module tt_um_Coline3003_spect_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire \clknet_leaf_0_top1.acquisition_clk ;
 wire \top1.PISO_ch1 ;
 wire \top1.PISO_time ;
 wire \top1.SL_ch ;
 wire \top1.SL_time ;
 wire \top1.acquisition_clk ;
 wire \top1.addr_in[0] ;
 wire \top1.addr_in[1] ;
 wire \top1.addr_in[2] ;
 wire \top1.addr_in[3] ;
 wire \top1.addr_in[4] ;
 wire \top1.addr_in[5] ;
 wire \top1.addr_in[6] ;
 wire \top1.addr_in[7] ;
 wire \top1.addr_in[8] ;
 wire \top1.addr_out[0] ;
 wire \top1.addr_out[1] ;
 wire \top1.addr_out[2] ;
 wire \top1.addr_out[3] ;
 wire \top1.addr_out[4] ;
 wire \top1.addr_out[5] ;
 wire \top1.addr_out[6] ;
 wire \top1.addr_out[7] ;
 wire \top1.addr_out[8] ;
 wire \top1.bank0_full ;
 wire \top1.bank1_full ;
 wire \top1.event_time[0] ;
 wire \top1.event_time[10] ;
 wire \top1.event_time[11] ;
 wire \top1.event_time[12] ;
 wire \top1.event_time[13] ;
 wire \top1.event_time[14] ;
 wire \top1.event_time[15] ;
 wire \top1.event_time[16] ;
 wire \top1.event_time[17] ;
 wire \top1.event_time[18] ;
 wire \top1.event_time[19] ;
 wire \top1.event_time[1] ;
 wire \top1.event_time[20] ;
 wire \top1.event_time[21] ;
 wire \top1.event_time[22] ;
 wire \top1.event_time[23] ;
 wire \top1.event_time[24] ;
 wire \top1.event_time[25] ;
 wire \top1.event_time[26] ;
 wire \top1.event_time[27] ;
 wire \top1.event_time[28] ;
 wire \top1.event_time[29] ;
 wire \top1.event_time[2] ;
 wire \top1.event_time[30] ;
 wire \top1.event_time[31] ;
 wire \top1.event_time[3] ;
 wire \top1.event_time[4] ;
 wire \top1.event_time[5] ;
 wire \top1.event_time[6] ;
 wire \top1.event_time[7] ;
 wire \top1.event_time[8] ;
 wire \top1.event_time[9] ;
 wire \top1.event_time_out[0] ;
 wire \top1.event_time_out[10] ;
 wire \top1.event_time_out[11] ;
 wire \top1.event_time_out[12] ;
 wire \top1.event_time_out[13] ;
 wire \top1.event_time_out[14] ;
 wire \top1.event_time_out[15] ;
 wire \top1.event_time_out[16] ;
 wire \top1.event_time_out[17] ;
 wire \top1.event_time_out[18] ;
 wire \top1.event_time_out[19] ;
 wire \top1.event_time_out[1] ;
 wire \top1.event_time_out[20] ;
 wire \top1.event_time_out[21] ;
 wire \top1.event_time_out[22] ;
 wire \top1.event_time_out[23] ;
 wire \top1.event_time_out[24] ;
 wire \top1.event_time_out[25] ;
 wire \top1.event_time_out[26] ;
 wire \top1.event_time_out[27] ;
 wire \top1.event_time_out[28] ;
 wire \top1.event_time_out[29] ;
 wire \top1.event_time_out[2] ;
 wire \top1.event_time_out[30] ;
 wire \top1.event_time_out[31] ;
 wire \top1.event_time_out[3] ;
 wire \top1.event_time_out[4] ;
 wire \top1.event_time_out[5] ;
 wire \top1.event_time_out[6] ;
 wire \top1.event_time_out[7] ;
 wire \top1.event_time_out[8] ;
 wire \top1.event_time_out[9] ;
 wire \top1.fsm.clk ;
 wire \top1.fsm.cpt[0] ;
 wire \top1.fsm.cpt[1] ;
 wire \top1.fsm.cpt[2] ;
 wire \top1.fsm.cpt[3] ;
 wire \top1.fsm.cpt[4] ;
 wire \top1.fsm.idx_final[0] ;
 wire \top1.fsm.idx_final[1] ;
 wire \top1.fsm.idx_final[2] ;
 wire \top1.fsm.idx_final[3] ;
 wire \top1.fsm.idx_final[4] ;
 wire \top1.fsm.idx_final[5] ;
 wire \top1.fsm.idx_final[6] ;
 wire \top1.fsm.idx_final[7] ;
 wire \top1.fsm.memorization_completed ;
 wire \top1.fsm.re ;
 wire \top1.fsm.reg_idx_final[0] ;
 wire \top1.fsm.reg_idx_final[1] ;
 wire \top1.fsm.reg_idx_final[2] ;
 wire \top1.fsm.reg_idx_final[3] ;
 wire \top1.fsm.reg_idx_final[4] ;
 wire \top1.fsm.reg_idx_final[5] ;
 wire \top1.fsm.reg_idx_final[6] ;
 wire \top1.fsm.reg_idx_final[7] ;
 wire \top1.fsm.sending_data ;
 wire \top1.fsm.sending_pending ;
 wire \top1.fsm.serial_readout ;
 wire \top1.fsm.signal_duration ;
 wire \top1.fsm.state_next[0] ;
 wire \top1.fsm.state_next[1] ;
 wire \top1.fsm.state_next[2] ;
 wire \top1.fsm.state_reg[0] ;
 wire \top1.fsm.state_reg[1] ;
 wire \top1.fsm.state_reg[2] ;
 wire \top1.mem_ctl.signal_detected ;
 wire \top1.mem_ctl.state_reg[0] ;
 wire \top1.mem_ctl.state_reg[1] ;
 wire \top1.memory1.data_out[0] ;
 wire \top1.memory1.data_out[1] ;
 wire \top1.memory1.data_out[2] ;
 wire \top1.memory1.mem1[0][0] ;
 wire \top1.memory1.mem1[0][1] ;
 wire \top1.memory1.mem1[0][2] ;
 wire \top1.memory1.mem1[100][0] ;
 wire \top1.memory1.mem1[100][1] ;
 wire \top1.memory1.mem1[100][2] ;
 wire \top1.memory1.mem1[101][0] ;
 wire \top1.memory1.mem1[101][1] ;
 wire \top1.memory1.mem1[101][2] ;
 wire \top1.memory1.mem1[102][0] ;
 wire \top1.memory1.mem1[102][1] ;
 wire \top1.memory1.mem1[102][2] ;
 wire \top1.memory1.mem1[103][0] ;
 wire \top1.memory1.mem1[103][1] ;
 wire \top1.memory1.mem1[103][2] ;
 wire \top1.memory1.mem1[104][0] ;
 wire \top1.memory1.mem1[104][1] ;
 wire \top1.memory1.mem1[104][2] ;
 wire \top1.memory1.mem1[105][0] ;
 wire \top1.memory1.mem1[105][1] ;
 wire \top1.memory1.mem1[105][2] ;
 wire \top1.memory1.mem1[106][0] ;
 wire \top1.memory1.mem1[106][1] ;
 wire \top1.memory1.mem1[106][2] ;
 wire \top1.memory1.mem1[107][0] ;
 wire \top1.memory1.mem1[107][1] ;
 wire \top1.memory1.mem1[107][2] ;
 wire \top1.memory1.mem1[108][0] ;
 wire \top1.memory1.mem1[108][1] ;
 wire \top1.memory1.mem1[108][2] ;
 wire \top1.memory1.mem1[109][0] ;
 wire \top1.memory1.mem1[109][1] ;
 wire \top1.memory1.mem1[109][2] ;
 wire \top1.memory1.mem1[10][0] ;
 wire \top1.memory1.mem1[10][1] ;
 wire \top1.memory1.mem1[10][2] ;
 wire \top1.memory1.mem1[110][0] ;
 wire \top1.memory1.mem1[110][1] ;
 wire \top1.memory1.mem1[110][2] ;
 wire \top1.memory1.mem1[111][0] ;
 wire \top1.memory1.mem1[111][1] ;
 wire \top1.memory1.mem1[111][2] ;
 wire \top1.memory1.mem1[112][0] ;
 wire \top1.memory1.mem1[112][1] ;
 wire \top1.memory1.mem1[112][2] ;
 wire \top1.memory1.mem1[113][0] ;
 wire \top1.memory1.mem1[113][1] ;
 wire \top1.memory1.mem1[113][2] ;
 wire \top1.memory1.mem1[114][0] ;
 wire \top1.memory1.mem1[114][1] ;
 wire \top1.memory1.mem1[114][2] ;
 wire \top1.memory1.mem1[115][0] ;
 wire \top1.memory1.mem1[115][1] ;
 wire \top1.memory1.mem1[115][2] ;
 wire \top1.memory1.mem1[116][0] ;
 wire \top1.memory1.mem1[116][1] ;
 wire \top1.memory1.mem1[116][2] ;
 wire \top1.memory1.mem1[117][0] ;
 wire \top1.memory1.mem1[117][1] ;
 wire \top1.memory1.mem1[117][2] ;
 wire \top1.memory1.mem1[118][0] ;
 wire \top1.memory1.mem1[118][1] ;
 wire \top1.memory1.mem1[118][2] ;
 wire \top1.memory1.mem1[119][0] ;
 wire \top1.memory1.mem1[119][1] ;
 wire \top1.memory1.mem1[119][2] ;
 wire \top1.memory1.mem1[11][0] ;
 wire \top1.memory1.mem1[11][1] ;
 wire \top1.memory1.mem1[11][2] ;
 wire \top1.memory1.mem1[120][0] ;
 wire \top1.memory1.mem1[120][1] ;
 wire \top1.memory1.mem1[120][2] ;
 wire \top1.memory1.mem1[121][0] ;
 wire \top1.memory1.mem1[121][1] ;
 wire \top1.memory1.mem1[121][2] ;
 wire \top1.memory1.mem1[122][0] ;
 wire \top1.memory1.mem1[122][1] ;
 wire \top1.memory1.mem1[122][2] ;
 wire \top1.memory1.mem1[123][0] ;
 wire \top1.memory1.mem1[123][1] ;
 wire \top1.memory1.mem1[123][2] ;
 wire \top1.memory1.mem1[124][0] ;
 wire \top1.memory1.mem1[124][1] ;
 wire \top1.memory1.mem1[124][2] ;
 wire \top1.memory1.mem1[125][0] ;
 wire \top1.memory1.mem1[125][1] ;
 wire \top1.memory1.mem1[125][2] ;
 wire \top1.memory1.mem1[126][0] ;
 wire \top1.memory1.mem1[126][1] ;
 wire \top1.memory1.mem1[126][2] ;
 wire \top1.memory1.mem1[127][0] ;
 wire \top1.memory1.mem1[127][1] ;
 wire \top1.memory1.mem1[127][2] ;
 wire \top1.memory1.mem1[128][0] ;
 wire \top1.memory1.mem1[128][1] ;
 wire \top1.memory1.mem1[128][2] ;
 wire \top1.memory1.mem1[129][0] ;
 wire \top1.memory1.mem1[129][1] ;
 wire \top1.memory1.mem1[129][2] ;
 wire \top1.memory1.mem1[12][0] ;
 wire \top1.memory1.mem1[12][1] ;
 wire \top1.memory1.mem1[12][2] ;
 wire \top1.memory1.mem1[130][0] ;
 wire \top1.memory1.mem1[130][1] ;
 wire \top1.memory1.mem1[130][2] ;
 wire \top1.memory1.mem1[131][0] ;
 wire \top1.memory1.mem1[131][1] ;
 wire \top1.memory1.mem1[131][2] ;
 wire \top1.memory1.mem1[132][0] ;
 wire \top1.memory1.mem1[132][1] ;
 wire \top1.memory1.mem1[132][2] ;
 wire \top1.memory1.mem1[133][0] ;
 wire \top1.memory1.mem1[133][1] ;
 wire \top1.memory1.mem1[133][2] ;
 wire \top1.memory1.mem1[134][0] ;
 wire \top1.memory1.mem1[134][1] ;
 wire \top1.memory1.mem1[134][2] ;
 wire \top1.memory1.mem1[135][0] ;
 wire \top1.memory1.mem1[135][1] ;
 wire \top1.memory1.mem1[135][2] ;
 wire \top1.memory1.mem1[136][0] ;
 wire \top1.memory1.mem1[136][1] ;
 wire \top1.memory1.mem1[136][2] ;
 wire \top1.memory1.mem1[137][0] ;
 wire \top1.memory1.mem1[137][1] ;
 wire \top1.memory1.mem1[137][2] ;
 wire \top1.memory1.mem1[138][0] ;
 wire \top1.memory1.mem1[138][1] ;
 wire \top1.memory1.mem1[138][2] ;
 wire \top1.memory1.mem1[139][0] ;
 wire \top1.memory1.mem1[139][1] ;
 wire \top1.memory1.mem1[139][2] ;
 wire \top1.memory1.mem1[13][0] ;
 wire \top1.memory1.mem1[13][1] ;
 wire \top1.memory1.mem1[13][2] ;
 wire \top1.memory1.mem1[140][0] ;
 wire \top1.memory1.mem1[140][1] ;
 wire \top1.memory1.mem1[140][2] ;
 wire \top1.memory1.mem1[141][0] ;
 wire \top1.memory1.mem1[141][1] ;
 wire \top1.memory1.mem1[141][2] ;
 wire \top1.memory1.mem1[142][0] ;
 wire \top1.memory1.mem1[142][1] ;
 wire \top1.memory1.mem1[142][2] ;
 wire \top1.memory1.mem1[143][0] ;
 wire \top1.memory1.mem1[143][1] ;
 wire \top1.memory1.mem1[143][2] ;
 wire \top1.memory1.mem1[144][0] ;
 wire \top1.memory1.mem1[144][1] ;
 wire \top1.memory1.mem1[144][2] ;
 wire \top1.memory1.mem1[145][0] ;
 wire \top1.memory1.mem1[145][1] ;
 wire \top1.memory1.mem1[145][2] ;
 wire \top1.memory1.mem1[146][0] ;
 wire \top1.memory1.mem1[146][1] ;
 wire \top1.memory1.mem1[146][2] ;
 wire \top1.memory1.mem1[147][0] ;
 wire \top1.memory1.mem1[147][1] ;
 wire \top1.memory1.mem1[147][2] ;
 wire \top1.memory1.mem1[148][0] ;
 wire \top1.memory1.mem1[148][1] ;
 wire \top1.memory1.mem1[148][2] ;
 wire \top1.memory1.mem1[149][0] ;
 wire \top1.memory1.mem1[149][1] ;
 wire \top1.memory1.mem1[149][2] ;
 wire \top1.memory1.mem1[14][0] ;
 wire \top1.memory1.mem1[14][1] ;
 wire \top1.memory1.mem1[14][2] ;
 wire \top1.memory1.mem1[150][0] ;
 wire \top1.memory1.mem1[150][1] ;
 wire \top1.memory1.mem1[150][2] ;
 wire \top1.memory1.mem1[151][0] ;
 wire \top1.memory1.mem1[151][1] ;
 wire \top1.memory1.mem1[151][2] ;
 wire \top1.memory1.mem1[152][0] ;
 wire \top1.memory1.mem1[152][1] ;
 wire \top1.memory1.mem1[152][2] ;
 wire \top1.memory1.mem1[153][0] ;
 wire \top1.memory1.mem1[153][1] ;
 wire \top1.memory1.mem1[153][2] ;
 wire \top1.memory1.mem1[154][0] ;
 wire \top1.memory1.mem1[154][1] ;
 wire \top1.memory1.mem1[154][2] ;
 wire \top1.memory1.mem1[155][0] ;
 wire \top1.memory1.mem1[155][1] ;
 wire \top1.memory1.mem1[155][2] ;
 wire \top1.memory1.mem1[156][0] ;
 wire \top1.memory1.mem1[156][1] ;
 wire \top1.memory1.mem1[156][2] ;
 wire \top1.memory1.mem1[157][0] ;
 wire \top1.memory1.mem1[157][1] ;
 wire \top1.memory1.mem1[157][2] ;
 wire \top1.memory1.mem1[158][0] ;
 wire \top1.memory1.mem1[158][1] ;
 wire \top1.memory1.mem1[158][2] ;
 wire \top1.memory1.mem1[159][0] ;
 wire \top1.memory1.mem1[159][1] ;
 wire \top1.memory1.mem1[159][2] ;
 wire \top1.memory1.mem1[15][0] ;
 wire \top1.memory1.mem1[15][1] ;
 wire \top1.memory1.mem1[15][2] ;
 wire \top1.memory1.mem1[160][0] ;
 wire \top1.memory1.mem1[160][1] ;
 wire \top1.memory1.mem1[160][2] ;
 wire \top1.memory1.mem1[161][0] ;
 wire \top1.memory1.mem1[161][1] ;
 wire \top1.memory1.mem1[161][2] ;
 wire \top1.memory1.mem1[162][0] ;
 wire \top1.memory1.mem1[162][1] ;
 wire \top1.memory1.mem1[162][2] ;
 wire \top1.memory1.mem1[163][0] ;
 wire \top1.memory1.mem1[163][1] ;
 wire \top1.memory1.mem1[163][2] ;
 wire \top1.memory1.mem1[164][0] ;
 wire \top1.memory1.mem1[164][1] ;
 wire \top1.memory1.mem1[164][2] ;
 wire \top1.memory1.mem1[165][0] ;
 wire \top1.memory1.mem1[165][1] ;
 wire \top1.memory1.mem1[165][2] ;
 wire \top1.memory1.mem1[166][0] ;
 wire \top1.memory1.mem1[166][1] ;
 wire \top1.memory1.mem1[166][2] ;
 wire \top1.memory1.mem1[167][0] ;
 wire \top1.memory1.mem1[167][1] ;
 wire \top1.memory1.mem1[167][2] ;
 wire \top1.memory1.mem1[168][0] ;
 wire \top1.memory1.mem1[168][1] ;
 wire \top1.memory1.mem1[168][2] ;
 wire \top1.memory1.mem1[169][0] ;
 wire \top1.memory1.mem1[169][1] ;
 wire \top1.memory1.mem1[169][2] ;
 wire \top1.memory1.mem1[16][0] ;
 wire \top1.memory1.mem1[16][1] ;
 wire \top1.memory1.mem1[16][2] ;
 wire \top1.memory1.mem1[170][0] ;
 wire \top1.memory1.mem1[170][1] ;
 wire \top1.memory1.mem1[170][2] ;
 wire \top1.memory1.mem1[171][0] ;
 wire \top1.memory1.mem1[171][1] ;
 wire \top1.memory1.mem1[171][2] ;
 wire \top1.memory1.mem1[172][0] ;
 wire \top1.memory1.mem1[172][1] ;
 wire \top1.memory1.mem1[172][2] ;
 wire \top1.memory1.mem1[173][0] ;
 wire \top1.memory1.mem1[173][1] ;
 wire \top1.memory1.mem1[173][2] ;
 wire \top1.memory1.mem1[174][0] ;
 wire \top1.memory1.mem1[174][1] ;
 wire \top1.memory1.mem1[174][2] ;
 wire \top1.memory1.mem1[175][0] ;
 wire \top1.memory1.mem1[175][1] ;
 wire \top1.memory1.mem1[175][2] ;
 wire \top1.memory1.mem1[176][0] ;
 wire \top1.memory1.mem1[176][1] ;
 wire \top1.memory1.mem1[176][2] ;
 wire \top1.memory1.mem1[177][0] ;
 wire \top1.memory1.mem1[177][1] ;
 wire \top1.memory1.mem1[177][2] ;
 wire \top1.memory1.mem1[178][0] ;
 wire \top1.memory1.mem1[178][1] ;
 wire \top1.memory1.mem1[178][2] ;
 wire \top1.memory1.mem1[179][0] ;
 wire \top1.memory1.mem1[179][1] ;
 wire \top1.memory1.mem1[179][2] ;
 wire \top1.memory1.mem1[17][0] ;
 wire \top1.memory1.mem1[17][1] ;
 wire \top1.memory1.mem1[17][2] ;
 wire \top1.memory1.mem1[180][0] ;
 wire \top1.memory1.mem1[180][1] ;
 wire \top1.memory1.mem1[180][2] ;
 wire \top1.memory1.mem1[181][0] ;
 wire \top1.memory1.mem1[181][1] ;
 wire \top1.memory1.mem1[181][2] ;
 wire \top1.memory1.mem1[182][0] ;
 wire \top1.memory1.mem1[182][1] ;
 wire \top1.memory1.mem1[182][2] ;
 wire \top1.memory1.mem1[183][0] ;
 wire \top1.memory1.mem1[183][1] ;
 wire \top1.memory1.mem1[183][2] ;
 wire \top1.memory1.mem1[184][0] ;
 wire \top1.memory1.mem1[184][1] ;
 wire \top1.memory1.mem1[184][2] ;
 wire \top1.memory1.mem1[185][0] ;
 wire \top1.memory1.mem1[185][1] ;
 wire \top1.memory1.mem1[185][2] ;
 wire \top1.memory1.mem1[186][0] ;
 wire \top1.memory1.mem1[186][1] ;
 wire \top1.memory1.mem1[186][2] ;
 wire \top1.memory1.mem1[187][0] ;
 wire \top1.memory1.mem1[187][1] ;
 wire \top1.memory1.mem1[187][2] ;
 wire \top1.memory1.mem1[188][0] ;
 wire \top1.memory1.mem1[188][1] ;
 wire \top1.memory1.mem1[188][2] ;
 wire \top1.memory1.mem1[189][0] ;
 wire \top1.memory1.mem1[189][1] ;
 wire \top1.memory1.mem1[189][2] ;
 wire \top1.memory1.mem1[18][0] ;
 wire \top1.memory1.mem1[18][1] ;
 wire \top1.memory1.mem1[18][2] ;
 wire \top1.memory1.mem1[190][0] ;
 wire \top1.memory1.mem1[190][1] ;
 wire \top1.memory1.mem1[190][2] ;
 wire \top1.memory1.mem1[191][0] ;
 wire \top1.memory1.mem1[191][1] ;
 wire \top1.memory1.mem1[191][2] ;
 wire \top1.memory1.mem1[192][0] ;
 wire \top1.memory1.mem1[192][1] ;
 wire \top1.memory1.mem1[192][2] ;
 wire \top1.memory1.mem1[193][0] ;
 wire \top1.memory1.mem1[193][1] ;
 wire \top1.memory1.mem1[193][2] ;
 wire \top1.memory1.mem1[194][0] ;
 wire \top1.memory1.mem1[194][1] ;
 wire \top1.memory1.mem1[194][2] ;
 wire \top1.memory1.mem1[195][0] ;
 wire \top1.memory1.mem1[195][1] ;
 wire \top1.memory1.mem1[195][2] ;
 wire \top1.memory1.mem1[196][0] ;
 wire \top1.memory1.mem1[196][1] ;
 wire \top1.memory1.mem1[196][2] ;
 wire \top1.memory1.mem1[197][0] ;
 wire \top1.memory1.mem1[197][1] ;
 wire \top1.memory1.mem1[197][2] ;
 wire \top1.memory1.mem1[198][0] ;
 wire \top1.memory1.mem1[198][1] ;
 wire \top1.memory1.mem1[198][2] ;
 wire \top1.memory1.mem1[199][0] ;
 wire \top1.memory1.mem1[199][1] ;
 wire \top1.memory1.mem1[199][2] ;
 wire \top1.memory1.mem1[19][0] ;
 wire \top1.memory1.mem1[19][1] ;
 wire \top1.memory1.mem1[19][2] ;
 wire \top1.memory1.mem1[1][0] ;
 wire \top1.memory1.mem1[1][1] ;
 wire \top1.memory1.mem1[1][2] ;
 wire \top1.memory1.mem1[20][0] ;
 wire \top1.memory1.mem1[20][1] ;
 wire \top1.memory1.mem1[20][2] ;
 wire \top1.memory1.mem1[21][0] ;
 wire \top1.memory1.mem1[21][1] ;
 wire \top1.memory1.mem1[21][2] ;
 wire \top1.memory1.mem1[22][0] ;
 wire \top1.memory1.mem1[22][1] ;
 wire \top1.memory1.mem1[22][2] ;
 wire \top1.memory1.mem1[23][0] ;
 wire \top1.memory1.mem1[23][1] ;
 wire \top1.memory1.mem1[23][2] ;
 wire \top1.memory1.mem1[24][0] ;
 wire \top1.memory1.mem1[24][1] ;
 wire \top1.memory1.mem1[24][2] ;
 wire \top1.memory1.mem1[25][0] ;
 wire \top1.memory1.mem1[25][1] ;
 wire \top1.memory1.mem1[25][2] ;
 wire \top1.memory1.mem1[26][0] ;
 wire \top1.memory1.mem1[26][1] ;
 wire \top1.memory1.mem1[26][2] ;
 wire \top1.memory1.mem1[27][0] ;
 wire \top1.memory1.mem1[27][1] ;
 wire \top1.memory1.mem1[27][2] ;
 wire \top1.memory1.mem1[28][0] ;
 wire \top1.memory1.mem1[28][1] ;
 wire \top1.memory1.mem1[28][2] ;
 wire \top1.memory1.mem1[29][0] ;
 wire \top1.memory1.mem1[29][1] ;
 wire \top1.memory1.mem1[29][2] ;
 wire \top1.memory1.mem1[2][0] ;
 wire \top1.memory1.mem1[2][1] ;
 wire \top1.memory1.mem1[2][2] ;
 wire \top1.memory1.mem1[30][0] ;
 wire \top1.memory1.mem1[30][1] ;
 wire \top1.memory1.mem1[30][2] ;
 wire \top1.memory1.mem1[31][0] ;
 wire \top1.memory1.mem1[31][1] ;
 wire \top1.memory1.mem1[31][2] ;
 wire \top1.memory1.mem1[32][0] ;
 wire \top1.memory1.mem1[32][1] ;
 wire \top1.memory1.mem1[32][2] ;
 wire \top1.memory1.mem1[33][0] ;
 wire \top1.memory1.mem1[33][1] ;
 wire \top1.memory1.mem1[33][2] ;
 wire \top1.memory1.mem1[34][0] ;
 wire \top1.memory1.mem1[34][1] ;
 wire \top1.memory1.mem1[34][2] ;
 wire \top1.memory1.mem1[35][0] ;
 wire \top1.memory1.mem1[35][1] ;
 wire \top1.memory1.mem1[35][2] ;
 wire \top1.memory1.mem1[36][0] ;
 wire \top1.memory1.mem1[36][1] ;
 wire \top1.memory1.mem1[36][2] ;
 wire \top1.memory1.mem1[37][0] ;
 wire \top1.memory1.mem1[37][1] ;
 wire \top1.memory1.mem1[37][2] ;
 wire \top1.memory1.mem1[38][0] ;
 wire \top1.memory1.mem1[38][1] ;
 wire \top1.memory1.mem1[38][2] ;
 wire \top1.memory1.mem1[39][0] ;
 wire \top1.memory1.mem1[39][1] ;
 wire \top1.memory1.mem1[39][2] ;
 wire \top1.memory1.mem1[3][0] ;
 wire \top1.memory1.mem1[3][1] ;
 wire \top1.memory1.mem1[3][2] ;
 wire \top1.memory1.mem1[40][0] ;
 wire \top1.memory1.mem1[40][1] ;
 wire \top1.memory1.mem1[40][2] ;
 wire \top1.memory1.mem1[41][0] ;
 wire \top1.memory1.mem1[41][1] ;
 wire \top1.memory1.mem1[41][2] ;
 wire \top1.memory1.mem1[42][0] ;
 wire \top1.memory1.mem1[42][1] ;
 wire \top1.memory1.mem1[42][2] ;
 wire \top1.memory1.mem1[43][0] ;
 wire \top1.memory1.mem1[43][1] ;
 wire \top1.memory1.mem1[43][2] ;
 wire \top1.memory1.mem1[44][0] ;
 wire \top1.memory1.mem1[44][1] ;
 wire \top1.memory1.mem1[44][2] ;
 wire \top1.memory1.mem1[45][0] ;
 wire \top1.memory1.mem1[45][1] ;
 wire \top1.memory1.mem1[45][2] ;
 wire \top1.memory1.mem1[46][0] ;
 wire \top1.memory1.mem1[46][1] ;
 wire \top1.memory1.mem1[46][2] ;
 wire \top1.memory1.mem1[47][0] ;
 wire \top1.memory1.mem1[47][1] ;
 wire \top1.memory1.mem1[47][2] ;
 wire \top1.memory1.mem1[48][0] ;
 wire \top1.memory1.mem1[48][1] ;
 wire \top1.memory1.mem1[48][2] ;
 wire \top1.memory1.mem1[49][0] ;
 wire \top1.memory1.mem1[49][1] ;
 wire \top1.memory1.mem1[49][2] ;
 wire \top1.memory1.mem1[4][0] ;
 wire \top1.memory1.mem1[4][1] ;
 wire \top1.memory1.mem1[4][2] ;
 wire \top1.memory1.mem1[50][0] ;
 wire \top1.memory1.mem1[50][1] ;
 wire \top1.memory1.mem1[50][2] ;
 wire \top1.memory1.mem1[51][0] ;
 wire \top1.memory1.mem1[51][1] ;
 wire \top1.memory1.mem1[51][2] ;
 wire \top1.memory1.mem1[52][0] ;
 wire \top1.memory1.mem1[52][1] ;
 wire \top1.memory1.mem1[52][2] ;
 wire \top1.memory1.mem1[53][0] ;
 wire \top1.memory1.mem1[53][1] ;
 wire \top1.memory1.mem1[53][2] ;
 wire \top1.memory1.mem1[54][0] ;
 wire \top1.memory1.mem1[54][1] ;
 wire \top1.memory1.mem1[54][2] ;
 wire \top1.memory1.mem1[55][0] ;
 wire \top1.memory1.mem1[55][1] ;
 wire \top1.memory1.mem1[55][2] ;
 wire \top1.memory1.mem1[56][0] ;
 wire \top1.memory1.mem1[56][1] ;
 wire \top1.memory1.mem1[56][2] ;
 wire \top1.memory1.mem1[57][0] ;
 wire \top1.memory1.mem1[57][1] ;
 wire \top1.memory1.mem1[57][2] ;
 wire \top1.memory1.mem1[58][0] ;
 wire \top1.memory1.mem1[58][1] ;
 wire \top1.memory1.mem1[58][2] ;
 wire \top1.memory1.mem1[59][0] ;
 wire \top1.memory1.mem1[59][1] ;
 wire \top1.memory1.mem1[59][2] ;
 wire \top1.memory1.mem1[5][0] ;
 wire \top1.memory1.mem1[5][1] ;
 wire \top1.memory1.mem1[5][2] ;
 wire \top1.memory1.mem1[60][0] ;
 wire \top1.memory1.mem1[60][1] ;
 wire \top1.memory1.mem1[60][2] ;
 wire \top1.memory1.mem1[61][0] ;
 wire \top1.memory1.mem1[61][1] ;
 wire \top1.memory1.mem1[61][2] ;
 wire \top1.memory1.mem1[62][0] ;
 wire \top1.memory1.mem1[62][1] ;
 wire \top1.memory1.mem1[62][2] ;
 wire \top1.memory1.mem1[63][0] ;
 wire \top1.memory1.mem1[63][1] ;
 wire \top1.memory1.mem1[63][2] ;
 wire \top1.memory1.mem1[64][0] ;
 wire \top1.memory1.mem1[64][1] ;
 wire \top1.memory1.mem1[64][2] ;
 wire \top1.memory1.mem1[65][0] ;
 wire \top1.memory1.mem1[65][1] ;
 wire \top1.memory1.mem1[65][2] ;
 wire \top1.memory1.mem1[66][0] ;
 wire \top1.memory1.mem1[66][1] ;
 wire \top1.memory1.mem1[66][2] ;
 wire \top1.memory1.mem1[67][0] ;
 wire \top1.memory1.mem1[67][1] ;
 wire \top1.memory1.mem1[67][2] ;
 wire \top1.memory1.mem1[68][0] ;
 wire \top1.memory1.mem1[68][1] ;
 wire \top1.memory1.mem1[68][2] ;
 wire \top1.memory1.mem1[69][0] ;
 wire \top1.memory1.mem1[69][1] ;
 wire \top1.memory1.mem1[69][2] ;
 wire \top1.memory1.mem1[6][0] ;
 wire \top1.memory1.mem1[6][1] ;
 wire \top1.memory1.mem1[6][2] ;
 wire \top1.memory1.mem1[70][0] ;
 wire \top1.memory1.mem1[70][1] ;
 wire \top1.memory1.mem1[70][2] ;
 wire \top1.memory1.mem1[71][0] ;
 wire \top1.memory1.mem1[71][1] ;
 wire \top1.memory1.mem1[71][2] ;
 wire \top1.memory1.mem1[72][0] ;
 wire \top1.memory1.mem1[72][1] ;
 wire \top1.memory1.mem1[72][2] ;
 wire \top1.memory1.mem1[73][0] ;
 wire \top1.memory1.mem1[73][1] ;
 wire \top1.memory1.mem1[73][2] ;
 wire \top1.memory1.mem1[74][0] ;
 wire \top1.memory1.mem1[74][1] ;
 wire \top1.memory1.mem1[74][2] ;
 wire \top1.memory1.mem1[75][0] ;
 wire \top1.memory1.mem1[75][1] ;
 wire \top1.memory1.mem1[75][2] ;
 wire \top1.memory1.mem1[76][0] ;
 wire \top1.memory1.mem1[76][1] ;
 wire \top1.memory1.mem1[76][2] ;
 wire \top1.memory1.mem1[77][0] ;
 wire \top1.memory1.mem1[77][1] ;
 wire \top1.memory1.mem1[77][2] ;
 wire \top1.memory1.mem1[78][0] ;
 wire \top1.memory1.mem1[78][1] ;
 wire \top1.memory1.mem1[78][2] ;
 wire \top1.memory1.mem1[79][0] ;
 wire \top1.memory1.mem1[79][1] ;
 wire \top1.memory1.mem1[79][2] ;
 wire \top1.memory1.mem1[7][0] ;
 wire \top1.memory1.mem1[7][1] ;
 wire \top1.memory1.mem1[7][2] ;
 wire \top1.memory1.mem1[80][0] ;
 wire \top1.memory1.mem1[80][1] ;
 wire \top1.memory1.mem1[80][2] ;
 wire \top1.memory1.mem1[81][0] ;
 wire \top1.memory1.mem1[81][1] ;
 wire \top1.memory1.mem1[81][2] ;
 wire \top1.memory1.mem1[82][0] ;
 wire \top1.memory1.mem1[82][1] ;
 wire \top1.memory1.mem1[82][2] ;
 wire \top1.memory1.mem1[83][0] ;
 wire \top1.memory1.mem1[83][1] ;
 wire \top1.memory1.mem1[83][2] ;
 wire \top1.memory1.mem1[84][0] ;
 wire \top1.memory1.mem1[84][1] ;
 wire \top1.memory1.mem1[84][2] ;
 wire \top1.memory1.mem1[85][0] ;
 wire \top1.memory1.mem1[85][1] ;
 wire \top1.memory1.mem1[85][2] ;
 wire \top1.memory1.mem1[86][0] ;
 wire \top1.memory1.mem1[86][1] ;
 wire \top1.memory1.mem1[86][2] ;
 wire \top1.memory1.mem1[87][0] ;
 wire \top1.memory1.mem1[87][1] ;
 wire \top1.memory1.mem1[87][2] ;
 wire \top1.memory1.mem1[88][0] ;
 wire \top1.memory1.mem1[88][1] ;
 wire \top1.memory1.mem1[88][2] ;
 wire \top1.memory1.mem1[89][0] ;
 wire \top1.memory1.mem1[89][1] ;
 wire \top1.memory1.mem1[89][2] ;
 wire \top1.memory1.mem1[8][0] ;
 wire \top1.memory1.mem1[8][1] ;
 wire \top1.memory1.mem1[8][2] ;
 wire \top1.memory1.mem1[90][0] ;
 wire \top1.memory1.mem1[90][1] ;
 wire \top1.memory1.mem1[90][2] ;
 wire \top1.memory1.mem1[91][0] ;
 wire \top1.memory1.mem1[91][1] ;
 wire \top1.memory1.mem1[91][2] ;
 wire \top1.memory1.mem1[92][0] ;
 wire \top1.memory1.mem1[92][1] ;
 wire \top1.memory1.mem1[92][2] ;
 wire \top1.memory1.mem1[93][0] ;
 wire \top1.memory1.mem1[93][1] ;
 wire \top1.memory1.mem1[93][2] ;
 wire \top1.memory1.mem1[94][0] ;
 wire \top1.memory1.mem1[94][1] ;
 wire \top1.memory1.mem1[94][2] ;
 wire \top1.memory1.mem1[95][0] ;
 wire \top1.memory1.mem1[95][1] ;
 wire \top1.memory1.mem1[95][2] ;
 wire \top1.memory1.mem1[96][0] ;
 wire \top1.memory1.mem1[96][1] ;
 wire \top1.memory1.mem1[96][2] ;
 wire \top1.memory1.mem1[97][0] ;
 wire \top1.memory1.mem1[97][1] ;
 wire \top1.memory1.mem1[97][2] ;
 wire \top1.memory1.mem1[98][0] ;
 wire \top1.memory1.mem1[98][1] ;
 wire \top1.memory1.mem1[98][2] ;
 wire \top1.memory1.mem1[99][0] ;
 wire \top1.memory1.mem1[99][1] ;
 wire \top1.memory1.mem1[99][2] ;
 wire \top1.memory1.mem1[9][0] ;
 wire \top1.memory1.mem1[9][1] ;
 wire \top1.memory1.mem1[9][2] ;
 wire \top1.memory1.mem2[0][0] ;
 wire \top1.memory1.mem2[0][1] ;
 wire \top1.memory1.mem2[0][2] ;
 wire \top1.memory1.mem2[100][0] ;
 wire \top1.memory1.mem2[100][1] ;
 wire \top1.memory1.mem2[100][2] ;
 wire \top1.memory1.mem2[101][0] ;
 wire \top1.memory1.mem2[101][1] ;
 wire \top1.memory1.mem2[101][2] ;
 wire \top1.memory1.mem2[102][0] ;
 wire \top1.memory1.mem2[102][1] ;
 wire \top1.memory1.mem2[102][2] ;
 wire \top1.memory1.mem2[103][0] ;
 wire \top1.memory1.mem2[103][1] ;
 wire \top1.memory1.mem2[103][2] ;
 wire \top1.memory1.mem2[104][0] ;
 wire \top1.memory1.mem2[104][1] ;
 wire \top1.memory1.mem2[104][2] ;
 wire \top1.memory1.mem2[105][0] ;
 wire \top1.memory1.mem2[105][1] ;
 wire \top1.memory1.mem2[105][2] ;
 wire \top1.memory1.mem2[106][0] ;
 wire \top1.memory1.mem2[106][1] ;
 wire \top1.memory1.mem2[106][2] ;
 wire \top1.memory1.mem2[107][0] ;
 wire \top1.memory1.mem2[107][1] ;
 wire \top1.memory1.mem2[107][2] ;
 wire \top1.memory1.mem2[108][0] ;
 wire \top1.memory1.mem2[108][1] ;
 wire \top1.memory1.mem2[108][2] ;
 wire \top1.memory1.mem2[109][0] ;
 wire \top1.memory1.mem2[109][1] ;
 wire \top1.memory1.mem2[109][2] ;
 wire \top1.memory1.mem2[10][0] ;
 wire \top1.memory1.mem2[10][1] ;
 wire \top1.memory1.mem2[10][2] ;
 wire \top1.memory1.mem2[110][0] ;
 wire \top1.memory1.mem2[110][1] ;
 wire \top1.memory1.mem2[110][2] ;
 wire \top1.memory1.mem2[111][0] ;
 wire \top1.memory1.mem2[111][1] ;
 wire \top1.memory1.mem2[111][2] ;
 wire \top1.memory1.mem2[112][0] ;
 wire \top1.memory1.mem2[112][1] ;
 wire \top1.memory1.mem2[112][2] ;
 wire \top1.memory1.mem2[113][0] ;
 wire \top1.memory1.mem2[113][1] ;
 wire \top1.memory1.mem2[113][2] ;
 wire \top1.memory1.mem2[114][0] ;
 wire \top1.memory1.mem2[114][1] ;
 wire \top1.memory1.mem2[114][2] ;
 wire \top1.memory1.mem2[115][0] ;
 wire \top1.memory1.mem2[115][1] ;
 wire \top1.memory1.mem2[115][2] ;
 wire \top1.memory1.mem2[116][0] ;
 wire \top1.memory1.mem2[116][1] ;
 wire \top1.memory1.mem2[116][2] ;
 wire \top1.memory1.mem2[117][0] ;
 wire \top1.memory1.mem2[117][1] ;
 wire \top1.memory1.mem2[117][2] ;
 wire \top1.memory1.mem2[118][0] ;
 wire \top1.memory1.mem2[118][1] ;
 wire \top1.memory1.mem2[118][2] ;
 wire \top1.memory1.mem2[119][0] ;
 wire \top1.memory1.mem2[119][1] ;
 wire \top1.memory1.mem2[119][2] ;
 wire \top1.memory1.mem2[11][0] ;
 wire \top1.memory1.mem2[11][1] ;
 wire \top1.memory1.mem2[11][2] ;
 wire \top1.memory1.mem2[120][0] ;
 wire \top1.memory1.mem2[120][1] ;
 wire \top1.memory1.mem2[120][2] ;
 wire \top1.memory1.mem2[121][0] ;
 wire \top1.memory1.mem2[121][1] ;
 wire \top1.memory1.mem2[121][2] ;
 wire \top1.memory1.mem2[122][0] ;
 wire \top1.memory1.mem2[122][1] ;
 wire \top1.memory1.mem2[122][2] ;
 wire \top1.memory1.mem2[123][0] ;
 wire \top1.memory1.mem2[123][1] ;
 wire \top1.memory1.mem2[123][2] ;
 wire \top1.memory1.mem2[124][0] ;
 wire \top1.memory1.mem2[124][1] ;
 wire \top1.memory1.mem2[124][2] ;
 wire \top1.memory1.mem2[125][0] ;
 wire \top1.memory1.mem2[125][1] ;
 wire \top1.memory1.mem2[125][2] ;
 wire \top1.memory1.mem2[126][0] ;
 wire \top1.memory1.mem2[126][1] ;
 wire \top1.memory1.mem2[126][2] ;
 wire \top1.memory1.mem2[127][0] ;
 wire \top1.memory1.mem2[127][1] ;
 wire \top1.memory1.mem2[127][2] ;
 wire \top1.memory1.mem2[128][0] ;
 wire \top1.memory1.mem2[128][1] ;
 wire \top1.memory1.mem2[128][2] ;
 wire \top1.memory1.mem2[129][0] ;
 wire \top1.memory1.mem2[129][1] ;
 wire \top1.memory1.mem2[129][2] ;
 wire \top1.memory1.mem2[12][0] ;
 wire \top1.memory1.mem2[12][1] ;
 wire \top1.memory1.mem2[12][2] ;
 wire \top1.memory1.mem2[130][0] ;
 wire \top1.memory1.mem2[130][1] ;
 wire \top1.memory1.mem2[130][2] ;
 wire \top1.memory1.mem2[131][0] ;
 wire \top1.memory1.mem2[131][1] ;
 wire \top1.memory1.mem2[131][2] ;
 wire \top1.memory1.mem2[132][0] ;
 wire \top1.memory1.mem2[132][1] ;
 wire \top1.memory1.mem2[132][2] ;
 wire \top1.memory1.mem2[133][0] ;
 wire \top1.memory1.mem2[133][1] ;
 wire \top1.memory1.mem2[133][2] ;
 wire \top1.memory1.mem2[134][0] ;
 wire \top1.memory1.mem2[134][1] ;
 wire \top1.memory1.mem2[134][2] ;
 wire \top1.memory1.mem2[135][0] ;
 wire \top1.memory1.mem2[135][1] ;
 wire \top1.memory1.mem2[135][2] ;
 wire \top1.memory1.mem2[136][0] ;
 wire \top1.memory1.mem2[136][1] ;
 wire \top1.memory1.mem2[136][2] ;
 wire \top1.memory1.mem2[137][0] ;
 wire \top1.memory1.mem2[137][1] ;
 wire \top1.memory1.mem2[137][2] ;
 wire \top1.memory1.mem2[138][0] ;
 wire \top1.memory1.mem2[138][1] ;
 wire \top1.memory1.mem2[138][2] ;
 wire \top1.memory1.mem2[139][0] ;
 wire \top1.memory1.mem2[139][1] ;
 wire \top1.memory1.mem2[139][2] ;
 wire \top1.memory1.mem2[13][0] ;
 wire \top1.memory1.mem2[13][1] ;
 wire \top1.memory1.mem2[13][2] ;
 wire \top1.memory1.mem2[140][0] ;
 wire \top1.memory1.mem2[140][1] ;
 wire \top1.memory1.mem2[140][2] ;
 wire \top1.memory1.mem2[141][0] ;
 wire \top1.memory1.mem2[141][1] ;
 wire \top1.memory1.mem2[141][2] ;
 wire \top1.memory1.mem2[142][0] ;
 wire \top1.memory1.mem2[142][1] ;
 wire \top1.memory1.mem2[142][2] ;
 wire \top1.memory1.mem2[143][0] ;
 wire \top1.memory1.mem2[143][1] ;
 wire \top1.memory1.mem2[143][2] ;
 wire \top1.memory1.mem2[144][0] ;
 wire \top1.memory1.mem2[144][1] ;
 wire \top1.memory1.mem2[144][2] ;
 wire \top1.memory1.mem2[145][0] ;
 wire \top1.memory1.mem2[145][1] ;
 wire \top1.memory1.mem2[145][2] ;
 wire \top1.memory1.mem2[146][0] ;
 wire \top1.memory1.mem2[146][1] ;
 wire \top1.memory1.mem2[146][2] ;
 wire \top1.memory1.mem2[147][0] ;
 wire \top1.memory1.mem2[147][1] ;
 wire \top1.memory1.mem2[147][2] ;
 wire \top1.memory1.mem2[148][0] ;
 wire \top1.memory1.mem2[148][1] ;
 wire \top1.memory1.mem2[148][2] ;
 wire \top1.memory1.mem2[149][0] ;
 wire \top1.memory1.mem2[149][1] ;
 wire \top1.memory1.mem2[149][2] ;
 wire \top1.memory1.mem2[14][0] ;
 wire \top1.memory1.mem2[14][1] ;
 wire \top1.memory1.mem2[14][2] ;
 wire \top1.memory1.mem2[150][0] ;
 wire \top1.memory1.mem2[150][1] ;
 wire \top1.memory1.mem2[150][2] ;
 wire \top1.memory1.mem2[151][0] ;
 wire \top1.memory1.mem2[151][1] ;
 wire \top1.memory1.mem2[151][2] ;
 wire \top1.memory1.mem2[152][0] ;
 wire \top1.memory1.mem2[152][1] ;
 wire \top1.memory1.mem2[152][2] ;
 wire \top1.memory1.mem2[153][0] ;
 wire \top1.memory1.mem2[153][1] ;
 wire \top1.memory1.mem2[153][2] ;
 wire \top1.memory1.mem2[154][0] ;
 wire \top1.memory1.mem2[154][1] ;
 wire \top1.memory1.mem2[154][2] ;
 wire \top1.memory1.mem2[155][0] ;
 wire \top1.memory1.mem2[155][1] ;
 wire \top1.memory1.mem2[155][2] ;
 wire \top1.memory1.mem2[156][0] ;
 wire \top1.memory1.mem2[156][1] ;
 wire \top1.memory1.mem2[156][2] ;
 wire \top1.memory1.mem2[157][0] ;
 wire \top1.memory1.mem2[157][1] ;
 wire \top1.memory1.mem2[157][2] ;
 wire \top1.memory1.mem2[158][0] ;
 wire \top1.memory1.mem2[158][1] ;
 wire \top1.memory1.mem2[158][2] ;
 wire \top1.memory1.mem2[159][0] ;
 wire \top1.memory1.mem2[159][1] ;
 wire \top1.memory1.mem2[159][2] ;
 wire \top1.memory1.mem2[15][0] ;
 wire \top1.memory1.mem2[15][1] ;
 wire \top1.memory1.mem2[15][2] ;
 wire \top1.memory1.mem2[160][0] ;
 wire \top1.memory1.mem2[160][1] ;
 wire \top1.memory1.mem2[160][2] ;
 wire \top1.memory1.mem2[161][0] ;
 wire \top1.memory1.mem2[161][1] ;
 wire \top1.memory1.mem2[161][2] ;
 wire \top1.memory1.mem2[162][0] ;
 wire \top1.memory1.mem2[162][1] ;
 wire \top1.memory1.mem2[162][2] ;
 wire \top1.memory1.mem2[163][0] ;
 wire \top1.memory1.mem2[163][1] ;
 wire \top1.memory1.mem2[163][2] ;
 wire \top1.memory1.mem2[164][0] ;
 wire \top1.memory1.mem2[164][1] ;
 wire \top1.memory1.mem2[164][2] ;
 wire \top1.memory1.mem2[165][0] ;
 wire \top1.memory1.mem2[165][1] ;
 wire \top1.memory1.mem2[165][2] ;
 wire \top1.memory1.mem2[166][0] ;
 wire \top1.memory1.mem2[166][1] ;
 wire \top1.memory1.mem2[166][2] ;
 wire \top1.memory1.mem2[167][0] ;
 wire \top1.memory1.mem2[167][1] ;
 wire \top1.memory1.mem2[167][2] ;
 wire \top1.memory1.mem2[168][0] ;
 wire \top1.memory1.mem2[168][1] ;
 wire \top1.memory1.mem2[168][2] ;
 wire \top1.memory1.mem2[169][0] ;
 wire \top1.memory1.mem2[169][1] ;
 wire \top1.memory1.mem2[169][2] ;
 wire \top1.memory1.mem2[16][0] ;
 wire \top1.memory1.mem2[16][1] ;
 wire \top1.memory1.mem2[16][2] ;
 wire \top1.memory1.mem2[170][0] ;
 wire \top1.memory1.mem2[170][1] ;
 wire \top1.memory1.mem2[170][2] ;
 wire \top1.memory1.mem2[171][0] ;
 wire \top1.memory1.mem2[171][1] ;
 wire \top1.memory1.mem2[171][2] ;
 wire \top1.memory1.mem2[172][0] ;
 wire \top1.memory1.mem2[172][1] ;
 wire \top1.memory1.mem2[172][2] ;
 wire \top1.memory1.mem2[173][0] ;
 wire \top1.memory1.mem2[173][1] ;
 wire \top1.memory1.mem2[173][2] ;
 wire \top1.memory1.mem2[174][0] ;
 wire \top1.memory1.mem2[174][1] ;
 wire \top1.memory1.mem2[174][2] ;
 wire \top1.memory1.mem2[175][0] ;
 wire \top1.memory1.mem2[175][1] ;
 wire \top1.memory1.mem2[175][2] ;
 wire \top1.memory1.mem2[176][0] ;
 wire \top1.memory1.mem2[176][1] ;
 wire \top1.memory1.mem2[176][2] ;
 wire \top1.memory1.mem2[177][0] ;
 wire \top1.memory1.mem2[177][1] ;
 wire \top1.memory1.mem2[177][2] ;
 wire \top1.memory1.mem2[178][0] ;
 wire \top1.memory1.mem2[178][1] ;
 wire \top1.memory1.mem2[178][2] ;
 wire \top1.memory1.mem2[179][0] ;
 wire \top1.memory1.mem2[179][1] ;
 wire \top1.memory1.mem2[179][2] ;
 wire \top1.memory1.mem2[17][0] ;
 wire \top1.memory1.mem2[17][1] ;
 wire \top1.memory1.mem2[17][2] ;
 wire \top1.memory1.mem2[180][0] ;
 wire \top1.memory1.mem2[180][1] ;
 wire \top1.memory1.mem2[180][2] ;
 wire \top1.memory1.mem2[181][0] ;
 wire \top1.memory1.mem2[181][1] ;
 wire \top1.memory1.mem2[181][2] ;
 wire \top1.memory1.mem2[182][0] ;
 wire \top1.memory1.mem2[182][1] ;
 wire \top1.memory1.mem2[182][2] ;
 wire \top1.memory1.mem2[183][0] ;
 wire \top1.memory1.mem2[183][1] ;
 wire \top1.memory1.mem2[183][2] ;
 wire \top1.memory1.mem2[184][0] ;
 wire \top1.memory1.mem2[184][1] ;
 wire \top1.memory1.mem2[184][2] ;
 wire \top1.memory1.mem2[185][0] ;
 wire \top1.memory1.mem2[185][1] ;
 wire \top1.memory1.mem2[185][2] ;
 wire \top1.memory1.mem2[186][0] ;
 wire \top1.memory1.mem2[186][1] ;
 wire \top1.memory1.mem2[186][2] ;
 wire \top1.memory1.mem2[187][0] ;
 wire \top1.memory1.mem2[187][1] ;
 wire \top1.memory1.mem2[187][2] ;
 wire \top1.memory1.mem2[188][0] ;
 wire \top1.memory1.mem2[188][1] ;
 wire \top1.memory1.mem2[188][2] ;
 wire \top1.memory1.mem2[189][0] ;
 wire \top1.memory1.mem2[189][1] ;
 wire \top1.memory1.mem2[189][2] ;
 wire \top1.memory1.mem2[18][0] ;
 wire \top1.memory1.mem2[18][1] ;
 wire \top1.memory1.mem2[18][2] ;
 wire \top1.memory1.mem2[190][0] ;
 wire \top1.memory1.mem2[190][1] ;
 wire \top1.memory1.mem2[190][2] ;
 wire \top1.memory1.mem2[191][0] ;
 wire \top1.memory1.mem2[191][1] ;
 wire \top1.memory1.mem2[191][2] ;
 wire \top1.memory1.mem2[192][0] ;
 wire \top1.memory1.mem2[192][1] ;
 wire \top1.memory1.mem2[192][2] ;
 wire \top1.memory1.mem2[193][0] ;
 wire \top1.memory1.mem2[193][1] ;
 wire \top1.memory1.mem2[193][2] ;
 wire \top1.memory1.mem2[194][0] ;
 wire \top1.memory1.mem2[194][1] ;
 wire \top1.memory1.mem2[194][2] ;
 wire \top1.memory1.mem2[195][0] ;
 wire \top1.memory1.mem2[195][1] ;
 wire \top1.memory1.mem2[195][2] ;
 wire \top1.memory1.mem2[196][0] ;
 wire \top1.memory1.mem2[196][1] ;
 wire \top1.memory1.mem2[196][2] ;
 wire \top1.memory1.mem2[197][0] ;
 wire \top1.memory1.mem2[197][1] ;
 wire \top1.memory1.mem2[197][2] ;
 wire \top1.memory1.mem2[198][0] ;
 wire \top1.memory1.mem2[198][1] ;
 wire \top1.memory1.mem2[198][2] ;
 wire \top1.memory1.mem2[199][0] ;
 wire \top1.memory1.mem2[199][1] ;
 wire \top1.memory1.mem2[199][2] ;
 wire \top1.memory1.mem2[19][0] ;
 wire \top1.memory1.mem2[19][1] ;
 wire \top1.memory1.mem2[19][2] ;
 wire \top1.memory1.mem2[1][0] ;
 wire \top1.memory1.mem2[1][1] ;
 wire \top1.memory1.mem2[1][2] ;
 wire \top1.memory1.mem2[20][0] ;
 wire \top1.memory1.mem2[20][1] ;
 wire \top1.memory1.mem2[20][2] ;
 wire \top1.memory1.mem2[21][0] ;
 wire \top1.memory1.mem2[21][1] ;
 wire \top1.memory1.mem2[21][2] ;
 wire \top1.memory1.mem2[22][0] ;
 wire \top1.memory1.mem2[22][1] ;
 wire \top1.memory1.mem2[22][2] ;
 wire \top1.memory1.mem2[23][0] ;
 wire \top1.memory1.mem2[23][1] ;
 wire \top1.memory1.mem2[23][2] ;
 wire \top1.memory1.mem2[24][0] ;
 wire \top1.memory1.mem2[24][1] ;
 wire \top1.memory1.mem2[24][2] ;
 wire \top1.memory1.mem2[25][0] ;
 wire \top1.memory1.mem2[25][1] ;
 wire \top1.memory1.mem2[25][2] ;
 wire \top1.memory1.mem2[26][0] ;
 wire \top1.memory1.mem2[26][1] ;
 wire \top1.memory1.mem2[26][2] ;
 wire \top1.memory1.mem2[27][0] ;
 wire \top1.memory1.mem2[27][1] ;
 wire \top1.memory1.mem2[27][2] ;
 wire \top1.memory1.mem2[28][0] ;
 wire \top1.memory1.mem2[28][1] ;
 wire \top1.memory1.mem2[28][2] ;
 wire \top1.memory1.mem2[29][0] ;
 wire \top1.memory1.mem2[29][1] ;
 wire \top1.memory1.mem2[29][2] ;
 wire \top1.memory1.mem2[2][0] ;
 wire \top1.memory1.mem2[2][1] ;
 wire \top1.memory1.mem2[2][2] ;
 wire \top1.memory1.mem2[30][0] ;
 wire \top1.memory1.mem2[30][1] ;
 wire \top1.memory1.mem2[30][2] ;
 wire \top1.memory1.mem2[31][0] ;
 wire \top1.memory1.mem2[31][1] ;
 wire \top1.memory1.mem2[31][2] ;
 wire \top1.memory1.mem2[32][0] ;
 wire \top1.memory1.mem2[32][1] ;
 wire \top1.memory1.mem2[32][2] ;
 wire \top1.memory1.mem2[33][0] ;
 wire \top1.memory1.mem2[33][1] ;
 wire \top1.memory1.mem2[33][2] ;
 wire \top1.memory1.mem2[34][0] ;
 wire \top1.memory1.mem2[34][1] ;
 wire \top1.memory1.mem2[34][2] ;
 wire \top1.memory1.mem2[35][0] ;
 wire \top1.memory1.mem2[35][1] ;
 wire \top1.memory1.mem2[35][2] ;
 wire \top1.memory1.mem2[36][0] ;
 wire \top1.memory1.mem2[36][1] ;
 wire \top1.memory1.mem2[36][2] ;
 wire \top1.memory1.mem2[37][0] ;
 wire \top1.memory1.mem2[37][1] ;
 wire \top1.memory1.mem2[37][2] ;
 wire \top1.memory1.mem2[38][0] ;
 wire \top1.memory1.mem2[38][1] ;
 wire \top1.memory1.mem2[38][2] ;
 wire \top1.memory1.mem2[39][0] ;
 wire \top1.memory1.mem2[39][1] ;
 wire \top1.memory1.mem2[39][2] ;
 wire \top1.memory1.mem2[3][0] ;
 wire \top1.memory1.mem2[3][1] ;
 wire \top1.memory1.mem2[3][2] ;
 wire \top1.memory1.mem2[40][0] ;
 wire \top1.memory1.mem2[40][1] ;
 wire \top1.memory1.mem2[40][2] ;
 wire \top1.memory1.mem2[41][0] ;
 wire \top1.memory1.mem2[41][1] ;
 wire \top1.memory1.mem2[41][2] ;
 wire \top1.memory1.mem2[42][0] ;
 wire \top1.memory1.mem2[42][1] ;
 wire \top1.memory1.mem2[42][2] ;
 wire \top1.memory1.mem2[43][0] ;
 wire \top1.memory1.mem2[43][1] ;
 wire \top1.memory1.mem2[43][2] ;
 wire \top1.memory1.mem2[44][0] ;
 wire \top1.memory1.mem2[44][1] ;
 wire \top1.memory1.mem2[44][2] ;
 wire \top1.memory1.mem2[45][0] ;
 wire \top1.memory1.mem2[45][1] ;
 wire \top1.memory1.mem2[45][2] ;
 wire \top1.memory1.mem2[46][0] ;
 wire \top1.memory1.mem2[46][1] ;
 wire \top1.memory1.mem2[46][2] ;
 wire \top1.memory1.mem2[47][0] ;
 wire \top1.memory1.mem2[47][1] ;
 wire \top1.memory1.mem2[47][2] ;
 wire \top1.memory1.mem2[48][0] ;
 wire \top1.memory1.mem2[48][1] ;
 wire \top1.memory1.mem2[48][2] ;
 wire \top1.memory1.mem2[49][0] ;
 wire \top1.memory1.mem2[49][1] ;
 wire \top1.memory1.mem2[49][2] ;
 wire \top1.memory1.mem2[4][0] ;
 wire \top1.memory1.mem2[4][1] ;
 wire \top1.memory1.mem2[4][2] ;
 wire \top1.memory1.mem2[50][0] ;
 wire \top1.memory1.mem2[50][1] ;
 wire \top1.memory1.mem2[50][2] ;
 wire \top1.memory1.mem2[51][0] ;
 wire \top1.memory1.mem2[51][1] ;
 wire \top1.memory1.mem2[51][2] ;
 wire \top1.memory1.mem2[52][0] ;
 wire \top1.memory1.mem2[52][1] ;
 wire \top1.memory1.mem2[52][2] ;
 wire \top1.memory1.mem2[53][0] ;
 wire \top1.memory1.mem2[53][1] ;
 wire \top1.memory1.mem2[53][2] ;
 wire \top1.memory1.mem2[54][0] ;
 wire \top1.memory1.mem2[54][1] ;
 wire \top1.memory1.mem2[54][2] ;
 wire \top1.memory1.mem2[55][0] ;
 wire \top1.memory1.mem2[55][1] ;
 wire \top1.memory1.mem2[55][2] ;
 wire \top1.memory1.mem2[56][0] ;
 wire \top1.memory1.mem2[56][1] ;
 wire \top1.memory1.mem2[56][2] ;
 wire \top1.memory1.mem2[57][0] ;
 wire \top1.memory1.mem2[57][1] ;
 wire \top1.memory1.mem2[57][2] ;
 wire \top1.memory1.mem2[58][0] ;
 wire \top1.memory1.mem2[58][1] ;
 wire \top1.memory1.mem2[58][2] ;
 wire \top1.memory1.mem2[59][0] ;
 wire \top1.memory1.mem2[59][1] ;
 wire \top1.memory1.mem2[59][2] ;
 wire \top1.memory1.mem2[5][0] ;
 wire \top1.memory1.mem2[5][1] ;
 wire \top1.memory1.mem2[5][2] ;
 wire \top1.memory1.mem2[60][0] ;
 wire \top1.memory1.mem2[60][1] ;
 wire \top1.memory1.mem2[60][2] ;
 wire \top1.memory1.mem2[61][0] ;
 wire \top1.memory1.mem2[61][1] ;
 wire \top1.memory1.mem2[61][2] ;
 wire \top1.memory1.mem2[62][0] ;
 wire \top1.memory1.mem2[62][1] ;
 wire \top1.memory1.mem2[62][2] ;
 wire \top1.memory1.mem2[63][0] ;
 wire \top1.memory1.mem2[63][1] ;
 wire \top1.memory1.mem2[63][2] ;
 wire \top1.memory1.mem2[64][0] ;
 wire \top1.memory1.mem2[64][1] ;
 wire \top1.memory1.mem2[64][2] ;
 wire \top1.memory1.mem2[65][0] ;
 wire \top1.memory1.mem2[65][1] ;
 wire \top1.memory1.mem2[65][2] ;
 wire \top1.memory1.mem2[66][0] ;
 wire \top1.memory1.mem2[66][1] ;
 wire \top1.memory1.mem2[66][2] ;
 wire \top1.memory1.mem2[67][0] ;
 wire \top1.memory1.mem2[67][1] ;
 wire \top1.memory1.mem2[67][2] ;
 wire \top1.memory1.mem2[68][0] ;
 wire \top1.memory1.mem2[68][1] ;
 wire \top1.memory1.mem2[68][2] ;
 wire \top1.memory1.mem2[69][0] ;
 wire \top1.memory1.mem2[69][1] ;
 wire \top1.memory1.mem2[69][2] ;
 wire \top1.memory1.mem2[6][0] ;
 wire \top1.memory1.mem2[6][1] ;
 wire \top1.memory1.mem2[6][2] ;
 wire \top1.memory1.mem2[70][0] ;
 wire \top1.memory1.mem2[70][1] ;
 wire \top1.memory1.mem2[70][2] ;
 wire \top1.memory1.mem2[71][0] ;
 wire \top1.memory1.mem2[71][1] ;
 wire \top1.memory1.mem2[71][2] ;
 wire \top1.memory1.mem2[72][0] ;
 wire \top1.memory1.mem2[72][1] ;
 wire \top1.memory1.mem2[72][2] ;
 wire \top1.memory1.mem2[73][0] ;
 wire \top1.memory1.mem2[73][1] ;
 wire \top1.memory1.mem2[73][2] ;
 wire \top1.memory1.mem2[74][0] ;
 wire \top1.memory1.mem2[74][1] ;
 wire \top1.memory1.mem2[74][2] ;
 wire \top1.memory1.mem2[75][0] ;
 wire \top1.memory1.mem2[75][1] ;
 wire \top1.memory1.mem2[75][2] ;
 wire \top1.memory1.mem2[76][0] ;
 wire \top1.memory1.mem2[76][1] ;
 wire \top1.memory1.mem2[76][2] ;
 wire \top1.memory1.mem2[77][0] ;
 wire \top1.memory1.mem2[77][1] ;
 wire \top1.memory1.mem2[77][2] ;
 wire \top1.memory1.mem2[78][0] ;
 wire \top1.memory1.mem2[78][1] ;
 wire \top1.memory1.mem2[78][2] ;
 wire \top1.memory1.mem2[79][0] ;
 wire \top1.memory1.mem2[79][1] ;
 wire \top1.memory1.mem2[79][2] ;
 wire \top1.memory1.mem2[7][0] ;
 wire \top1.memory1.mem2[7][1] ;
 wire \top1.memory1.mem2[7][2] ;
 wire \top1.memory1.mem2[80][0] ;
 wire \top1.memory1.mem2[80][1] ;
 wire \top1.memory1.mem2[80][2] ;
 wire \top1.memory1.mem2[81][0] ;
 wire \top1.memory1.mem2[81][1] ;
 wire \top1.memory1.mem2[81][2] ;
 wire \top1.memory1.mem2[82][0] ;
 wire \top1.memory1.mem2[82][1] ;
 wire \top1.memory1.mem2[82][2] ;
 wire \top1.memory1.mem2[83][0] ;
 wire \top1.memory1.mem2[83][1] ;
 wire \top1.memory1.mem2[83][2] ;
 wire \top1.memory1.mem2[84][0] ;
 wire \top1.memory1.mem2[84][1] ;
 wire \top1.memory1.mem2[84][2] ;
 wire \top1.memory1.mem2[85][0] ;
 wire \top1.memory1.mem2[85][1] ;
 wire \top1.memory1.mem2[85][2] ;
 wire \top1.memory1.mem2[86][0] ;
 wire \top1.memory1.mem2[86][1] ;
 wire \top1.memory1.mem2[86][2] ;
 wire \top1.memory1.mem2[87][0] ;
 wire \top1.memory1.mem2[87][1] ;
 wire \top1.memory1.mem2[87][2] ;
 wire \top1.memory1.mem2[88][0] ;
 wire \top1.memory1.mem2[88][1] ;
 wire \top1.memory1.mem2[88][2] ;
 wire \top1.memory1.mem2[89][0] ;
 wire \top1.memory1.mem2[89][1] ;
 wire \top1.memory1.mem2[89][2] ;
 wire \top1.memory1.mem2[8][0] ;
 wire \top1.memory1.mem2[8][1] ;
 wire \top1.memory1.mem2[8][2] ;
 wire \top1.memory1.mem2[90][0] ;
 wire \top1.memory1.mem2[90][1] ;
 wire \top1.memory1.mem2[90][2] ;
 wire \top1.memory1.mem2[91][0] ;
 wire \top1.memory1.mem2[91][1] ;
 wire \top1.memory1.mem2[91][2] ;
 wire \top1.memory1.mem2[92][0] ;
 wire \top1.memory1.mem2[92][1] ;
 wire \top1.memory1.mem2[92][2] ;
 wire \top1.memory1.mem2[93][0] ;
 wire \top1.memory1.mem2[93][1] ;
 wire \top1.memory1.mem2[93][2] ;
 wire \top1.memory1.mem2[94][0] ;
 wire \top1.memory1.mem2[94][1] ;
 wire \top1.memory1.mem2[94][2] ;
 wire \top1.memory1.mem2[95][0] ;
 wire \top1.memory1.mem2[95][1] ;
 wire \top1.memory1.mem2[95][2] ;
 wire \top1.memory1.mem2[96][0] ;
 wire \top1.memory1.mem2[96][1] ;
 wire \top1.memory1.mem2[96][2] ;
 wire \top1.memory1.mem2[97][0] ;
 wire \top1.memory1.mem2[97][1] ;
 wire \top1.memory1.mem2[97][2] ;
 wire \top1.memory1.mem2[98][0] ;
 wire \top1.memory1.mem2[98][1] ;
 wire \top1.memory1.mem2[98][2] ;
 wire \top1.memory1.mem2[99][0] ;
 wire \top1.memory1.mem2[99][1] ;
 wire \top1.memory1.mem2[99][2] ;
 wire \top1.memory1.mem2[9][0] ;
 wire \top1.memory1.mem2[9][1] ;
 wire \top1.memory1.mem2[9][2] ;
 wire \top1.memory2.data_out[0] ;
 wire \top1.memory2.data_out[1] ;
 wire \top1.memory2.data_out[2] ;
 wire \top1.memory2.mem1[0][0] ;
 wire \top1.memory2.mem1[0][1] ;
 wire \top1.memory2.mem1[0][2] ;
 wire \top1.memory2.mem1[100][0] ;
 wire \top1.memory2.mem1[100][1] ;
 wire \top1.memory2.mem1[100][2] ;
 wire \top1.memory2.mem1[101][0] ;
 wire \top1.memory2.mem1[101][1] ;
 wire \top1.memory2.mem1[101][2] ;
 wire \top1.memory2.mem1[102][0] ;
 wire \top1.memory2.mem1[102][1] ;
 wire \top1.memory2.mem1[102][2] ;
 wire \top1.memory2.mem1[103][0] ;
 wire \top1.memory2.mem1[103][1] ;
 wire \top1.memory2.mem1[103][2] ;
 wire \top1.memory2.mem1[104][0] ;
 wire \top1.memory2.mem1[104][1] ;
 wire \top1.memory2.mem1[104][2] ;
 wire \top1.memory2.mem1[105][0] ;
 wire \top1.memory2.mem1[105][1] ;
 wire \top1.memory2.mem1[105][2] ;
 wire \top1.memory2.mem1[106][0] ;
 wire \top1.memory2.mem1[106][1] ;
 wire \top1.memory2.mem1[106][2] ;
 wire \top1.memory2.mem1[107][0] ;
 wire \top1.memory2.mem1[107][1] ;
 wire \top1.memory2.mem1[107][2] ;
 wire \top1.memory2.mem1[108][0] ;
 wire \top1.memory2.mem1[108][1] ;
 wire \top1.memory2.mem1[108][2] ;
 wire \top1.memory2.mem1[109][0] ;
 wire \top1.memory2.mem1[109][1] ;
 wire \top1.memory2.mem1[109][2] ;
 wire \top1.memory2.mem1[10][0] ;
 wire \top1.memory2.mem1[10][1] ;
 wire \top1.memory2.mem1[10][2] ;
 wire \top1.memory2.mem1[110][0] ;
 wire \top1.memory2.mem1[110][1] ;
 wire \top1.memory2.mem1[110][2] ;
 wire \top1.memory2.mem1[111][0] ;
 wire \top1.memory2.mem1[111][1] ;
 wire \top1.memory2.mem1[111][2] ;
 wire \top1.memory2.mem1[112][0] ;
 wire \top1.memory2.mem1[112][1] ;
 wire \top1.memory2.mem1[112][2] ;
 wire \top1.memory2.mem1[113][0] ;
 wire \top1.memory2.mem1[113][1] ;
 wire \top1.memory2.mem1[113][2] ;
 wire \top1.memory2.mem1[114][0] ;
 wire \top1.memory2.mem1[114][1] ;
 wire \top1.memory2.mem1[114][2] ;
 wire \top1.memory2.mem1[115][0] ;
 wire \top1.memory2.mem1[115][1] ;
 wire \top1.memory2.mem1[115][2] ;
 wire \top1.memory2.mem1[116][0] ;
 wire \top1.memory2.mem1[116][1] ;
 wire \top1.memory2.mem1[116][2] ;
 wire \top1.memory2.mem1[117][0] ;
 wire \top1.memory2.mem1[117][1] ;
 wire \top1.memory2.mem1[117][2] ;
 wire \top1.memory2.mem1[118][0] ;
 wire \top1.memory2.mem1[118][1] ;
 wire \top1.memory2.mem1[118][2] ;
 wire \top1.memory2.mem1[119][0] ;
 wire \top1.memory2.mem1[119][1] ;
 wire \top1.memory2.mem1[119][2] ;
 wire \top1.memory2.mem1[11][0] ;
 wire \top1.memory2.mem1[11][1] ;
 wire \top1.memory2.mem1[11][2] ;
 wire \top1.memory2.mem1[120][0] ;
 wire \top1.memory2.mem1[120][1] ;
 wire \top1.memory2.mem1[120][2] ;
 wire \top1.memory2.mem1[121][0] ;
 wire \top1.memory2.mem1[121][1] ;
 wire \top1.memory2.mem1[121][2] ;
 wire \top1.memory2.mem1[122][0] ;
 wire \top1.memory2.mem1[122][1] ;
 wire \top1.memory2.mem1[122][2] ;
 wire \top1.memory2.mem1[123][0] ;
 wire \top1.memory2.mem1[123][1] ;
 wire \top1.memory2.mem1[123][2] ;
 wire \top1.memory2.mem1[124][0] ;
 wire \top1.memory2.mem1[124][1] ;
 wire \top1.memory2.mem1[124][2] ;
 wire \top1.memory2.mem1[125][0] ;
 wire \top1.memory2.mem1[125][1] ;
 wire \top1.memory2.mem1[125][2] ;
 wire \top1.memory2.mem1[126][0] ;
 wire \top1.memory2.mem1[126][1] ;
 wire \top1.memory2.mem1[126][2] ;
 wire \top1.memory2.mem1[127][0] ;
 wire \top1.memory2.mem1[127][1] ;
 wire \top1.memory2.mem1[127][2] ;
 wire \top1.memory2.mem1[128][0] ;
 wire \top1.memory2.mem1[128][1] ;
 wire \top1.memory2.mem1[128][2] ;
 wire \top1.memory2.mem1[129][0] ;
 wire \top1.memory2.mem1[129][1] ;
 wire \top1.memory2.mem1[129][2] ;
 wire \top1.memory2.mem1[12][0] ;
 wire \top1.memory2.mem1[12][1] ;
 wire \top1.memory2.mem1[12][2] ;
 wire \top1.memory2.mem1[130][0] ;
 wire \top1.memory2.mem1[130][1] ;
 wire \top1.memory2.mem1[130][2] ;
 wire \top1.memory2.mem1[131][0] ;
 wire \top1.memory2.mem1[131][1] ;
 wire \top1.memory2.mem1[131][2] ;
 wire \top1.memory2.mem1[132][0] ;
 wire \top1.memory2.mem1[132][1] ;
 wire \top1.memory2.mem1[132][2] ;
 wire \top1.memory2.mem1[133][0] ;
 wire \top1.memory2.mem1[133][1] ;
 wire \top1.memory2.mem1[133][2] ;
 wire \top1.memory2.mem1[134][0] ;
 wire \top1.memory2.mem1[134][1] ;
 wire \top1.memory2.mem1[134][2] ;
 wire \top1.memory2.mem1[135][0] ;
 wire \top1.memory2.mem1[135][1] ;
 wire \top1.memory2.mem1[135][2] ;
 wire \top1.memory2.mem1[136][0] ;
 wire \top1.memory2.mem1[136][1] ;
 wire \top1.memory2.mem1[136][2] ;
 wire \top1.memory2.mem1[137][0] ;
 wire \top1.memory2.mem1[137][1] ;
 wire \top1.memory2.mem1[137][2] ;
 wire \top1.memory2.mem1[138][0] ;
 wire \top1.memory2.mem1[138][1] ;
 wire \top1.memory2.mem1[138][2] ;
 wire \top1.memory2.mem1[139][0] ;
 wire \top1.memory2.mem1[139][1] ;
 wire \top1.memory2.mem1[139][2] ;
 wire \top1.memory2.mem1[13][0] ;
 wire \top1.memory2.mem1[13][1] ;
 wire \top1.memory2.mem1[13][2] ;
 wire \top1.memory2.mem1[140][0] ;
 wire \top1.memory2.mem1[140][1] ;
 wire \top1.memory2.mem1[140][2] ;
 wire \top1.memory2.mem1[141][0] ;
 wire \top1.memory2.mem1[141][1] ;
 wire \top1.memory2.mem1[141][2] ;
 wire \top1.memory2.mem1[142][0] ;
 wire \top1.memory2.mem1[142][1] ;
 wire \top1.memory2.mem1[142][2] ;
 wire \top1.memory2.mem1[143][0] ;
 wire \top1.memory2.mem1[143][1] ;
 wire \top1.memory2.mem1[143][2] ;
 wire \top1.memory2.mem1[144][0] ;
 wire \top1.memory2.mem1[144][1] ;
 wire \top1.memory2.mem1[144][2] ;
 wire \top1.memory2.mem1[145][0] ;
 wire \top1.memory2.mem1[145][1] ;
 wire \top1.memory2.mem1[145][2] ;
 wire \top1.memory2.mem1[146][0] ;
 wire \top1.memory2.mem1[146][1] ;
 wire \top1.memory2.mem1[146][2] ;
 wire \top1.memory2.mem1[147][0] ;
 wire \top1.memory2.mem1[147][1] ;
 wire \top1.memory2.mem1[147][2] ;
 wire \top1.memory2.mem1[148][0] ;
 wire \top1.memory2.mem1[148][1] ;
 wire \top1.memory2.mem1[148][2] ;
 wire \top1.memory2.mem1[149][0] ;
 wire \top1.memory2.mem1[149][1] ;
 wire \top1.memory2.mem1[149][2] ;
 wire \top1.memory2.mem1[14][0] ;
 wire \top1.memory2.mem1[14][1] ;
 wire \top1.memory2.mem1[14][2] ;
 wire \top1.memory2.mem1[150][0] ;
 wire \top1.memory2.mem1[150][1] ;
 wire \top1.memory2.mem1[150][2] ;
 wire \top1.memory2.mem1[151][0] ;
 wire \top1.memory2.mem1[151][1] ;
 wire \top1.memory2.mem1[151][2] ;
 wire \top1.memory2.mem1[152][0] ;
 wire \top1.memory2.mem1[152][1] ;
 wire \top1.memory2.mem1[152][2] ;
 wire \top1.memory2.mem1[153][0] ;
 wire \top1.memory2.mem1[153][1] ;
 wire \top1.memory2.mem1[153][2] ;
 wire \top1.memory2.mem1[154][0] ;
 wire \top1.memory2.mem1[154][1] ;
 wire \top1.memory2.mem1[154][2] ;
 wire \top1.memory2.mem1[155][0] ;
 wire \top1.memory2.mem1[155][1] ;
 wire \top1.memory2.mem1[155][2] ;
 wire \top1.memory2.mem1[156][0] ;
 wire \top1.memory2.mem1[156][1] ;
 wire \top1.memory2.mem1[156][2] ;
 wire \top1.memory2.mem1[157][0] ;
 wire \top1.memory2.mem1[157][1] ;
 wire \top1.memory2.mem1[157][2] ;
 wire \top1.memory2.mem1[158][0] ;
 wire \top1.memory2.mem1[158][1] ;
 wire \top1.memory2.mem1[158][2] ;
 wire \top1.memory2.mem1[159][0] ;
 wire \top1.memory2.mem1[159][1] ;
 wire \top1.memory2.mem1[159][2] ;
 wire \top1.memory2.mem1[15][0] ;
 wire \top1.memory2.mem1[15][1] ;
 wire \top1.memory2.mem1[15][2] ;
 wire \top1.memory2.mem1[160][0] ;
 wire \top1.memory2.mem1[160][1] ;
 wire \top1.memory2.mem1[160][2] ;
 wire \top1.memory2.mem1[161][0] ;
 wire \top1.memory2.mem1[161][1] ;
 wire \top1.memory2.mem1[161][2] ;
 wire \top1.memory2.mem1[162][0] ;
 wire \top1.memory2.mem1[162][1] ;
 wire \top1.memory2.mem1[162][2] ;
 wire \top1.memory2.mem1[163][0] ;
 wire \top1.memory2.mem1[163][1] ;
 wire \top1.memory2.mem1[163][2] ;
 wire \top1.memory2.mem1[164][0] ;
 wire \top1.memory2.mem1[164][1] ;
 wire \top1.memory2.mem1[164][2] ;
 wire \top1.memory2.mem1[165][0] ;
 wire \top1.memory2.mem1[165][1] ;
 wire \top1.memory2.mem1[165][2] ;
 wire \top1.memory2.mem1[166][0] ;
 wire \top1.memory2.mem1[166][1] ;
 wire \top1.memory2.mem1[166][2] ;
 wire \top1.memory2.mem1[167][0] ;
 wire \top1.memory2.mem1[167][1] ;
 wire \top1.memory2.mem1[167][2] ;
 wire \top1.memory2.mem1[168][0] ;
 wire \top1.memory2.mem1[168][1] ;
 wire \top1.memory2.mem1[168][2] ;
 wire \top1.memory2.mem1[169][0] ;
 wire \top1.memory2.mem1[169][1] ;
 wire \top1.memory2.mem1[169][2] ;
 wire \top1.memory2.mem1[16][0] ;
 wire \top1.memory2.mem1[16][1] ;
 wire \top1.memory2.mem1[16][2] ;
 wire \top1.memory2.mem1[170][0] ;
 wire \top1.memory2.mem1[170][1] ;
 wire \top1.memory2.mem1[170][2] ;
 wire \top1.memory2.mem1[171][0] ;
 wire \top1.memory2.mem1[171][1] ;
 wire \top1.memory2.mem1[171][2] ;
 wire \top1.memory2.mem1[172][0] ;
 wire \top1.memory2.mem1[172][1] ;
 wire \top1.memory2.mem1[172][2] ;
 wire \top1.memory2.mem1[173][0] ;
 wire \top1.memory2.mem1[173][1] ;
 wire \top1.memory2.mem1[173][2] ;
 wire \top1.memory2.mem1[174][0] ;
 wire \top1.memory2.mem1[174][1] ;
 wire \top1.memory2.mem1[174][2] ;
 wire \top1.memory2.mem1[175][0] ;
 wire \top1.memory2.mem1[175][1] ;
 wire \top1.memory2.mem1[175][2] ;
 wire \top1.memory2.mem1[176][0] ;
 wire \top1.memory2.mem1[176][1] ;
 wire \top1.memory2.mem1[176][2] ;
 wire \top1.memory2.mem1[177][0] ;
 wire \top1.memory2.mem1[177][1] ;
 wire \top1.memory2.mem1[177][2] ;
 wire \top1.memory2.mem1[178][0] ;
 wire \top1.memory2.mem1[178][1] ;
 wire \top1.memory2.mem1[178][2] ;
 wire \top1.memory2.mem1[179][0] ;
 wire \top1.memory2.mem1[179][1] ;
 wire \top1.memory2.mem1[179][2] ;
 wire \top1.memory2.mem1[17][0] ;
 wire \top1.memory2.mem1[17][1] ;
 wire \top1.memory2.mem1[17][2] ;
 wire \top1.memory2.mem1[180][0] ;
 wire \top1.memory2.mem1[180][1] ;
 wire \top1.memory2.mem1[180][2] ;
 wire \top1.memory2.mem1[181][0] ;
 wire \top1.memory2.mem1[181][1] ;
 wire \top1.memory2.mem1[181][2] ;
 wire \top1.memory2.mem1[182][0] ;
 wire \top1.memory2.mem1[182][1] ;
 wire \top1.memory2.mem1[182][2] ;
 wire \top1.memory2.mem1[183][0] ;
 wire \top1.memory2.mem1[183][1] ;
 wire \top1.memory2.mem1[183][2] ;
 wire \top1.memory2.mem1[184][0] ;
 wire \top1.memory2.mem1[184][1] ;
 wire \top1.memory2.mem1[184][2] ;
 wire \top1.memory2.mem1[185][0] ;
 wire \top1.memory2.mem1[185][1] ;
 wire \top1.memory2.mem1[185][2] ;
 wire \top1.memory2.mem1[186][0] ;
 wire \top1.memory2.mem1[186][1] ;
 wire \top1.memory2.mem1[186][2] ;
 wire \top1.memory2.mem1[187][0] ;
 wire \top1.memory2.mem1[187][1] ;
 wire \top1.memory2.mem1[187][2] ;
 wire \top1.memory2.mem1[188][0] ;
 wire \top1.memory2.mem1[188][1] ;
 wire \top1.memory2.mem1[188][2] ;
 wire \top1.memory2.mem1[189][0] ;
 wire \top1.memory2.mem1[189][1] ;
 wire \top1.memory2.mem1[189][2] ;
 wire \top1.memory2.mem1[18][0] ;
 wire \top1.memory2.mem1[18][1] ;
 wire \top1.memory2.mem1[18][2] ;
 wire \top1.memory2.mem1[190][0] ;
 wire \top1.memory2.mem1[190][1] ;
 wire \top1.memory2.mem1[190][2] ;
 wire \top1.memory2.mem1[191][0] ;
 wire \top1.memory2.mem1[191][1] ;
 wire \top1.memory2.mem1[191][2] ;
 wire \top1.memory2.mem1[192][0] ;
 wire \top1.memory2.mem1[192][1] ;
 wire \top1.memory2.mem1[192][2] ;
 wire \top1.memory2.mem1[193][0] ;
 wire \top1.memory2.mem1[193][1] ;
 wire \top1.memory2.mem1[193][2] ;
 wire \top1.memory2.mem1[194][0] ;
 wire \top1.memory2.mem1[194][1] ;
 wire \top1.memory2.mem1[194][2] ;
 wire \top1.memory2.mem1[195][0] ;
 wire \top1.memory2.mem1[195][1] ;
 wire \top1.memory2.mem1[195][2] ;
 wire \top1.memory2.mem1[196][0] ;
 wire \top1.memory2.mem1[196][1] ;
 wire \top1.memory2.mem1[196][2] ;
 wire \top1.memory2.mem1[197][0] ;
 wire \top1.memory2.mem1[197][1] ;
 wire \top1.memory2.mem1[197][2] ;
 wire \top1.memory2.mem1[198][0] ;
 wire \top1.memory2.mem1[198][1] ;
 wire \top1.memory2.mem1[198][2] ;
 wire \top1.memory2.mem1[199][0] ;
 wire \top1.memory2.mem1[199][1] ;
 wire \top1.memory2.mem1[199][2] ;
 wire \top1.memory2.mem1[19][0] ;
 wire \top1.memory2.mem1[19][1] ;
 wire \top1.memory2.mem1[19][2] ;
 wire \top1.memory2.mem1[1][0] ;
 wire \top1.memory2.mem1[1][1] ;
 wire \top1.memory2.mem1[1][2] ;
 wire \top1.memory2.mem1[20][0] ;
 wire \top1.memory2.mem1[20][1] ;
 wire \top1.memory2.mem1[20][2] ;
 wire \top1.memory2.mem1[21][0] ;
 wire \top1.memory2.mem1[21][1] ;
 wire \top1.memory2.mem1[21][2] ;
 wire \top1.memory2.mem1[22][0] ;
 wire \top1.memory2.mem1[22][1] ;
 wire \top1.memory2.mem1[22][2] ;
 wire \top1.memory2.mem1[23][0] ;
 wire \top1.memory2.mem1[23][1] ;
 wire \top1.memory2.mem1[23][2] ;
 wire \top1.memory2.mem1[24][0] ;
 wire \top1.memory2.mem1[24][1] ;
 wire \top1.memory2.mem1[24][2] ;
 wire \top1.memory2.mem1[25][0] ;
 wire \top1.memory2.mem1[25][1] ;
 wire \top1.memory2.mem1[25][2] ;
 wire \top1.memory2.mem1[26][0] ;
 wire \top1.memory2.mem1[26][1] ;
 wire \top1.memory2.mem1[26][2] ;
 wire \top1.memory2.mem1[27][0] ;
 wire \top1.memory2.mem1[27][1] ;
 wire \top1.memory2.mem1[27][2] ;
 wire \top1.memory2.mem1[28][0] ;
 wire \top1.memory2.mem1[28][1] ;
 wire \top1.memory2.mem1[28][2] ;
 wire \top1.memory2.mem1[29][0] ;
 wire \top1.memory2.mem1[29][1] ;
 wire \top1.memory2.mem1[29][2] ;
 wire \top1.memory2.mem1[2][0] ;
 wire \top1.memory2.mem1[2][1] ;
 wire \top1.memory2.mem1[2][2] ;
 wire \top1.memory2.mem1[30][0] ;
 wire \top1.memory2.mem1[30][1] ;
 wire \top1.memory2.mem1[30][2] ;
 wire \top1.memory2.mem1[31][0] ;
 wire \top1.memory2.mem1[31][1] ;
 wire \top1.memory2.mem1[31][2] ;
 wire \top1.memory2.mem1[32][0] ;
 wire \top1.memory2.mem1[32][1] ;
 wire \top1.memory2.mem1[32][2] ;
 wire \top1.memory2.mem1[33][0] ;
 wire \top1.memory2.mem1[33][1] ;
 wire \top1.memory2.mem1[33][2] ;
 wire \top1.memory2.mem1[34][0] ;
 wire \top1.memory2.mem1[34][1] ;
 wire \top1.memory2.mem1[34][2] ;
 wire \top1.memory2.mem1[35][0] ;
 wire \top1.memory2.mem1[35][1] ;
 wire \top1.memory2.mem1[35][2] ;
 wire \top1.memory2.mem1[36][0] ;
 wire \top1.memory2.mem1[36][1] ;
 wire \top1.memory2.mem1[36][2] ;
 wire \top1.memory2.mem1[37][0] ;
 wire \top1.memory2.mem1[37][1] ;
 wire \top1.memory2.mem1[37][2] ;
 wire \top1.memory2.mem1[38][0] ;
 wire \top1.memory2.mem1[38][1] ;
 wire \top1.memory2.mem1[38][2] ;
 wire \top1.memory2.mem1[39][0] ;
 wire \top1.memory2.mem1[39][1] ;
 wire \top1.memory2.mem1[39][2] ;
 wire \top1.memory2.mem1[3][0] ;
 wire \top1.memory2.mem1[3][1] ;
 wire \top1.memory2.mem1[3][2] ;
 wire \top1.memory2.mem1[40][0] ;
 wire \top1.memory2.mem1[40][1] ;
 wire \top1.memory2.mem1[40][2] ;
 wire \top1.memory2.mem1[41][0] ;
 wire \top1.memory2.mem1[41][1] ;
 wire \top1.memory2.mem1[41][2] ;
 wire \top1.memory2.mem1[42][0] ;
 wire \top1.memory2.mem1[42][1] ;
 wire \top1.memory2.mem1[42][2] ;
 wire \top1.memory2.mem1[43][0] ;
 wire \top1.memory2.mem1[43][1] ;
 wire \top1.memory2.mem1[43][2] ;
 wire \top1.memory2.mem1[44][0] ;
 wire \top1.memory2.mem1[44][1] ;
 wire \top1.memory2.mem1[44][2] ;
 wire \top1.memory2.mem1[45][0] ;
 wire \top1.memory2.mem1[45][1] ;
 wire \top1.memory2.mem1[45][2] ;
 wire \top1.memory2.mem1[46][0] ;
 wire \top1.memory2.mem1[46][1] ;
 wire \top1.memory2.mem1[46][2] ;
 wire \top1.memory2.mem1[47][0] ;
 wire \top1.memory2.mem1[47][1] ;
 wire \top1.memory2.mem1[47][2] ;
 wire \top1.memory2.mem1[48][0] ;
 wire \top1.memory2.mem1[48][1] ;
 wire \top1.memory2.mem1[48][2] ;
 wire \top1.memory2.mem1[49][0] ;
 wire \top1.memory2.mem1[49][1] ;
 wire \top1.memory2.mem1[49][2] ;
 wire \top1.memory2.mem1[4][0] ;
 wire \top1.memory2.mem1[4][1] ;
 wire \top1.memory2.mem1[4][2] ;
 wire \top1.memory2.mem1[50][0] ;
 wire \top1.memory2.mem1[50][1] ;
 wire \top1.memory2.mem1[50][2] ;
 wire \top1.memory2.mem1[51][0] ;
 wire \top1.memory2.mem1[51][1] ;
 wire \top1.memory2.mem1[51][2] ;
 wire \top1.memory2.mem1[52][0] ;
 wire \top1.memory2.mem1[52][1] ;
 wire \top1.memory2.mem1[52][2] ;
 wire \top1.memory2.mem1[53][0] ;
 wire \top1.memory2.mem1[53][1] ;
 wire \top1.memory2.mem1[53][2] ;
 wire \top1.memory2.mem1[54][0] ;
 wire \top1.memory2.mem1[54][1] ;
 wire \top1.memory2.mem1[54][2] ;
 wire \top1.memory2.mem1[55][0] ;
 wire \top1.memory2.mem1[55][1] ;
 wire \top1.memory2.mem1[55][2] ;
 wire \top1.memory2.mem1[56][0] ;
 wire \top1.memory2.mem1[56][1] ;
 wire \top1.memory2.mem1[56][2] ;
 wire \top1.memory2.mem1[57][0] ;
 wire \top1.memory2.mem1[57][1] ;
 wire \top1.memory2.mem1[57][2] ;
 wire \top1.memory2.mem1[58][0] ;
 wire \top1.memory2.mem1[58][1] ;
 wire \top1.memory2.mem1[58][2] ;
 wire \top1.memory2.mem1[59][0] ;
 wire \top1.memory2.mem1[59][1] ;
 wire \top1.memory2.mem1[59][2] ;
 wire \top1.memory2.mem1[5][0] ;
 wire \top1.memory2.mem1[5][1] ;
 wire \top1.memory2.mem1[5][2] ;
 wire \top1.memory2.mem1[60][0] ;
 wire \top1.memory2.mem1[60][1] ;
 wire \top1.memory2.mem1[60][2] ;
 wire \top1.memory2.mem1[61][0] ;
 wire \top1.memory2.mem1[61][1] ;
 wire \top1.memory2.mem1[61][2] ;
 wire \top1.memory2.mem1[62][0] ;
 wire \top1.memory2.mem1[62][1] ;
 wire \top1.memory2.mem1[62][2] ;
 wire \top1.memory2.mem1[63][0] ;
 wire \top1.memory2.mem1[63][1] ;
 wire \top1.memory2.mem1[63][2] ;
 wire \top1.memory2.mem1[64][0] ;
 wire \top1.memory2.mem1[64][1] ;
 wire \top1.memory2.mem1[64][2] ;
 wire \top1.memory2.mem1[65][0] ;
 wire \top1.memory2.mem1[65][1] ;
 wire \top1.memory2.mem1[65][2] ;
 wire \top1.memory2.mem1[66][0] ;
 wire \top1.memory2.mem1[66][1] ;
 wire \top1.memory2.mem1[66][2] ;
 wire \top1.memory2.mem1[67][0] ;
 wire \top1.memory2.mem1[67][1] ;
 wire \top1.memory2.mem1[67][2] ;
 wire \top1.memory2.mem1[68][0] ;
 wire \top1.memory2.mem1[68][1] ;
 wire \top1.memory2.mem1[68][2] ;
 wire \top1.memory2.mem1[69][0] ;
 wire \top1.memory2.mem1[69][1] ;
 wire \top1.memory2.mem1[69][2] ;
 wire \top1.memory2.mem1[6][0] ;
 wire \top1.memory2.mem1[6][1] ;
 wire \top1.memory2.mem1[6][2] ;
 wire \top1.memory2.mem1[70][0] ;
 wire \top1.memory2.mem1[70][1] ;
 wire \top1.memory2.mem1[70][2] ;
 wire \top1.memory2.mem1[71][0] ;
 wire \top1.memory2.mem1[71][1] ;
 wire \top1.memory2.mem1[71][2] ;
 wire \top1.memory2.mem1[72][0] ;
 wire \top1.memory2.mem1[72][1] ;
 wire \top1.memory2.mem1[72][2] ;
 wire \top1.memory2.mem1[73][0] ;
 wire \top1.memory2.mem1[73][1] ;
 wire \top1.memory2.mem1[73][2] ;
 wire \top1.memory2.mem1[74][0] ;
 wire \top1.memory2.mem1[74][1] ;
 wire \top1.memory2.mem1[74][2] ;
 wire \top1.memory2.mem1[75][0] ;
 wire \top1.memory2.mem1[75][1] ;
 wire \top1.memory2.mem1[75][2] ;
 wire \top1.memory2.mem1[76][0] ;
 wire \top1.memory2.mem1[76][1] ;
 wire \top1.memory2.mem1[76][2] ;
 wire \top1.memory2.mem1[77][0] ;
 wire \top1.memory2.mem1[77][1] ;
 wire \top1.memory2.mem1[77][2] ;
 wire \top1.memory2.mem1[78][0] ;
 wire \top1.memory2.mem1[78][1] ;
 wire \top1.memory2.mem1[78][2] ;
 wire \top1.memory2.mem1[79][0] ;
 wire \top1.memory2.mem1[79][1] ;
 wire \top1.memory2.mem1[79][2] ;
 wire \top1.memory2.mem1[7][0] ;
 wire \top1.memory2.mem1[7][1] ;
 wire \top1.memory2.mem1[7][2] ;
 wire \top1.memory2.mem1[80][0] ;
 wire \top1.memory2.mem1[80][1] ;
 wire \top1.memory2.mem1[80][2] ;
 wire \top1.memory2.mem1[81][0] ;
 wire \top1.memory2.mem1[81][1] ;
 wire \top1.memory2.mem1[81][2] ;
 wire \top1.memory2.mem1[82][0] ;
 wire \top1.memory2.mem1[82][1] ;
 wire \top1.memory2.mem1[82][2] ;
 wire \top1.memory2.mem1[83][0] ;
 wire \top1.memory2.mem1[83][1] ;
 wire \top1.memory2.mem1[83][2] ;
 wire \top1.memory2.mem1[84][0] ;
 wire \top1.memory2.mem1[84][1] ;
 wire \top1.memory2.mem1[84][2] ;
 wire \top1.memory2.mem1[85][0] ;
 wire \top1.memory2.mem1[85][1] ;
 wire \top1.memory2.mem1[85][2] ;
 wire \top1.memory2.mem1[86][0] ;
 wire \top1.memory2.mem1[86][1] ;
 wire \top1.memory2.mem1[86][2] ;
 wire \top1.memory2.mem1[87][0] ;
 wire \top1.memory2.mem1[87][1] ;
 wire \top1.memory2.mem1[87][2] ;
 wire \top1.memory2.mem1[88][0] ;
 wire \top1.memory2.mem1[88][1] ;
 wire \top1.memory2.mem1[88][2] ;
 wire \top1.memory2.mem1[89][0] ;
 wire \top1.memory2.mem1[89][1] ;
 wire \top1.memory2.mem1[89][2] ;
 wire \top1.memory2.mem1[8][0] ;
 wire \top1.memory2.mem1[8][1] ;
 wire \top1.memory2.mem1[8][2] ;
 wire \top1.memory2.mem1[90][0] ;
 wire \top1.memory2.mem1[90][1] ;
 wire \top1.memory2.mem1[90][2] ;
 wire \top1.memory2.mem1[91][0] ;
 wire \top1.memory2.mem1[91][1] ;
 wire \top1.memory2.mem1[91][2] ;
 wire \top1.memory2.mem1[92][0] ;
 wire \top1.memory2.mem1[92][1] ;
 wire \top1.memory2.mem1[92][2] ;
 wire \top1.memory2.mem1[93][0] ;
 wire \top1.memory2.mem1[93][1] ;
 wire \top1.memory2.mem1[93][2] ;
 wire \top1.memory2.mem1[94][0] ;
 wire \top1.memory2.mem1[94][1] ;
 wire \top1.memory2.mem1[94][2] ;
 wire \top1.memory2.mem1[95][0] ;
 wire \top1.memory2.mem1[95][1] ;
 wire \top1.memory2.mem1[95][2] ;
 wire \top1.memory2.mem1[96][0] ;
 wire \top1.memory2.mem1[96][1] ;
 wire \top1.memory2.mem1[96][2] ;
 wire \top1.memory2.mem1[97][0] ;
 wire \top1.memory2.mem1[97][1] ;
 wire \top1.memory2.mem1[97][2] ;
 wire \top1.memory2.mem1[98][0] ;
 wire \top1.memory2.mem1[98][1] ;
 wire \top1.memory2.mem1[98][2] ;
 wire \top1.memory2.mem1[99][0] ;
 wire \top1.memory2.mem1[99][1] ;
 wire \top1.memory2.mem1[99][2] ;
 wire \top1.memory2.mem1[9][0] ;
 wire \top1.memory2.mem1[9][1] ;
 wire \top1.memory2.mem1[9][2] ;
 wire \top1.memory2.mem2[0][0] ;
 wire \top1.memory2.mem2[0][1] ;
 wire \top1.memory2.mem2[0][2] ;
 wire \top1.memory2.mem2[100][0] ;
 wire \top1.memory2.mem2[100][1] ;
 wire \top1.memory2.mem2[100][2] ;
 wire \top1.memory2.mem2[101][0] ;
 wire \top1.memory2.mem2[101][1] ;
 wire \top1.memory2.mem2[101][2] ;
 wire \top1.memory2.mem2[102][0] ;
 wire \top1.memory2.mem2[102][1] ;
 wire \top1.memory2.mem2[102][2] ;
 wire \top1.memory2.mem2[103][0] ;
 wire \top1.memory2.mem2[103][1] ;
 wire \top1.memory2.mem2[103][2] ;
 wire \top1.memory2.mem2[104][0] ;
 wire \top1.memory2.mem2[104][1] ;
 wire \top1.memory2.mem2[104][2] ;
 wire \top1.memory2.mem2[105][0] ;
 wire \top1.memory2.mem2[105][1] ;
 wire \top1.memory2.mem2[105][2] ;
 wire \top1.memory2.mem2[106][0] ;
 wire \top1.memory2.mem2[106][1] ;
 wire \top1.memory2.mem2[106][2] ;
 wire \top1.memory2.mem2[107][0] ;
 wire \top1.memory2.mem2[107][1] ;
 wire \top1.memory2.mem2[107][2] ;
 wire \top1.memory2.mem2[108][0] ;
 wire \top1.memory2.mem2[108][1] ;
 wire \top1.memory2.mem2[108][2] ;
 wire \top1.memory2.mem2[109][0] ;
 wire \top1.memory2.mem2[109][1] ;
 wire \top1.memory2.mem2[109][2] ;
 wire \top1.memory2.mem2[10][0] ;
 wire \top1.memory2.mem2[10][1] ;
 wire \top1.memory2.mem2[10][2] ;
 wire \top1.memory2.mem2[110][0] ;
 wire \top1.memory2.mem2[110][1] ;
 wire \top1.memory2.mem2[110][2] ;
 wire \top1.memory2.mem2[111][0] ;
 wire \top1.memory2.mem2[111][1] ;
 wire \top1.memory2.mem2[111][2] ;
 wire \top1.memory2.mem2[112][0] ;
 wire \top1.memory2.mem2[112][1] ;
 wire \top1.memory2.mem2[112][2] ;
 wire \top1.memory2.mem2[113][0] ;
 wire \top1.memory2.mem2[113][1] ;
 wire \top1.memory2.mem2[113][2] ;
 wire \top1.memory2.mem2[114][0] ;
 wire \top1.memory2.mem2[114][1] ;
 wire \top1.memory2.mem2[114][2] ;
 wire \top1.memory2.mem2[115][0] ;
 wire \top1.memory2.mem2[115][1] ;
 wire \top1.memory2.mem2[115][2] ;
 wire \top1.memory2.mem2[116][0] ;
 wire \top1.memory2.mem2[116][1] ;
 wire \top1.memory2.mem2[116][2] ;
 wire \top1.memory2.mem2[117][0] ;
 wire \top1.memory2.mem2[117][1] ;
 wire \top1.memory2.mem2[117][2] ;
 wire \top1.memory2.mem2[118][0] ;
 wire \top1.memory2.mem2[118][1] ;
 wire \top1.memory2.mem2[118][2] ;
 wire \top1.memory2.mem2[119][0] ;
 wire \top1.memory2.mem2[119][1] ;
 wire \top1.memory2.mem2[119][2] ;
 wire \top1.memory2.mem2[11][0] ;
 wire \top1.memory2.mem2[11][1] ;
 wire \top1.memory2.mem2[11][2] ;
 wire \top1.memory2.mem2[120][0] ;
 wire \top1.memory2.mem2[120][1] ;
 wire \top1.memory2.mem2[120][2] ;
 wire \top1.memory2.mem2[121][0] ;
 wire \top1.memory2.mem2[121][1] ;
 wire \top1.memory2.mem2[121][2] ;
 wire \top1.memory2.mem2[122][0] ;
 wire \top1.memory2.mem2[122][1] ;
 wire \top1.memory2.mem2[122][2] ;
 wire \top1.memory2.mem2[123][0] ;
 wire \top1.memory2.mem2[123][1] ;
 wire \top1.memory2.mem2[123][2] ;
 wire \top1.memory2.mem2[124][0] ;
 wire \top1.memory2.mem2[124][1] ;
 wire \top1.memory2.mem2[124][2] ;
 wire \top1.memory2.mem2[125][0] ;
 wire \top1.memory2.mem2[125][1] ;
 wire \top1.memory2.mem2[125][2] ;
 wire \top1.memory2.mem2[126][0] ;
 wire \top1.memory2.mem2[126][1] ;
 wire \top1.memory2.mem2[126][2] ;
 wire \top1.memory2.mem2[127][0] ;
 wire \top1.memory2.mem2[127][1] ;
 wire \top1.memory2.mem2[127][2] ;
 wire \top1.memory2.mem2[128][0] ;
 wire \top1.memory2.mem2[128][1] ;
 wire \top1.memory2.mem2[128][2] ;
 wire \top1.memory2.mem2[129][0] ;
 wire \top1.memory2.mem2[129][1] ;
 wire \top1.memory2.mem2[129][2] ;
 wire \top1.memory2.mem2[12][0] ;
 wire \top1.memory2.mem2[12][1] ;
 wire \top1.memory2.mem2[12][2] ;
 wire \top1.memory2.mem2[130][0] ;
 wire \top1.memory2.mem2[130][1] ;
 wire \top1.memory2.mem2[130][2] ;
 wire \top1.memory2.mem2[131][0] ;
 wire \top1.memory2.mem2[131][1] ;
 wire \top1.memory2.mem2[131][2] ;
 wire \top1.memory2.mem2[132][0] ;
 wire \top1.memory2.mem2[132][1] ;
 wire \top1.memory2.mem2[132][2] ;
 wire \top1.memory2.mem2[133][0] ;
 wire \top1.memory2.mem2[133][1] ;
 wire \top1.memory2.mem2[133][2] ;
 wire \top1.memory2.mem2[134][0] ;
 wire \top1.memory2.mem2[134][1] ;
 wire \top1.memory2.mem2[134][2] ;
 wire \top1.memory2.mem2[135][0] ;
 wire \top1.memory2.mem2[135][1] ;
 wire \top1.memory2.mem2[135][2] ;
 wire \top1.memory2.mem2[136][0] ;
 wire \top1.memory2.mem2[136][1] ;
 wire \top1.memory2.mem2[136][2] ;
 wire \top1.memory2.mem2[137][0] ;
 wire \top1.memory2.mem2[137][1] ;
 wire \top1.memory2.mem2[137][2] ;
 wire \top1.memory2.mem2[138][0] ;
 wire \top1.memory2.mem2[138][1] ;
 wire \top1.memory2.mem2[138][2] ;
 wire \top1.memory2.mem2[139][0] ;
 wire \top1.memory2.mem2[139][1] ;
 wire \top1.memory2.mem2[139][2] ;
 wire \top1.memory2.mem2[13][0] ;
 wire \top1.memory2.mem2[13][1] ;
 wire \top1.memory2.mem2[13][2] ;
 wire \top1.memory2.mem2[140][0] ;
 wire \top1.memory2.mem2[140][1] ;
 wire \top1.memory2.mem2[140][2] ;
 wire \top1.memory2.mem2[141][0] ;
 wire \top1.memory2.mem2[141][1] ;
 wire \top1.memory2.mem2[141][2] ;
 wire \top1.memory2.mem2[142][0] ;
 wire \top1.memory2.mem2[142][1] ;
 wire \top1.memory2.mem2[142][2] ;
 wire \top1.memory2.mem2[143][0] ;
 wire \top1.memory2.mem2[143][1] ;
 wire \top1.memory2.mem2[143][2] ;
 wire \top1.memory2.mem2[144][0] ;
 wire \top1.memory2.mem2[144][1] ;
 wire \top1.memory2.mem2[144][2] ;
 wire \top1.memory2.mem2[145][0] ;
 wire \top1.memory2.mem2[145][1] ;
 wire \top1.memory2.mem2[145][2] ;
 wire \top1.memory2.mem2[146][0] ;
 wire \top1.memory2.mem2[146][1] ;
 wire \top1.memory2.mem2[146][2] ;
 wire \top1.memory2.mem2[147][0] ;
 wire \top1.memory2.mem2[147][1] ;
 wire \top1.memory2.mem2[147][2] ;
 wire \top1.memory2.mem2[148][0] ;
 wire \top1.memory2.mem2[148][1] ;
 wire \top1.memory2.mem2[148][2] ;
 wire \top1.memory2.mem2[149][0] ;
 wire \top1.memory2.mem2[149][1] ;
 wire \top1.memory2.mem2[149][2] ;
 wire \top1.memory2.mem2[14][0] ;
 wire \top1.memory2.mem2[14][1] ;
 wire \top1.memory2.mem2[14][2] ;
 wire \top1.memory2.mem2[150][0] ;
 wire \top1.memory2.mem2[150][1] ;
 wire \top1.memory2.mem2[150][2] ;
 wire \top1.memory2.mem2[151][0] ;
 wire \top1.memory2.mem2[151][1] ;
 wire \top1.memory2.mem2[151][2] ;
 wire \top1.memory2.mem2[152][0] ;
 wire \top1.memory2.mem2[152][1] ;
 wire \top1.memory2.mem2[152][2] ;
 wire \top1.memory2.mem2[153][0] ;
 wire \top1.memory2.mem2[153][1] ;
 wire \top1.memory2.mem2[153][2] ;
 wire \top1.memory2.mem2[154][0] ;
 wire \top1.memory2.mem2[154][1] ;
 wire \top1.memory2.mem2[154][2] ;
 wire \top1.memory2.mem2[155][0] ;
 wire \top1.memory2.mem2[155][1] ;
 wire \top1.memory2.mem2[155][2] ;
 wire \top1.memory2.mem2[156][0] ;
 wire \top1.memory2.mem2[156][1] ;
 wire \top1.memory2.mem2[156][2] ;
 wire \top1.memory2.mem2[157][0] ;
 wire \top1.memory2.mem2[157][1] ;
 wire \top1.memory2.mem2[157][2] ;
 wire \top1.memory2.mem2[158][0] ;
 wire \top1.memory2.mem2[158][1] ;
 wire \top1.memory2.mem2[158][2] ;
 wire \top1.memory2.mem2[159][0] ;
 wire \top1.memory2.mem2[159][1] ;
 wire \top1.memory2.mem2[159][2] ;
 wire \top1.memory2.mem2[15][0] ;
 wire \top1.memory2.mem2[15][1] ;
 wire \top1.memory2.mem2[15][2] ;
 wire \top1.memory2.mem2[160][0] ;
 wire \top1.memory2.mem2[160][1] ;
 wire \top1.memory2.mem2[160][2] ;
 wire \top1.memory2.mem2[161][0] ;
 wire \top1.memory2.mem2[161][1] ;
 wire \top1.memory2.mem2[161][2] ;
 wire \top1.memory2.mem2[162][0] ;
 wire \top1.memory2.mem2[162][1] ;
 wire \top1.memory2.mem2[162][2] ;
 wire \top1.memory2.mem2[163][0] ;
 wire \top1.memory2.mem2[163][1] ;
 wire \top1.memory2.mem2[163][2] ;
 wire \top1.memory2.mem2[164][0] ;
 wire \top1.memory2.mem2[164][1] ;
 wire \top1.memory2.mem2[164][2] ;
 wire \top1.memory2.mem2[165][0] ;
 wire \top1.memory2.mem2[165][1] ;
 wire \top1.memory2.mem2[165][2] ;
 wire \top1.memory2.mem2[166][0] ;
 wire \top1.memory2.mem2[166][1] ;
 wire \top1.memory2.mem2[166][2] ;
 wire \top1.memory2.mem2[167][0] ;
 wire \top1.memory2.mem2[167][1] ;
 wire \top1.memory2.mem2[167][2] ;
 wire \top1.memory2.mem2[168][0] ;
 wire \top1.memory2.mem2[168][1] ;
 wire \top1.memory2.mem2[168][2] ;
 wire \top1.memory2.mem2[169][0] ;
 wire \top1.memory2.mem2[169][1] ;
 wire \top1.memory2.mem2[169][2] ;
 wire \top1.memory2.mem2[16][0] ;
 wire \top1.memory2.mem2[16][1] ;
 wire \top1.memory2.mem2[16][2] ;
 wire \top1.memory2.mem2[170][0] ;
 wire \top1.memory2.mem2[170][1] ;
 wire \top1.memory2.mem2[170][2] ;
 wire \top1.memory2.mem2[171][0] ;
 wire \top1.memory2.mem2[171][1] ;
 wire \top1.memory2.mem2[171][2] ;
 wire \top1.memory2.mem2[172][0] ;
 wire \top1.memory2.mem2[172][1] ;
 wire \top1.memory2.mem2[172][2] ;
 wire \top1.memory2.mem2[173][0] ;
 wire \top1.memory2.mem2[173][1] ;
 wire \top1.memory2.mem2[173][2] ;
 wire \top1.memory2.mem2[174][0] ;
 wire \top1.memory2.mem2[174][1] ;
 wire \top1.memory2.mem2[174][2] ;
 wire \top1.memory2.mem2[175][0] ;
 wire \top1.memory2.mem2[175][1] ;
 wire \top1.memory2.mem2[175][2] ;
 wire \top1.memory2.mem2[176][0] ;
 wire \top1.memory2.mem2[176][1] ;
 wire \top1.memory2.mem2[176][2] ;
 wire \top1.memory2.mem2[177][0] ;
 wire \top1.memory2.mem2[177][1] ;
 wire \top1.memory2.mem2[177][2] ;
 wire \top1.memory2.mem2[178][0] ;
 wire \top1.memory2.mem2[178][1] ;
 wire \top1.memory2.mem2[178][2] ;
 wire \top1.memory2.mem2[179][0] ;
 wire \top1.memory2.mem2[179][1] ;
 wire \top1.memory2.mem2[179][2] ;
 wire \top1.memory2.mem2[17][0] ;
 wire \top1.memory2.mem2[17][1] ;
 wire \top1.memory2.mem2[17][2] ;
 wire \top1.memory2.mem2[180][0] ;
 wire \top1.memory2.mem2[180][1] ;
 wire \top1.memory2.mem2[180][2] ;
 wire \top1.memory2.mem2[181][0] ;
 wire \top1.memory2.mem2[181][1] ;
 wire \top1.memory2.mem2[181][2] ;
 wire \top1.memory2.mem2[182][0] ;
 wire \top1.memory2.mem2[182][1] ;
 wire \top1.memory2.mem2[182][2] ;
 wire \top1.memory2.mem2[183][0] ;
 wire \top1.memory2.mem2[183][1] ;
 wire \top1.memory2.mem2[183][2] ;
 wire \top1.memory2.mem2[184][0] ;
 wire \top1.memory2.mem2[184][1] ;
 wire \top1.memory2.mem2[184][2] ;
 wire \top1.memory2.mem2[185][0] ;
 wire \top1.memory2.mem2[185][1] ;
 wire \top1.memory2.mem2[185][2] ;
 wire \top1.memory2.mem2[186][0] ;
 wire \top1.memory2.mem2[186][1] ;
 wire \top1.memory2.mem2[186][2] ;
 wire \top1.memory2.mem2[187][0] ;
 wire \top1.memory2.mem2[187][1] ;
 wire \top1.memory2.mem2[187][2] ;
 wire \top1.memory2.mem2[188][0] ;
 wire \top1.memory2.mem2[188][1] ;
 wire \top1.memory2.mem2[188][2] ;
 wire \top1.memory2.mem2[189][0] ;
 wire \top1.memory2.mem2[189][1] ;
 wire \top1.memory2.mem2[189][2] ;
 wire \top1.memory2.mem2[18][0] ;
 wire \top1.memory2.mem2[18][1] ;
 wire \top1.memory2.mem2[18][2] ;
 wire \top1.memory2.mem2[190][0] ;
 wire \top1.memory2.mem2[190][1] ;
 wire \top1.memory2.mem2[190][2] ;
 wire \top1.memory2.mem2[191][0] ;
 wire \top1.memory2.mem2[191][1] ;
 wire \top1.memory2.mem2[191][2] ;
 wire \top1.memory2.mem2[192][0] ;
 wire \top1.memory2.mem2[192][1] ;
 wire \top1.memory2.mem2[192][2] ;
 wire \top1.memory2.mem2[193][0] ;
 wire \top1.memory2.mem2[193][1] ;
 wire \top1.memory2.mem2[193][2] ;
 wire \top1.memory2.mem2[194][0] ;
 wire \top1.memory2.mem2[194][1] ;
 wire \top1.memory2.mem2[194][2] ;
 wire \top1.memory2.mem2[195][0] ;
 wire \top1.memory2.mem2[195][1] ;
 wire \top1.memory2.mem2[195][2] ;
 wire \top1.memory2.mem2[196][0] ;
 wire \top1.memory2.mem2[196][1] ;
 wire \top1.memory2.mem2[196][2] ;
 wire \top1.memory2.mem2[197][0] ;
 wire \top1.memory2.mem2[197][1] ;
 wire \top1.memory2.mem2[197][2] ;
 wire \top1.memory2.mem2[198][0] ;
 wire \top1.memory2.mem2[198][1] ;
 wire \top1.memory2.mem2[198][2] ;
 wire \top1.memory2.mem2[199][0] ;
 wire \top1.memory2.mem2[199][1] ;
 wire \top1.memory2.mem2[199][2] ;
 wire \top1.memory2.mem2[19][0] ;
 wire \top1.memory2.mem2[19][1] ;
 wire \top1.memory2.mem2[19][2] ;
 wire \top1.memory2.mem2[1][0] ;
 wire \top1.memory2.mem2[1][1] ;
 wire \top1.memory2.mem2[1][2] ;
 wire \top1.memory2.mem2[20][0] ;
 wire \top1.memory2.mem2[20][1] ;
 wire \top1.memory2.mem2[20][2] ;
 wire \top1.memory2.mem2[21][0] ;
 wire \top1.memory2.mem2[21][1] ;
 wire \top1.memory2.mem2[21][2] ;
 wire \top1.memory2.mem2[22][0] ;
 wire \top1.memory2.mem2[22][1] ;
 wire \top1.memory2.mem2[22][2] ;
 wire \top1.memory2.mem2[23][0] ;
 wire \top1.memory2.mem2[23][1] ;
 wire \top1.memory2.mem2[23][2] ;
 wire \top1.memory2.mem2[24][0] ;
 wire \top1.memory2.mem2[24][1] ;
 wire \top1.memory2.mem2[24][2] ;
 wire \top1.memory2.mem2[25][0] ;
 wire \top1.memory2.mem2[25][1] ;
 wire \top1.memory2.mem2[25][2] ;
 wire \top1.memory2.mem2[26][0] ;
 wire \top1.memory2.mem2[26][1] ;
 wire \top1.memory2.mem2[26][2] ;
 wire \top1.memory2.mem2[27][0] ;
 wire \top1.memory2.mem2[27][1] ;
 wire \top1.memory2.mem2[27][2] ;
 wire \top1.memory2.mem2[28][0] ;
 wire \top1.memory2.mem2[28][1] ;
 wire \top1.memory2.mem2[28][2] ;
 wire \top1.memory2.mem2[29][0] ;
 wire \top1.memory2.mem2[29][1] ;
 wire \top1.memory2.mem2[29][2] ;
 wire \top1.memory2.mem2[2][0] ;
 wire \top1.memory2.mem2[2][1] ;
 wire \top1.memory2.mem2[2][2] ;
 wire \top1.memory2.mem2[30][0] ;
 wire \top1.memory2.mem2[30][1] ;
 wire \top1.memory2.mem2[30][2] ;
 wire \top1.memory2.mem2[31][0] ;
 wire \top1.memory2.mem2[31][1] ;
 wire \top1.memory2.mem2[31][2] ;
 wire \top1.memory2.mem2[32][0] ;
 wire \top1.memory2.mem2[32][1] ;
 wire \top1.memory2.mem2[32][2] ;
 wire \top1.memory2.mem2[33][0] ;
 wire \top1.memory2.mem2[33][1] ;
 wire \top1.memory2.mem2[33][2] ;
 wire \top1.memory2.mem2[34][0] ;
 wire \top1.memory2.mem2[34][1] ;
 wire \top1.memory2.mem2[34][2] ;
 wire \top1.memory2.mem2[35][0] ;
 wire \top1.memory2.mem2[35][1] ;
 wire \top1.memory2.mem2[35][2] ;
 wire \top1.memory2.mem2[36][0] ;
 wire \top1.memory2.mem2[36][1] ;
 wire \top1.memory2.mem2[36][2] ;
 wire \top1.memory2.mem2[37][0] ;
 wire \top1.memory2.mem2[37][1] ;
 wire \top1.memory2.mem2[37][2] ;
 wire \top1.memory2.mem2[38][0] ;
 wire \top1.memory2.mem2[38][1] ;
 wire \top1.memory2.mem2[38][2] ;
 wire \top1.memory2.mem2[39][0] ;
 wire \top1.memory2.mem2[39][1] ;
 wire \top1.memory2.mem2[39][2] ;
 wire \top1.memory2.mem2[3][0] ;
 wire \top1.memory2.mem2[3][1] ;
 wire \top1.memory2.mem2[3][2] ;
 wire \top1.memory2.mem2[40][0] ;
 wire \top1.memory2.mem2[40][1] ;
 wire \top1.memory2.mem2[40][2] ;
 wire \top1.memory2.mem2[41][0] ;
 wire \top1.memory2.mem2[41][1] ;
 wire \top1.memory2.mem2[41][2] ;
 wire \top1.memory2.mem2[42][0] ;
 wire \top1.memory2.mem2[42][1] ;
 wire \top1.memory2.mem2[42][2] ;
 wire \top1.memory2.mem2[43][0] ;
 wire \top1.memory2.mem2[43][1] ;
 wire \top1.memory2.mem2[43][2] ;
 wire \top1.memory2.mem2[44][0] ;
 wire \top1.memory2.mem2[44][1] ;
 wire \top1.memory2.mem2[44][2] ;
 wire \top1.memory2.mem2[45][0] ;
 wire \top1.memory2.mem2[45][1] ;
 wire \top1.memory2.mem2[45][2] ;
 wire \top1.memory2.mem2[46][0] ;
 wire \top1.memory2.mem2[46][1] ;
 wire \top1.memory2.mem2[46][2] ;
 wire \top1.memory2.mem2[47][0] ;
 wire \top1.memory2.mem2[47][1] ;
 wire \top1.memory2.mem2[47][2] ;
 wire \top1.memory2.mem2[48][0] ;
 wire \top1.memory2.mem2[48][1] ;
 wire \top1.memory2.mem2[48][2] ;
 wire \top1.memory2.mem2[49][0] ;
 wire \top1.memory2.mem2[49][1] ;
 wire \top1.memory2.mem2[49][2] ;
 wire \top1.memory2.mem2[4][0] ;
 wire \top1.memory2.mem2[4][1] ;
 wire \top1.memory2.mem2[4][2] ;
 wire \top1.memory2.mem2[50][0] ;
 wire \top1.memory2.mem2[50][1] ;
 wire \top1.memory2.mem2[50][2] ;
 wire \top1.memory2.mem2[51][0] ;
 wire \top1.memory2.mem2[51][1] ;
 wire \top1.memory2.mem2[51][2] ;
 wire \top1.memory2.mem2[52][0] ;
 wire \top1.memory2.mem2[52][1] ;
 wire \top1.memory2.mem2[52][2] ;
 wire \top1.memory2.mem2[53][0] ;
 wire \top1.memory2.mem2[53][1] ;
 wire \top1.memory2.mem2[53][2] ;
 wire \top1.memory2.mem2[54][0] ;
 wire \top1.memory2.mem2[54][1] ;
 wire \top1.memory2.mem2[54][2] ;
 wire \top1.memory2.mem2[55][0] ;
 wire \top1.memory2.mem2[55][1] ;
 wire \top1.memory2.mem2[55][2] ;
 wire \top1.memory2.mem2[56][0] ;
 wire \top1.memory2.mem2[56][1] ;
 wire \top1.memory2.mem2[56][2] ;
 wire \top1.memory2.mem2[57][0] ;
 wire \top1.memory2.mem2[57][1] ;
 wire \top1.memory2.mem2[57][2] ;
 wire \top1.memory2.mem2[58][0] ;
 wire \top1.memory2.mem2[58][1] ;
 wire \top1.memory2.mem2[58][2] ;
 wire \top1.memory2.mem2[59][0] ;
 wire \top1.memory2.mem2[59][1] ;
 wire \top1.memory2.mem2[59][2] ;
 wire \top1.memory2.mem2[5][0] ;
 wire \top1.memory2.mem2[5][1] ;
 wire \top1.memory2.mem2[5][2] ;
 wire \top1.memory2.mem2[60][0] ;
 wire \top1.memory2.mem2[60][1] ;
 wire \top1.memory2.mem2[60][2] ;
 wire \top1.memory2.mem2[61][0] ;
 wire \top1.memory2.mem2[61][1] ;
 wire \top1.memory2.mem2[61][2] ;
 wire \top1.memory2.mem2[62][0] ;
 wire \top1.memory2.mem2[62][1] ;
 wire \top1.memory2.mem2[62][2] ;
 wire \top1.memory2.mem2[63][0] ;
 wire \top1.memory2.mem2[63][1] ;
 wire \top1.memory2.mem2[63][2] ;
 wire \top1.memory2.mem2[64][0] ;
 wire \top1.memory2.mem2[64][1] ;
 wire \top1.memory2.mem2[64][2] ;
 wire \top1.memory2.mem2[65][0] ;
 wire \top1.memory2.mem2[65][1] ;
 wire \top1.memory2.mem2[65][2] ;
 wire \top1.memory2.mem2[66][0] ;
 wire \top1.memory2.mem2[66][1] ;
 wire \top1.memory2.mem2[66][2] ;
 wire \top1.memory2.mem2[67][0] ;
 wire \top1.memory2.mem2[67][1] ;
 wire \top1.memory2.mem2[67][2] ;
 wire \top1.memory2.mem2[68][0] ;
 wire \top1.memory2.mem2[68][1] ;
 wire \top1.memory2.mem2[68][2] ;
 wire \top1.memory2.mem2[69][0] ;
 wire \top1.memory2.mem2[69][1] ;
 wire \top1.memory2.mem2[69][2] ;
 wire \top1.memory2.mem2[6][0] ;
 wire \top1.memory2.mem2[6][1] ;
 wire \top1.memory2.mem2[6][2] ;
 wire \top1.memory2.mem2[70][0] ;
 wire \top1.memory2.mem2[70][1] ;
 wire \top1.memory2.mem2[70][2] ;
 wire \top1.memory2.mem2[71][0] ;
 wire \top1.memory2.mem2[71][1] ;
 wire \top1.memory2.mem2[71][2] ;
 wire \top1.memory2.mem2[72][0] ;
 wire \top1.memory2.mem2[72][1] ;
 wire \top1.memory2.mem2[72][2] ;
 wire \top1.memory2.mem2[73][0] ;
 wire \top1.memory2.mem2[73][1] ;
 wire \top1.memory2.mem2[73][2] ;
 wire \top1.memory2.mem2[74][0] ;
 wire \top1.memory2.mem2[74][1] ;
 wire \top1.memory2.mem2[74][2] ;
 wire \top1.memory2.mem2[75][0] ;
 wire \top1.memory2.mem2[75][1] ;
 wire \top1.memory2.mem2[75][2] ;
 wire \top1.memory2.mem2[76][0] ;
 wire \top1.memory2.mem2[76][1] ;
 wire \top1.memory2.mem2[76][2] ;
 wire \top1.memory2.mem2[77][0] ;
 wire \top1.memory2.mem2[77][1] ;
 wire \top1.memory2.mem2[77][2] ;
 wire \top1.memory2.mem2[78][0] ;
 wire \top1.memory2.mem2[78][1] ;
 wire \top1.memory2.mem2[78][2] ;
 wire \top1.memory2.mem2[79][0] ;
 wire \top1.memory2.mem2[79][1] ;
 wire \top1.memory2.mem2[79][2] ;
 wire \top1.memory2.mem2[7][0] ;
 wire \top1.memory2.mem2[7][1] ;
 wire \top1.memory2.mem2[7][2] ;
 wire \top1.memory2.mem2[80][0] ;
 wire \top1.memory2.mem2[80][1] ;
 wire \top1.memory2.mem2[80][2] ;
 wire \top1.memory2.mem2[81][0] ;
 wire \top1.memory2.mem2[81][1] ;
 wire \top1.memory2.mem2[81][2] ;
 wire \top1.memory2.mem2[82][0] ;
 wire \top1.memory2.mem2[82][1] ;
 wire \top1.memory2.mem2[82][2] ;
 wire \top1.memory2.mem2[83][0] ;
 wire \top1.memory2.mem2[83][1] ;
 wire \top1.memory2.mem2[83][2] ;
 wire \top1.memory2.mem2[84][0] ;
 wire \top1.memory2.mem2[84][1] ;
 wire \top1.memory2.mem2[84][2] ;
 wire \top1.memory2.mem2[85][0] ;
 wire \top1.memory2.mem2[85][1] ;
 wire \top1.memory2.mem2[85][2] ;
 wire \top1.memory2.mem2[86][0] ;
 wire \top1.memory2.mem2[86][1] ;
 wire \top1.memory2.mem2[86][2] ;
 wire \top1.memory2.mem2[87][0] ;
 wire \top1.memory2.mem2[87][1] ;
 wire \top1.memory2.mem2[87][2] ;
 wire \top1.memory2.mem2[88][0] ;
 wire \top1.memory2.mem2[88][1] ;
 wire \top1.memory2.mem2[88][2] ;
 wire \top1.memory2.mem2[89][0] ;
 wire \top1.memory2.mem2[89][1] ;
 wire \top1.memory2.mem2[89][2] ;
 wire \top1.memory2.mem2[8][0] ;
 wire \top1.memory2.mem2[8][1] ;
 wire \top1.memory2.mem2[8][2] ;
 wire \top1.memory2.mem2[90][0] ;
 wire \top1.memory2.mem2[90][1] ;
 wire \top1.memory2.mem2[90][2] ;
 wire \top1.memory2.mem2[91][0] ;
 wire \top1.memory2.mem2[91][1] ;
 wire \top1.memory2.mem2[91][2] ;
 wire \top1.memory2.mem2[92][0] ;
 wire \top1.memory2.mem2[92][1] ;
 wire \top1.memory2.mem2[92][2] ;
 wire \top1.memory2.mem2[93][0] ;
 wire \top1.memory2.mem2[93][1] ;
 wire \top1.memory2.mem2[93][2] ;
 wire \top1.memory2.mem2[94][0] ;
 wire \top1.memory2.mem2[94][1] ;
 wire \top1.memory2.mem2[94][2] ;
 wire \top1.memory2.mem2[95][0] ;
 wire \top1.memory2.mem2[95][1] ;
 wire \top1.memory2.mem2[95][2] ;
 wire \top1.memory2.mem2[96][0] ;
 wire \top1.memory2.mem2[96][1] ;
 wire \top1.memory2.mem2[96][2] ;
 wire \top1.memory2.mem2[97][0] ;
 wire \top1.memory2.mem2[97][1] ;
 wire \top1.memory2.mem2[97][2] ;
 wire \top1.memory2.mem2[98][0] ;
 wire \top1.memory2.mem2[98][1] ;
 wire \top1.memory2.mem2[98][2] ;
 wire \top1.memory2.mem2[99][0] ;
 wire \top1.memory2.mem2[99][1] ;
 wire \top1.memory2.mem2[99][2] ;
 wire \top1.memory2.mem2[9][0] ;
 wire \top1.memory2.mem2[9][1] ;
 wire \top1.memory2.mem2[9][2] ;
 wire \top1.mux.data_out ;
 wire \top1.piso_time_reg.register[0] ;
 wire \top1.piso_time_reg.register[10] ;
 wire \top1.piso_time_reg.register[11] ;
 wire \top1.piso_time_reg.register[12] ;
 wire \top1.piso_time_reg.register[13] ;
 wire \top1.piso_time_reg.register[14] ;
 wire \top1.piso_time_reg.register[15] ;
 wire \top1.piso_time_reg.register[16] ;
 wire \top1.piso_time_reg.register[17] ;
 wire \top1.piso_time_reg.register[18] ;
 wire \top1.piso_time_reg.register[19] ;
 wire \top1.piso_time_reg.register[1] ;
 wire \top1.piso_time_reg.register[20] ;
 wire \top1.piso_time_reg.register[21] ;
 wire \top1.piso_time_reg.register[22] ;
 wire \top1.piso_time_reg.register[23] ;
 wire \top1.piso_time_reg.register[24] ;
 wire \top1.piso_time_reg.register[25] ;
 wire \top1.piso_time_reg.register[26] ;
 wire \top1.piso_time_reg.register[27] ;
 wire \top1.piso_time_reg.register[28] ;
 wire \top1.piso_time_reg.register[29] ;
 wire \top1.piso_time_reg.register[2] ;
 wire \top1.piso_time_reg.register[30] ;
 wire \top1.piso_time_reg.register[3] ;
 wire \top1.piso_time_reg.register[4] ;
 wire \top1.piso_time_reg.register[5] ;
 wire \top1.piso_time_reg.register[6] ;
 wire \top1.piso_time_reg.register[7] ;
 wire \top1.piso_time_reg.register[8] ;
 wire \top1.piso_time_reg.register[9] ;
 wire \top1.reg1.register[0] ;
 wire \top1.reg1.register[1] ;
 wire \top1.reg2.register[0] ;
 wire \top1.reg2.register[1] ;
 wire \top1.reg2.serial_out ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6203;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net6319;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6325;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;
 wire net6619;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6623;
 wire net6624;
 wire net6625;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6629;
 wire net6630;
 wire net6631;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6638;
 wire net6639;
 wire net6640;
 wire net6641;
 wire net6642;
 wire net6643;
 wire net6644;
 wire net6645;
 wire net6646;
 wire net6647;
 wire net6648;
 wire net6649;
 wire net6650;
 wire net6651;
 wire net6652;
 wire net6653;
 wire net6654;
 wire net6655;
 wire net6656;
 wire net6657;
 wire net6658;
 wire net6659;
 wire net6660;
 wire net6661;
 wire net6662;
 wire net6663;
 wire net6664;
 wire net6665;
 wire net6666;
 wire net6667;
 wire net6668;
 wire net6669;
 wire net6670;
 wire net6671;
 wire net6672;
 wire net6673;
 wire net6674;
 wire net6675;
 wire net6676;
 wire net6677;
 wire net6678;
 wire net6679;
 wire net6680;
 wire net6681;
 wire net6682;
 wire net6683;
 wire net6684;
 wire net6685;
 wire net6686;
 wire net6687;
 wire net6688;
 wire net6689;
 wire net6690;
 wire net6691;
 wire net6692;
 wire net6693;
 wire net6694;
 wire net6695;
 wire net6696;
 wire net6697;
 wire net6698;
 wire net6699;
 wire net6700;
 wire net6701;
 wire net6702;
 wire net6703;
 wire net6704;
 wire net6705;
 wire net6706;
 wire net6707;
 wire net6708;
 wire net6709;
 wire net6710;
 wire net6711;
 wire net6712;
 wire net6713;
 wire net6714;
 wire net6715;
 wire net6716;
 wire net6717;
 wire net6718;
 wire net6719;
 wire net6720;
 wire net6721;
 wire net6722;
 wire net6723;
 wire net6724;
 wire net6725;
 wire net6726;
 wire net6727;
 wire net6728;
 wire net6729;
 wire net6730;
 wire net6731;
 wire net6732;
 wire net6733;
 wire net6734;
 wire net6735;
 wire net6736;
 wire net6737;
 wire net6738;
 wire net6739;
 wire net6740;
 wire net6741;
 wire net6742;
 wire net6743;
 wire net6744;
 wire net6745;
 wire net6746;
 wire net6747;
 wire net6748;
 wire net6749;
 wire net6750;
 wire net6751;
 wire net6752;
 wire net6753;
 wire net6754;
 wire net6755;
 wire net6756;
 wire net6757;
 wire net6758;
 wire net6759;
 wire net6760;
 wire net6761;
 wire net6762;
 wire net6763;
 wire net6764;
 wire net6765;
 wire net6766;
 wire net6767;
 wire net6768;
 wire net6769;
 wire net6770;
 wire net6771;
 wire net6772;
 wire net6773;
 wire net6774;
 wire net6775;
 wire net6776;
 wire net6777;
 wire net6778;
 wire net6779;
 wire net6780;
 wire net6781;
 wire net6782;
 wire net6783;
 wire net6784;
 wire net6785;
 wire net6786;
 wire net6787;
 wire net6788;
 wire net6789;
 wire net6790;
 wire net6791;
 wire net6792;
 wire net6793;
 wire net6794;
 wire net6795;
 wire net6796;
 wire net6797;
 wire net6798;
 wire net6799;
 wire net6800;
 wire net6801;
 wire net6802;
 wire net6803;
 wire net6804;
 wire net6805;
 wire net6806;
 wire net6807;
 wire net6808;
 wire net6809;
 wire net6810;
 wire net6811;
 wire net6812;
 wire net6813;
 wire net6814;
 wire net6815;
 wire net6816;
 wire net6817;
 wire net6818;
 wire net6819;
 wire net6820;
 wire net6821;
 wire net6822;
 wire net6823;
 wire net6824;
 wire net6825;
 wire net6826;
 wire net6827;
 wire net6828;
 wire net6829;
 wire net6830;
 wire net6831;
 wire net6832;
 wire net6833;
 wire net6834;
 wire net6835;
 wire net6836;
 wire net6837;
 wire net6838;
 wire net6839;
 wire net6840;
 wire net6841;
 wire net6842;
 wire net6843;
 wire net6844;
 wire net6845;
 wire net6846;
 wire net6847;
 wire net6848;
 wire net6849;
 wire net6850;
 wire net6851;
 wire net6852;
 wire net6853;
 wire net6854;
 wire net6855;
 wire net6856;
 wire net6857;
 wire net6858;
 wire net6859;
 wire net6860;
 wire net6861;
 wire net6862;
 wire net6863;
 wire net6864;
 wire net6865;
 wire net6866;
 wire net6867;
 wire net6868;
 wire net6869;
 wire net6870;
 wire net6871;
 wire net6872;
 wire net6873;
 wire net6874;
 wire net6875;
 wire net6876;
 wire net6877;
 wire net6878;
 wire net6879;
 wire net6880;
 wire net6881;
 wire net6882;
 wire net6883;
 wire net6884;
 wire net6885;
 wire net6886;
 wire net6887;
 wire net6888;
 wire net6889;
 wire net6890;
 wire net6891;
 wire net6892;
 wire net6893;
 wire net6894;
 wire net6895;
 wire net6896;
 wire net6897;
 wire net6898;
 wire net6899;
 wire net6900;
 wire net6901;
 wire net6902;
 wire net6903;
 wire net6904;
 wire net6905;
 wire net6906;
 wire net6907;
 wire net6908;
 wire net6909;
 wire net6910;
 wire net6911;
 wire net6912;
 wire net6913;
 wire net6914;
 wire net6915;
 wire net6916;
 wire net6917;
 wire net6918;
 wire net6919;
 wire net6920;
 wire net6921;
 wire net6922;
 wire net6923;
 wire net6924;
 wire net6925;
 wire net6926;
 wire net6927;
 wire net6928;
 wire net6929;
 wire net6930;
 wire net6931;
 wire net6932;
 wire net6933;
 wire net6934;
 wire net6935;
 wire net6936;
 wire net6937;
 wire net6938;
 wire net6939;
 wire net6940;
 wire net6941;
 wire net6942;
 wire net6943;
 wire net6944;
 wire net6945;
 wire net6946;
 wire net6947;
 wire net6948;
 wire net6949;
 wire net6950;
 wire net6951;
 wire net6952;
 wire net6953;
 wire net6954;
 wire net6955;
 wire net6956;
 wire net6957;
 wire net6958;
 wire net6959;
 wire net6960;
 wire net6961;
 wire net6962;
 wire net6963;
 wire net6964;
 wire net6965;
 wire net6966;
 wire net6967;
 wire net6968;
 wire net6969;
 wire net6970;
 wire net6971;
 wire net6972;
 wire net6973;
 wire net6974;
 wire net6975;
 wire net6976;
 wire net6977;
 wire net6978;
 wire net6979;
 wire net6980;
 wire net6981;
 wire net6982;
 wire net6983;
 wire net6984;
 wire net6985;
 wire net6986;
 wire net6987;
 wire net6988;
 wire net6989;
 wire net6990;
 wire net6991;
 wire net6992;
 wire net6993;
 wire net6994;
 wire net6995;
 wire net6996;
 wire net6997;
 wire net6998;
 wire net6999;
 wire net7000;
 wire net7001;
 wire net7002;
 wire net7003;
 wire net7004;
 wire net7005;
 wire net7006;
 wire net7007;
 wire net7008;
 wire net7009;
 wire net7010;
 wire net7011;
 wire net7012;
 wire net7013;
 wire net7014;
 wire net7015;
 wire net7016;
 wire net7017;
 wire net7018;
 wire net7019;
 wire net7020;
 wire net7021;
 wire net7022;
 wire net7023;
 wire net7024;
 wire net7025;
 wire net7026;
 wire net7027;
 wire net7028;
 wire net7029;
 wire net7030;
 wire net7031;
 wire net7032;
 wire net7033;
 wire net7034;
 wire net7035;
 wire net7036;
 wire net7037;
 wire net7038;
 wire net7039;
 wire net7040;
 wire net7041;
 wire net7042;
 wire net7043;
 wire net7044;
 wire net7045;
 wire net7046;
 wire net7047;
 wire net7048;
 wire net7049;
 wire net7050;
 wire net7051;
 wire net7052;
 wire net7053;
 wire net7054;
 wire net7055;
 wire net7056;
 wire net7057;
 wire net7058;
 wire net7059;
 wire net7060;
 wire net7061;
 wire net7062;
 wire net7063;
 wire net7064;
 wire net7065;
 wire net7066;
 wire net7067;
 wire net7068;
 wire net7069;
 wire net7070;
 wire net7071;
 wire net7072;
 wire net7073;
 wire net7074;
 wire net7075;
 wire net7076;
 wire net7077;
 wire net7078;
 wire net7079;
 wire net7080;
 wire net7081;
 wire net7082;
 wire net7083;
 wire net7084;
 wire net7085;
 wire net7086;
 wire net7087;
 wire net7088;
 wire net7089;
 wire net7090;
 wire net7091;
 wire net7092;
 wire net7093;
 wire net7094;
 wire net7095;
 wire net7096;
 wire net7097;
 wire net7098;
 wire net7099;
 wire net7100;
 wire net7101;
 wire net7102;
 wire net7103;
 wire net7104;
 wire net7105;
 wire net7106;
 wire net7107;
 wire net7108;
 wire net7109;
 wire net7110;
 wire net7111;
 wire net7112;
 wire net7113;
 wire net7114;
 wire net7115;
 wire net7116;
 wire net7117;
 wire net7118;
 wire net7119;
 wire net7120;
 wire net7121;
 wire net7122;
 wire net7123;
 wire net7124;
 wire net7125;
 wire net7126;
 wire net7127;
 wire net7128;
 wire net7129;
 wire net7130;
 wire net7131;
 wire net7132;
 wire net7133;
 wire net7134;
 wire net7135;
 wire net7136;
 wire net7137;
 wire net7138;
 wire net7139;
 wire net7140;
 wire net7141;
 wire net7142;
 wire net7143;
 wire net7144;
 wire net7145;
 wire net7146;
 wire net7147;
 wire net7148;
 wire net7149;
 wire net7150;
 wire net7151;
 wire net7152;
 wire net7153;
 wire net7154;
 wire net7155;
 wire net7156;
 wire net7157;
 wire net7158;
 wire net7159;
 wire net7160;
 wire net7161;
 wire net7162;
 wire net7163;
 wire net7164;
 wire net7165;
 wire net7166;
 wire net7167;
 wire net7168;
 wire net7169;
 wire net7170;
 wire net7171;
 wire net7172;
 wire net7173;
 wire net7174;
 wire net7175;
 wire net7176;
 wire net7177;
 wire net7178;
 wire net7179;
 wire net7180;
 wire net7181;
 wire net7182;
 wire net7183;
 wire net7184;
 wire net7185;
 wire net7186;
 wire net7187;
 wire net7188;
 wire net7189;
 wire net7190;
 wire net7191;
 wire net7192;
 wire net7193;
 wire net7194;
 wire net7195;
 wire net7196;
 wire net7197;
 wire net7198;
 wire net7199;
 wire net7200;
 wire net7201;
 wire net7202;
 wire net7203;
 wire net7204;
 wire net7205;
 wire net7206;
 wire net7207;
 wire net7208;
 wire net7209;
 wire net7210;
 wire net7211;
 wire net7212;
 wire net7213;
 wire net7214;
 wire net7215;
 wire net7216;
 wire net7217;
 wire net7218;
 wire net7219;
 wire net7220;
 wire net7221;
 wire net7222;
 wire net7223;
 wire net7224;
 wire net7225;
 wire net7226;
 wire net7227;
 wire net7228;
 wire net7229;
 wire net7230;
 wire net7231;
 wire net7232;
 wire net7233;
 wire net7234;
 wire net7235;
 wire net7236;
 wire net7237;
 wire net7238;
 wire net7239;
 wire net7240;
 wire net7241;
 wire net7242;
 wire net7243;
 wire net7244;
 wire net7245;
 wire net7246;
 wire net7247;
 wire net7248;
 wire net7249;
 wire net7250;
 wire net7251;
 wire net7252;
 wire net7253;
 wire net7254;
 wire net7255;
 wire net7256;
 wire net7257;
 wire net7258;
 wire net7259;
 wire net7260;
 wire net7261;
 wire net7262;
 wire net7263;
 wire net7264;
 wire net7265;
 wire net7266;
 wire net7267;
 wire net7268;
 wire net7269;
 wire net7270;
 wire net7271;
 wire net7272;
 wire net7273;
 wire net7274;
 wire net7275;
 wire net7276;
 wire net7277;
 wire net7278;
 wire net7279;
 wire net7280;
 wire net7281;
 wire net7282;
 wire net7283;
 wire net7284;
 wire net7285;
 wire net7286;
 wire net7287;
 wire net7288;
 wire net7289;
 wire net7290;
 wire net7291;
 wire net7292;
 wire net7293;
 wire net7294;
 wire net7295;
 wire net7296;
 wire net7297;
 wire net7298;
 wire net7299;
 wire net7300;
 wire net7301;
 wire net7302;
 wire net7303;
 wire net7304;
 wire net7305;
 wire net7306;
 wire net7307;
 wire net7308;
 wire net7309;
 wire net7310;
 wire net7311;
 wire net7312;
 wire net7313;
 wire net7314;
 wire net7315;
 wire net7316;
 wire net7317;
 wire net7318;
 wire net7319;
 wire net7320;
 wire net7321;
 wire net7322;
 wire net7323;
 wire net7324;
 wire net7325;
 wire net7326;
 wire net7327;
 wire net7328;
 wire net7329;
 wire net7330;
 wire net7331;
 wire net7332;
 wire net7333;
 wire net7334;
 wire net7335;
 wire net7336;
 wire net7337;
 wire net7338;
 wire net7339;
 wire net7340;
 wire net7341;
 wire net7342;
 wire net7343;
 wire net7344;
 wire net7345;
 wire net7346;
 wire net7347;
 wire net7348;
 wire net7349;
 wire net7350;
 wire net7351;
 wire net7352;
 wire net7353;
 wire net7354;
 wire net7355;
 wire net7356;
 wire net7357;
 wire net7358;
 wire net7359;
 wire net7360;
 wire net7361;
 wire net7362;
 wire net7363;
 wire net7364;
 wire net7365;
 wire net7366;
 wire net7367;
 wire net7368;
 wire net7369;
 wire net7370;
 wire net7371;
 wire net7372;
 wire net7373;
 wire net7374;
 wire net7375;
 wire net7376;
 wire net7377;
 wire net7378;
 wire net7379;
 wire net7380;
 wire net7381;
 wire net7382;
 wire net7383;
 wire net7384;
 wire net7385;
 wire net7386;
 wire net7387;
 wire net7388;
 wire net7389;
 wire net7390;
 wire net7391;
 wire net7392;
 wire net7393;
 wire net7394;
 wire net7395;
 wire net7396;
 wire net7397;
 wire net7398;
 wire net7399;
 wire net7400;
 wire net7401;
 wire net7402;
 wire net7403;
 wire net7404;
 wire net7405;
 wire net7406;
 wire net7407;
 wire net7408;
 wire net7409;
 wire net7410;
 wire net7411;
 wire net7412;
 wire net7413;
 wire net7414;
 wire net7415;
 wire net7416;
 wire net7417;
 wire net7418;
 wire net7419;
 wire net7420;
 wire net7421;
 wire net7422;
 wire net7423;
 wire net7424;
 wire net7425;
 wire net7426;
 wire net7427;
 wire net7428;
 wire net7429;
 wire net7430;
 wire net7431;
 wire net7432;
 wire net7433;
 wire net7434;
 wire net7435;
 wire net7436;
 wire net7437;
 wire net7438;
 wire net7439;
 wire net7440;
 wire net7441;
 wire net7442;
 wire net7443;
 wire net7444;
 wire net7445;
 wire net7446;
 wire net7447;
 wire net7448;
 wire net7449;
 wire net7450;
 wire net7451;
 wire net7452;
 wire net7453;
 wire net7454;
 wire net7455;
 wire net7456;
 wire net7457;
 wire net7458;
 wire net7459;
 wire net7460;
 wire net7461;
 wire net7462;
 wire net7463;
 wire net7464;
 wire net7465;
 wire net7466;
 wire net7467;
 wire net7468;
 wire net7469;
 wire net7470;
 wire net7471;
 wire net7472;
 wire net7473;
 wire net7474;
 wire net7475;
 wire net7476;
 wire net7477;
 wire net7478;
 wire net7479;
 wire net7480;
 wire net7481;
 wire net7482;
 wire net7483;
 wire net7484;
 wire net7485;
 wire net7486;
 wire net7487;
 wire net7488;
 wire net7489;
 wire net7490;
 wire net7491;
 wire net7492;
 wire net7493;
 wire net7494;
 wire net7495;
 wire net7496;
 wire net7497;
 wire net7498;
 wire net7499;
 wire net7500;
 wire net7501;
 wire net7502;
 wire net7503;
 wire net7504;
 wire net7505;
 wire net7506;
 wire net7507;
 wire net7508;
 wire net7509;
 wire net7510;
 wire net7511;
 wire net7512;
 wire net7513;
 wire net7514;
 wire net7515;
 wire net7516;
 wire net7517;
 wire net7518;
 wire net7519;
 wire net7520;
 wire net7521;
 wire net7522;
 wire net7523;
 wire net7524;
 wire net7525;
 wire net7526;
 wire net7527;
 wire net7528;
 wire net7529;
 wire net7530;
 wire net7531;
 wire net7532;
 wire net7533;
 wire net7534;
 wire net7535;
 wire net7536;
 wire net7537;
 wire net7538;
 wire net7539;
 wire net7540;
 wire net7541;
 wire net7542;
 wire net7543;
 wire net7544;
 wire net7545;
 wire net7546;
 wire net7547;
 wire net7548;
 wire net7549;
 wire net7550;
 wire net7551;
 wire net7552;
 wire net7553;
 wire net7554;
 wire net7555;
 wire net7556;
 wire net7557;
 wire net7558;
 wire net7559;
 wire net7560;
 wire net7561;
 wire net7562;
 wire net7563;
 wire net7564;
 wire net7565;
 wire net7566;
 wire net7567;
 wire net7568;
 wire net7569;
 wire net7570;
 wire net7571;
 wire net7572;
 wire net7573;
 wire net7574;
 wire net7575;
 wire net7576;
 wire net7577;
 wire net7578;
 wire net7579;
 wire net7580;
 wire net7581;
 wire net7582;
 wire net7583;
 wire net7584;
 wire net7585;
 wire net7586;
 wire net7587;
 wire net7588;
 wire net7589;
 wire net7590;
 wire net7591;
 wire net7592;
 wire net7593;
 wire net7594;
 wire net7595;
 wire net7596;
 wire net7597;
 wire net7598;
 wire net7599;
 wire net7600;
 wire net7601;
 wire net7602;
 wire net7603;
 wire net7604;
 wire net7605;
 wire net7606;
 wire net7607;
 wire net7608;
 wire net7609;
 wire net7610;
 wire net7611;
 wire net7612;
 wire net7613;
 wire net7614;
 wire net7615;
 wire net7616;
 wire net7617;
 wire net7618;
 wire net7619;
 wire net7620;
 wire net7621;
 wire net7622;
 wire net7623;
 wire net7624;
 wire net7625;
 wire net7626;
 wire net7627;
 wire net7628;
 wire net7629;
 wire net7630;
 wire net7631;
 wire net7632;
 wire net7633;
 wire net7634;
 wire net7635;
 wire net7636;
 wire net7637;
 wire net7638;
 wire net7639;
 wire net7640;
 wire net7641;
 wire net7642;
 wire net7643;
 wire net7644;
 wire net7645;
 wire net7646;
 wire net7647;
 wire net7648;
 wire net7649;
 wire net7650;
 wire net7651;
 wire net7652;
 wire net7653;
 wire net7654;
 wire net7655;
 wire net7656;
 wire net7657;
 wire net7658;
 wire net7659;
 wire net7660;
 wire net7661;
 wire net7662;
 wire net7663;
 wire net7664;
 wire net7665;
 wire net7666;
 wire net7667;
 wire net7668;
 wire net7669;
 wire net7670;
 wire net7671;
 wire net7672;
 wire net7673;
 wire net7674;
 wire net7675;
 wire net7676;
 wire net7677;
 wire net7678;
 wire net7679;
 wire net7680;
 wire net7681;
 wire net7682;
 wire net7683;
 wire net7684;
 wire net7685;
 wire net7686;
 wire net7687;
 wire net7688;
 wire net7689;
 wire net7690;
 wire net7691;
 wire net7692;
 wire net7693;
 wire net7694;
 wire net7695;
 wire net7696;
 wire net7697;
 wire net7698;
 wire net7699;
 wire net7700;
 wire net7701;
 wire net7702;
 wire net7703;
 wire net7704;
 wire net7705;
 wire net7706;
 wire net7707;
 wire net7708;
 wire net7709;
 wire net7710;
 wire net7711;
 wire net7712;
 wire net7713;
 wire net7714;
 wire net7715;
 wire net7716;
 wire net7717;
 wire net7718;
 wire net7719;
 wire net7720;
 wire net7721;
 wire net7722;
 wire net7723;
 wire net7724;
 wire net7725;
 wire net7726;
 wire net7727;
 wire net7728;
 wire net7729;
 wire net7730;
 wire net7731;
 wire net7732;
 wire net7733;
 wire net7734;
 wire net7735;
 wire net7736;
 wire net7737;
 wire net7738;
 wire net7739;
 wire net7740;
 wire net7741;
 wire net7742;
 wire net7743;
 wire net7744;
 wire net7745;
 wire net7746;
 wire net7747;
 wire net7748;
 wire net7749;
 wire net7750;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire \clknet_leaf_1_top1.acquisition_clk ;
 wire \clknet_leaf_2_top1.acquisition_clk ;
 wire \clknet_leaf_3_top1.acquisition_clk ;
 wire \clknet_leaf_4_top1.acquisition_clk ;
 wire \clknet_leaf_5_top1.acquisition_clk ;
 wire \clknet_leaf_6_top1.acquisition_clk ;
 wire \clknet_leaf_7_top1.acquisition_clk ;
 wire \clknet_leaf_8_top1.acquisition_clk ;
 wire \clknet_leaf_9_top1.acquisition_clk ;
 wire \clknet_leaf_10_top1.acquisition_clk ;
 wire \clknet_leaf_11_top1.acquisition_clk ;
 wire \clknet_leaf_12_top1.acquisition_clk ;
 wire \clknet_leaf_13_top1.acquisition_clk ;
 wire \clknet_leaf_14_top1.acquisition_clk ;
 wire \clknet_leaf_15_top1.acquisition_clk ;
 wire \clknet_leaf_16_top1.acquisition_clk ;
 wire \clknet_leaf_17_top1.acquisition_clk ;
 wire \clknet_leaf_18_top1.acquisition_clk ;
 wire \clknet_leaf_19_top1.acquisition_clk ;
 wire \clknet_leaf_20_top1.acquisition_clk ;
 wire \clknet_leaf_21_top1.acquisition_clk ;
 wire \clknet_leaf_22_top1.acquisition_clk ;
 wire \clknet_leaf_23_top1.acquisition_clk ;
 wire \clknet_leaf_24_top1.acquisition_clk ;
 wire \clknet_leaf_25_top1.acquisition_clk ;
 wire \clknet_leaf_26_top1.acquisition_clk ;
 wire \clknet_leaf_27_top1.acquisition_clk ;
 wire \clknet_leaf_28_top1.acquisition_clk ;
 wire \clknet_leaf_29_top1.acquisition_clk ;
 wire \clknet_leaf_30_top1.acquisition_clk ;
 wire \clknet_leaf_31_top1.acquisition_clk ;
 wire \clknet_leaf_32_top1.acquisition_clk ;
 wire \clknet_leaf_33_top1.acquisition_clk ;
 wire \clknet_leaf_34_top1.acquisition_clk ;
 wire \clknet_leaf_35_top1.acquisition_clk ;
 wire \clknet_leaf_36_top1.acquisition_clk ;
 wire \clknet_leaf_37_top1.acquisition_clk ;
 wire \clknet_leaf_38_top1.acquisition_clk ;
 wire \clknet_leaf_39_top1.acquisition_clk ;
 wire \clknet_leaf_40_top1.acquisition_clk ;
 wire \clknet_leaf_41_top1.acquisition_clk ;
 wire \clknet_leaf_42_top1.acquisition_clk ;
 wire \clknet_leaf_43_top1.acquisition_clk ;
 wire \clknet_leaf_44_top1.acquisition_clk ;
 wire \clknet_leaf_45_top1.acquisition_clk ;
 wire \clknet_leaf_46_top1.acquisition_clk ;
 wire \clknet_leaf_47_top1.acquisition_clk ;
 wire \clknet_leaf_48_top1.acquisition_clk ;
 wire \clknet_leaf_49_top1.acquisition_clk ;
 wire \clknet_leaf_50_top1.acquisition_clk ;
 wire \clknet_leaf_51_top1.acquisition_clk ;
 wire \clknet_leaf_52_top1.acquisition_clk ;
 wire \clknet_leaf_53_top1.acquisition_clk ;
 wire \clknet_leaf_54_top1.acquisition_clk ;
 wire \clknet_leaf_55_top1.acquisition_clk ;
 wire \clknet_leaf_56_top1.acquisition_clk ;
 wire \clknet_leaf_57_top1.acquisition_clk ;
 wire \clknet_leaf_58_top1.acquisition_clk ;
 wire \clknet_leaf_59_top1.acquisition_clk ;
 wire \clknet_leaf_60_top1.acquisition_clk ;
 wire \clknet_leaf_61_top1.acquisition_clk ;
 wire \clknet_leaf_62_top1.acquisition_clk ;
 wire \clknet_leaf_63_top1.acquisition_clk ;
 wire \clknet_leaf_64_top1.acquisition_clk ;
 wire \clknet_leaf_65_top1.acquisition_clk ;
 wire \clknet_leaf_66_top1.acquisition_clk ;
 wire \clknet_leaf_67_top1.acquisition_clk ;
 wire \clknet_leaf_68_top1.acquisition_clk ;
 wire \clknet_leaf_69_top1.acquisition_clk ;
 wire \clknet_leaf_70_top1.acquisition_clk ;
 wire \clknet_leaf_71_top1.acquisition_clk ;
 wire \clknet_leaf_72_top1.acquisition_clk ;
 wire \clknet_leaf_73_top1.acquisition_clk ;
 wire \clknet_leaf_74_top1.acquisition_clk ;
 wire \clknet_leaf_75_top1.acquisition_clk ;
 wire \clknet_leaf_76_top1.acquisition_clk ;
 wire \clknet_leaf_77_top1.acquisition_clk ;
 wire \clknet_leaf_78_top1.acquisition_clk ;
 wire \clknet_leaf_79_top1.acquisition_clk ;
 wire \clknet_leaf_80_top1.acquisition_clk ;
 wire \clknet_leaf_81_top1.acquisition_clk ;
 wire \clknet_leaf_82_top1.acquisition_clk ;
 wire \clknet_leaf_83_top1.acquisition_clk ;
 wire \clknet_leaf_84_top1.acquisition_clk ;
 wire \clknet_leaf_85_top1.acquisition_clk ;
 wire \clknet_leaf_86_top1.acquisition_clk ;
 wire \clknet_leaf_87_top1.acquisition_clk ;
 wire \clknet_leaf_88_top1.acquisition_clk ;
 wire \clknet_leaf_89_top1.acquisition_clk ;
 wire \clknet_leaf_90_top1.acquisition_clk ;
 wire \clknet_leaf_91_top1.acquisition_clk ;
 wire \clknet_leaf_92_top1.acquisition_clk ;
 wire \clknet_leaf_93_top1.acquisition_clk ;
 wire \clknet_leaf_94_top1.acquisition_clk ;
 wire \clknet_leaf_95_top1.acquisition_clk ;
 wire \clknet_leaf_96_top1.acquisition_clk ;
 wire \clknet_leaf_97_top1.acquisition_clk ;
 wire \clknet_leaf_98_top1.acquisition_clk ;
 wire \clknet_leaf_99_top1.acquisition_clk ;
 wire \clknet_leaf_100_top1.acquisition_clk ;
 wire \clknet_leaf_101_top1.acquisition_clk ;
 wire \clknet_leaf_102_top1.acquisition_clk ;
 wire \clknet_leaf_103_top1.acquisition_clk ;
 wire \clknet_leaf_104_top1.acquisition_clk ;
 wire \clknet_leaf_105_top1.acquisition_clk ;
 wire \clknet_leaf_106_top1.acquisition_clk ;
 wire \clknet_leaf_107_top1.acquisition_clk ;
 wire \clknet_leaf_108_top1.acquisition_clk ;
 wire \clknet_leaf_109_top1.acquisition_clk ;
 wire \clknet_leaf_110_top1.acquisition_clk ;
 wire \clknet_leaf_111_top1.acquisition_clk ;
 wire \clknet_leaf_112_top1.acquisition_clk ;
 wire \clknet_leaf_113_top1.acquisition_clk ;
 wire \clknet_leaf_114_top1.acquisition_clk ;
 wire \clknet_leaf_115_top1.acquisition_clk ;
 wire \clknet_leaf_116_top1.acquisition_clk ;
 wire \clknet_leaf_117_top1.acquisition_clk ;
 wire \clknet_leaf_118_top1.acquisition_clk ;
 wire \clknet_leaf_119_top1.acquisition_clk ;
 wire \clknet_leaf_120_top1.acquisition_clk ;
 wire \clknet_leaf_121_top1.acquisition_clk ;
 wire \clknet_leaf_122_top1.acquisition_clk ;
 wire \clknet_leaf_123_top1.acquisition_clk ;
 wire \clknet_leaf_124_top1.acquisition_clk ;
 wire \clknet_leaf_125_top1.acquisition_clk ;
 wire \clknet_leaf_126_top1.acquisition_clk ;
 wire \clknet_leaf_127_top1.acquisition_clk ;
 wire \clknet_leaf_128_top1.acquisition_clk ;
 wire \clknet_leaf_129_top1.acquisition_clk ;
 wire \clknet_leaf_130_top1.acquisition_clk ;
 wire \clknet_leaf_131_top1.acquisition_clk ;
 wire \clknet_leaf_132_top1.acquisition_clk ;
 wire \clknet_leaf_133_top1.acquisition_clk ;
 wire \clknet_leaf_134_top1.acquisition_clk ;
 wire \clknet_leaf_135_top1.acquisition_clk ;
 wire \clknet_leaf_136_top1.acquisition_clk ;
 wire \clknet_leaf_137_top1.acquisition_clk ;
 wire \clknet_leaf_138_top1.acquisition_clk ;
 wire \clknet_leaf_139_top1.acquisition_clk ;
 wire \clknet_leaf_140_top1.acquisition_clk ;
 wire \clknet_leaf_141_top1.acquisition_clk ;
 wire \clknet_leaf_142_top1.acquisition_clk ;
 wire \clknet_leaf_143_top1.acquisition_clk ;
 wire \clknet_leaf_144_top1.acquisition_clk ;
 wire \clknet_leaf_145_top1.acquisition_clk ;
 wire \clknet_leaf_146_top1.acquisition_clk ;
 wire \clknet_leaf_147_top1.acquisition_clk ;
 wire \clknet_leaf_148_top1.acquisition_clk ;
 wire \clknet_leaf_149_top1.acquisition_clk ;
 wire \clknet_leaf_150_top1.acquisition_clk ;
 wire \clknet_leaf_151_top1.acquisition_clk ;
 wire \clknet_leaf_152_top1.acquisition_clk ;
 wire \clknet_leaf_153_top1.acquisition_clk ;
 wire \clknet_leaf_154_top1.acquisition_clk ;
 wire \clknet_leaf_155_top1.acquisition_clk ;
 wire \clknet_leaf_156_top1.acquisition_clk ;
 wire \clknet_leaf_157_top1.acquisition_clk ;
 wire \clknet_leaf_158_top1.acquisition_clk ;
 wire \clknet_leaf_159_top1.acquisition_clk ;
 wire \clknet_leaf_160_top1.acquisition_clk ;
 wire \clknet_leaf_161_top1.acquisition_clk ;
 wire \clknet_leaf_162_top1.acquisition_clk ;
 wire \clknet_leaf_163_top1.acquisition_clk ;
 wire \clknet_leaf_164_top1.acquisition_clk ;
 wire \clknet_leaf_165_top1.acquisition_clk ;
 wire \clknet_leaf_166_top1.acquisition_clk ;
 wire \clknet_leaf_167_top1.acquisition_clk ;
 wire \clknet_leaf_168_top1.acquisition_clk ;
 wire \clknet_leaf_169_top1.acquisition_clk ;
 wire \clknet_leaf_170_top1.acquisition_clk ;
 wire \clknet_leaf_171_top1.acquisition_clk ;
 wire \clknet_leaf_172_top1.acquisition_clk ;
 wire \clknet_leaf_173_top1.acquisition_clk ;
 wire \clknet_leaf_174_top1.acquisition_clk ;
 wire \clknet_leaf_175_top1.acquisition_clk ;
 wire \clknet_leaf_176_top1.acquisition_clk ;
 wire \clknet_leaf_177_top1.acquisition_clk ;
 wire \clknet_leaf_178_top1.acquisition_clk ;
 wire \clknet_leaf_179_top1.acquisition_clk ;
 wire \clknet_leaf_180_top1.acquisition_clk ;
 wire \clknet_leaf_181_top1.acquisition_clk ;
 wire \clknet_leaf_182_top1.acquisition_clk ;
 wire \clknet_leaf_183_top1.acquisition_clk ;
 wire \clknet_leaf_184_top1.acquisition_clk ;
 wire \clknet_leaf_185_top1.acquisition_clk ;
 wire \clknet_leaf_186_top1.acquisition_clk ;
 wire \clknet_leaf_187_top1.acquisition_clk ;
 wire \clknet_leaf_188_top1.acquisition_clk ;
 wire \clknet_leaf_189_top1.acquisition_clk ;
 wire \clknet_leaf_190_top1.acquisition_clk ;
 wire \clknet_leaf_191_top1.acquisition_clk ;
 wire \clknet_leaf_192_top1.acquisition_clk ;
 wire \clknet_leaf_193_top1.acquisition_clk ;
 wire \clknet_leaf_194_top1.acquisition_clk ;
 wire \clknet_leaf_195_top1.acquisition_clk ;
 wire \clknet_leaf_196_top1.acquisition_clk ;
 wire \clknet_leaf_197_top1.acquisition_clk ;
 wire \clknet_leaf_198_top1.acquisition_clk ;
 wire \clknet_leaf_199_top1.acquisition_clk ;
 wire \clknet_leaf_200_top1.acquisition_clk ;
 wire \clknet_leaf_201_top1.acquisition_clk ;
 wire \clknet_leaf_202_top1.acquisition_clk ;
 wire \clknet_leaf_203_top1.acquisition_clk ;
 wire \clknet_leaf_204_top1.acquisition_clk ;
 wire \clknet_leaf_205_top1.acquisition_clk ;
 wire \clknet_leaf_206_top1.acquisition_clk ;
 wire \clknet_leaf_207_top1.acquisition_clk ;
 wire \clknet_leaf_208_top1.acquisition_clk ;
 wire \clknet_leaf_209_top1.acquisition_clk ;
 wire \clknet_leaf_210_top1.acquisition_clk ;
 wire \clknet_leaf_211_top1.acquisition_clk ;
 wire \clknet_leaf_212_top1.acquisition_clk ;
 wire \clknet_leaf_213_top1.acquisition_clk ;
 wire \clknet_leaf_214_top1.acquisition_clk ;
 wire \clknet_leaf_215_top1.acquisition_clk ;
 wire \clknet_leaf_216_top1.acquisition_clk ;
 wire \clknet_leaf_217_top1.acquisition_clk ;
 wire \clknet_leaf_218_top1.acquisition_clk ;
 wire \clknet_leaf_219_top1.acquisition_clk ;
 wire \clknet_leaf_220_top1.acquisition_clk ;
 wire \clknet_leaf_221_top1.acquisition_clk ;
 wire \clknet_leaf_222_top1.acquisition_clk ;
 wire \clknet_leaf_223_top1.acquisition_clk ;
 wire \clknet_leaf_224_top1.acquisition_clk ;
 wire \clknet_leaf_225_top1.acquisition_clk ;
 wire \clknet_leaf_226_top1.acquisition_clk ;
 wire \clknet_leaf_227_top1.acquisition_clk ;
 wire \clknet_leaf_228_top1.acquisition_clk ;
 wire \clknet_leaf_229_top1.acquisition_clk ;
 wire \clknet_leaf_230_top1.acquisition_clk ;
 wire \clknet_leaf_231_top1.acquisition_clk ;
 wire \clknet_leaf_232_top1.acquisition_clk ;
 wire \clknet_leaf_233_top1.acquisition_clk ;
 wire \clknet_leaf_234_top1.acquisition_clk ;
 wire \clknet_leaf_235_top1.acquisition_clk ;
 wire \clknet_leaf_236_top1.acquisition_clk ;
 wire \clknet_leaf_237_top1.acquisition_clk ;
 wire \clknet_leaf_238_top1.acquisition_clk ;
 wire \clknet_leaf_239_top1.acquisition_clk ;
 wire \clknet_leaf_240_top1.acquisition_clk ;
 wire \clknet_leaf_241_top1.acquisition_clk ;
 wire \clknet_leaf_242_top1.acquisition_clk ;
 wire \clknet_leaf_243_top1.acquisition_clk ;
 wire \clknet_leaf_244_top1.acquisition_clk ;
 wire \clknet_leaf_245_top1.acquisition_clk ;
 wire \clknet_leaf_246_top1.acquisition_clk ;
 wire \clknet_leaf_247_top1.acquisition_clk ;
 wire \clknet_leaf_248_top1.acquisition_clk ;
 wire \clknet_leaf_249_top1.acquisition_clk ;
 wire \clknet_leaf_250_top1.acquisition_clk ;
 wire \clknet_leaf_251_top1.acquisition_clk ;
 wire \clknet_leaf_252_top1.acquisition_clk ;
 wire \clknet_leaf_253_top1.acquisition_clk ;
 wire \clknet_leaf_254_top1.acquisition_clk ;
 wire \clknet_leaf_255_top1.acquisition_clk ;
 wire \clknet_leaf_256_top1.acquisition_clk ;
 wire \clknet_leaf_257_top1.acquisition_clk ;
 wire \clknet_leaf_258_top1.acquisition_clk ;
 wire \clknet_leaf_259_top1.acquisition_clk ;
 wire \clknet_leaf_260_top1.acquisition_clk ;
 wire \clknet_leaf_261_top1.acquisition_clk ;
 wire \clknet_leaf_262_top1.acquisition_clk ;
 wire \clknet_leaf_263_top1.acquisition_clk ;
 wire \clknet_leaf_264_top1.acquisition_clk ;
 wire \clknet_leaf_265_top1.acquisition_clk ;
 wire \clknet_leaf_266_top1.acquisition_clk ;
 wire \clknet_leaf_267_top1.acquisition_clk ;
 wire \clknet_leaf_268_top1.acquisition_clk ;
 wire \clknet_leaf_269_top1.acquisition_clk ;
 wire \clknet_leaf_270_top1.acquisition_clk ;
 wire \clknet_leaf_271_top1.acquisition_clk ;
 wire \clknet_leaf_272_top1.acquisition_clk ;
 wire \clknet_leaf_273_top1.acquisition_clk ;
 wire \clknet_leaf_274_top1.acquisition_clk ;
 wire \clknet_leaf_275_top1.acquisition_clk ;
 wire \clknet_leaf_276_top1.acquisition_clk ;
 wire \clknet_leaf_277_top1.acquisition_clk ;
 wire \clknet_leaf_278_top1.acquisition_clk ;
 wire \clknet_leaf_279_top1.acquisition_clk ;
 wire \clknet_leaf_280_top1.acquisition_clk ;
 wire \clknet_leaf_281_top1.acquisition_clk ;
 wire \clknet_leaf_282_top1.acquisition_clk ;
 wire \clknet_leaf_283_top1.acquisition_clk ;
 wire \clknet_leaf_284_top1.acquisition_clk ;
 wire \clknet_leaf_285_top1.acquisition_clk ;
 wire \clknet_leaf_286_top1.acquisition_clk ;
 wire \clknet_leaf_287_top1.acquisition_clk ;
 wire \clknet_leaf_288_top1.acquisition_clk ;
 wire \clknet_leaf_289_top1.acquisition_clk ;
 wire \clknet_leaf_290_top1.acquisition_clk ;
 wire \clknet_leaf_291_top1.acquisition_clk ;
 wire \clknet_leaf_292_top1.acquisition_clk ;
 wire \clknet_leaf_293_top1.acquisition_clk ;
 wire \clknet_leaf_294_top1.acquisition_clk ;
 wire \clknet_leaf_295_top1.acquisition_clk ;
 wire \clknet_leaf_296_top1.acquisition_clk ;
 wire \clknet_leaf_297_top1.acquisition_clk ;
 wire \clknet_leaf_298_top1.acquisition_clk ;
 wire \clknet_leaf_299_top1.acquisition_clk ;
 wire \clknet_leaf_300_top1.acquisition_clk ;
 wire \clknet_leaf_301_top1.acquisition_clk ;
 wire \clknet_leaf_302_top1.acquisition_clk ;
 wire \clknet_0_top1.acquisition_clk ;
 wire \clknet_3_0_0_top1.acquisition_clk ;
 wire \clknet_3_1_0_top1.acquisition_clk ;
 wire \clknet_3_2_0_top1.acquisition_clk ;
 wire \clknet_3_3_0_top1.acquisition_clk ;
 wire \clknet_3_4_0_top1.acquisition_clk ;
 wire \clknet_3_5_0_top1.acquisition_clk ;
 wire \clknet_3_6_0_top1.acquisition_clk ;
 wire \clknet_3_7_0_top1.acquisition_clk ;
 wire \clknet_6_0_0_top1.acquisition_clk ;
 wire \clknet_6_1_0_top1.acquisition_clk ;
 wire \clknet_6_2_0_top1.acquisition_clk ;
 wire \clknet_6_3_0_top1.acquisition_clk ;
 wire \clknet_6_4_0_top1.acquisition_clk ;
 wire \clknet_6_5_0_top1.acquisition_clk ;
 wire \clknet_6_6_0_top1.acquisition_clk ;
 wire \clknet_6_7_0_top1.acquisition_clk ;
 wire \clknet_6_8_0_top1.acquisition_clk ;
 wire \clknet_6_9_0_top1.acquisition_clk ;
 wire \clknet_6_10_0_top1.acquisition_clk ;
 wire \clknet_6_11_0_top1.acquisition_clk ;
 wire \clknet_6_12_0_top1.acquisition_clk ;
 wire \clknet_6_13_0_top1.acquisition_clk ;
 wire \clknet_6_14_0_top1.acquisition_clk ;
 wire \clknet_6_15_0_top1.acquisition_clk ;
 wire \clknet_6_16_0_top1.acquisition_clk ;
 wire \clknet_6_17_0_top1.acquisition_clk ;
 wire \clknet_6_18_0_top1.acquisition_clk ;
 wire \clknet_6_19_0_top1.acquisition_clk ;
 wire \clknet_6_20_0_top1.acquisition_clk ;
 wire \clknet_6_21_0_top1.acquisition_clk ;
 wire \clknet_6_22_0_top1.acquisition_clk ;
 wire \clknet_6_23_0_top1.acquisition_clk ;
 wire \clknet_6_24_0_top1.acquisition_clk ;
 wire \clknet_6_25_0_top1.acquisition_clk ;
 wire \clknet_6_26_0_top1.acquisition_clk ;
 wire \clknet_6_27_0_top1.acquisition_clk ;
 wire \clknet_6_28_0_top1.acquisition_clk ;
 wire \clknet_6_29_0_top1.acquisition_clk ;
 wire \clknet_6_30_0_top1.acquisition_clk ;
 wire \clknet_6_31_0_top1.acquisition_clk ;
 wire \clknet_6_32_0_top1.acquisition_clk ;
 wire \clknet_6_33_0_top1.acquisition_clk ;
 wire \clknet_6_34_0_top1.acquisition_clk ;
 wire \clknet_6_35_0_top1.acquisition_clk ;
 wire \clknet_6_36_0_top1.acquisition_clk ;
 wire \clknet_6_37_0_top1.acquisition_clk ;
 wire \clknet_6_38_0_top1.acquisition_clk ;
 wire \clknet_6_39_0_top1.acquisition_clk ;
 wire \clknet_6_40_0_top1.acquisition_clk ;
 wire \clknet_6_41_0_top1.acquisition_clk ;
 wire \clknet_6_42_0_top1.acquisition_clk ;
 wire \clknet_6_43_0_top1.acquisition_clk ;
 wire \clknet_6_44_0_top1.acquisition_clk ;
 wire \clknet_6_45_0_top1.acquisition_clk ;
 wire \clknet_6_46_0_top1.acquisition_clk ;
 wire \clknet_6_47_0_top1.acquisition_clk ;
 wire \clknet_6_48_0_top1.acquisition_clk ;
 wire \clknet_6_49_0_top1.acquisition_clk ;
 wire \clknet_6_50_0_top1.acquisition_clk ;
 wire \clknet_6_51_0_top1.acquisition_clk ;
 wire \clknet_6_52_0_top1.acquisition_clk ;
 wire \clknet_6_53_0_top1.acquisition_clk ;
 wire \clknet_6_54_0_top1.acquisition_clk ;
 wire \clknet_6_55_0_top1.acquisition_clk ;
 wire \clknet_6_56_0_top1.acquisition_clk ;
 wire \clknet_6_57_0_top1.acquisition_clk ;
 wire \clknet_6_58_0_top1.acquisition_clk ;
 wire \clknet_6_59_0_top1.acquisition_clk ;
 wire \clknet_6_60_0_top1.acquisition_clk ;
 wire \clknet_6_61_0_top1.acquisition_clk ;
 wire \clknet_6_62_0_top1.acquisition_clk ;
 wire \clknet_6_63_0_top1.acquisition_clk ;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;

 sg13g2_inv_2 _12413_ (.Y(_03826_),
    .A(\top1.fsm.state_reg[1] ));
 sg13g2_inv_4 _12414_ (.A(net6131),
    .Y(_03827_));
 sg13g2_inv_1 _12415_ (.Y(_03828_),
    .A(net6125));
 sg13g2_inv_4 _12416_ (.A(net6117),
    .Y(_03829_));
 sg13g2_inv_4 _12417_ (.A(net6115),
    .Y(_03830_));
 sg13g2_inv_2 _12418_ (.Y(_03831_),
    .A(net6111));
 sg13g2_inv_1 _12419_ (.Y(_03832_),
    .A(\top1.fsm.re ));
 sg13g2_inv_1 _12420_ (.Y(_03833_),
    .A(\top1.fsm.signal_duration ));
 sg13g2_inv_1 _12421_ (.Y(_03834_),
    .A(\top1.event_time[25] ));
 sg13g2_inv_1 _12422_ (.Y(_03835_),
    .A(\top1.event_time[11] ));
 sg13g2_inv_1 _12423_ (.Y(_03836_),
    .A(\top1.event_time[10] ));
 sg13g2_inv_1 _12424_ (.Y(_03837_),
    .A(\top1.event_time[12] ));
 sg13g2_inv_1 _12425_ (.Y(_03838_),
    .A(\top1.event_time[13] ));
 sg13g2_inv_1 _12426_ (.Y(_03839_),
    .A(\top1.event_time[19] ));
 sg13g2_inv_1 _12427_ (.Y(_03840_),
    .A(\top1.event_time[18] ));
 sg13g2_inv_1 _12428_ (.Y(_00053_),
    .A(\top1.event_time[0] ));
 sg13g2_inv_1 _12429_ (.Y(_03841_),
    .A(\top1.event_time[3] ));
 sg13g2_inv_1 _12430_ (.Y(_03842_),
    .A(\top1.event_time[28] ));
 sg13g2_inv_1 _12431_ (.Y(_03843_),
    .A(\top1.event_time[27] ));
 sg13g2_inv_1 _12432_ (.Y(_03844_),
    .A(\top1.event_time[31] ));
 sg13g2_inv_2 _12433_ (.Y(_03845_),
    .A(net4864));
 sg13g2_inv_2 _12434_ (.Y(_03846_),
    .A(\top1.addr_in[4] ));
 sg13g2_inv_2 _12435_ (.Y(_03847_),
    .A(net7562));
 sg13g2_inv_4 _12436_ (.A(net7561),
    .Y(_03848_));
 sg13g2_inv_1 _12437_ (.Y(_03849_),
    .A(\top1.memory2.data_out[0] ));
 sg13g2_inv_1 _12438_ (.Y(_03850_),
    .A(\top1.memory2.data_out[1] ));
 sg13g2_inv_1 _12439_ (.Y(_03851_),
    .A(\top1.memory1.data_out[0] ));
 sg13g2_inv_1 _12440_ (.Y(_03852_),
    .A(\top1.memory1.data_out[1] ));
 sg13g2_inv_1 _12441_ (.Y(_03853_),
    .A(\top1.memory1.data_out[2] ));
 sg13g2_inv_1 _12442_ (.Y(_03854_),
    .A(\top1.memory2.mem2[69][0] ));
 sg13g2_inv_1 _12443_ (.Y(_03855_),
    .A(\top1.memory2.mem2[70][0] ));
 sg13g2_inv_1 _12444_ (.Y(_03856_),
    .A(\top1.memory2.mem2[71][0] ));
 sg13g2_inv_1 _12445_ (.Y(_03857_),
    .A(\top1.memory2.mem2[148][0] ));
 sg13g2_inv_1 _12446_ (.Y(_03858_),
    .A(\top1.memory2.mem2[149][0] ));
 sg13g2_inv_1 _12447_ (.Y(_03859_),
    .A(\top1.memory2.mem2[150][0] ));
 sg13g2_inv_1 _12448_ (.Y(_03860_),
    .A(\top1.memory2.mem2[151][0] ));
 sg13g2_inv_1 _12449_ (.Y(_03861_),
    .A(\top1.memory2.mem1[20][1] ));
 sg13g2_inv_1 _12450_ (.Y(_03862_),
    .A(\top1.memory2.mem1[21][1] ));
 sg13g2_inv_1 _12451_ (.Y(_03863_),
    .A(\top1.memory2.mem1[22][1] ));
 sg13g2_inv_1 _12452_ (.Y(_03864_),
    .A(\top1.memory2.mem1[23][1] ));
 sg13g2_inv_1 _12453_ (.Y(_03865_),
    .A(\top1.memory2.mem2[5][1] ));
 sg13g2_inv_1 _12454_ (.Y(_03866_),
    .A(\top1.memory2.mem2[6][1] ));
 sg13g2_inv_1 _12455_ (.Y(_03867_),
    .A(\top1.memory2.mem2[7][1] ));
 sg13g2_inv_1 _12456_ (.Y(_03868_),
    .A(\top1.memory2.mem2[20][1] ));
 sg13g2_inv_1 _12457_ (.Y(_03869_),
    .A(\top1.memory2.mem2[21][1] ));
 sg13g2_inv_1 _12458_ (.Y(_03870_),
    .A(\top1.memory2.mem2[22][1] ));
 sg13g2_inv_1 _12459_ (.Y(_03871_),
    .A(\top1.memory2.mem2[23][1] ));
 sg13g2_inv_1 _12460_ (.Y(_03872_),
    .A(\top1.memory2.mem1[21][2] ));
 sg13g2_inv_1 _12461_ (.Y(_03873_),
    .A(\top1.memory2.mem1[22][2] ));
 sg13g2_inv_1 _12462_ (.Y(_03874_),
    .A(\top1.memory2.mem1[23][2] ));
 sg13g2_inv_1 _12463_ (.Y(_03875_),
    .A(\top1.memory2.mem2[133][2] ));
 sg13g2_inv_1 _12464_ (.Y(_03876_),
    .A(\top1.memory2.mem2[134][2] ));
 sg13g2_inv_1 _12465_ (.Y(_03877_),
    .A(\top1.memory2.mem2[135][2] ));
 sg13g2_inv_1 _12466_ (.Y(_03878_),
    .A(\top1.memory1.mem1[21][0] ));
 sg13g2_inv_1 _12467_ (.Y(_03879_),
    .A(\top1.memory1.mem1[22][0] ));
 sg13g2_inv_1 _12468_ (.Y(_03880_),
    .A(\top1.memory1.mem1[23][0] ));
 sg13g2_inv_1 _12469_ (.Y(_03881_),
    .A(\top1.memory1.mem2[68][0] ));
 sg13g2_inv_1 _12470_ (.Y(_03882_),
    .A(\top1.memory1.mem2[69][0] ));
 sg13g2_inv_1 _12471_ (.Y(_03883_),
    .A(\top1.memory1.mem2[70][0] ));
 sg13g2_inv_1 _12472_ (.Y(_03884_),
    .A(\top1.memory1.mem2[71][0] ));
 sg13g2_inv_1 _12473_ (.Y(_03885_),
    .A(\top1.memory1.mem1[4][1] ));
 sg13g2_inv_1 _12474_ (.Y(_03886_),
    .A(\top1.memory1.mem1[5][1] ));
 sg13g2_inv_1 _12475_ (.Y(_03887_),
    .A(\top1.memory1.mem1[6][1] ));
 sg13g2_inv_1 _12476_ (.Y(_03888_),
    .A(\top1.memory1.mem1[7][1] ));
 sg13g2_inv_1 _12477_ (.Y(_03889_),
    .A(\top1.memory1.mem1[20][1] ));
 sg13g2_inv_1 _12478_ (.Y(_03890_),
    .A(\top1.memory1.mem1[21][1] ));
 sg13g2_inv_1 _12479_ (.Y(_03891_),
    .A(\top1.memory1.mem1[22][1] ));
 sg13g2_inv_1 _12480_ (.Y(_03892_),
    .A(\top1.memory1.mem1[23][1] ));
 sg13g2_inv_1 _12481_ (.Y(_03893_),
    .A(\top1.memory1.mem1[68][1] ));
 sg13g2_inv_1 _12482_ (.Y(_03894_),
    .A(\top1.memory1.mem1[69][1] ));
 sg13g2_inv_1 _12483_ (.Y(_03895_),
    .A(\top1.memory1.mem1[70][1] ));
 sg13g2_inv_1 _12484_ (.Y(_03896_),
    .A(\top1.memory1.mem1[71][1] ));
 sg13g2_inv_1 _12485_ (.Y(_03897_),
    .A(\top1.memory1.mem2[5][1] ));
 sg13g2_inv_1 _12486_ (.Y(_03898_),
    .A(\top1.memory1.mem2[6][1] ));
 sg13g2_inv_1 _12487_ (.Y(_03899_),
    .A(\top1.memory1.mem2[7][1] ));
 sg13g2_inv_1 _12488_ (.Y(_03900_),
    .A(\top1.memory1.mem2[69][1] ));
 sg13g2_inv_1 _12489_ (.Y(_03901_),
    .A(\top1.memory1.mem2[70][1] ));
 sg13g2_inv_1 _12490_ (.Y(_03902_),
    .A(\top1.memory1.mem2[71][1] ));
 sg13g2_inv_1 _12491_ (.Y(_03903_),
    .A(\top1.memory1.mem1[8][2] ));
 sg13g2_inv_1 _12492_ (.Y(_03904_),
    .A(\top1.memory1.mem1[9][2] ));
 sg13g2_inv_1 _12493_ (.Y(_03905_),
    .A(\top1.memory1.mem1[24][2] ));
 sg13g2_inv_1 _12494_ (.Y(_03906_),
    .A(\top1.memory1.mem1[25][2] ));
 sg13g2_inv_1 _12495_ (.Y(_03907_),
    .A(\top1.memory1.mem1[26][2] ));
 sg13g2_inv_1 _12496_ (.Y(_03908_),
    .A(\top1.memory1.mem1[27][2] ));
 sg13g2_inv_1 _12497_ (.Y(_03909_),
    .A(\top1.memory1.mem1[88][2] ));
 sg13g2_inv_1 _12498_ (.Y(_03910_),
    .A(\top1.memory1.mem1[89][2] ));
 sg13g2_inv_1 _12499_ (.Y(_03911_),
    .A(\top1.memory1.mem1[90][2] ));
 sg13g2_inv_1 _12500_ (.Y(_03912_),
    .A(\top1.memory1.mem1[91][2] ));
 sg13g2_inv_1 _12501_ (.Y(_03913_),
    .A(\top1.memory1.mem2[9][2] ));
 sg13g2_inv_1 _12502_ (.Y(_03914_),
    .A(\top1.memory1.mem2[10][2] ));
 sg13g2_inv_1 _12503_ (.Y(_03915_),
    .A(\top1.memory1.mem2[11][2] ));
 sg13g2_inv_1 _12504_ (.Y(_03916_),
    .A(\top1.memory1.mem2[25][2] ));
 sg13g2_inv_1 _12505_ (.Y(_03917_),
    .A(\top1.memory1.mem2[26][2] ));
 sg13g2_inv_1 _12506_ (.Y(_03918_),
    .A(\top1.memory1.mem2[27][2] ));
 sg13g2_inv_1 _12507_ (.Y(_03919_),
    .A(\top1.memory1.mem2[72][2] ));
 sg13g2_inv_1 _12508_ (.Y(_03920_),
    .A(\top1.memory1.mem2[73][2] ));
 sg13g2_inv_1 _12509_ (.Y(_03921_),
    .A(\top1.memory1.mem2[74][2] ));
 sg13g2_inv_1 _12510_ (.Y(_03922_),
    .A(\top1.memory1.mem2[75][2] ));
 sg13g2_inv_1 _12511_ (.Y(_03923_),
    .A(\top1.memory1.mem2[194][2] ));
 sg13g2_inv_1 _12512_ (.Y(_03924_),
    .A(net10));
 sg13g2_inv_1 _12513_ (.Y(_03925_),
    .A(net13));
 sg13g2_inv_1 _12514_ (.Y(_03926_),
    .A(net14));
 sg13g2_inv_1 _12515_ (.Y(_03927_),
    .A(net2));
 sg13g2_inv_1 _12516_ (.Y(_03928_),
    .A(net5));
 sg13g2_inv_1 _12517_ (.Y(_03929_),
    .A(net6));
 sg13g2_xnor2_1 _12518_ (.Y(_03930_),
    .A(\top1.fsm.reg_idx_final[2] ),
    .B(net6129));
 sg13g2_xnor2_1 _12519_ (.Y(_03931_),
    .A(\top1.fsm.reg_idx_final[5] ),
    .B(net6117));
 sg13g2_xnor2_1 _12520_ (.Y(_03932_),
    .A(\top1.fsm.reg_idx_final[1] ),
    .B(net6153));
 sg13g2_xnor2_1 _12521_ (.Y(_03933_),
    .A(\top1.fsm.reg_idx_final[6] ),
    .B(net6114));
 sg13g2_xnor2_1 _12522_ (.Y(_03934_),
    .A(\top1.fsm.reg_idx_final[3] ),
    .B(\top1.addr_out[3] ));
 sg13g2_xnor2_1 _12523_ (.Y(_03935_),
    .A(\top1.fsm.reg_idx_final[7] ),
    .B(net6112));
 sg13g2_xnor2_1 _12524_ (.Y(_03936_),
    .A(\top1.fsm.reg_idx_final[4] ),
    .B(net6123));
 sg13g2_xor2_1 _12525_ (.B(net6205),
    .A(\top1.fsm.reg_idx_final[0] ),
    .X(_03937_));
 sg13g2_nand4_1 _12526_ (.B(_03934_),
    .C(_03935_),
    .A(_03932_),
    .Y(_03938_),
    .D(_03936_));
 sg13g2_nand3_1 _12527_ (.B(_03931_),
    .C(_03933_),
    .A(_03930_),
    .Y(_03939_));
 sg13g2_nor3_2 _12528_ (.A(_03937_),
    .B(_03938_),
    .C(_03939_),
    .Y(_03940_));
 sg13g2_nor2_1 _12529_ (.A(\top1.fsm.cpt[2] ),
    .B(\top1.fsm.cpt[3] ),
    .Y(_03941_));
 sg13g2_nand2_1 _12530_ (.Y(_03942_),
    .A(_00064_),
    .B(_03941_));
 sg13g2_nor2b_1 _12531_ (.A(\top1.fsm.cpt[1] ),
    .B_N(\top1.fsm.cpt[0] ),
    .Y(_03943_));
 sg13g2_nand3_1 _12532_ (.B(_03941_),
    .C(_03943_),
    .A(_00064_),
    .Y(_03944_));
 sg13g2_nand3_1 _12533_ (.B(net6110),
    .C(\top1.fsm.state_reg[2] ),
    .A(\top1.fsm.state_reg[1] ),
    .Y(_03945_));
 sg13g2_nor2_1 _12534_ (.A(_03940_),
    .B(_03945_),
    .Y(_03946_));
 sg13g2_nand2b_1 _12535_ (.Y(_03947_),
    .B(\top1.fsm.cpt[1] ),
    .A_N(\top1.fsm.cpt[0] ));
 sg13g2_nor2_1 _12536_ (.A(_03942_),
    .B(_03947_),
    .Y(_03948_));
 sg13g2_a21oi_2 _12537_ (.B1(_03945_),
    .Y(_03949_),
    .A2(_03948_),
    .A1(_03940_));
 sg13g2_o21ai_1 _12538_ (.B1(_03949_),
    .Y(_03950_),
    .A1(_03940_),
    .A2(_03944_));
 sg13g2_and2_1 _12539_ (.A(\top1.fsm.state_reg[1] ),
    .B(_00063_),
    .X(_03951_));
 sg13g2_nand2b_2 _12540_ (.Y(_03952_),
    .B(_00063_),
    .A_N(net6110));
 sg13g2_nor2_2 _12541_ (.A(_03826_),
    .B(_03952_),
    .Y(_03953_));
 sg13g2_nand2_1 _12542_ (.Y(_03954_),
    .A(\top1.fsm.cpt[2] ),
    .B(\top1.fsm.cpt[3] ));
 sg13g2_nor3_1 _12543_ (.A(_00064_),
    .B(_03947_),
    .C(_03954_),
    .Y(_03955_));
 sg13g2_and2_1 _12544_ (.A(_03953_),
    .B(_03955_),
    .X(_03956_));
 sg13g2_nand2_1 _12545_ (.Y(_03957_),
    .A(\top1.fsm.signal_duration ),
    .B(_03956_));
 sg13g2_nor2b_1 _12546_ (.A(\top1.fsm.state_reg[1] ),
    .B_N(net6110),
    .Y(_03958_));
 sg13g2_a21oi_1 _12547_ (.A1(_00063_),
    .A2(_03958_),
    .Y(_03959_),
    .B1(_03953_));
 sg13g2_nor2_2 _12548_ (.A(\top1.bank0_full ),
    .B(\top1.bank1_full ),
    .Y(_03960_));
 sg13g2_nand2b_1 _12549_ (.Y(_03961_),
    .B(_03960_),
    .A_N(\top1.fsm.sending_pending ));
 sg13g2_and2_2 _12550_ (.A(net6110),
    .B(_03951_),
    .X(_03962_));
 sg13g2_nor2_1 _12551_ (.A(\top1.fsm.state_reg[2] ),
    .B(_03962_),
    .Y(_03963_));
 sg13g2_nand3_1 _12552_ (.B(_03961_),
    .C(_03963_),
    .A(_03959_),
    .Y(_03964_));
 sg13g2_nor2b_1 _12553_ (.A(net6110),
    .B_N(\top1.fsm.state_reg[2] ),
    .Y(_03965_));
 sg13g2_inv_1 _12554_ (.Y(_03966_),
    .A(_03965_));
 sg13g2_nor2_1 _12555_ (.A(\top1.fsm.state_reg[1] ),
    .B(net6110),
    .Y(_03967_));
 sg13g2_nor2_1 _12556_ (.A(\top1.fsm.state_reg[1] ),
    .B(_03966_),
    .Y(_03968_));
 sg13g2_nand2_1 _12557_ (.Y(_03969_),
    .A(_03826_),
    .B(_03965_));
 sg13g2_nor2_1 _12558_ (.A(_03944_),
    .B(_03969_),
    .Y(_03970_));
 sg13g2_nor2_2 _12559_ (.A(_03826_),
    .B(_03966_),
    .Y(_03971_));
 sg13g2_nand2_2 _12560_ (.Y(_03972_),
    .A(\top1.fsm.state_reg[2] ),
    .B(_03958_));
 sg13g2_a21oi_1 _12561_ (.A1(\top1.fsm.sending_pending ),
    .A2(\top1.fsm.re ),
    .Y(_03973_),
    .B1(_03972_));
 sg13g2_nor3_1 _12562_ (.A(_03970_),
    .B(_03971_),
    .C(_03973_),
    .Y(_03974_));
 sg13g2_nand4_1 _12563_ (.B(_03957_),
    .C(_03964_),
    .A(_03950_),
    .Y(\top1.fsm.state_next[0] ),
    .D(_03974_));
 sg13g2_nor2_1 _12564_ (.A(_03949_),
    .B(_03971_),
    .Y(_03975_));
 sg13g2_nor2_2 _12565_ (.A(net6124),
    .B(net6118),
    .Y(_03976_));
 sg13g2_or2_2 _12566_ (.X(_03977_),
    .B(net6117),
    .A(net6121));
 sg13g2_nor2_2 _12567_ (.A(net6102),
    .B(_03831_),
    .Y(_03978_));
 sg13g2_nand2_2 _12568_ (.Y(_03979_),
    .A(net6114),
    .B(net6112));
 sg13g2_nor2_2 _12569_ (.A(_03977_),
    .B(_03979_),
    .Y(_03980_));
 sg13g2_nor2b_1 _12570_ (.A(net6128),
    .B_N(net6127),
    .Y(_03981_));
 sg13g2_nand2b_2 _12571_ (.Y(_03982_),
    .B(net6127),
    .A_N(net6128));
 sg13g2_nor2_1 _12572_ (.A(net6218),
    .B(net6150),
    .Y(_03983_));
 sg13g2_or2_2 _12573_ (.X(_03984_),
    .B(net6138),
    .A(net6202));
 sg13g2_nand3_1 _12574_ (.B(net6084),
    .C(net6050),
    .A(_03980_),
    .Y(_03985_));
 sg13g2_nand2b_1 _12575_ (.Y(_03986_),
    .B(_03985_),
    .A_N(_03944_));
 sg13g2_nor2_1 _12576_ (.A(_00066_),
    .B(_03960_),
    .Y(_03987_));
 sg13g2_a21oi_1 _12577_ (.A1(_00065_),
    .A2(_03987_),
    .Y(_03988_),
    .B1(_03972_));
 sg13g2_or2_1 _12578_ (.X(_03989_),
    .B(_03988_),
    .A(_03962_));
 sg13g2_a221oi_1 _12579_ (.B2(_03986_),
    .C1(_03989_),
    .B1(_03968_),
    .A1(_03833_),
    .Y(_03990_),
    .A2(_03956_));
 sg13g2_nand2_1 _12580_ (.Y(\top1.fsm.state_next[2] ),
    .A(_03975_),
    .B(_03990_));
 sg13g2_nor2b_1 _12581_ (.A(\top1.mem_ctl.state_reg[0] ),
    .B_N(\top1.mem_ctl.state_reg[1] ),
    .Y(\top1.fsm.memorization_completed ));
 sg13g2_nor2_2 _12582_ (.A(net9),
    .B(net1),
    .Y(_03991_));
 sg13g2_inv_4 _12583_ (.A(_03991_),
    .Y(\top1.mem_ctl.signal_detected ));
 sg13g2_nand2b_1 _12584_ (.Y(_03992_),
    .B(_03961_),
    .A_N(_03972_));
 sg13g2_o21ai_1 _12585_ (.B1(_03959_),
    .Y(_03993_),
    .A1(_00066_),
    .A2(_03992_));
 sg13g2_a21oi_1 _12586_ (.A1(_03970_),
    .A2(_03985_),
    .Y(_03994_),
    .B1(_03993_));
 sg13g2_nand2_1 _12587_ (.Y(\top1.fsm.state_next[1] ),
    .A(_03975_),
    .B(_03994_));
 sg13g2_or2_1 _12588_ (.X(\top1.fsm.serial_readout ),
    .B(_03951_),
    .A(\top1.fsm.state_reg[2] ));
 sg13g2_nor2_1 _12589_ (.A(net4870),
    .B(\top1.mem_ctl.signal_detected ),
    .Y(_03995_));
 sg13g2_nand2b_2 _12590_ (.Y(_03996_),
    .B(_03995_),
    .A_N(\top1.mem_ctl.state_reg[0] ));
 sg13g2_nor4_1 _12591_ (.A(\top1.fsm.state_reg[1] ),
    .B(\top1.fsm.state_reg[2] ),
    .C(_03952_),
    .D(_03996_),
    .Y(_03997_));
 sg13g2_nor2b_1 _12592_ (.A(_03997_),
    .B_N(net16),
    .Y(\top1.fsm.clk ));
 sg13g2_and2_1 _12593_ (.A(clk),
    .B(_03996_),
    .X(\top1.acquisition_clk ));
 sg13g2_nor2_1 _12594_ (.A(_03967_),
    .B(\top1.fsm.serial_readout ),
    .Y(\top1.SL_time ));
 sg13g2_mux2_1 _12595_ (.A0(\top1.piso_time_reg.register[0] ),
    .A1(\top1.event_time_out[0] ),
    .S(net5829),
    .X(_00046_));
 sg13g2_mux2_1 _12596_ (.A0(\top1.piso_time_reg.register[1] ),
    .A1(\top1.event_time_out[1] ),
    .S(net5829),
    .X(_00015_));
 sg13g2_mux2_1 _12597_ (.A0(\top1.piso_time_reg.register[2] ),
    .A1(\top1.event_time_out[2] ),
    .S(net5829),
    .X(_00026_));
 sg13g2_mux2_1 _12598_ (.A0(\top1.piso_time_reg.register[3] ),
    .A1(\top1.event_time_out[3] ),
    .S(net5829),
    .X(_00037_));
 sg13g2_mux2_1 _12599_ (.A0(\top1.piso_time_reg.register[4] ),
    .A1(\top1.event_time_out[4] ),
    .S(net5829),
    .X(_00039_));
 sg13g2_mux2_1 _12600_ (.A0(\top1.piso_time_reg.register[5] ),
    .A1(\top1.event_time_out[5] ),
    .S(net5827),
    .X(_00040_));
 sg13g2_mux2_1 _12601_ (.A0(\top1.piso_time_reg.register[6] ),
    .A1(\top1.event_time_out[6] ),
    .S(net5827),
    .X(_00041_));
 sg13g2_mux2_1 _12602_ (.A0(\top1.piso_time_reg.register[7] ),
    .A1(\top1.event_time_out[7] ),
    .S(net5827),
    .X(_00042_));
 sg13g2_mux2_1 _12603_ (.A0(\top1.piso_time_reg.register[8] ),
    .A1(\top1.event_time_out[8] ),
    .S(net5827),
    .X(_00043_));
 sg13g2_mux2_1 _12604_ (.A0(\top1.piso_time_reg.register[9] ),
    .A1(\top1.event_time_out[9] ),
    .S(net5828),
    .X(_00044_));
 sg13g2_mux2_1 _12605_ (.A0(\top1.piso_time_reg.register[10] ),
    .A1(\top1.event_time_out[10] ),
    .S(net5827),
    .X(_00045_));
 sg13g2_mux2_1 _12606_ (.A0(\top1.piso_time_reg.register[11] ),
    .A1(\top1.event_time_out[11] ),
    .S(net5827),
    .X(_00016_));
 sg13g2_mux2_1 _12607_ (.A0(\top1.piso_time_reg.register[12] ),
    .A1(\top1.event_time_out[12] ),
    .S(net5827),
    .X(_00017_));
 sg13g2_mux2_1 _12608_ (.A0(\top1.piso_time_reg.register[13] ),
    .A1(\top1.event_time_out[13] ),
    .S(net5827),
    .X(_00018_));
 sg13g2_mux2_1 _12609_ (.A0(\top1.piso_time_reg.register[14] ),
    .A1(\top1.event_time_out[14] ),
    .S(net5828),
    .X(_00019_));
 sg13g2_mux2_1 _12610_ (.A0(\top1.piso_time_reg.register[15] ),
    .A1(\top1.event_time_out[15] ),
    .S(net5828),
    .X(_00020_));
 sg13g2_mux2_1 _12611_ (.A0(\top1.piso_time_reg.register[16] ),
    .A1(\top1.event_time_out[16] ),
    .S(net5826),
    .X(_00021_));
 sg13g2_mux2_1 _12612_ (.A0(\top1.piso_time_reg.register[17] ),
    .A1(\top1.event_time_out[17] ),
    .S(net5830),
    .X(_00022_));
 sg13g2_mux2_1 _12613_ (.A0(\top1.piso_time_reg.register[18] ),
    .A1(\top1.event_time_out[18] ),
    .S(net5826),
    .X(_00023_));
 sg13g2_mux2_1 _12614_ (.A0(\top1.piso_time_reg.register[19] ),
    .A1(\top1.event_time_out[19] ),
    .S(net5826),
    .X(_00024_));
 sg13g2_mux2_1 _12615_ (.A0(\top1.piso_time_reg.register[20] ),
    .A1(\top1.event_time_out[20] ),
    .S(net5826),
    .X(_00025_));
 sg13g2_mux2_1 _12616_ (.A0(\top1.piso_time_reg.register[21] ),
    .A1(\top1.event_time_out[21] ),
    .S(net5826),
    .X(_00027_));
 sg13g2_mux2_1 _12617_ (.A0(\top1.piso_time_reg.register[22] ),
    .A1(\top1.event_time_out[22] ),
    .S(net5830),
    .X(_00028_));
 sg13g2_mux2_1 _12618_ (.A0(\top1.piso_time_reg.register[23] ),
    .A1(\top1.event_time_out[23] ),
    .S(net5825),
    .X(_00029_));
 sg13g2_mux2_1 _12619_ (.A0(\top1.piso_time_reg.register[24] ),
    .A1(\top1.event_time_out[24] ),
    .S(net5825),
    .X(_00030_));
 sg13g2_mux2_1 _12620_ (.A0(\top1.piso_time_reg.register[25] ),
    .A1(\top1.event_time_out[25] ),
    .S(net5825),
    .X(_00031_));
 sg13g2_mux2_1 _12621_ (.A0(\top1.piso_time_reg.register[26] ),
    .A1(\top1.event_time_out[26] ),
    .S(net5825),
    .X(_00032_));
 sg13g2_mux2_1 _12622_ (.A0(\top1.piso_time_reg.register[27] ),
    .A1(\top1.event_time_out[27] ),
    .S(net5825),
    .X(_00033_));
 sg13g2_mux2_1 _12623_ (.A0(\top1.piso_time_reg.register[28] ),
    .A1(\top1.event_time_out[28] ),
    .S(net5825),
    .X(_00034_));
 sg13g2_mux2_1 _12624_ (.A0(\top1.piso_time_reg.register[29] ),
    .A1(\top1.event_time_out[29] ),
    .S(net5826),
    .X(_00035_));
 sg13g2_mux2_1 _12625_ (.A0(\top1.piso_time_reg.register[30] ),
    .A1(\top1.event_time_out[30] ),
    .S(net5825),
    .X(_00036_));
 sg13g2_and2_1 _12626_ (.A(\top1.event_time_out[31] ),
    .B(net5825),
    .X(_00038_));
 sg13g2_xor2_1 _12627_ (.B(\top1.event_time[0] ),
    .A(\top1.event_time[1] ),
    .X(_00054_));
 sg13g2_nand3_1 _12628_ (.B(\top1.event_time[0] ),
    .C(\top1.event_time[2] ),
    .A(\top1.event_time[1] ),
    .Y(_03998_));
 sg13g2_a21o_1 _12629_ (.A2(\top1.event_time[0] ),
    .A1(\top1.event_time[1] ),
    .B1(\top1.event_time[2] ),
    .X(_03999_));
 sg13g2_and2_1 _12630_ (.A(_03998_),
    .B(_03999_),
    .X(_00055_));
 sg13g2_nand3_1 _12631_ (.B(\top1.event_time[8] ),
    .C(\top1.event_time[9] ),
    .A(\top1.event_time[6] ),
    .Y(_04000_));
 sg13g2_or2_1 _12632_ (.X(_04001_),
    .B(\top1.event_time[4] ),
    .A(\top1.event_time[3] ));
 sg13g2_nand2_1 _12633_ (.Y(_04002_),
    .A(\top1.event_time[5] ),
    .B(\top1.event_time[7] ));
 sg13g2_nor4_2 _12634_ (.A(_03998_),
    .B(_04000_),
    .C(_04001_),
    .Y(_04003_),
    .D(_04002_));
 sg13g2_or4_2 _12635_ (.A(_03998_),
    .B(_04000_),
    .C(_04001_),
    .D(_04002_),
    .X(_04004_));
 sg13g2_and2_1 _12636_ (.A(_03841_),
    .B(_03998_),
    .X(_04005_));
 sg13g2_nor2_1 _12637_ (.A(_03841_),
    .B(_03998_),
    .Y(_04006_));
 sg13g2_nor3_1 _12638_ (.A(_04003_),
    .B(_04005_),
    .C(_04006_),
    .Y(_00056_));
 sg13g2_and2_1 _12639_ (.A(\top1.event_time[4] ),
    .B(_04006_),
    .X(_04007_));
 sg13g2_xor2_1 _12640_ (.B(_04006_),
    .A(\top1.event_time[4] ),
    .X(_00057_));
 sg13g2_nor2_1 _12641_ (.A(\top1.event_time[5] ),
    .B(_04007_),
    .Y(_04008_));
 sg13g2_and2_1 _12642_ (.A(\top1.event_time[5] ),
    .B(_04007_),
    .X(_04009_));
 sg13g2_nor3_1 _12643_ (.A(_04003_),
    .B(_04008_),
    .C(_04009_),
    .Y(_00058_));
 sg13g2_nor2_1 _12644_ (.A(\top1.event_time[6] ),
    .B(_04009_),
    .Y(_04010_));
 sg13g2_and2_1 _12645_ (.A(\top1.event_time[6] ),
    .B(_04009_),
    .X(_04011_));
 sg13g2_nor3_1 _12646_ (.A(_04003_),
    .B(_04010_),
    .C(_04011_),
    .Y(_00059_));
 sg13g2_nor2_1 _12647_ (.A(\top1.event_time[7] ),
    .B(_04011_),
    .Y(_04012_));
 sg13g2_and2_1 _12648_ (.A(\top1.event_time[7] ),
    .B(_04011_),
    .X(_04013_));
 sg13g2_nor3_1 _12649_ (.A(_04003_),
    .B(_04012_),
    .C(_04013_),
    .Y(_00060_));
 sg13g2_a21o_1 _12650_ (.A2(_04013_),
    .A1(\top1.event_time[8] ),
    .B1(_04003_),
    .X(_04014_));
 sg13g2_nor2_1 _12651_ (.A(\top1.event_time[8] ),
    .B(_04013_),
    .Y(_04015_));
 sg13g2_nor2_1 _12652_ (.A(_04014_),
    .B(_04015_),
    .Y(_00061_));
 sg13g2_a21oi_1 _12653_ (.A1(\top1.event_time[8] ),
    .A2(_04013_),
    .Y(_04016_),
    .B1(\top1.event_time[9] ));
 sg13g2_a21oi_1 _12654_ (.A1(\top1.event_time[9] ),
    .A2(_04014_),
    .Y(_00062_),
    .B1(_04016_));
 sg13g2_mux2_1 _12655_ (.A0(\top1.PISO_ch1 ),
    .A1(\top1.PISO_time ),
    .S(_03963_),
    .X(\top1.mux.data_out ));
 sg13g2_nand2_1 _12656_ (.Y(_04017_),
    .A(_03945_),
    .B(_03969_));
 sg13g2_nor2_2 _12657_ (.A(_03953_),
    .B(_04017_),
    .Y(_04018_));
 sg13g2_nand2_1 _12658_ (.Y(_04019_),
    .A(_03972_),
    .B(_04018_));
 sg13g2_a21oi_1 _12659_ (.A1(_03826_),
    .A2(_00063_),
    .Y(\top1.SL_ch ),
    .B1(_04019_));
 sg13g2_nor2_1 _12660_ (.A(\top1.reg2.register[0] ),
    .B(net5823),
    .Y(_04020_));
 sg13g2_a21oi_2 _12661_ (.B1(_04020_),
    .Y(_00052_),
    .A2(net5823),
    .A1(_03849_));
 sg13g2_nor2_1 _12662_ (.A(\top1.reg2.register[1] ),
    .B(net5822),
    .Y(_04021_));
 sg13g2_a21oi_1 _12663_ (.A1(_03850_),
    .A2(net5822),
    .Y(_00050_),
    .B1(_04021_));
 sg13g2_and2_1 _12664_ (.A(\top1.memory2.data_out[2] ),
    .B(net5822),
    .X(_00051_));
 sg13g2_nor2_1 _12665_ (.A(\top1.reg1.register[0] ),
    .B(net5822),
    .Y(_04022_));
 sg13g2_a21oi_2 _12666_ (.B1(_04022_),
    .Y(_00049_),
    .A2(net5822),
    .A1(_03851_));
 sg13g2_nor2_1 _12667_ (.A(\top1.reg1.register[1] ),
    .B(net5822),
    .Y(_04023_));
 sg13g2_a21oi_1 _12668_ (.A1(_03852_),
    .A2(net5822),
    .Y(_00047_),
    .B1(_04023_));
 sg13g2_and2_1 _12669_ (.A(\top1.memory1.data_out[2] ),
    .B(net5822),
    .X(_00048_));
 sg13g2_nor2_1 _12670_ (.A(\top1.fsm.cpt[0] ),
    .B(_04018_),
    .Y(_00001_));
 sg13g2_and2_1 _12671_ (.A(\top1.fsm.cpt[1] ),
    .B(\top1.fsm.cpt[0] ),
    .X(_04024_));
 sg13g2_nor2_1 _12672_ (.A(\top1.fsm.cpt[1] ),
    .B(\top1.fsm.cpt[0] ),
    .Y(_04025_));
 sg13g2_nor3_1 _12673_ (.A(_04018_),
    .B(_04024_),
    .C(_04025_),
    .Y(_00002_));
 sg13g2_xnor2_1 _12674_ (.Y(_04026_),
    .A(\top1.fsm.cpt[2] ),
    .B(_04024_));
 sg13g2_nor2_1 _12675_ (.A(_04018_),
    .B(_04026_),
    .Y(_00003_));
 sg13g2_nor2b_1 _12676_ (.A(_03954_),
    .B_N(_04024_),
    .Y(_04027_));
 sg13g2_a21oi_1 _12677_ (.A1(\top1.fsm.cpt[2] ),
    .A2(_04024_),
    .Y(_04028_),
    .B1(\top1.fsm.cpt[3] ));
 sg13g2_nor3_1 _12678_ (.A(_04018_),
    .B(_04027_),
    .C(_04028_),
    .Y(_00004_));
 sg13g2_xnor2_1 _12679_ (.Y(_04029_),
    .A(\top1.fsm.cpt[4] ),
    .B(_04027_));
 sg13g2_nor2_1 _12680_ (.A(_04018_),
    .B(_04029_),
    .Y(_00005_));
 sg13g2_nor2b_1 _12681_ (.A(net7565),
    .B_N(net7566),
    .Y(_00007_));
 sg13g2_and2_2 _12682_ (.A(net4863),
    .B(net7564),
    .X(_04030_));
 sg13g2_nand2_2 _12683_ (.Y(_04031_),
    .A(net7565),
    .B(net7564));
 sg13g2_nor2_2 _12684_ (.A(\top1.addr_in[0] ),
    .B(\top1.addr_in[1] ),
    .Y(_04032_));
 sg13g2_or2_2 _12685_ (.X(_04033_),
    .B(net7564),
    .A(net7565));
 sg13g2_and3_1 _12686_ (.X(_00008_),
    .A(net7566),
    .B(_04031_),
    .C(_04033_));
 sg13g2_o21ai_1 _12687_ (.B1(net7566),
    .Y(_04034_),
    .A1(_03845_),
    .A2(_04031_));
 sg13g2_a21oi_1 _12688_ (.A1(_03845_),
    .A2(_04031_),
    .Y(_00009_),
    .B1(_04034_));
 sg13g2_nor2_2 _12689_ (.A(net7563),
    .B(\top1.addr_in[4] ),
    .Y(_04035_));
 sg13g2_nor4_1 _12690_ (.A(\top1.addr_in[5] ),
    .B(\top1.addr_in[4] ),
    .C(_03847_),
    .D(_03848_),
    .Y(_04036_));
 sg13g2_nor2_2 _12691_ (.A(_03845_),
    .B(\top1.addr_in[3] ),
    .Y(_04037_));
 sg13g2_nand2b_2 _12692_ (.Y(_04038_),
    .B(\top1.addr_in[2] ),
    .A_N(\top1.addr_in[3] ));
 sg13g2_nor2_1 _12693_ (.A(_04031_),
    .B(_04038_),
    .Y(_04039_));
 sg13g2_nand2_2 _12694_ (.Y(_04040_),
    .A(_04030_),
    .B(_04037_));
 sg13g2_nand2_2 _12695_ (.Y(_04041_),
    .A(net7412),
    .B(net7406));
 sg13g2_o21ai_1 _12696_ (.B1(net7566),
    .Y(_04042_),
    .A1(\top1.mem_ctl.state_reg[1] ),
    .A2(_04041_));
 sg13g2_nand2_2 _12697_ (.Y(_04043_),
    .A(\top1.addr_in[2] ),
    .B(\top1.addr_in[3] ));
 sg13g2_nor2_2 _12698_ (.A(_04031_),
    .B(_04043_),
    .Y(_04044_));
 sg13g2_or2_2 _12699_ (.X(_04045_),
    .B(_04043_),
    .A(_04031_));
 sg13g2_a21oi_1 _12700_ (.A1(net4864),
    .A2(_04030_),
    .Y(_04046_),
    .B1(\top1.addr_in[3] ));
 sg13g2_nor3_1 _12701_ (.A(_04042_),
    .B(net7403),
    .C(net4865),
    .Y(_00010_));
 sg13g2_o21ai_1 _12702_ (.B1(net7566),
    .Y(_04047_),
    .A1(_03846_),
    .A2(_04045_));
 sg13g2_a21oi_1 _12703_ (.A1(net4867),
    .A2(net7402),
    .Y(_00011_),
    .B1(_04047_));
 sg13g2_a21oi_1 _12704_ (.A1(net4866),
    .A2(net7403),
    .Y(_04048_),
    .B1(net7563));
 sg13g2_nand2_2 _12705_ (.Y(_04049_),
    .A(\top1.addr_in[5] ),
    .B(\top1.addr_in[4] ));
 sg13g2_or2_1 _12706_ (.X(_04050_),
    .B(_04049_),
    .A(net7402));
 sg13g2_nand2_1 _12707_ (.Y(_04051_),
    .A(net7566),
    .B(_04050_));
 sg13g2_nor2_1 _12708_ (.A(_04048_),
    .B(_04051_),
    .Y(_00012_));
 sg13g2_xnor2_1 _12709_ (.Y(_04052_),
    .A(_03847_),
    .B(_04050_));
 sg13g2_nor2_1 _12710_ (.A(_04042_),
    .B(_04052_),
    .Y(_00013_));
 sg13g2_o21ai_1 _12711_ (.B1(net7561),
    .Y(_04053_),
    .A1(_03847_),
    .A2(_04050_));
 sg13g2_nor2_2 _12712_ (.A(_03847_),
    .B(net7561),
    .Y(_04054_));
 sg13g2_nand2_2 _12713_ (.Y(_04055_),
    .A(\top1.addr_in[6] ),
    .B(_03848_));
 sg13g2_nand4_1 _12714_ (.B(\top1.addr_in[4] ),
    .C(net7403),
    .A(\top1.addr_in[5] ),
    .Y(_04056_),
    .D(_04054_));
 sg13g2_nor2_2 _12715_ (.A(_04049_),
    .B(_04055_),
    .Y(_04057_));
 sg13g2_a21oi_1 _12716_ (.A1(_04053_),
    .A2(_04056_),
    .Y(_00014_),
    .B1(_04042_));
 sg13g2_nor2b_2 _12717_ (.A(\top1.mem_ctl.state_reg[1] ),
    .B_N(net7566),
    .Y(_04058_));
 sg13g2_nand2b_1 _12718_ (.Y(_04059_),
    .B(net7566),
    .A_N(\top1.mem_ctl.state_reg[1] ));
 sg13g2_nor2_1 _12719_ (.A(_00000_),
    .B(_04059_),
    .Y(_04060_));
 sg13g2_nand2b_2 _12720_ (.Y(_04061_),
    .B(_04058_),
    .A_N(_00000_));
 sg13g2_nor2b_2 _12721_ (.A(net7564),
    .B_N(net7565),
    .Y(_04062_));
 sg13g2_nand2b_1 _12722_ (.Y(_04063_),
    .B(net7565),
    .A_N(net7564));
 sg13g2_nor2_1 _12723_ (.A(_04038_),
    .B(_04063_),
    .Y(_04064_));
 sg13g2_nand2_2 _12724_ (.Y(_04065_),
    .A(_04037_),
    .B(_04062_));
 sg13g2_nand3_1 _12725_ (.B(net7380),
    .C(net7361),
    .A(net7410),
    .Y(_04066_));
 sg13g2_a21oi_1 _12726_ (.A1(net1),
    .A2(_03927_),
    .Y(_04067_),
    .B1(net3));
 sg13g2_o21ai_1 _12727_ (.B1(_03928_),
    .Y(_04068_),
    .A1(net4),
    .A2(_04067_));
 sg13g2_a21oi_2 _12728_ (.B1(net7),
    .Y(_04069_),
    .A2(_04068_),
    .A1(_03929_));
 sg13g2_nand2_1 _12729_ (.Y(_04070_),
    .A(net2658),
    .B(net7113));
 sg13g2_o21ai_1 _12730_ (.B1(_04070_),
    .Y(_00074_),
    .A1(net7112),
    .A2(net7316));
 sg13g2_nor2_1 _12731_ (.A(net2),
    .B(net3),
    .Y(_04071_));
 sg13g2_nor3_1 _12732_ (.A(net4),
    .B(net5),
    .C(_04071_),
    .Y(_04072_));
 sg13g2_nor3_2 _12733_ (.A(net6),
    .B(net7),
    .C(_04072_),
    .Y(_04073_));
 sg13g2_nand2_1 _12734_ (.Y(_04074_),
    .A(net3905),
    .B(net7112));
 sg13g2_o21ai_1 _12735_ (.B1(_04074_),
    .Y(_00075_),
    .A1(net7113),
    .A2(net7516));
 sg13g2_nor4_2 _12736_ (.A(net4),
    .B(net5),
    .C(net6),
    .Y(_04075_),
    .D(net7));
 sg13g2_nand2_1 _12737_ (.Y(_04076_),
    .A(net3014),
    .B(net7113));
 sg13g2_o21ai_1 _12738_ (.B1(_04076_),
    .Y(_00076_),
    .A1(net7113),
    .A2(net7670));
 sg13g2_nor2_2 _12739_ (.A(\top1.addr_in[2] ),
    .B(\top1.addr_in[3] ),
    .Y(_04077_));
 sg13g2_and2_2 _12740_ (.A(_04030_),
    .B(_04077_),
    .X(_04078_));
 sg13g2_nand2_2 _12741_ (.Y(_04079_),
    .A(_04030_),
    .B(_04077_));
 sg13g2_nand3_1 _12742_ (.B(net7379),
    .C(net7285),
    .A(net7410),
    .Y(_04080_));
 sg13g2_nand2_1 _12743_ (.Y(_04081_),
    .A(net3590),
    .B(net7111));
 sg13g2_o21ai_1 _12744_ (.B1(_04081_),
    .Y(_00077_),
    .A1(net7316),
    .A2(net7111));
 sg13g2_nand2_1 _12745_ (.Y(_04082_),
    .A(net3326),
    .B(net7111));
 sg13g2_o21ai_1 _12746_ (.B1(_04082_),
    .Y(_00078_),
    .A1(net7516),
    .A2(net7111));
 sg13g2_nand2_1 _12747_ (.Y(_04083_),
    .A(net2451),
    .B(net7110));
 sg13g2_o21ai_1 _12748_ (.B1(_04083_),
    .Y(_00079_),
    .A1(net7670),
    .A2(net7110));
 sg13g2_nor2b_2 _12749_ (.A(net7565),
    .B_N(net7564),
    .Y(_04084_));
 sg13g2_nand2b_1 _12750_ (.Y(_04085_),
    .B(net7564),
    .A_N(net7565));
 sg13g2_nor2_1 _12751_ (.A(_04038_),
    .B(_04085_),
    .Y(_04086_));
 sg13g2_nand2_2 _12752_ (.Y(_04087_),
    .A(_04037_),
    .B(_04084_));
 sg13g2_nand3_1 _12753_ (.B(net7380),
    .C(net7281),
    .A(net7411),
    .Y(_04088_));
 sg13g2_nand2_1 _12754_ (.Y(_04089_),
    .A(net2803),
    .B(net7109));
 sg13g2_o21ai_1 _12755_ (.B1(_04089_),
    .Y(_00080_),
    .A1(net7316),
    .A2(net7109));
 sg13g2_nand2_1 _12756_ (.Y(_04090_),
    .A(net3483),
    .B(net7109));
 sg13g2_o21ai_1 _12757_ (.B1(_04090_),
    .Y(_00081_),
    .A1(net7516),
    .A2(net7108));
 sg13g2_nand2_1 _12758_ (.Y(_04091_),
    .A(net2755),
    .B(net7109));
 sg13g2_o21ai_1 _12759_ (.B1(_04091_),
    .Y(_00082_),
    .A1(net7670),
    .A2(net7108));
 sg13g2_nor2_2 _12760_ (.A(_04033_),
    .B(_04038_),
    .Y(_04092_));
 sg13g2_nand2_2 _12761_ (.Y(_04093_),
    .A(_04032_),
    .B(_04037_));
 sg13g2_nand3_1 _12762_ (.B(net7379),
    .C(net7280),
    .A(net7411),
    .Y(_04094_));
 sg13g2_nand2_1 _12763_ (.Y(_04095_),
    .A(net3700),
    .B(net7105));
 sg13g2_o21ai_1 _12764_ (.B1(_04095_),
    .Y(_00083_),
    .A1(net7316),
    .A2(net7105));
 sg13g2_nand2_1 _12765_ (.Y(_04096_),
    .A(net3147),
    .B(net7106));
 sg13g2_o21ai_1 _12766_ (.B1(_04096_),
    .Y(_00084_),
    .A1(net7516),
    .A2(net7106));
 sg13g2_nand2_1 _12767_ (.Y(_04097_),
    .A(net3691),
    .B(net7106));
 sg13g2_o21ai_1 _12768_ (.B1(_04097_),
    .Y(_00085_),
    .A1(net7670),
    .A2(net7105));
 sg13g2_nor2b_2 _12769_ (.A(\top1.addr_in[2] ),
    .B_N(\top1.addr_in[3] ),
    .Y(_04098_));
 sg13g2_nand2_2 _12770_ (.Y(_04099_),
    .A(_03845_),
    .B(\top1.addr_in[3] ));
 sg13g2_nor2_1 _12771_ (.A(_04085_),
    .B(_04099_),
    .Y(_04100_));
 sg13g2_nand2_2 _12772_ (.Y(_04101_),
    .A(_04084_),
    .B(_04098_));
 sg13g2_nand3_1 _12773_ (.B(net7391),
    .C(net7103),
    .A(net7115),
    .Y(_04102_));
 sg13g2_nand2_1 _12774_ (.Y(_04103_),
    .A(net2793),
    .B(net6734));
 sg13g2_o21ai_1 _12775_ (.B1(_04103_),
    .Y(_00086_),
    .A1(net7344),
    .A2(net6734));
 sg13g2_nand2_1 _12776_ (.Y(_04104_),
    .A(net2707),
    .B(net6734));
 sg13g2_o21ai_1 _12777_ (.B1(_04104_),
    .Y(_00087_),
    .A1(net7542),
    .A2(net6734));
 sg13g2_nand2_1 _12778_ (.Y(_04105_),
    .A(net2852),
    .B(net6735));
 sg13g2_o21ai_1 _12779_ (.B1(_04105_),
    .Y(_00088_),
    .A1(net7708),
    .A2(net6735));
 sg13g2_and2_2 _12780_ (.A(_04062_),
    .B(_04077_),
    .X(_04106_));
 sg13g2_nand2_2 _12781_ (.Y(_04107_),
    .A(_04062_),
    .B(_04077_));
 sg13g2_nand2_2 _12782_ (.Y(_04108_),
    .A(net7563),
    .B(_03846_));
 sg13g2_nor2_2 _12783_ (.A(_04055_),
    .B(_04108_),
    .Y(_04109_));
 sg13g2_nand3_1 _12784_ (.B(_03846_),
    .C(_04054_),
    .A(net7563),
    .Y(_04110_));
 sg13g2_nor3_1 _12785_ (.A(net7374),
    .B(net7276),
    .C(net7097),
    .Y(_04111_));
 sg13g2_nor2_1 _12786_ (.A(net4362),
    .B(net6732),
    .Y(_04112_));
 sg13g2_a21oi_1 _12787_ (.A1(net7328),
    .A2(net6732),
    .Y(_00089_),
    .B1(_04112_));
 sg13g2_nor2_1 _12788_ (.A(net4809),
    .B(net6732),
    .Y(_04113_));
 sg13g2_a21oi_1 _12789_ (.A1(net7526),
    .A2(net6732),
    .Y(_00090_),
    .B1(_04113_));
 sg13g2_nor2_1 _12790_ (.A(net4533),
    .B(net6733),
    .Y(_04114_));
 sg13g2_a21oi_1 _12791_ (.A1(net7684),
    .A2(net6732),
    .Y(_00091_),
    .B1(_04114_));
 sg13g2_and2_2 _12792_ (.A(_04077_),
    .B(_04084_),
    .X(_04115_));
 sg13g2_nand2_2 _12793_ (.Y(_04116_),
    .A(_04077_),
    .B(_04084_));
 sg13g2_nand2b_2 _12794_ (.Y(_04117_),
    .B(\top1.addr_in[4] ),
    .A_N(net7563));
 sg13g2_nor2_2 _12795_ (.A(_04055_),
    .B(_04117_),
    .Y(_04118_));
 sg13g2_or2_1 _12796_ (.X(_04119_),
    .B(_04117_),
    .A(_04055_));
 sg13g2_nor3_1 _12797_ (.A(net7369),
    .B(net7271),
    .C(net7092),
    .Y(_04120_));
 sg13g2_nor2_1 _12798_ (.A(net4724),
    .B(net6730),
    .Y(_04121_));
 sg13g2_a21oi_1 _12799_ (.A1(net7292),
    .A2(net6730),
    .Y(_00092_),
    .B1(_04121_));
 sg13g2_nor2_1 _12800_ (.A(net4395),
    .B(net6730),
    .Y(_04122_));
 sg13g2_a21oi_1 _12801_ (.A1(net7491),
    .A2(net6730),
    .Y(_00093_),
    .B1(_04122_));
 sg13g2_nor2_1 _12802_ (.A(net4797),
    .B(net6731),
    .Y(_04123_));
 sg13g2_a21oi_1 _12803_ (.A1(net7650),
    .A2(net6731),
    .Y(_00094_),
    .B1(_04123_));
 sg13g2_nor3_1 _12804_ (.A(net7369),
    .B(net7275),
    .C(net7092),
    .Y(_04124_));
 sg13g2_nor2_1 _12805_ (.A(net4822),
    .B(net6728),
    .Y(_04125_));
 sg13g2_a21oi_1 _12806_ (.A1(net7292),
    .A2(net6728),
    .Y(_00095_),
    .B1(_04125_));
 sg13g2_nor2_1 _12807_ (.A(net4610),
    .B(net6728),
    .Y(_04126_));
 sg13g2_a21oi_1 _12808_ (.A1(net7491),
    .A2(net6728),
    .Y(_00096_),
    .B1(_04126_));
 sg13g2_nor2_1 _12809_ (.A(net4591),
    .B(net6729),
    .Y(_04127_));
 sg13g2_a21oi_1 _12810_ (.A1(net7650),
    .A2(net6729),
    .Y(_00097_),
    .B1(_04127_));
 sg13g2_nor3_2 _12811_ (.A(net7563),
    .B(\top1.addr_in[4] ),
    .C(net7562),
    .Y(_04128_));
 sg13g2_and2_2 _12812_ (.A(_03848_),
    .B(_04128_),
    .X(_04129_));
 sg13g2_nand2_2 _12813_ (.Y(_04130_),
    .A(_03848_),
    .B(_04128_));
 sg13g2_nor3_2 _12814_ (.A(net7372),
    .B(net7276),
    .C(net7270),
    .Y(_04131_));
 sg13g2_nor2_1 _12815_ (.A(net4572),
    .B(net7090),
    .Y(_04132_));
 sg13g2_a21oi_1 _12816_ (.A1(net7319),
    .A2(net7090),
    .Y(_00098_),
    .B1(_04132_));
 sg13g2_nor2_1 _12817_ (.A(net4756),
    .B(net7091),
    .Y(_04133_));
 sg13g2_a21oi_1 _12818_ (.A1(net7520),
    .A2(net7091),
    .Y(_00099_),
    .B1(_04133_));
 sg13g2_nor2_1 _12819_ (.A(net3959),
    .B(net7090),
    .Y(_04134_));
 sg13g2_a21oi_1 _12820_ (.A1(net7676),
    .A2(net7090),
    .Y(_00100_),
    .B1(_04134_));
 sg13g2_nand3_1 _12821_ (.B(net7406),
    .C(_04058_),
    .A(net7412),
    .Y(_04135_));
 sg13g2_nor2_1 _12822_ (.A(_04041_),
    .B(net7370),
    .Y(_04136_));
 sg13g2_nor2_1 _12823_ (.A(net4621),
    .B(net6727),
    .Y(_04137_));
 sg13g2_a21oi_1 _12824_ (.A1(net7316),
    .A2(net6726),
    .Y(_00101_),
    .B1(_04137_));
 sg13g2_nor2_1 _12825_ (.A(net4355),
    .B(net6727),
    .Y(_04138_));
 sg13g2_a21oi_1 _12826_ (.A1(net7516),
    .A2(net6726),
    .Y(_00102_),
    .B1(_04138_));
 sg13g2_nor2_1 _12827_ (.A(net4842),
    .B(net6726),
    .Y(_04139_));
 sg13g2_a21oi_1 _12828_ (.A1(net7670),
    .A2(net6726),
    .Y(_00103_),
    .B1(_04139_));
 sg13g2_nor2_1 _12829_ (.A(_04043_),
    .B(_04063_),
    .Y(_04140_));
 sg13g2_nand2b_2 _12830_ (.Y(_04141_),
    .B(_04062_),
    .A_N(_04043_));
 sg13g2_nor3_2 _12831_ (.A(net7562),
    .B(_03848_),
    .C(_04049_),
    .Y(_04142_));
 sg13g2_nand3_1 _12832_ (.B(net7265),
    .C(net7262),
    .A(net7386),
    .Y(_04143_));
 sg13g2_nand2_1 _12833_ (.Y(_04144_),
    .A(net3428),
    .B(net7088));
 sg13g2_o21ai_1 _12834_ (.B1(_04144_),
    .Y(_00104_),
    .A1(net7338),
    .A2(net7088));
 sg13g2_nand2_1 _12835_ (.Y(_04145_),
    .A(net4052),
    .B(net7088));
 sg13g2_o21ai_1 _12836_ (.B1(_04145_),
    .Y(_00105_),
    .A1(net7536),
    .A2(net7088));
 sg13g2_nand2_1 _12837_ (.Y(_04146_),
    .A(net4492),
    .B(net7088));
 sg13g2_o21ai_1 _12838_ (.B1(_04146_),
    .Y(_00106_),
    .A1(net7694),
    .A2(net7088));
 sg13g2_nand3_1 _12839_ (.B(net7286),
    .C(net7261),
    .A(net7386),
    .Y(_04147_));
 sg13g2_nand2_1 _12840_ (.Y(_04148_),
    .A(net3376),
    .B(net7087));
 sg13g2_o21ai_1 _12841_ (.B1(_04148_),
    .Y(_00107_),
    .A1(net7338),
    .A2(net7087));
 sg13g2_nand2_1 _12842_ (.Y(_04149_),
    .A(net2769),
    .B(net7086));
 sg13g2_o21ai_1 _12843_ (.B1(_04149_),
    .Y(_00108_),
    .A1(net7537),
    .A2(net7086));
 sg13g2_nand2_1 _12844_ (.Y(_04150_),
    .A(net3659),
    .B(net7086));
 sg13g2_o21ai_1 _12845_ (.B1(_04150_),
    .Y(_00109_),
    .A1(net7696),
    .A2(net7086));
 sg13g2_nor2_1 _12846_ (.A(_04063_),
    .B(_04099_),
    .Y(_04151_));
 sg13g2_nand2_2 _12847_ (.Y(_04152_),
    .A(_04062_),
    .B(_04098_));
 sg13g2_nor3_2 _12848_ (.A(net7562),
    .B(_03848_),
    .C(_04108_),
    .Y(_04153_));
 sg13g2_nand4_1 _12849_ (.B(_03846_),
    .C(_03847_),
    .A(net7563),
    .Y(_04154_),
    .D(net7561));
 sg13g2_nand3_1 _12850_ (.B(net7085),
    .C(net7082),
    .A(net7382),
    .Y(_04155_));
 sg13g2_nand2_1 _12851_ (.Y(_04156_),
    .A(net2813),
    .B(net6724));
 sg13g2_o21ai_1 _12852_ (.B1(_04156_),
    .Y(_00110_),
    .A1(net7317),
    .A2(net6724));
 sg13g2_nand2_1 _12853_ (.Y(_04157_),
    .A(net3030),
    .B(net6724));
 sg13g2_o21ai_1 _12854_ (.B1(_04157_),
    .Y(_00111_),
    .A1(net7517),
    .A2(net6724));
 sg13g2_nand2_1 _12855_ (.Y(_04158_),
    .A(net3615),
    .B(net6725));
 sg13g2_o21ai_1 _12856_ (.B1(_04158_),
    .Y(_00112_),
    .A1(net7689),
    .A2(net6725));
 sg13g2_nor3_2 _12857_ (.A(net7562),
    .B(net7561),
    .C(_04108_),
    .Y(_04159_));
 sg13g2_nand3_1 _12858_ (.B(net7279),
    .C(net7072),
    .A(net7387),
    .Y(_04160_));
 sg13g2_nand2_1 _12859_ (.Y(_04161_),
    .A(net3132),
    .B(net6722));
 sg13g2_o21ai_1 _12860_ (.B1(_04161_),
    .Y(_00113_),
    .A1(net7339),
    .A2(net6722));
 sg13g2_nand2_1 _12861_ (.Y(_04162_),
    .A(net3386),
    .B(net6723));
 sg13g2_o21ai_1 _12862_ (.B1(_04162_),
    .Y(_00114_),
    .A1(net7537),
    .A2(net6723));
 sg13g2_nand2_1 _12863_ (.Y(_04163_),
    .A(net3029),
    .B(net6722));
 sg13g2_o21ai_1 _12864_ (.B1(_04163_),
    .Y(_00115_),
    .A1(net7697),
    .A2(net6722));
 sg13g2_nor3_2 _12865_ (.A(net7562),
    .B(_03848_),
    .C(_04117_),
    .Y(_04164_));
 sg13g2_nand3b_1 _12866_ (.B(_03847_),
    .C(net7561),
    .Y(_04165_),
    .A_N(_04117_));
 sg13g2_nand3_1 _12867_ (.B(net7377),
    .C(net7254),
    .A(net7403),
    .Y(_04166_));
 sg13g2_nand2_1 _12868_ (.Y(_04167_),
    .A(net2764),
    .B(net7070));
 sg13g2_o21ai_1 _12869_ (.B1(_04167_),
    .Y(_00116_),
    .A1(net7305),
    .A2(net7070));
 sg13g2_nand2_1 _12870_ (.Y(_04168_),
    .A(net2515),
    .B(net7070));
 sg13g2_o21ai_1 _12871_ (.B1(_04168_),
    .Y(_00117_),
    .A1(net7503),
    .A2(net7070));
 sg13g2_nand2_1 _12872_ (.Y(_04169_),
    .A(net3545),
    .B(net7071));
 sg13g2_o21ai_1 _12873_ (.B1(_04169_),
    .Y(_00118_),
    .A1(net7672),
    .A2(net7071));
 sg13g2_nand3_1 _12874_ (.B(net7286),
    .C(net7073),
    .A(net7395),
    .Y(_04170_));
 sg13g2_nand2_1 _12875_ (.Y(_04171_),
    .A(net2824),
    .B(net6720));
 sg13g2_o21ai_1 _12876_ (.B1(_04171_),
    .Y(_00119_),
    .A1(net7340),
    .A2(net6720));
 sg13g2_nand2_1 _12877_ (.Y(_04172_),
    .A(net2923),
    .B(net6720));
 sg13g2_o21ai_1 _12878_ (.B1(_04172_),
    .Y(_00120_),
    .A1(net7534),
    .A2(net6720));
 sg13g2_nand2_1 _12879_ (.Y(_04173_),
    .A(net4185),
    .B(net6721));
 sg13g2_o21ai_1 _12880_ (.B1(_04173_),
    .Y(_00121_),
    .A1(net7695),
    .A2(net6721));
 sg13g2_nand3_1 _12881_ (.B(net7361),
    .C(net7256),
    .A(net7377),
    .Y(_04174_));
 sg13g2_nand2_1 _12882_ (.Y(_04175_),
    .A(net3844),
    .B(net7068));
 sg13g2_o21ai_1 _12883_ (.B1(_04175_),
    .Y(_00122_),
    .A1(net7303),
    .A2(net7068));
 sg13g2_nand2_1 _12884_ (.Y(_04176_),
    .A(net3037),
    .B(net7068));
 sg13g2_o21ai_1 _12885_ (.B1(_04176_),
    .Y(_00123_),
    .A1(net7501),
    .A2(net7068));
 sg13g2_nand2_1 _12886_ (.Y(_04177_),
    .A(net2547),
    .B(net7069));
 sg13g2_o21ai_1 _12887_ (.B1(_04177_),
    .Y(_00124_),
    .A1(net7671),
    .A2(net7069));
 sg13g2_nand3_1 _12888_ (.B(net7274),
    .C(net7073),
    .A(net7395),
    .Y(_04178_));
 sg13g2_nand2_1 _12889_ (.Y(_04179_),
    .A(net2497),
    .B(net6718));
 sg13g2_o21ai_1 _12890_ (.B1(_04179_),
    .Y(_00125_),
    .A1(net7337),
    .A2(net6718));
 sg13g2_nand2_1 _12891_ (.Y(_04180_),
    .A(net3589),
    .B(net6718));
 sg13g2_o21ai_1 _12892_ (.B1(_04180_),
    .Y(_00126_),
    .A1(net7534),
    .A2(net6718));
 sg13g2_nand2_1 _12893_ (.Y(_04181_),
    .A(net3656),
    .B(net6719));
 sg13g2_o21ai_1 _12894_ (.B1(_04181_),
    .Y(_00127_),
    .A1(net7695),
    .A2(net6719));
 sg13g2_nand2_2 _12895_ (.Y(_04182_),
    .A(net7561),
    .B(_04128_));
 sg13g2_nor2_1 _12896_ (.A(_04031_),
    .B(_04099_),
    .Y(_04183_));
 sg13g2_nand2_2 _12897_ (.Y(_04184_),
    .A(_04030_),
    .B(_04098_));
 sg13g2_nor3_2 _12898_ (.A(net7367),
    .B(net7252),
    .C(_04184_),
    .Y(_04185_));
 sg13g2_nor2_1 _12899_ (.A(net3523),
    .B(net7064),
    .Y(_04186_));
 sg13g2_a21oi_1 _12900_ (.A1(net7304),
    .A2(net7064),
    .Y(_00128_),
    .B1(_04186_));
 sg13g2_nor2_1 _12901_ (.A(net4393),
    .B(net7064),
    .Y(_04187_));
 sg13g2_a21oi_1 _12902_ (.A1(net7502),
    .A2(net7064),
    .Y(_00129_),
    .B1(_04187_));
 sg13g2_nor2_1 _12903_ (.A(net4476),
    .B(net7063),
    .Y(_04188_));
 sg13g2_a21oi_1 _12904_ (.A1(net7658),
    .A2(net7063),
    .Y(_00130_),
    .B1(_04188_));
 sg13g2_nand3_1 _12905_ (.B(net7278),
    .C(net7073),
    .A(net7395),
    .Y(_04189_));
 sg13g2_nand2_1 _12906_ (.Y(_04190_),
    .A(net3765),
    .B(net6716));
 sg13g2_o21ai_1 _12907_ (.B1(_04190_),
    .Y(_00131_),
    .A1(net7337),
    .A2(net6716));
 sg13g2_nand2_1 _12908_ (.Y(_04191_),
    .A(net2905),
    .B(net6716));
 sg13g2_o21ai_1 _12909_ (.B1(_04191_),
    .Y(_00132_),
    .A1(net7535),
    .A2(net6716));
 sg13g2_nand2_1 _12910_ (.Y(_04192_),
    .A(net3953),
    .B(net6717));
 sg13g2_o21ai_1 _12911_ (.B1(_04192_),
    .Y(_00133_),
    .A1(net7695),
    .A2(net6717));
 sg13g2_nor3_2 _12912_ (.A(net7366),
    .B(net7275),
    .C(net7251),
    .Y(_04193_));
 sg13g2_nor2_1 _12913_ (.A(net4192),
    .B(net7061),
    .Y(_04194_));
 sg13g2_a21oi_1 _12914_ (.A1(net7298),
    .A2(net7061),
    .Y(_00134_),
    .B1(_04194_));
 sg13g2_nor2_1 _12915_ (.A(net3980),
    .B(net7062),
    .Y(_04195_));
 sg13g2_a21oi_1 _12916_ (.A1(net7497),
    .A2(net7062),
    .Y(_00135_),
    .B1(_04195_));
 sg13g2_nor2_1 _12917_ (.A(net4410),
    .B(net7062),
    .Y(_04196_));
 sg13g2_a21oi_1 _12918_ (.A1(net7657),
    .A2(net7062),
    .Y(_00136_),
    .B1(_04196_));
 sg13g2_and2_2 _12919_ (.A(_04032_),
    .B(_04077_),
    .X(_04197_));
 sg13g2_nand2_2 _12920_ (.Y(_04198_),
    .A(_04032_),
    .B(_04077_));
 sg13g2_nand3_1 _12921_ (.B(net7073),
    .C(net7248),
    .A(net7395),
    .Y(_04199_));
 sg13g2_nand2_1 _12922_ (.Y(_04200_),
    .A(net2617),
    .B(net6714));
 sg13g2_o21ai_1 _12923_ (.B1(_04200_),
    .Y(_00137_),
    .A1(net7337),
    .A2(net6714));
 sg13g2_nand2_1 _12924_ (.Y(_04201_),
    .A(net3808),
    .B(net6714));
 sg13g2_o21ai_1 _12925_ (.B1(_04201_),
    .Y(_00138_),
    .A1(net7535),
    .A2(net6714));
 sg13g2_nand2_1 _12926_ (.Y(_04202_),
    .A(net2916),
    .B(net6715));
 sg13g2_o21ai_1 _12927_ (.B1(_04202_),
    .Y(_00139_),
    .A1(net7695),
    .A2(net6715));
 sg13g2_nand3_1 _12928_ (.B(net7114),
    .C(net7391),
    .A(net7409),
    .Y(_04203_));
 sg13g2_nand2_1 _12929_ (.Y(_04204_),
    .A(net4041),
    .B(net6712));
 sg13g2_o21ai_1 _12930_ (.B1(_04204_),
    .Y(_00140_),
    .A1(net7346),
    .A2(net6712));
 sg13g2_nand2_1 _12931_ (.Y(_04205_),
    .A(net2951),
    .B(net6713));
 sg13g2_o21ai_1 _12932_ (.B1(_04205_),
    .Y(_00141_),
    .A1(net7544),
    .A2(net6713));
 sg13g2_nand2_1 _12933_ (.Y(_04206_),
    .A(net3869),
    .B(net6712));
 sg13g2_o21ai_1 _12934_ (.B1(_04206_),
    .Y(_00142_),
    .A1(net7703),
    .A2(net6712));
 sg13g2_nor3_2 _12935_ (.A(net7562),
    .B(\top1.addr_in[7] ),
    .C(_04117_),
    .Y(_04207_));
 sg13g2_nand3_1 _12936_ (.B(net7381),
    .C(net7244),
    .A(net7403),
    .Y(_04208_));
 sg13g2_nand2_1 _12937_ (.Y(_04209_),
    .A(net3258),
    .B(net7059));
 sg13g2_o21ai_1 _12938_ (.B1(_04209_),
    .Y(_00143_),
    .A1(net7334),
    .A2(net7059));
 sg13g2_nand2_1 _12939_ (.Y(_04210_),
    .A(net3358),
    .B(net7059));
 sg13g2_o21ai_1 _12940_ (.B1(_04210_),
    .Y(_00144_),
    .A1(net7519),
    .A2(net7059));
 sg13g2_nand2_1 _12941_ (.Y(_04211_),
    .A(net2757),
    .B(net7060));
 sg13g2_o21ai_1 _12942_ (.B1(_04211_),
    .Y(_00145_),
    .A1(net7676),
    .A2(net7060));
 sg13g2_nand3_1 _12943_ (.B(net7101),
    .C(net7266),
    .A(net7390),
    .Y(_04212_));
 sg13g2_nand2_1 _12944_ (.Y(_04213_),
    .A(net3895),
    .B(net6711));
 sg13g2_o21ai_1 _12945_ (.B1(_04213_),
    .Y(_00146_),
    .A1(net7341),
    .A2(net6710));
 sg13g2_nand2_1 _12946_ (.Y(_04214_),
    .A(net3811),
    .B(net6710));
 sg13g2_o21ai_1 _12947_ (.B1(_04214_),
    .Y(_00147_),
    .A1(net7539),
    .A2(net6710));
 sg13g2_nand2_1 _12948_ (.Y(_04215_),
    .A(net3525),
    .B(net6710));
 sg13g2_o21ai_1 _12949_ (.B1(_04215_),
    .Y(_00148_),
    .A1(net7700),
    .A2(net6711));
 sg13g2_nor2_1 _12950_ (.A(_04043_),
    .B(_04085_),
    .Y(_04216_));
 sg13g2_nand2b_2 _12951_ (.Y(_04217_),
    .B(_04084_),
    .A_N(_04043_));
 sg13g2_nand3_1 _12952_ (.B(net7243),
    .C(net7237),
    .A(net7381),
    .Y(_04218_));
 sg13g2_nand2_1 _12953_ (.Y(_04219_),
    .A(net2584),
    .B(net7058));
 sg13g2_o21ai_1 _12954_ (.B1(_04219_),
    .Y(_00149_),
    .A1(net7334),
    .A2(net7058));
 sg13g2_nand2_1 _12955_ (.Y(_04220_),
    .A(net3084),
    .B(net7057));
 sg13g2_o21ai_1 _12956_ (.B1(_04220_),
    .Y(_00150_),
    .A1(net7519),
    .A2(net7057));
 sg13g2_nand2_1 _12957_ (.Y(_04221_),
    .A(net3399),
    .B(net7057));
 sg13g2_o21ai_1 _12958_ (.B1(_04221_),
    .Y(_00151_),
    .A1(net7676),
    .A2(net7057));
 sg13g2_nor3_1 _12959_ (.A(net7374),
    .B(net7284),
    .C(net7097),
    .Y(_04222_));
 sg13g2_nor2_1 _12960_ (.A(net4356),
    .B(net6708),
    .Y(_04223_));
 sg13g2_a21oi_1 _12961_ (.A1(net7328),
    .A2(net6708),
    .Y(_00152_),
    .B1(_04223_));
 sg13g2_nor2_1 _12962_ (.A(net4664),
    .B(net6708),
    .Y(_04224_));
 sg13g2_a21oi_1 _12963_ (.A1(net7526),
    .A2(net6708),
    .Y(_00153_),
    .B1(_04224_));
 sg13g2_nor2_1 _12964_ (.A(net4244),
    .B(net6709),
    .Y(_04225_));
 sg13g2_a21oi_1 _12965_ (.A1(net7684),
    .A2(net6708),
    .Y(_00154_),
    .B1(_04225_));
 sg13g2_nor3_2 _12966_ (.A(net7372),
    .B(net7272),
    .C(net7270),
    .Y(_04226_));
 sg13g2_nor2_1 _12967_ (.A(net4742),
    .B(net7055),
    .Y(_04227_));
 sg13g2_a21oi_1 _12968_ (.A1(net7319),
    .A2(net7055),
    .Y(_00155_),
    .B1(_04227_));
 sg13g2_nor2_1 _12969_ (.A(net4466),
    .B(net7056),
    .Y(_04228_));
 sg13g2_a21oi_1 _12970_ (.A1(net7520),
    .A2(net7056),
    .Y(_00156_),
    .B1(_04228_));
 sg13g2_nor2_1 _12971_ (.A(net4156),
    .B(net7056),
    .Y(_04229_));
 sg13g2_a21oi_1 _12972_ (.A1(net7676),
    .A2(net7055),
    .Y(_00157_),
    .B1(_04229_));
 sg13g2_nand3_1 _12973_ (.B(net7094),
    .C(net7085),
    .A(net7375),
    .Y(_04230_));
 sg13g2_nand2_1 _12974_ (.Y(_04231_),
    .A(net3017),
    .B(net6707));
 sg13g2_o21ai_1 _12975_ (.B1(_04231_),
    .Y(_00158_),
    .A1(net7293),
    .A2(net6707));
 sg13g2_nand2_1 _12976_ (.Y(_04232_),
    .A(net3825),
    .B(net6706));
 sg13g2_o21ai_1 _12977_ (.B1(_04232_),
    .Y(_00159_),
    .A1(net7492),
    .A2(net6706));
 sg13g2_nand2_1 _12978_ (.Y(_04233_),
    .A(net2939),
    .B(net6707));
 sg13g2_o21ai_1 _12979_ (.B1(_04233_),
    .Y(_00160_),
    .A1(net7651),
    .A2(net6707));
 sg13g2_nor2_2 _12980_ (.A(_04033_),
    .B(_04043_),
    .Y(_04234_));
 sg13g2_or2_2 _12981_ (.X(_04235_),
    .B(_04043_),
    .A(_04033_));
 sg13g2_nand3_1 _12982_ (.B(net7243),
    .C(net7236),
    .A(net7381),
    .Y(_04236_));
 sg13g2_nand2_1 _12983_ (.Y(_04237_),
    .A(net2448),
    .B(net7054));
 sg13g2_o21ai_1 _12984_ (.B1(_04237_),
    .Y(_00161_),
    .A1(net7334),
    .A2(net7054));
 sg13g2_nand2_1 _12985_ (.Y(_04238_),
    .A(net2444),
    .B(net7053));
 sg13g2_o21ai_1 _12986_ (.B1(_04238_),
    .Y(_00162_),
    .A1(net7519),
    .A2(net7053));
 sg13g2_nand2_1 _12987_ (.Y(_04239_),
    .A(net2936),
    .B(net7053));
 sg13g2_o21ai_1 _12988_ (.B1(_04239_),
    .Y(_00163_),
    .A1(net7676),
    .A2(net7053));
 sg13g2_and2_1 _12989_ (.A(_04035_),
    .B(_04054_),
    .X(_04240_));
 sg13g2_nand2_1 _12990_ (.Y(_04241_),
    .A(_04035_),
    .B(_04054_));
 sg13g2_nor3_1 _12991_ (.A(net7402),
    .B(net7364),
    .C(net7048),
    .Y(_04242_));
 sg13g2_nor2_1 _12992_ (.A(net4757),
    .B(net6705),
    .Y(_04243_));
 sg13g2_a21oi_1 _12993_ (.A1(net7287),
    .A2(net6705),
    .Y(_00164_),
    .B1(_04243_));
 sg13g2_nor2_1 _12994_ (.A(net4059),
    .B(net6704),
    .Y(_04244_));
 sg13g2_a21oi_1 _12995_ (.A1(net7488),
    .A2(net6704),
    .Y(_00165_),
    .B1(_04244_));
 sg13g2_nor2_1 _12996_ (.A(net4854),
    .B(net6705),
    .Y(_04245_));
 sg13g2_a21oi_1 _12997_ (.A1(net7646),
    .A2(net6705),
    .Y(_00166_),
    .B1(_04245_));
 sg13g2_nand3_1 _12998_ (.B(net7065),
    .C(_04207_),
    .A(net7385),
    .Y(_04246_));
 sg13g2_nand2_1 _12999_ (.Y(_04247_),
    .A(net3423),
    .B(net6702));
 sg13g2_o21ai_1 _13000_ (.B1(_04247_),
    .Y(_00167_),
    .A1(net7334),
    .A2(net6702));
 sg13g2_nand2_1 _13001_ (.Y(_04248_),
    .A(net3956),
    .B(net6702));
 sg13g2_o21ai_1 _13002_ (.B1(_04248_),
    .Y(_00168_),
    .A1(net7530),
    .A2(net6702));
 sg13g2_nand2_1 _13003_ (.Y(_04249_),
    .A(net2950),
    .B(net6703));
 sg13g2_o21ai_1 _13004_ (.B1(_04249_),
    .Y(_00169_),
    .A1(net7691),
    .A2(net6703));
 sg13g2_nor3_2 _13005_ (.A(net7372),
    .B(_04079_),
    .C(net7270),
    .Y(_04250_));
 sg13g2_nor2_1 _13006_ (.A(net4595),
    .B(net7046),
    .Y(_04251_));
 sg13g2_a21oi_1 _13007_ (.A1(net7319),
    .A2(net7046),
    .Y(_00170_),
    .B1(_04251_));
 sg13g2_nor2_1 _13008_ (.A(net4157),
    .B(net7047),
    .Y(_04252_));
 sg13g2_a21oi_1 _13009_ (.A1(net7520),
    .A2(net7047),
    .Y(_00171_),
    .B1(_04252_));
 sg13g2_nor2_1 _13010_ (.A(net3657),
    .B(net7047),
    .Y(_04253_));
 sg13g2_a21oi_1 _13011_ (.A1(net7676),
    .A2(net7046),
    .Y(_00172_),
    .B1(_04253_));
 sg13g2_nand3_1 _13012_ (.B(net7265),
    .C(net7073),
    .A(net7395),
    .Y(_04254_));
 sg13g2_nand2_1 _13013_ (.Y(_04255_),
    .A(net3738),
    .B(net6701));
 sg13g2_o21ai_1 _13014_ (.B1(_04255_),
    .Y(_00173_),
    .A1(net7352),
    .A2(net6701));
 sg13g2_nand2_1 _13015_ (.Y(_04256_),
    .A(net3047),
    .B(net6701));
 sg13g2_o21ai_1 _13016_ (.B1(_04256_),
    .Y(_00174_),
    .A1(net7550),
    .A2(net6701));
 sg13g2_nand2_1 _13017_ (.Y(_04257_),
    .A(net3480),
    .B(net6700));
 sg13g2_o21ai_1 _13018_ (.B1(_04257_),
    .Y(_00175_),
    .A1(net7696),
    .A2(net6700));
 sg13g2_nor3_1 _13019_ (.A(net7369),
    .B(net7092),
    .C(net7245),
    .Y(_04258_));
 sg13g2_nor2_1 _13020_ (.A(net4285),
    .B(net6698),
    .Y(_04259_));
 sg13g2_a21oi_1 _13021_ (.A1(net7292),
    .A2(net6698),
    .Y(_00176_),
    .B1(_04259_));
 sg13g2_nor2_1 _13022_ (.A(net4378),
    .B(net6698),
    .Y(_04260_));
 sg13g2_a21oi_1 _13023_ (.A1(net7491),
    .A2(net6698),
    .Y(_00177_),
    .B1(_04260_));
 sg13g2_nor2_1 _13024_ (.A(net4835),
    .B(net6699),
    .Y(_04261_));
 sg13g2_a21oi_1 _13025_ (.A1(net7650),
    .A2(net6699),
    .Y(_00178_),
    .B1(_04261_));
 sg13g2_nand3_1 _13026_ (.B(net7383),
    .C(_04129_),
    .A(net7407),
    .Y(_04262_));
 sg13g2_nand2_1 _13027_ (.Y(_04263_),
    .A(net2788),
    .B(net7044));
 sg13g2_o21ai_1 _13028_ (.B1(_04263_),
    .Y(_00179_),
    .A1(net7320),
    .A2(net7044));
 sg13g2_nand2_1 _13029_ (.Y(_04264_),
    .A(net3625),
    .B(net7045));
 sg13g2_o21ai_1 _13030_ (.B1(_04264_),
    .Y(_00180_),
    .A1(net7519),
    .A2(net7045));
 sg13g2_nand2_1 _13031_ (.Y(_04265_),
    .A(net2832),
    .B(net7044));
 sg13g2_o21ai_1 _13032_ (.B1(_04265_),
    .Y(_00181_),
    .A1(net7675),
    .A2(net7044));
 sg13g2_nor3_1 _13033_ (.A(net7364),
    .B(_04217_),
    .C(net7048),
    .Y(_04266_));
 sg13g2_nor2_1 _13034_ (.A(net4637),
    .B(net6697),
    .Y(_04267_));
 sg13g2_a21oi_1 _13035_ (.A1(net7287),
    .A2(net6697),
    .Y(_00182_),
    .B1(_04267_));
 sg13g2_nor2_1 _13036_ (.A(net4778),
    .B(net6696),
    .Y(_04268_));
 sg13g2_a21oi_1 _13037_ (.A1(net7488),
    .A2(net6696),
    .Y(_00183_),
    .B1(_04268_));
 sg13g2_nor2_1 _13038_ (.A(net3873),
    .B(net6697),
    .Y(_04269_));
 sg13g2_a21oi_1 _13039_ (.A1(net7646),
    .A2(net6697),
    .Y(_00184_),
    .B1(_04269_));
 sg13g2_nor3_1 _13040_ (.A(net7364),
    .B(_04141_),
    .C(net7048),
    .Y(_04270_));
 sg13g2_nor2_1 _13041_ (.A(net3903),
    .B(net6695),
    .Y(_04271_));
 sg13g2_a21oi_1 _13042_ (.A1(net7287),
    .A2(net6695),
    .Y(_00185_),
    .B1(_04271_));
 sg13g2_nor2_1 _13043_ (.A(net4795),
    .B(net6694),
    .Y(_04272_));
 sg13g2_a21oi_1 _13044_ (.A1(net7488),
    .A2(net6694),
    .Y(_00186_),
    .B1(_04272_));
 sg13g2_nor2_1 _13045_ (.A(net4856),
    .B(net6695),
    .Y(_04273_));
 sg13g2_a21oi_1 _13046_ (.A1(net7646),
    .A2(net6695),
    .Y(_00187_),
    .B1(_04273_));
 sg13g2_nor3_1 _13047_ (.A(net7364),
    .B(_04235_),
    .C(net7048),
    .Y(_04274_));
 sg13g2_nor2_1 _13048_ (.A(net4314),
    .B(net6693),
    .Y(_04275_));
 sg13g2_a21oi_1 _13049_ (.A1(net7287),
    .A2(net6693),
    .Y(_00188_),
    .B1(_04275_));
 sg13g2_nor2_1 _13050_ (.A(net4814),
    .B(net6692),
    .Y(_04276_));
 sg13g2_a21oi_1 _13051_ (.A1(net7488),
    .A2(net6692),
    .Y(_00189_),
    .B1(_04276_));
 sg13g2_nor2_1 _13052_ (.A(net4550),
    .B(net6693),
    .Y(_04277_));
 sg13g2_a21oi_1 _13053_ (.A1(net7646),
    .A2(net6693),
    .Y(_00190_),
    .B1(_04277_));
 sg13g2_nor3_2 _13054_ (.A(net7365),
    .B(_04184_),
    .C(net7051),
    .Y(_04278_));
 sg13g2_nor2_1 _13055_ (.A(net3914),
    .B(net6691),
    .Y(_04279_));
 sg13g2_a21oi_1 _13056_ (.A1(net7294),
    .A2(net6690),
    .Y(_00191_),
    .B1(_04279_));
 sg13g2_nor2_1 _13057_ (.A(net4377),
    .B(net6690),
    .Y(_04280_));
 sg13g2_a21oi_1 _13058_ (.A1(net7492),
    .A2(net6691),
    .Y(_00192_),
    .B1(_04280_));
 sg13g2_nor2_1 _13059_ (.A(net4029),
    .B(net6691),
    .Y(_04281_));
 sg13g2_a21oi_1 _13060_ (.A1(net7649),
    .A2(net6691),
    .Y(_00193_),
    .B1(_04281_));
 sg13g2_nor3_2 _13061_ (.A(net7365),
    .B(_04101_),
    .C(net7051),
    .Y(_04282_));
 sg13g2_nor2_1 _13062_ (.A(net4163),
    .B(net6689),
    .Y(_04283_));
 sg13g2_a21oi_1 _13063_ (.A1(net7294),
    .A2(net6689),
    .Y(_00194_),
    .B1(_04283_));
 sg13g2_nor2_1 _13064_ (.A(net3871),
    .B(net6688),
    .Y(_04284_));
 sg13g2_a21oi_1 _13065_ (.A1(net7492),
    .A2(net6688),
    .Y(_00195_),
    .B1(_04284_));
 sg13g2_nor2_1 _13066_ (.A(net4434),
    .B(net6689),
    .Y(_04285_));
 sg13g2_a21oi_1 _13067_ (.A1(net7645),
    .A2(net6689),
    .Y(_00196_),
    .B1(_04285_));
 sg13g2_nor3_2 _13068_ (.A(net7365),
    .B(_04152_),
    .C(net7051),
    .Y(_04286_));
 sg13g2_nor2_1 _13069_ (.A(net4441),
    .B(net6686),
    .Y(_04287_));
 sg13g2_a21oi_1 _13070_ (.A1(net7294),
    .A2(net6686),
    .Y(_00197_),
    .B1(_04287_));
 sg13g2_nor2_1 _13071_ (.A(net4738),
    .B(net6687),
    .Y(_04288_));
 sg13g2_a21oi_1 _13072_ (.A1(net7492),
    .A2(net6687),
    .Y(_00198_),
    .B1(_04288_));
 sg13g2_nor2_1 _13073_ (.A(net4390),
    .B(net6687),
    .Y(_04289_));
 sg13g2_a21oi_1 _13074_ (.A1(net7645),
    .A2(net6687),
    .Y(_00199_),
    .B1(_04289_));
 sg13g2_nor2_1 _13075_ (.A(_04033_),
    .B(_04099_),
    .Y(_04290_));
 sg13g2_nand2_2 _13076_ (.Y(_04291_),
    .A(_04032_),
    .B(_04098_));
 sg13g2_nor3_2 _13077_ (.A(net7365),
    .B(net7051),
    .C(net7234),
    .Y(_04292_));
 sg13g2_nor2_1 _13078_ (.A(net4654),
    .B(net6684),
    .Y(_04293_));
 sg13g2_a21oi_1 _13079_ (.A1(net7294),
    .A2(net6684),
    .Y(_00200_),
    .B1(_04293_));
 sg13g2_nor2_1 _13080_ (.A(net4342),
    .B(net6685),
    .Y(_04294_));
 sg13g2_a21oi_1 _13081_ (.A1(net7492),
    .A2(net6685),
    .Y(_00201_),
    .B1(_04294_));
 sg13g2_nor2_1 _13082_ (.A(net4406),
    .B(net6685),
    .Y(_04295_));
 sg13g2_a21oi_1 _13083_ (.A1(net7645),
    .A2(net6685),
    .Y(_00202_),
    .B1(_04295_));
 sg13g2_nand3_1 _13084_ (.B(net7376),
    .C(_04240_),
    .A(net7406),
    .Y(_04296_));
 sg13g2_nand2_1 _13085_ (.Y(_04297_),
    .A(net3649),
    .B(net6682));
 sg13g2_o21ai_1 _13086_ (.B1(_04297_),
    .Y(_00203_),
    .A1(net7294),
    .A2(net6682));
 sg13g2_nand2_1 _13087_ (.Y(_04298_),
    .A(net3299),
    .B(net6682));
 sg13g2_o21ai_1 _13088_ (.B1(_04298_),
    .Y(_00204_),
    .A1(net7493),
    .A2(net6682));
 sg13g2_nand2_1 _13089_ (.Y(_04299_),
    .A(net2853),
    .B(net6682));
 sg13g2_o21ai_1 _13090_ (.B1(_04299_),
    .Y(_00205_),
    .A1(net7649),
    .A2(net6682));
 sg13g2_nor3_1 _13091_ (.A(net7374),
    .B(net7097),
    .C(net7246),
    .Y(_04300_));
 sg13g2_nor2_1 _13092_ (.A(net4848),
    .B(net6680),
    .Y(_04301_));
 sg13g2_a21oi_1 _13093_ (.A1(net7328),
    .A2(net6680),
    .Y(_00206_),
    .B1(_04301_));
 sg13g2_nor2_1 _13094_ (.A(net4514),
    .B(net6680),
    .Y(_04302_));
 sg13g2_a21oi_1 _13095_ (.A1(net7526),
    .A2(net6680),
    .Y(_00207_),
    .B1(_04302_));
 sg13g2_nor2_1 _13096_ (.A(net4820),
    .B(net6681),
    .Y(_04303_));
 sg13g2_a21oi_1 _13097_ (.A1(net7684),
    .A2(net6680),
    .Y(_00208_),
    .B1(_04303_));
 sg13g2_nor3_1 _13098_ (.A(net7365),
    .B(_04087_),
    .C(net7051),
    .Y(_04304_));
 sg13g2_nor2_1 _13099_ (.A(net4178),
    .B(net6678),
    .Y(_04305_));
 sg13g2_a21oi_1 _13100_ (.A1(net7294),
    .A2(net6678),
    .Y(_00209_),
    .B1(_04305_));
 sg13g2_nor2_1 _13101_ (.A(net4417),
    .B(net6678),
    .Y(_04306_));
 sg13g2_a21oi_1 _13102_ (.A1(net7492),
    .A2(net6678),
    .Y(_00210_),
    .B1(_04306_));
 sg13g2_nor2_1 _13103_ (.A(net4167),
    .B(net6678),
    .Y(_04307_));
 sg13g2_a21oi_1 _13104_ (.A1(net7649),
    .A2(net6678),
    .Y(_00211_),
    .B1(_04307_));
 sg13g2_nand3_1 _13105_ (.B(net7375),
    .C(net7094),
    .A(net7403),
    .Y(_04308_));
 sg13g2_nand2_1 _13106_ (.Y(_04309_),
    .A(net2656),
    .B(net6676));
 sg13g2_o21ai_1 _13107_ (.B1(_04309_),
    .Y(_00212_),
    .A1(net7292),
    .A2(net6676));
 sg13g2_nand2_1 _13108_ (.Y(_04310_),
    .A(net3056),
    .B(net6676));
 sg13g2_o21ai_1 _13109_ (.B1(_04310_),
    .Y(_00213_),
    .A1(net7504),
    .A2(net6676));
 sg13g2_nand2_1 _13110_ (.Y(_04311_),
    .A(net2632),
    .B(net6676));
 sg13g2_o21ai_1 _13111_ (.B1(_04311_),
    .Y(_00214_),
    .A1(net7650),
    .A2(net6676));
 sg13g2_nor3_1 _13112_ (.A(net7373),
    .B(_04087_),
    .C(net7269),
    .Y(_04312_));
 sg13g2_nor2_1 _13113_ (.A(net4617),
    .B(net6675),
    .Y(_04313_));
 sg13g2_a21oi_1 _13114_ (.A1(net7320),
    .A2(net6675),
    .Y(_00215_),
    .B1(_04313_));
 sg13g2_nor2_1 _13115_ (.A(net4798),
    .B(net6675),
    .Y(_04314_));
 sg13g2_a21oi_1 _13116_ (.A1(net7519),
    .A2(net6675),
    .Y(_00216_),
    .B1(_04314_));
 sg13g2_nor2_1 _13117_ (.A(net4667),
    .B(net6674),
    .Y(_04315_));
 sg13g2_a21oi_1 _13118_ (.A1(net7675),
    .A2(net6674),
    .Y(_00217_),
    .B1(_04315_));
 sg13g2_nand3_1 _13119_ (.B(net7391),
    .C(net7084),
    .A(net7115),
    .Y(_04316_));
 sg13g2_nand2_1 _13120_ (.Y(_04317_),
    .A(net2587),
    .B(net6672));
 sg13g2_o21ai_1 _13121_ (.B1(_04317_),
    .Y(_00218_),
    .A1(net7344),
    .A2(net6672));
 sg13g2_nand2_1 _13122_ (.Y(_04318_),
    .A(net3417),
    .B(net6672));
 sg13g2_o21ai_1 _13123_ (.B1(_04318_),
    .Y(_00219_),
    .A1(net7542),
    .A2(net6672));
 sg13g2_nand2_1 _13124_ (.Y(_04319_),
    .A(net3069),
    .B(net6673));
 sg13g2_o21ai_1 _13125_ (.B1(_04319_),
    .Y(_00220_),
    .A1(net7708),
    .A2(net6673));
 sg13g2_nand3_1 _13126_ (.B(net7391),
    .C(net7043),
    .A(net7115),
    .Y(_04320_));
 sg13g2_nand2_1 _13127_ (.Y(_04321_),
    .A(net3566),
    .B(net6670));
 sg13g2_o21ai_1 _13128_ (.B1(_04321_),
    .Y(_00221_),
    .A1(net7344),
    .A2(net6670));
 sg13g2_nand2_1 _13129_ (.Y(_04322_),
    .A(net3228),
    .B(net6670));
 sg13g2_o21ai_1 _13130_ (.B1(_04322_),
    .Y(_00222_),
    .A1(net7542),
    .A2(net6670));
 sg13g2_nand2_1 _13131_ (.Y(_04323_),
    .A(net3367),
    .B(net6671));
 sg13g2_o21ai_1 _13132_ (.B1(_04323_),
    .Y(_00223_),
    .A1(net7702),
    .A2(net6671));
 sg13g2_nand3_1 _13133_ (.B(_04129_),
    .C(net7067),
    .A(net7383),
    .Y(_04324_));
 sg13g2_nand2_1 _13134_ (.Y(_04325_),
    .A(net4076),
    .B(net6668));
 sg13g2_o21ai_1 _13135_ (.B1(_04325_),
    .Y(_00224_),
    .A1(net7319),
    .A2(net6668));
 sg13g2_nand2_1 _13136_ (.Y(_04326_),
    .A(net3353),
    .B(net6668));
 sg13g2_o21ai_1 _13137_ (.B1(_04326_),
    .Y(_00225_),
    .A1(net7520),
    .A2(net6668));
 sg13g2_nand2_1 _13138_ (.Y(_04327_),
    .A(net3707),
    .B(net6669));
 sg13g2_o21ai_1 _13139_ (.B1(_04327_),
    .Y(_00226_),
    .A1(net7675),
    .A2(net6669));
 sg13g2_nand3_1 _13140_ (.B(net7391),
    .C(net7283),
    .A(net7114),
    .Y(_04328_));
 sg13g2_nand2_1 _13141_ (.Y(_04329_),
    .A(net3349),
    .B(net6666));
 sg13g2_o21ai_1 _13142_ (.B1(_04329_),
    .Y(_00227_),
    .A1(net7346),
    .A2(net6666));
 sg13g2_nand2_1 _13143_ (.Y(_04330_),
    .A(net2945),
    .B(net6667));
 sg13g2_o21ai_1 _13144_ (.B1(_04330_),
    .Y(_00228_),
    .A1(net7544),
    .A2(net6667));
 sg13g2_nand2_1 _13145_ (.Y(_04331_),
    .A(net3343),
    .B(net6666));
 sg13g2_o21ai_1 _13146_ (.B1(_04331_),
    .Y(_00229_),
    .A1(net7703),
    .A2(net6666));
 sg13g2_nand3_1 _13147_ (.B(net7391),
    .C(net7363),
    .A(net7114),
    .Y(_04332_));
 sg13g2_nand2_1 _13148_ (.Y(_04333_),
    .A(net3732),
    .B(net6664));
 sg13g2_o21ai_1 _13149_ (.B1(_04333_),
    .Y(_00230_),
    .A1(net7346),
    .A2(net6664));
 sg13g2_nand2_1 _13150_ (.Y(_04334_),
    .A(net3107),
    .B(net6665));
 sg13g2_o21ai_1 _13151_ (.B1(_04334_),
    .Y(_00231_),
    .A1(net7544),
    .A2(net6665));
 sg13g2_nand2_1 _13152_ (.Y(_04335_),
    .A(net3557),
    .B(net6664));
 sg13g2_o21ai_1 _13153_ (.B1(_04335_),
    .Y(_00232_),
    .A1(net7703),
    .A2(net6664));
 sg13g2_nand3_1 _13154_ (.B(net7379),
    .C(net7273),
    .A(net7411),
    .Y(_04336_));
 sg13g2_nand2_1 _13155_ (.Y(_04337_),
    .A(net2601),
    .B(net7040));
 sg13g2_o21ai_1 _13156_ (.B1(_04337_),
    .Y(_00233_),
    .A1(net7316),
    .A2(net7040));
 sg13g2_nand2_1 _13157_ (.Y(_04338_),
    .A(net3058),
    .B(net7041));
 sg13g2_o21ai_1 _13158_ (.B1(_04338_),
    .Y(_00234_),
    .A1(net7516),
    .A2(net7040));
 sg13g2_nand2_1 _13159_ (.Y(_04339_),
    .A(net3586),
    .B(net7041));
 sg13g2_o21ai_1 _13160_ (.B1(_04339_),
    .Y(_00235_),
    .A1(net7674),
    .A2(net7041));
 sg13g2_nand3_1 _13161_ (.B(net7379),
    .C(net7277),
    .A(net7411),
    .Y(_04340_));
 sg13g2_nand2_1 _13162_ (.Y(_04341_),
    .A(net2959),
    .B(net7038));
 sg13g2_o21ai_1 _13163_ (.B1(_04341_),
    .Y(_00236_),
    .A1(net7315),
    .A2(net7038));
 sg13g2_nand2_1 _13164_ (.Y(_04342_),
    .A(net2693),
    .B(net7039));
 sg13g2_o21ai_1 _13165_ (.B1(_04342_),
    .Y(_00237_),
    .A1(net7516),
    .A2(net7039));
 sg13g2_nand2_1 _13166_ (.Y(_04343_),
    .A(net3008),
    .B(net7038));
 sg13g2_o21ai_1 _13167_ (.B1(_04343_),
    .Y(_00238_),
    .A1(net7670),
    .A2(net7038));
 sg13g2_nand3_1 _13168_ (.B(net7379),
    .C(net7247),
    .A(net7411),
    .Y(_04344_));
 sg13g2_nand2_1 _13169_ (.Y(_04345_),
    .A(net2563),
    .B(net7036));
 sg13g2_o21ai_1 _13170_ (.B1(_04345_),
    .Y(_00239_),
    .A1(net7316),
    .A2(net7036));
 sg13g2_nand2_1 _13171_ (.Y(_04346_),
    .A(net3240),
    .B(net7036));
 sg13g2_o21ai_1 _13172_ (.B1(_04346_),
    .Y(_00240_),
    .A1(net7516),
    .A2(net7036));
 sg13g2_nand2_1 _13173_ (.Y(_04347_),
    .A(net4332),
    .B(net7036));
 sg13g2_o21ai_1 _13174_ (.B1(_04347_),
    .Y(_00241_),
    .A1(net7674),
    .A2(net7036));
 sg13g2_nand3_1 _13175_ (.B(net7386),
    .C(net7262),
    .A(net7404),
    .Y(_04348_));
 sg13g2_nand2_1 _13176_ (.Y(_04349_),
    .A(net2445),
    .B(net7034));
 sg13g2_o21ai_1 _13177_ (.B1(_04349_),
    .Y(_00242_),
    .A1(net7338),
    .A2(net7034));
 sg13g2_nand2_1 _13178_ (.Y(_04350_),
    .A(net2870),
    .B(net7035));
 sg13g2_o21ai_1 _13179_ (.B1(_04350_),
    .Y(_00243_),
    .A1(net7536),
    .A2(net7034));
 sg13g2_nand2_1 _13180_ (.Y(_04351_),
    .A(net3734),
    .B(net7034));
 sg13g2_o21ai_1 _13181_ (.B1(_04351_),
    .Y(_00244_),
    .A1(net7694),
    .A2(net7034));
 sg13g2_nand3_1 _13182_ (.B(net7262),
    .C(net7238),
    .A(net7386),
    .Y(_04352_));
 sg13g2_nand2_1 _13183_ (.Y(_04353_),
    .A(net3522),
    .B(net7032));
 sg13g2_o21ai_1 _13184_ (.B1(_04353_),
    .Y(_00245_),
    .A1(net7338),
    .A2(net7032));
 sg13g2_nand2_1 _13185_ (.Y(_04354_),
    .A(net3932),
    .B(net7033));
 sg13g2_o21ai_1 _13186_ (.B1(_04354_),
    .Y(_00246_),
    .A1(net7536),
    .A2(net7033));
 sg13g2_nand2_1 _13187_ (.Y(_04355_),
    .A(net3896),
    .B(net7032));
 sg13g2_o21ai_1 _13188_ (.B1(_04355_),
    .Y(_00247_),
    .A1(net7694),
    .A2(net7032));
 sg13g2_nand3_1 _13189_ (.B(net7273),
    .C(net7244),
    .A(net7385),
    .Y(_04356_));
 sg13g2_nand2_1 _13190_ (.Y(_04357_),
    .A(net3797),
    .B(net7030));
 sg13g2_o21ai_1 _13191_ (.B1(_04357_),
    .Y(_00248_),
    .A1(net7335),
    .A2(net7030));
 sg13g2_nand2_1 _13192_ (.Y(_04358_),
    .A(net3698),
    .B(net7031));
 sg13g2_o21ai_1 _13193_ (.B1(_04358_),
    .Y(_00249_),
    .A1(net7531),
    .A2(net7031));
 sg13g2_nand2_1 _13194_ (.Y(_04359_),
    .A(net4027),
    .B(net7031));
 sg13g2_o21ai_1 _13195_ (.B1(_04359_),
    .Y(_00250_),
    .A1(net7691),
    .A2(net7031));
 sg13g2_nand3_1 _13196_ (.B(net7262),
    .C(net7235),
    .A(net7386),
    .Y(_04360_));
 sg13g2_nand2_1 _13197_ (.Y(_04361_),
    .A(net3210),
    .B(net7028));
 sg13g2_o21ai_1 _13198_ (.B1(_04361_),
    .Y(_00251_),
    .A1(net7338),
    .A2(net7028));
 sg13g2_nand2_1 _13199_ (.Y(_04362_),
    .A(net3341),
    .B(net7028));
 sg13g2_o21ai_1 _13200_ (.B1(_04362_),
    .Y(_00252_),
    .A1(net7536),
    .A2(net7028));
 sg13g2_nand2_1 _13201_ (.Y(_04363_),
    .A(net3908),
    .B(net7028));
 sg13g2_o21ai_1 _13202_ (.B1(_04363_),
    .Y(_00253_),
    .A1(net7694),
    .A2(net7028));
 sg13g2_nand3_1 _13203_ (.B(net7261),
    .C(net7066),
    .A(net7389),
    .Y(_04364_));
 sg13g2_nand2_1 _13204_ (.Y(_04365_),
    .A(net3291),
    .B(net6662));
 sg13g2_o21ai_1 _13205_ (.B1(_04365_),
    .Y(_00254_),
    .A1(net7335),
    .A2(net6662));
 sg13g2_nand2_1 _13206_ (.Y(_04366_),
    .A(net2501),
    .B(net6662));
 sg13g2_o21ai_1 _13207_ (.B1(_04366_),
    .Y(_00255_),
    .A1(net7536),
    .A2(net6662));
 sg13g2_nand2_1 _13208_ (.Y(_04367_),
    .A(net3032),
    .B(net6662));
 sg13g2_o21ai_1 _13209_ (.B1(_04367_),
    .Y(_00256_),
    .A1(net7692),
    .A2(net6663));
 sg13g2_nand3_1 _13210_ (.B(net7102),
    .C(net7261),
    .A(net7389),
    .Y(_04368_));
 sg13g2_nand2_1 _13211_ (.Y(_04369_),
    .A(net2810),
    .B(net6660));
 sg13g2_o21ai_1 _13212_ (.B1(_04369_),
    .Y(_00257_),
    .A1(net7335),
    .A2(net6660));
 sg13g2_nand2_1 _13213_ (.Y(_04370_),
    .A(net3374),
    .B(net6660));
 sg13g2_o21ai_1 _13214_ (.B1(_04370_),
    .Y(_00258_),
    .A1(net7536),
    .A2(net6660));
 sg13g2_nand2_1 _13215_ (.Y(_04371_),
    .A(net3517),
    .B(net6660));
 sg13g2_o21ai_1 _13216_ (.B1(_04371_),
    .Y(_00259_),
    .A1(net7691),
    .A2(net6661));
 sg13g2_nand3_1 _13217_ (.B(net7261),
    .C(net7083),
    .A(net7385),
    .Y(_04372_));
 sg13g2_nand2_1 _13218_ (.Y(_04373_),
    .A(net3697),
    .B(net6658));
 sg13g2_o21ai_1 _13219_ (.B1(_04373_),
    .Y(_00260_),
    .A1(net7335),
    .A2(net6658));
 sg13g2_nand2_1 _13220_ (.Y(_04374_),
    .A(net3801),
    .B(net6658));
 sg13g2_o21ai_1 _13221_ (.B1(_04374_),
    .Y(_00261_),
    .A1(net7532),
    .A2(net6658));
 sg13g2_nand2_1 _13222_ (.Y(_04375_),
    .A(net3713),
    .B(net6658));
 sg13g2_o21ai_1 _13223_ (.B1(_04375_),
    .Y(_00262_),
    .A1(net7691),
    .A2(net6659));
 sg13g2_nand3_1 _13224_ (.B(net7261),
    .C(net7042),
    .A(net7385),
    .Y(_04376_));
 sg13g2_nand2_1 _13225_ (.Y(_04377_),
    .A(net2447),
    .B(net6656));
 sg13g2_o21ai_1 _13226_ (.B1(_04377_),
    .Y(_00263_),
    .A1(net7335),
    .A2(net6656));
 sg13g2_nand2_1 _13227_ (.Y(_04378_),
    .A(net2718),
    .B(net6656));
 sg13g2_o21ai_1 _13228_ (.B1(_04378_),
    .Y(_00264_),
    .A1(net7532),
    .A2(net6656));
 sg13g2_nand2_1 _13229_ (.Y(_04379_),
    .A(net3043),
    .B(net6656));
 sg13g2_o21ai_1 _13230_ (.B1(_04379_),
    .Y(_00265_),
    .A1(net7691),
    .A2(net6657));
 sg13g2_nand3_1 _13231_ (.B(net7388),
    .C(net7263),
    .A(net7408),
    .Y(_04380_));
 sg13g2_nand2_1 _13232_ (.Y(_04381_),
    .A(net2833),
    .B(net7026));
 sg13g2_o21ai_1 _13233_ (.B1(_04381_),
    .Y(_00266_),
    .A1(net7337),
    .A2(net7026));
 sg13g2_nand2_1 _13234_ (.Y(_04382_),
    .A(net3179),
    .B(net7026));
 sg13g2_o21ai_1 _13235_ (.B1(_04382_),
    .Y(_00267_),
    .A1(net7534),
    .A2(net7026));
 sg13g2_nand2_1 _13236_ (.Y(_04383_),
    .A(net2676),
    .B(net7027));
 sg13g2_o21ai_1 _13237_ (.B1(_04383_),
    .Y(_00268_),
    .A1(net7694),
    .A2(net7027));
 sg13g2_nand3_1 _13238_ (.B(net7282),
    .C(net7263),
    .A(net7388),
    .Y(_04384_));
 sg13g2_nand2_1 _13239_ (.Y(_04385_),
    .A(net3856),
    .B(net7024));
 sg13g2_o21ai_1 _13240_ (.B1(_04385_),
    .Y(_00269_),
    .A1(net7337),
    .A2(net7024));
 sg13g2_nand2_1 _13241_ (.Y(_04386_),
    .A(net2780),
    .B(net7024));
 sg13g2_o21ai_1 _13242_ (.B1(_04386_),
    .Y(_00270_),
    .A1(net7534),
    .A2(net7024));
 sg13g2_nand2_1 _13243_ (.Y(_04387_),
    .A(net3264),
    .B(net7025));
 sg13g2_o21ai_1 _13244_ (.B1(_04387_),
    .Y(_00271_),
    .A1(net7694),
    .A2(net7024));
 sg13g2_nand3_1 _13245_ (.B(net7362),
    .C(net7263),
    .A(net7388),
    .Y(_04388_));
 sg13g2_nand2_1 _13246_ (.Y(_04389_),
    .A(net3693),
    .B(net7022));
 sg13g2_o21ai_1 _13247_ (.B1(_04389_),
    .Y(_00272_),
    .A1(net7337),
    .A2(net7022));
 sg13g2_nand2_1 _13248_ (.Y(_04390_),
    .A(net3500),
    .B(net7022));
 sg13g2_o21ai_1 _13249_ (.B1(_04390_),
    .Y(_00273_),
    .A1(net7533),
    .A2(net7022));
 sg13g2_nand2_1 _13250_ (.Y(_04391_),
    .A(net3110),
    .B(net7023));
 sg13g2_o21ai_1 _13251_ (.B1(_04391_),
    .Y(_00274_),
    .A1(net7694),
    .A2(net7023));
 sg13g2_nand3_1 _13252_ (.B(net7279),
    .C(net7263),
    .A(net7388),
    .Y(_04392_));
 sg13g2_nand2_1 _13253_ (.Y(_04393_),
    .A(net3231),
    .B(net7020));
 sg13g2_o21ai_1 _13254_ (.B1(_04393_),
    .Y(_00275_),
    .A1(net7337),
    .A2(net7020));
 sg13g2_nand2_1 _13255_ (.Y(_04394_),
    .A(net2992),
    .B(net7020));
 sg13g2_o21ai_1 _13256_ (.B1(_04394_),
    .Y(_00276_),
    .A1(net7533),
    .A2(net7020));
 sg13g2_nand2_1 _13257_ (.Y(_04395_),
    .A(net3252),
    .B(net7021));
 sg13g2_o21ai_1 _13258_ (.B1(_04395_),
    .Y(_00277_),
    .A1(net7694),
    .A2(net7021));
 sg13g2_nand3_1 _13259_ (.B(net7277),
    .C(net7244),
    .A(net7385),
    .Y(_04396_));
 sg13g2_nand2_1 _13260_ (.Y(_04397_),
    .A(net3105),
    .B(net7018));
 sg13g2_o21ai_1 _13261_ (.B1(_04397_),
    .Y(_00278_),
    .A1(net7335),
    .A2(net7018));
 sg13g2_nand2_1 _13262_ (.Y(_04398_),
    .A(net2993),
    .B(net7019));
 sg13g2_o21ai_1 _13263_ (.B1(_04398_),
    .Y(_00279_),
    .A1(net7530),
    .A2(net7019));
 sg13g2_nand2_1 _13264_ (.Y(_04399_),
    .A(net2820),
    .B(net7019));
 sg13g2_o21ai_1 _13265_ (.B1(_04399_),
    .Y(_00280_),
    .A1(net7691),
    .A2(net7019));
 sg13g2_nand3_1 _13266_ (.B(net7273),
    .C(net7261),
    .A(net7386),
    .Y(_04400_));
 sg13g2_nand2_1 _13267_ (.Y(_04401_),
    .A(net2882),
    .B(net7017));
 sg13g2_o21ai_1 _13268_ (.B1(_04401_),
    .Y(_00281_),
    .A1(net7338),
    .A2(net7017));
 sg13g2_nand2_1 _13269_ (.Y(_04402_),
    .A(net3930),
    .B(net7016));
 sg13g2_o21ai_1 _13270_ (.B1(_04402_),
    .Y(_00282_),
    .A1(net7537),
    .A2(net7016));
 sg13g2_nand2_1 _13271_ (.Y(_04403_),
    .A(net3770),
    .B(net7016));
 sg13g2_o21ai_1 _13272_ (.B1(_04403_),
    .Y(_00283_),
    .A1(net7696),
    .A2(net7016));
 sg13g2_nand3_1 _13273_ (.B(net7277),
    .C(net7261),
    .A(net7386),
    .Y(_04404_));
 sg13g2_nand2_1 _13274_ (.Y(_04405_),
    .A(net2627),
    .B(net7014));
 sg13g2_o21ai_1 _13275_ (.B1(_04405_),
    .Y(_00284_),
    .A1(net7338),
    .A2(net7014));
 sg13g2_nand2_1 _13276_ (.Y(_04406_),
    .A(net3813),
    .B(net7014));
 sg13g2_o21ai_1 _13277_ (.B1(_04406_),
    .Y(_00285_),
    .A1(net7536),
    .A2(net7014));
 sg13g2_nand2_1 _13278_ (.Y(_04407_),
    .A(net2766),
    .B(net7014));
 sg13g2_o21ai_1 _13279_ (.B1(_04407_),
    .Y(_00286_),
    .A1(net7696),
    .A2(net7014));
 sg13g2_nand3_1 _13280_ (.B(net7261),
    .C(net7247),
    .A(net7386),
    .Y(_04408_));
 sg13g2_nand2_1 _13281_ (.Y(_04409_),
    .A(net2744),
    .B(net7012));
 sg13g2_o21ai_1 _13282_ (.B1(_04409_),
    .Y(_00287_),
    .A1(net7338),
    .A2(net7012));
 sg13g2_nand2_1 _13283_ (.Y(_04410_),
    .A(net3235),
    .B(net7012));
 sg13g2_o21ai_1 _13284_ (.B1(_04410_),
    .Y(_00288_),
    .A1(net7536),
    .A2(net7012));
 sg13g2_nand2_1 _13285_ (.Y(_04411_),
    .A(net2912),
    .B(net7012));
 sg13g2_o21ai_1 _13286_ (.B1(_04411_),
    .Y(_00289_),
    .A1(net7696),
    .A2(net7012));
 sg13g2_nand3_1 _13287_ (.B(net7384),
    .C(net7079),
    .A(net7404),
    .Y(_04412_));
 sg13g2_nand2_1 _13288_ (.Y(_04413_),
    .A(net4172),
    .B(net6654));
 sg13g2_o21ai_1 _13289_ (.B1(_04413_),
    .Y(_00290_),
    .A1(net7313),
    .A2(net6654));
 sg13g2_nand2_1 _13290_ (.Y(_04414_),
    .A(net2471),
    .B(net6655));
 sg13g2_o21ai_1 _13291_ (.B1(_04414_),
    .Y(_00291_),
    .A1(net7511),
    .A2(net6654));
 sg13g2_nand2_1 _13292_ (.Y(_04415_),
    .A(net3159),
    .B(net6655));
 sg13g2_o21ai_1 _13293_ (.B1(_04415_),
    .Y(_00292_),
    .A1(net7682),
    .A2(net6655));
 sg13g2_nand3_1 _13294_ (.B(net7078),
    .C(net7237),
    .A(net7384),
    .Y(_04416_));
 sg13g2_nand2_1 _13295_ (.Y(_04417_),
    .A(net3279),
    .B(net6652));
 sg13g2_o21ai_1 _13296_ (.B1(_04417_),
    .Y(_00293_),
    .A1(net7312),
    .A2(net6652));
 sg13g2_nand2_1 _13297_ (.Y(_04418_),
    .A(net3378),
    .B(net6653));
 sg13g2_o21ai_1 _13298_ (.B1(_04418_),
    .Y(_00294_),
    .A1(net7510),
    .A2(net6653));
 sg13g2_nand2_1 _13299_ (.Y(_04419_),
    .A(net3843),
    .B(net6652));
 sg13g2_o21ai_1 _13300_ (.B1(_04419_),
    .Y(_00295_),
    .A1(net7669),
    .A2(net6653));
 sg13g2_nand3_1 _13301_ (.B(net7264),
    .C(net7078),
    .A(net7384),
    .Y(_04420_));
 sg13g2_nand2_1 _13302_ (.Y(_04421_),
    .A(net3310),
    .B(net6650));
 sg13g2_o21ai_1 _13303_ (.B1(_04421_),
    .Y(_00296_),
    .A1(net7312),
    .A2(net6650));
 sg13g2_nand2_1 _13304_ (.Y(_04422_),
    .A(net3140),
    .B(net6650));
 sg13g2_o21ai_1 _13305_ (.B1(_04422_),
    .Y(_00297_),
    .A1(net7512),
    .A2(net6650));
 sg13g2_nand2_1 _13306_ (.Y(_04423_),
    .A(net3634),
    .B(net6651));
 sg13g2_o21ai_1 _13307_ (.B1(_04423_),
    .Y(_00298_),
    .A1(net7669),
    .A2(net6651));
 sg13g2_nand3_1 _13308_ (.B(net7078),
    .C(net7236),
    .A(net7384),
    .Y(_04424_));
 sg13g2_nand2_1 _13309_ (.Y(_04425_),
    .A(net3194),
    .B(net6648));
 sg13g2_o21ai_1 _13310_ (.B1(_04425_),
    .Y(_00299_),
    .A1(net7312),
    .A2(net6648));
 sg13g2_nand2_1 _13311_ (.Y(_04426_),
    .A(net2456),
    .B(net6648));
 sg13g2_o21ai_1 _13312_ (.B1(_04426_),
    .Y(_00300_),
    .A1(net7512),
    .A2(net6648));
 sg13g2_nand2_1 _13313_ (.Y(_04427_),
    .A(net2507),
    .B(net6649));
 sg13g2_o21ai_1 _13314_ (.B1(_04427_),
    .Y(_00301_),
    .A1(net7669),
    .A2(net6649));
 sg13g2_nand3_1 _13315_ (.B(net7082),
    .C(net7065),
    .A(net7382),
    .Y(_04428_));
 sg13g2_nand2_1 _13316_ (.Y(_04429_),
    .A(net3034),
    .B(net6646));
 sg13g2_o21ai_1 _13317_ (.B1(_04429_),
    .Y(_00302_),
    .A1(net7317),
    .A2(net6646));
 sg13g2_nand2_1 _13318_ (.Y(_04430_),
    .A(net3087),
    .B(net6646));
 sg13g2_o21ai_1 _13319_ (.B1(_04430_),
    .Y(_00303_),
    .A1(net7517),
    .A2(net6646));
 sg13g2_nand2_1 _13320_ (.Y(_04431_),
    .A(net3883),
    .B(net6647));
 sg13g2_o21ai_1 _13321_ (.B1(_04431_),
    .Y(_00304_),
    .A1(net7689),
    .A2(net6647));
 sg13g2_nand3_1 _13322_ (.B(net7104),
    .C(net7082),
    .A(net7382),
    .Y(_04432_));
 sg13g2_nand2_1 _13323_ (.Y(_04433_),
    .A(net2980),
    .B(net6644));
 sg13g2_o21ai_1 _13324_ (.B1(_04433_),
    .Y(_00305_),
    .A1(net7317),
    .A2(net6644));
 sg13g2_nand2_1 _13325_ (.Y(_04434_),
    .A(net3702),
    .B(net6644));
 sg13g2_o21ai_1 _13326_ (.B1(_04434_),
    .Y(_00306_),
    .A1(net7517),
    .A2(net6644));
 sg13g2_nand2_1 _13327_ (.Y(_04435_),
    .A(net2537),
    .B(net6645));
 sg13g2_o21ai_1 _13328_ (.B1(_04435_),
    .Y(_00307_),
    .A1(net7689),
    .A2(net6645));
 sg13g2_nand3_1 _13329_ (.B(net7247),
    .C(net7244),
    .A(net7385),
    .Y(_04436_));
 sg13g2_nand2_1 _13330_ (.Y(_04437_),
    .A(net3342),
    .B(net7010));
 sg13g2_o21ai_1 _13331_ (.B1(_04437_),
    .Y(_00308_),
    .A1(net7335),
    .A2(net7010));
 sg13g2_nand2_1 _13332_ (.Y(_04438_),
    .A(net2546),
    .B(net7011));
 sg13g2_o21ai_1 _13333_ (.B1(_04438_),
    .Y(_00309_),
    .A1(net7530),
    .A2(net7011));
 sg13g2_nand2_1 _13334_ (.Y(_04439_),
    .A(net2775),
    .B(net7011));
 sg13g2_o21ai_1 _13335_ (.B1(_04439_),
    .Y(_00310_),
    .A1(net7691),
    .A2(net7011));
 sg13g2_nand3_1 _13336_ (.B(net7078),
    .C(net7043),
    .A(net7382),
    .Y(_04440_));
 sg13g2_nand2_1 _13337_ (.Y(_04441_),
    .A(net3013),
    .B(net6642));
 sg13g2_o21ai_1 _13338_ (.B1(_04441_),
    .Y(_00311_),
    .A1(net7317),
    .A2(net6642));
 sg13g2_nand2_1 _13339_ (.Y(_04442_),
    .A(net2748),
    .B(net6642));
 sg13g2_o21ai_1 _13340_ (.B1(_04442_),
    .Y(_00312_),
    .A1(net7517),
    .A2(net6642));
 sg13g2_nand2_1 _13341_ (.Y(_04443_),
    .A(net2717),
    .B(net6643));
 sg13g2_o21ai_1 _13342_ (.B1(_04443_),
    .Y(_00313_),
    .A1(net7689),
    .A2(net6643));
 sg13g2_nand3_1 _13343_ (.B(net7382),
    .C(net7079),
    .A(net7407),
    .Y(_04444_));
 sg13g2_nand2_1 _13344_ (.Y(_04445_),
    .A(net2800),
    .B(net6640));
 sg13g2_o21ai_1 _13345_ (.B1(_04445_),
    .Y(_00314_),
    .A1(net7318),
    .A2(net6640));
 sg13g2_nand2_1 _13346_ (.Y(_04446_),
    .A(net3427),
    .B(net6640));
 sg13g2_o21ai_1 _13347_ (.B1(_04446_),
    .Y(_00315_),
    .A1(net7517),
    .A2(net6640));
 sg13g2_nand2_1 _13348_ (.Y(_04447_),
    .A(net3227),
    .B(net6641));
 sg13g2_o21ai_1 _13349_ (.B1(_04447_),
    .Y(_00316_),
    .A1(net7677),
    .A2(net6641));
 sg13g2_nand3_1 _13350_ (.B(net7283),
    .C(net7078),
    .A(net7382),
    .Y(_04448_));
 sg13g2_nand2_1 _13351_ (.Y(_04449_),
    .A(net3854),
    .B(net6638));
 sg13g2_o21ai_1 _13352_ (.B1(_04449_),
    .Y(_00317_),
    .A1(net7318),
    .A2(net6638));
 sg13g2_nand2_1 _13353_ (.Y(_04450_),
    .A(net2855),
    .B(net6638));
 sg13g2_o21ai_1 _13354_ (.B1(_04450_),
    .Y(_00318_),
    .A1(net7518),
    .A2(net6638));
 sg13g2_nand2_1 _13355_ (.Y(_04451_),
    .A(net3706),
    .B(net6639));
 sg13g2_o21ai_1 _13356_ (.B1(_04451_),
    .Y(_00319_),
    .A1(net7677),
    .A2(net6639));
 sg13g2_nand3_1 _13357_ (.B(net7361),
    .C(net7078),
    .A(net7382),
    .Y(_04452_));
 sg13g2_nand2_1 _13358_ (.Y(_04453_),
    .A(net3302),
    .B(net6636));
 sg13g2_o21ai_1 _13359_ (.B1(_04453_),
    .Y(_00320_),
    .A1(net7318),
    .A2(net6636));
 sg13g2_nand2_1 _13360_ (.Y(_04454_),
    .A(net3599),
    .B(net6636));
 sg13g2_o21ai_1 _13361_ (.B1(_04454_),
    .Y(_00321_),
    .A1(net7517),
    .A2(net6636));
 sg13g2_nand2_1 _13362_ (.Y(_04455_),
    .A(net3790),
    .B(net6637));
 sg13g2_o21ai_1 _13363_ (.B1(_04455_),
    .Y(_00322_),
    .A1(net7677),
    .A2(net6637));
 sg13g2_nand3_1 _13364_ (.B(net7280),
    .C(net7078),
    .A(net7382),
    .Y(_04456_));
 sg13g2_nand2_1 _13365_ (.Y(_04457_),
    .A(net2667),
    .B(net6634));
 sg13g2_o21ai_1 _13366_ (.B1(_04457_),
    .Y(_00323_),
    .A1(net7318),
    .A2(net6634));
 sg13g2_nand2_1 _13367_ (.Y(_04458_),
    .A(net2602),
    .B(net6634));
 sg13g2_o21ai_1 _13368_ (.B1(_04458_),
    .Y(_00324_),
    .A1(net7517),
    .A2(net6634));
 sg13g2_nand2_1 _13369_ (.Y(_04459_),
    .A(net3263),
    .B(net6635));
 sg13g2_o21ai_1 _13370_ (.B1(_04459_),
    .Y(_00325_),
    .A1(net7677),
    .A2(net6635));
 sg13g2_nand3_1 _13371_ (.B(net7285),
    .C(net7078),
    .A(net7383),
    .Y(_04460_));
 sg13g2_nand2_1 _13372_ (.Y(_04461_),
    .A(net3133),
    .B(net6632));
 sg13g2_o21ai_1 _13373_ (.B1(_04461_),
    .Y(_00326_),
    .A1(net7317),
    .A2(net6632));
 sg13g2_nand2_1 _13374_ (.Y(_04462_),
    .A(net3548),
    .B(net6632));
 sg13g2_o21ai_1 _13375_ (.B1(_04462_),
    .Y(_00327_),
    .A1(net7518),
    .A2(net6632));
 sg13g2_nand2_1 _13376_ (.Y(_04463_),
    .A(net2920),
    .B(net6633));
 sg13g2_o21ai_1 _13377_ (.B1(_04463_),
    .Y(_00328_),
    .A1(net7677),
    .A2(net6633));
 sg13g2_nor3_1 _13378_ (.A(net7372),
    .B(net7272),
    .C(_04154_),
    .Y(_04464_));
 sg13g2_nor2_1 _13379_ (.A(net4728),
    .B(net7008),
    .Y(_04465_));
 sg13g2_a21oi_1 _13380_ (.A1(net7317),
    .A2(net7008),
    .Y(_00329_),
    .B1(_04465_));
 sg13g2_nor2_1 _13381_ (.A(net3802),
    .B(net7008),
    .Y(_04466_));
 sg13g2_a21oi_1 _13382_ (.A1(net7517),
    .A2(net7008),
    .Y(_00330_),
    .B1(_04466_));
 sg13g2_nor2_1 _13383_ (.A(net4114),
    .B(net7009),
    .Y(_04467_));
 sg13g2_a21oi_1 _13384_ (.A1(net7677),
    .A2(net7009),
    .Y(_00331_),
    .B1(_04467_));
 sg13g2_nor3_1 _13385_ (.A(net7372),
    .B(net7276),
    .C(_04154_),
    .Y(_04468_));
 sg13g2_nor2_1 _13386_ (.A(net4203),
    .B(net7006),
    .Y(_04469_));
 sg13g2_a21oi_1 _13387_ (.A1(net7317),
    .A2(net7006),
    .Y(_00332_),
    .B1(_04469_));
 sg13g2_nor2_1 _13388_ (.A(net4307),
    .B(net7006),
    .Y(_04470_));
 sg13g2_a21oi_1 _13389_ (.A1(net7518),
    .A2(net7006),
    .Y(_00333_),
    .B1(_04470_));
 sg13g2_nor2_1 _13390_ (.A(net4120),
    .B(net7007),
    .Y(_04471_));
 sg13g2_a21oi_1 _13391_ (.A1(net7677),
    .A2(net7007),
    .Y(_00334_),
    .B1(_04471_));
 sg13g2_nor3_1 _13392_ (.A(net7372),
    .B(_04154_),
    .C(net7246),
    .Y(_04472_));
 sg13g2_nor2_1 _13393_ (.A(net3542),
    .B(net7004),
    .Y(_04473_));
 sg13g2_a21oi_1 _13394_ (.A1(net7317),
    .A2(net7004),
    .Y(_00335_),
    .B1(_04473_));
 sg13g2_nor2_1 _13395_ (.A(net4329),
    .B(net7004),
    .Y(_04474_));
 sg13g2_a21oi_1 _13396_ (.A1(net7518),
    .A2(net7004),
    .Y(_00336_),
    .B1(_04474_));
 sg13g2_nor2_1 _13397_ (.A(net4598),
    .B(net7005),
    .Y(_04475_));
 sg13g2_a21oi_1 _13398_ (.A1(net7677),
    .A2(net7005),
    .Y(_00337_),
    .B1(_04475_));
 sg13g2_nor3_2 _13399_ (.A(net7402),
    .B(net7370),
    .C(net7269),
    .Y(_04476_));
 sg13g2_nor2_1 _13400_ (.A(net4833),
    .B(net7002),
    .Y(_04477_));
 sg13g2_a21oi_1 _13401_ (.A1(net7322),
    .A2(net7003),
    .Y(_00338_),
    .B1(_04477_));
 sg13g2_nor2_1 _13402_ (.A(net4030),
    .B(net7002),
    .Y(_04478_));
 sg13g2_a21oi_1 _13403_ (.A1(net7515),
    .A2(net7002),
    .Y(_00339_),
    .B1(_04478_));
 sg13g2_nor2_1 _13404_ (.A(net4473),
    .B(net7003),
    .Y(_04479_));
 sg13g2_a21oi_1 _13405_ (.A1(net7673),
    .A2(net7003),
    .Y(_00340_),
    .B1(_04479_));
 sg13g2_nand3_1 _13406_ (.B(net7255),
    .C(net7237),
    .A(net7377),
    .Y(_04480_));
 sg13g2_nand2_1 _13407_ (.Y(_04481_),
    .A(net2561),
    .B(net7000));
 sg13g2_o21ai_1 _13408_ (.B1(_04481_),
    .Y(_00341_),
    .A1(net7305),
    .A2(net7000));
 sg13g2_nand2_1 _13409_ (.Y(_04482_),
    .A(net2782),
    .B(net7000));
 sg13g2_o21ai_1 _13410_ (.B1(_04482_),
    .Y(_00342_),
    .A1(net7503),
    .A2(net7000));
 sg13g2_nand2_1 _13411_ (.Y(_04483_),
    .A(net2490),
    .B(net7001));
 sg13g2_o21ai_1 _13412_ (.B1(_04483_),
    .Y(_00343_),
    .A1(net7661),
    .A2(net7001));
 sg13g2_nand3_1 _13413_ (.B(net7264),
    .C(net7254),
    .A(net7377),
    .Y(_04484_));
 sg13g2_nand2_1 _13414_ (.Y(_04485_),
    .A(net2840),
    .B(net6998));
 sg13g2_o21ai_1 _13415_ (.B1(_04485_),
    .Y(_00344_),
    .A1(net7303),
    .A2(net6998));
 sg13g2_nand2_1 _13416_ (.Y(_04486_),
    .A(net3313),
    .B(net6998));
 sg13g2_o21ai_1 _13417_ (.B1(_04486_),
    .Y(_00345_),
    .A1(net7501),
    .A2(net6998));
 sg13g2_nand2_1 _13418_ (.Y(_04487_),
    .A(net2506),
    .B(net6999));
 sg13g2_o21ai_1 _13419_ (.B1(_04487_),
    .Y(_00346_),
    .A1(net7672),
    .A2(net6999));
 sg13g2_nand3_1 _13420_ (.B(net7254),
    .C(net7236),
    .A(net7378),
    .Y(_04488_));
 sg13g2_nand2_1 _13421_ (.Y(_04489_),
    .A(net3070),
    .B(net6996));
 sg13g2_o21ai_1 _13422_ (.B1(_04489_),
    .Y(_00347_),
    .A1(net7303),
    .A2(net6996));
 sg13g2_nand2_1 _13423_ (.Y(_04490_),
    .A(net2523),
    .B(net6996));
 sg13g2_o21ai_1 _13424_ (.B1(_04490_),
    .Y(_00348_),
    .A1(net7501),
    .A2(net6996));
 sg13g2_nand2_1 _13425_ (.Y(_04491_),
    .A(net3184),
    .B(net6997));
 sg13g2_o21ai_1 _13426_ (.B1(_04491_),
    .Y(_00349_),
    .A1(net7661),
    .A2(net6997));
 sg13g2_nand3_1 _13427_ (.B(net7256),
    .C(net7065),
    .A(net7378),
    .Y(_04492_));
 sg13g2_nand2_1 _13428_ (.Y(_04493_),
    .A(net2635),
    .B(net6630));
 sg13g2_o21ai_1 _13429_ (.B1(_04493_),
    .Y(_00350_),
    .A1(net7315),
    .A2(net6630));
 sg13g2_nand2_1 _13430_ (.Y(_04494_),
    .A(net3031),
    .B(net6631));
 sg13g2_o21ai_1 _13431_ (.B1(_04494_),
    .Y(_00351_),
    .A1(net7514),
    .A2(net6631));
 sg13g2_nand2_1 _13432_ (.Y(_04495_),
    .A(net2607),
    .B(net6630));
 sg13g2_o21ai_1 _13433_ (.B1(_04495_),
    .Y(_00352_),
    .A1(net7671),
    .A2(net6630));
 sg13g2_nand3_1 _13434_ (.B(net7104),
    .C(net7256),
    .A(net7378),
    .Y(_04496_));
 sg13g2_nand2_1 _13435_ (.Y(_04497_),
    .A(net2608),
    .B(net6628));
 sg13g2_o21ai_1 _13436_ (.B1(_04497_),
    .Y(_00353_),
    .A1(net7315),
    .A2(net6628));
 sg13g2_nand2_1 _13437_ (.Y(_04498_),
    .A(net2868),
    .B(net6629));
 sg13g2_o21ai_1 _13438_ (.B1(_04498_),
    .Y(_00354_),
    .A1(net7514),
    .A2(net6629));
 sg13g2_nand2_1 _13439_ (.Y(_04499_),
    .A(net3446),
    .B(net6628));
 sg13g2_o21ai_1 _13440_ (.B1(_04499_),
    .Y(_00355_),
    .A1(net7672),
    .A2(net6628));
 sg13g2_nand3_1 _13441_ (.B(net7085),
    .C(net7256),
    .A(net7378),
    .Y(_04500_));
 sg13g2_nand2_1 _13442_ (.Y(_04501_),
    .A(net4036),
    .B(net6627));
 sg13g2_o21ai_1 _13443_ (.B1(_04501_),
    .Y(_00356_),
    .A1(net7315),
    .A2(net6627));
 sg13g2_nand2_1 _13444_ (.Y(_04502_),
    .A(net3119),
    .B(net6626));
 sg13g2_o21ai_1 _13445_ (.B1(_04502_),
    .Y(_00357_),
    .A1(net7514),
    .A2(net6626));
 sg13g2_nand2_1 _13446_ (.Y(_04503_),
    .A(net4144),
    .B(net6626));
 sg13g2_o21ai_1 _13447_ (.B1(_04503_),
    .Y(_00358_),
    .A1(net7672),
    .A2(net6626));
 sg13g2_nand3_1 _13448_ (.B(net7256),
    .C(net7043),
    .A(net7378),
    .Y(_04504_));
 sg13g2_nand2_1 _13449_ (.Y(_04505_),
    .A(net4287),
    .B(net6625));
 sg13g2_o21ai_1 _13450_ (.B1(_04505_),
    .Y(_00359_),
    .A1(net7315),
    .A2(net6625));
 sg13g2_nand2_1 _13451_ (.Y(_04506_),
    .A(net2726),
    .B(net6624));
 sg13g2_o21ai_1 _13452_ (.B1(_04506_),
    .Y(_00360_),
    .A1(net7514),
    .A2(net6624));
 sg13g2_nand2_1 _13453_ (.Y(_04507_),
    .A(net4035),
    .B(net6624));
 sg13g2_o21ai_1 _13454_ (.B1(_04507_),
    .Y(_00361_),
    .A1(net7672),
    .A2(net6624));
 sg13g2_nand3_1 _13455_ (.B(net7377),
    .C(net7255),
    .A(net7406),
    .Y(_04508_));
 sg13g2_nand2_1 _13456_ (.Y(_04509_),
    .A(net3063),
    .B(net6994));
 sg13g2_o21ai_1 _13457_ (.B1(_04509_),
    .Y(_00362_),
    .A1(net7303),
    .A2(net6994));
 sg13g2_nand2_1 _13458_ (.Y(_04510_),
    .A(net4160),
    .B(net6994));
 sg13g2_o21ai_1 _13459_ (.B1(_04510_),
    .Y(_00363_),
    .A1(net7501),
    .A2(net6994));
 sg13g2_nand2_1 _13460_ (.Y(_04511_),
    .A(net2441),
    .B(net6995));
 sg13g2_o21ai_1 _13461_ (.B1(_04511_),
    .Y(_00364_),
    .A1(net7671),
    .A2(net6995));
 sg13g2_nand3_1 _13462_ (.B(net7281),
    .C(net7256),
    .A(net7377),
    .Y(_04512_));
 sg13g2_nand2_1 _13463_ (.Y(_04513_),
    .A(net2742),
    .B(net6992));
 sg13g2_o21ai_1 _13464_ (.B1(_04513_),
    .Y(_00365_),
    .A1(net7302),
    .A2(net6992));
 sg13g2_nand2_1 _13465_ (.Y(_04514_),
    .A(net2941),
    .B(net6992));
 sg13g2_o21ai_1 _13466_ (.B1(_04514_),
    .Y(_00366_),
    .A1(net7503),
    .A2(net6992));
 sg13g2_nand2_1 _13467_ (.Y(_04515_),
    .A(net2651),
    .B(net6993));
 sg13g2_o21ai_1 _13468_ (.B1(_04515_),
    .Y(_00367_),
    .A1(net7670),
    .A2(net6993));
 sg13g2_nand3_1 _13469_ (.B(_04129_),
    .C(net7237),
    .A(net7379),
    .Y(_04516_));
 sg13g2_nand2_1 _13470_ (.Y(_04517_),
    .A(net3778),
    .B(net6990));
 sg13g2_o21ai_1 _13471_ (.B1(_04517_),
    .Y(_00368_),
    .A1(net7322),
    .A2(net6990));
 sg13g2_nand2_1 _13472_ (.Y(_04518_),
    .A(net2901),
    .B(net6990));
 sg13g2_o21ai_1 _13473_ (.B1(_04518_),
    .Y(_00369_),
    .A1(net7515),
    .A2(net6990));
 sg13g2_nand2_1 _13474_ (.Y(_04519_),
    .A(net3533),
    .B(net6990));
 sg13g2_o21ai_1 _13475_ (.B1(_04519_),
    .Y(_00370_),
    .A1(net7673),
    .A2(net6990));
 sg13g2_nand3_1 _13476_ (.B(net7280),
    .C(net7256),
    .A(net7377),
    .Y(_04520_));
 sg13g2_nand2_1 _13477_ (.Y(_04521_),
    .A(net3682),
    .B(net6988));
 sg13g2_o21ai_1 _13478_ (.B1(_04521_),
    .Y(_00371_),
    .A1(net7315),
    .A2(net6988));
 sg13g2_nand2_1 _13479_ (.Y(_04522_),
    .A(net4115),
    .B(net6988));
 sg13g2_o21ai_1 _13480_ (.B1(_04522_),
    .Y(_00372_),
    .A1(net7514),
    .A2(net6988));
 sg13g2_nand2_1 _13481_ (.Y(_04523_),
    .A(net3435),
    .B(net6989));
 sg13g2_o21ai_1 _13482_ (.B1(_04523_),
    .Y(_00373_),
    .A1(net7671),
    .A2(net6989));
 sg13g2_nand3_1 _13483_ (.B(net7285),
    .C(net7254),
    .A(net7377),
    .Y(_04524_));
 sg13g2_nand2_1 _13484_ (.Y(_04525_),
    .A(net3518),
    .B(net6986));
 sg13g2_o21ai_1 _13485_ (.B1(_04525_),
    .Y(_00374_),
    .A1(net7303),
    .A2(net6986));
 sg13g2_nand2_1 _13486_ (.Y(_04526_),
    .A(net3827),
    .B(net6986));
 sg13g2_o21ai_1 _13487_ (.B1(_04526_),
    .Y(_00375_),
    .A1(net7501),
    .A2(net6986));
 sg13g2_nand2_1 _13488_ (.Y(_04527_),
    .A(net3139),
    .B(net6987));
 sg13g2_o21ai_1 _13489_ (.B1(_04527_),
    .Y(_00376_),
    .A1(net7671),
    .A2(net6987));
 sg13g2_nor3_1 _13490_ (.A(net7370),
    .B(net7271),
    .C(_04165_),
    .Y(_04528_));
 sg13g2_nor2_1 _13491_ (.A(net4709),
    .B(net6984),
    .Y(_04529_));
 sg13g2_a21oi_1 _13492_ (.A1(net7303),
    .A2(net6984),
    .Y(_00377_),
    .B1(_04529_));
 sg13g2_nor2_1 _13493_ (.A(net3820),
    .B(net6984),
    .Y(_04530_));
 sg13g2_a21oi_1 _13494_ (.A1(net7501),
    .A2(net6984),
    .Y(_00378_),
    .B1(_04530_));
 sg13g2_nor2_1 _13495_ (.A(net4556),
    .B(net6985),
    .Y(_04531_));
 sg13g2_a21oi_1 _13496_ (.A1(net7671),
    .A2(net6985),
    .Y(_00379_),
    .B1(_04531_));
 sg13g2_nor3_1 _13497_ (.A(net7370),
    .B(net7275),
    .C(_04165_),
    .Y(_04532_));
 sg13g2_nor2_1 _13498_ (.A(net4451),
    .B(net6982),
    .Y(_04533_));
 sg13g2_a21oi_1 _13499_ (.A1(net7303),
    .A2(net6982),
    .Y(_00380_),
    .B1(_04533_));
 sg13g2_nor2_1 _13500_ (.A(net4372),
    .B(net6982),
    .Y(_04534_));
 sg13g2_a21oi_1 _13501_ (.A1(net7501),
    .A2(net6982),
    .Y(_00381_),
    .B1(_04534_));
 sg13g2_nor2_1 _13502_ (.A(net4305),
    .B(net6983),
    .Y(_04535_));
 sg13g2_a21oi_1 _13503_ (.A1(net7671),
    .A2(net6983),
    .Y(_00382_),
    .B1(_04535_));
 sg13g2_nor3_1 _13504_ (.A(net7370),
    .B(_04165_),
    .C(net7245),
    .Y(_04536_));
 sg13g2_nor2_1 _13505_ (.A(net4646),
    .B(net6980),
    .Y(_04537_));
 sg13g2_a21oi_1 _13506_ (.A1(net7303),
    .A2(net6980),
    .Y(_00383_),
    .B1(_04537_));
 sg13g2_nor2_1 _13507_ (.A(net4311),
    .B(net6980),
    .Y(_04538_));
 sg13g2_a21oi_1 _13508_ (.A1(net7501),
    .A2(net6980),
    .Y(_00384_),
    .B1(_04538_));
 sg13g2_nor2_1 _13509_ (.A(net4328),
    .B(net6981),
    .Y(_04539_));
 sg13g2_a21oi_1 _13510_ (.A1(net7671),
    .A2(net6981),
    .Y(_00385_),
    .B1(_04539_));
 sg13g2_nor3_1 _13511_ (.A(net7402),
    .B(net7366),
    .C(net7251),
    .Y(_04540_));
 sg13g2_nor2_1 _13512_ (.A(net4238),
    .B(net6978),
    .Y(_04541_));
 sg13g2_a21oi_1 _13513_ (.A1(net7299),
    .A2(net6978),
    .Y(_00386_),
    .B1(_04541_));
 sg13g2_nor2_1 _13514_ (.A(net4486),
    .B(net6979),
    .Y(_04542_));
 sg13g2_a21oi_1 _13515_ (.A1(net7497),
    .A2(net6979),
    .Y(_00387_),
    .B1(_04542_));
 sg13g2_nor2_1 _13516_ (.A(net3476),
    .B(net6978),
    .Y(_04543_));
 sg13g2_a21oi_1 _13517_ (.A1(net7657),
    .A2(net6978),
    .Y(_00388_),
    .B1(_04543_));
 sg13g2_nor3_1 _13518_ (.A(net7366),
    .B(net7251),
    .C(_04217_),
    .Y(_04544_));
 sg13g2_nor2_1 _13519_ (.A(net4606),
    .B(net6977),
    .Y(_04545_));
 sg13g2_a21oi_1 _13520_ (.A1(net7298),
    .A2(net6977),
    .Y(_00389_),
    .B1(_04545_));
 sg13g2_nor2_1 _13521_ (.A(net4519),
    .B(net6976),
    .Y(_04546_));
 sg13g2_a21oi_1 _13522_ (.A1(net7497),
    .A2(net6976),
    .Y(_00390_),
    .B1(_04546_));
 sg13g2_nor2_1 _13523_ (.A(net4063),
    .B(net6976),
    .Y(_04547_));
 sg13g2_a21oi_1 _13524_ (.A1(net7657),
    .A2(net6976),
    .Y(_00391_),
    .B1(_04547_));
 sg13g2_nor3_1 _13525_ (.A(net7366),
    .B(_04141_),
    .C(net7251),
    .Y(_04548_));
 sg13g2_nor2_1 _13526_ (.A(net4805),
    .B(net6975),
    .Y(_04549_));
 sg13g2_a21oi_1 _13527_ (.A1(net7298),
    .A2(net6975),
    .Y(_00392_),
    .B1(_04549_));
 sg13g2_nor2_1 _13528_ (.A(net4146),
    .B(net6974),
    .Y(_04550_));
 sg13g2_a21oi_1 _13529_ (.A1(net7497),
    .A2(net6974),
    .Y(_00393_),
    .B1(_04550_));
 sg13g2_nor2_1 _13530_ (.A(net4784),
    .B(net6974),
    .Y(_04551_));
 sg13g2_a21oi_1 _13531_ (.A1(net7657),
    .A2(net6974),
    .Y(_00394_),
    .B1(_04551_));
 sg13g2_nor3_1 _13532_ (.A(net7366),
    .B(net7251),
    .C(_04235_),
    .Y(_04552_));
 sg13g2_nor2_1 _13533_ (.A(net4695),
    .B(net6973),
    .Y(_04553_));
 sg13g2_a21oi_1 _13534_ (.A1(net7298),
    .A2(net6973),
    .Y(_00395_),
    .B1(_04553_));
 sg13g2_nor2_1 _13535_ (.A(net3436),
    .B(net6972),
    .Y(_04554_));
 sg13g2_a21oi_1 _13536_ (.A1(net7497),
    .A2(net6972),
    .Y(_00396_),
    .B1(_04554_));
 sg13g2_nor2_1 _13537_ (.A(net4385),
    .B(net6972),
    .Y(_04555_));
 sg13g2_a21oi_1 _13538_ (.A1(net7657),
    .A2(net6972),
    .Y(_00397_),
    .B1(_04555_));
 sg13g2_nand3_1 _13539_ (.B(_04129_),
    .C(net7264),
    .A(net7379),
    .Y(_04556_));
 sg13g2_nand2_1 _13540_ (.Y(_04557_),
    .A(net3460),
    .B(net6971));
 sg13g2_o21ai_1 _13541_ (.B1(_04557_),
    .Y(_00398_),
    .A1(net7315),
    .A2(net6971));
 sg13g2_nand2_1 _13542_ (.Y(_04558_),
    .A(net2559),
    .B(net6970));
 sg13g2_o21ai_1 _13543_ (.B1(_04558_),
    .Y(_00399_),
    .A1(net7515),
    .A2(net6970));
 sg13g2_nand2_1 _13544_ (.Y(_04559_),
    .A(net3247),
    .B(net6971));
 sg13g2_o21ai_1 _13545_ (.B1(_04559_),
    .Y(_00400_),
    .A1(net7673),
    .A2(net6971));
 sg13g2_nor3_2 _13546_ (.A(net7367),
    .B(_04101_),
    .C(net7252),
    .Y(_04560_));
 sg13g2_nor2_1 _13547_ (.A(net4286),
    .B(net6969),
    .Y(_04561_));
 sg13g2_a21oi_1 _13548_ (.A1(net7304),
    .A2(net6969),
    .Y(_00401_),
    .B1(_04561_));
 sg13g2_nor2_1 _13549_ (.A(net4249),
    .B(net6969),
    .Y(_04562_));
 sg13g2_a21oi_1 _13550_ (.A1(net7502),
    .A2(net6969),
    .Y(_00402_),
    .B1(_04562_));
 sg13g2_nor2_1 _13551_ (.A(net4648),
    .B(net6968),
    .Y(_04563_));
 sg13g2_a21oi_1 _13552_ (.A1(net7658),
    .A2(net6968),
    .Y(_00403_),
    .B1(_04563_));
 sg13g2_nor3_2 _13553_ (.A(net7367),
    .B(_04152_),
    .C(net7252),
    .Y(_04564_));
 sg13g2_nor2_1 _13554_ (.A(net4484),
    .B(net6967),
    .Y(_04565_));
 sg13g2_a21oi_1 _13555_ (.A1(net7304),
    .A2(net6967),
    .Y(_00404_),
    .B1(_04565_));
 sg13g2_nor2_1 _13556_ (.A(net4616),
    .B(net6967),
    .Y(_04566_));
 sg13g2_a21oi_1 _13557_ (.A1(net7502),
    .A2(net6967),
    .Y(_00405_),
    .B1(_04566_));
 sg13g2_nor2_1 _13558_ (.A(net4456),
    .B(net6966),
    .Y(_04567_));
 sg13g2_a21oi_1 _13559_ (.A1(net7658),
    .A2(net6966),
    .Y(_00406_),
    .B1(_04567_));
 sg13g2_nor3_1 _13560_ (.A(net7367),
    .B(net7252),
    .C(net7234),
    .Y(_04568_));
 sg13g2_nor2_1 _13561_ (.A(net3893),
    .B(net6965),
    .Y(_04569_));
 sg13g2_a21oi_1 _13562_ (.A1(net7304),
    .A2(net6965),
    .Y(_00407_),
    .B1(_04569_));
 sg13g2_nor2_1 _13563_ (.A(net3863),
    .B(net6964),
    .Y(_04570_));
 sg13g2_a21oi_1 _13564_ (.A1(net7498),
    .A2(net6965),
    .Y(_00408_),
    .B1(_04570_));
 sg13g2_nor2_1 _13565_ (.A(net4442),
    .B(net6965),
    .Y(_04571_));
 sg13g2_a21oi_1 _13566_ (.A1(net7658),
    .A2(net6964),
    .Y(_00409_),
    .B1(_04571_));
 sg13g2_nor3_1 _13567_ (.A(_04040_),
    .B(net7368),
    .C(net7252),
    .Y(_04572_));
 sg13g2_nor2_1 _13568_ (.A(net4554),
    .B(net6622),
    .Y(_04573_));
 sg13g2_a21oi_1 _13569_ (.A1(net7299),
    .A2(net6622),
    .Y(_00410_),
    .B1(_04573_));
 sg13g2_nor2_1 _13570_ (.A(net4113),
    .B(net6622),
    .Y(_04574_));
 sg13g2_a21oi_1 _13571_ (.A1(net7498),
    .A2(net6622),
    .Y(_00411_),
    .B1(_04574_));
 sg13g2_nor2_1 _13572_ (.A(net4025),
    .B(net6623),
    .Y(_04575_));
 sg13g2_a21oi_1 _13573_ (.A1(net7658),
    .A2(net6623),
    .Y(_00412_),
    .B1(_04575_));
 sg13g2_nand3_1 _13574_ (.B(net7391),
    .C(_04092_),
    .A(net7114),
    .Y(_04576_));
 sg13g2_nand2_1 _13575_ (.Y(_04577_),
    .A(net3502),
    .B(net6620));
 sg13g2_o21ai_1 _13576_ (.B1(_04577_),
    .Y(_00413_),
    .A1(net7346),
    .A2(net6620));
 sg13g2_nand2_1 _13577_ (.Y(_04578_),
    .A(net2875),
    .B(net6621));
 sg13g2_o21ai_1 _13578_ (.B1(_04578_),
    .Y(_00414_),
    .A1(net7544),
    .A2(net6621));
 sg13g2_nand2_1 _13579_ (.Y(_04579_),
    .A(net3661),
    .B(net6620));
 sg13g2_o21ai_1 _13580_ (.B1(_04579_),
    .Y(_00415_),
    .A1(net7703),
    .A2(net6620));
 sg13g2_nor3_2 _13581_ (.A(net7370),
    .B(net7269),
    .C(_04235_),
    .Y(_04580_));
 sg13g2_nor2_1 _13582_ (.A(net4803),
    .B(net6963),
    .Y(_04581_));
 sg13g2_a21oi_1 _13583_ (.A1(net7315),
    .A2(net6963),
    .Y(_00416_),
    .B1(_04581_));
 sg13g2_nor2_1 _13584_ (.A(net3982),
    .B(net6962),
    .Y(_04582_));
 sg13g2_a21oi_1 _13585_ (.A1(net7515),
    .A2(net6962),
    .Y(_00417_),
    .B1(_04582_));
 sg13g2_nor2_1 _13586_ (.A(net4642),
    .B(net6963),
    .Y(_04583_));
 sg13g2_a21oi_1 _13587_ (.A1(net7673),
    .A2(net6963),
    .Y(_00418_),
    .B1(_04583_));
 sg13g2_nand3_1 _13588_ (.B(net7392),
    .C(net7286),
    .A(net7115),
    .Y(_04584_));
 sg13g2_nand2_1 _13589_ (.Y(_04585_),
    .A(net3403),
    .B(net6618));
 sg13g2_o21ai_1 _13590_ (.B1(_04585_),
    .Y(_00419_),
    .A1(net7346),
    .A2(net6618));
 sg13g2_nand2_1 _13591_ (.Y(_04586_),
    .A(net3720),
    .B(net6618));
 sg13g2_o21ai_1 _13592_ (.B1(_04586_),
    .Y(_00420_),
    .A1(net7546),
    .A2(net6618));
 sg13g2_nand2_1 _13593_ (.Y(_04587_),
    .A(net4179),
    .B(net6619));
 sg13g2_o21ai_1 _13594_ (.B1(_04587_),
    .Y(_00421_),
    .A1(net7707),
    .A2(net6619));
 sg13g2_nand3_1 _13595_ (.B(net7393),
    .C(net7274),
    .A(net7115),
    .Y(_04588_));
 sg13g2_nand2_1 _13596_ (.Y(_04589_),
    .A(net3246),
    .B(net6616));
 sg13g2_o21ai_1 _13597_ (.B1(_04589_),
    .Y(_00422_),
    .A1(net7346),
    .A2(net6616));
 sg13g2_nand2_1 _13598_ (.Y(_04590_),
    .A(net4104),
    .B(net6616));
 sg13g2_o21ai_1 _13599_ (.B1(_04590_),
    .Y(_00423_),
    .A1(net7546),
    .A2(net6616));
 sg13g2_nand2_1 _13600_ (.Y(_04591_),
    .A(net2729),
    .B(net6617));
 sg13g2_o21ai_1 _13601_ (.B1(_04591_),
    .Y(_00424_),
    .A1(net7707),
    .A2(net6617));
 sg13g2_nor3_2 _13602_ (.A(net7366),
    .B(net7251),
    .C(net7245),
    .Y(_04592_));
 sg13g2_nor2_1 _13603_ (.A(net4117),
    .B(net6960),
    .Y(_04593_));
 sg13g2_a21oi_1 _13604_ (.A1(net7298),
    .A2(net6960),
    .Y(_00425_),
    .B1(_04593_));
 sg13g2_nor2_1 _13605_ (.A(net3864),
    .B(net6960),
    .Y(_04594_));
 sg13g2_a21oi_1 _13606_ (.A1(net7497),
    .A2(net6960),
    .Y(_00426_),
    .B1(_04594_));
 sg13g2_nor2_1 _13607_ (.A(net4277),
    .B(net6961),
    .Y(_04595_));
 sg13g2_a21oi_1 _13608_ (.A1(net7657),
    .A2(net6961),
    .Y(_00427_),
    .B1(_04595_));
 sg13g2_nand3_1 _13609_ (.B(net7393),
    .C(net7278),
    .A(net7115),
    .Y(_04596_));
 sg13g2_nand2_1 _13610_ (.Y(_04597_),
    .A(net2739),
    .B(net6614));
 sg13g2_o21ai_1 _13611_ (.B1(_04597_),
    .Y(_00428_),
    .A1(net7346),
    .A2(net6614));
 sg13g2_nand2_1 _13612_ (.Y(_04598_),
    .A(net3796),
    .B(net6614));
 sg13g2_o21ai_1 _13613_ (.B1(_04598_),
    .Y(_00429_),
    .A1(net7546),
    .A2(net6614));
 sg13g2_nand2_1 _13614_ (.Y(_04599_),
    .A(net3572),
    .B(net6615));
 sg13g2_o21ai_1 _13615_ (.B1(_04599_),
    .Y(_00430_),
    .A1(net7707),
    .A2(net6615));
 sg13g2_nand3_1 _13616_ (.B(net7393),
    .C(net7248),
    .A(net7115),
    .Y(_04600_));
 sg13g2_nand2_1 _13617_ (.Y(_04601_),
    .A(net3389),
    .B(net6612));
 sg13g2_o21ai_1 _13618_ (.B1(_04601_),
    .Y(_00431_),
    .A1(net7346),
    .A2(net6612));
 sg13g2_nand2_1 _13619_ (.Y(_04602_),
    .A(net3348),
    .B(net6612));
 sg13g2_o21ai_1 _13620_ (.B1(_04602_),
    .Y(_00432_),
    .A1(net7546),
    .A2(net6612));
 sg13g2_nand2_1 _13621_ (.Y(_04603_),
    .A(net4069),
    .B(net6613));
 sg13g2_o21ai_1 _13622_ (.B1(_04603_),
    .Y(_00433_),
    .A1(net7707),
    .A2(net6613));
 sg13g2_nor2_2 _13623_ (.A(_04056_),
    .B(net7374),
    .Y(_04604_));
 sg13g2_nor2_1 _13624_ (.A(net4551),
    .B(net6610),
    .Y(_04605_));
 sg13g2_a21oi_1 _13625_ (.A1(net7342),
    .A2(net6610),
    .Y(_00434_),
    .B1(_04605_));
 sg13g2_nor2_1 _13626_ (.A(net4638),
    .B(net6611),
    .Y(_04606_));
 sg13g2_a21oi_1 _13627_ (.A1(net7540),
    .A2(net6611),
    .Y(_00435_),
    .B1(_04606_));
 sg13g2_nor2_1 _13628_ (.A(net4467),
    .B(net6610),
    .Y(_04607_));
 sg13g2_a21oi_1 _13629_ (.A1(net7700),
    .A2(net6610),
    .Y(_00436_),
    .B1(_04607_));
 sg13g2_nand3_1 _13630_ (.B(net7390),
    .C(net7101),
    .A(net7405),
    .Y(_04608_));
 sg13g2_nand2_1 _13631_ (.Y(_04609_),
    .A(net2723),
    .B(net6609));
 sg13g2_o21ai_1 _13632_ (.B1(_04609_),
    .Y(_00437_),
    .A1(net7341),
    .A2(net6608));
 sg13g2_nand2_1 _13633_ (.Y(_04610_),
    .A(net3122),
    .B(net6608));
 sg13g2_o21ai_1 _13634_ (.B1(_04610_),
    .Y(_00438_),
    .A1(net7539),
    .A2(net6608));
 sg13g2_nand2_1 _13635_ (.Y(_04611_),
    .A(net4234),
    .B(net6608));
 sg13g2_o21ai_1 _13636_ (.B1(_04611_),
    .Y(_00439_),
    .A1(net7701),
    .A2(net6609));
 sg13g2_nand3_1 _13637_ (.B(net7099),
    .C(net7239),
    .A(net7390),
    .Y(_04612_));
 sg13g2_nand2_1 _13638_ (.Y(_04613_),
    .A(net2960),
    .B(net6607));
 sg13g2_o21ai_1 _13639_ (.B1(_04613_),
    .Y(_00440_),
    .A1(net7341),
    .A2(net6606));
 sg13g2_nand2_1 _13640_ (.Y(_04614_),
    .A(net4640),
    .B(net6606));
 sg13g2_o21ai_1 _13641_ (.B1(_04614_),
    .Y(_00441_),
    .A1(net7539),
    .A2(net6606));
 sg13g2_nand2_1 _13642_ (.Y(_04615_),
    .A(net2735),
    .B(net6606));
 sg13g2_o21ai_1 _13643_ (.B1(_04615_),
    .Y(_00442_),
    .A1(net7700),
    .A2(net6607));
 sg13g2_nand3_1 _13644_ (.B(net7392),
    .C(net7239),
    .A(net7114),
    .Y(_04616_));
 sg13g2_nand2_1 _13645_ (.Y(_04617_),
    .A(net3369),
    .B(net6605));
 sg13g2_o21ai_1 _13646_ (.B1(_04617_),
    .Y(_00443_),
    .A1(net7342),
    .A2(net6605));
 sg13g2_nand2_1 _13647_ (.Y(_04618_),
    .A(net4047),
    .B(net6604));
 sg13g2_o21ai_1 _13648_ (.B1(_04618_),
    .Y(_00444_),
    .A1(net7540),
    .A2(net6604));
 sg13g2_nand2_1 _13649_ (.Y(_04619_),
    .A(net3226),
    .B(net6604));
 sg13g2_o21ai_1 _13650_ (.B1(_04619_),
    .Y(_00445_),
    .A1(net7700),
    .A2(net6604));
 sg13g2_nor3_2 _13651_ (.A(net7369),
    .B(_04101_),
    .C(net7269),
    .Y(_04620_));
 sg13g2_nor2_1 _13652_ (.A(net4766),
    .B(net6958),
    .Y(_04621_));
 sg13g2_a21oi_1 _13653_ (.A1(net7319),
    .A2(net6958),
    .Y(_00446_),
    .B1(_04621_));
 sg13g2_nor2_1 _13654_ (.A(net4421),
    .B(net6958),
    .Y(_04622_));
 sg13g2_a21oi_1 _13655_ (.A1(net7514),
    .A2(net6958),
    .Y(_00447_),
    .B1(_04622_));
 sg13g2_nor2_1 _13656_ (.A(net3793),
    .B(net6958),
    .Y(_04623_));
 sg13g2_a21oi_1 _13657_ (.A1(net7675),
    .A2(net6958),
    .Y(_00448_),
    .B1(_04623_));
 sg13g2_nand3_1 _13658_ (.B(net7099),
    .C(_04234_),
    .A(net7390),
    .Y(_04624_));
 sg13g2_nand2_1 _13659_ (.Y(_04625_),
    .A(net2517),
    .B(net6602));
 sg13g2_o21ai_1 _13660_ (.B1(_04625_),
    .Y(_00449_),
    .A1(net7341),
    .A2(net6603));
 sg13g2_nand2_1 _13661_ (.Y(_04626_),
    .A(net2926),
    .B(net6602));
 sg13g2_o21ai_1 _13662_ (.B1(_04626_),
    .Y(_00450_),
    .A1(net7539),
    .A2(net6602));
 sg13g2_nand2_1 _13663_ (.Y(_04627_),
    .A(net2527),
    .B(net6602));
 sg13g2_o21ai_1 _13664_ (.B1(_04627_),
    .Y(_00451_),
    .A1(net7700),
    .A2(net6603));
 sg13g2_nand3_1 _13665_ (.B(net7392),
    .C(net7266),
    .A(net7114),
    .Y(_04628_));
 sg13g2_nand2_1 _13666_ (.Y(_04629_),
    .A(net4195),
    .B(net6601));
 sg13g2_o21ai_1 _13667_ (.B1(_04629_),
    .Y(_00452_),
    .A1(net7342),
    .A2(net6601));
 sg13g2_nand2_1 _13668_ (.Y(_04630_),
    .A(net4322),
    .B(net6600));
 sg13g2_o21ai_1 _13669_ (.B1(_04630_),
    .Y(_00453_),
    .A1(net7540),
    .A2(net6600));
 sg13g2_nand2_1 _13670_ (.Y(_04631_),
    .A(net2869),
    .B(net6600));
 sg13g2_o21ai_1 _13671_ (.B1(_04631_),
    .Y(_00454_),
    .A1(net7700),
    .A2(net6600));
 sg13g2_nand3_1 _13672_ (.B(net7099),
    .C(net7067),
    .A(net7394),
    .Y(_04632_));
 sg13g2_nand2_1 _13673_ (.Y(_04633_),
    .A(net2703),
    .B(net6599));
 sg13g2_o21ai_1 _13674_ (.B1(_04633_),
    .Y(_00455_),
    .A1(net7341),
    .A2(net6599));
 sg13g2_nand2_1 _13675_ (.Y(_04634_),
    .A(net3290),
    .B(net6598));
 sg13g2_o21ai_1 _13676_ (.B1(_04634_),
    .Y(_00456_),
    .A1(net7539),
    .A2(net6598));
 sg13g2_nand2_1 _13677_ (.Y(_04635_),
    .A(net4101),
    .B(net6598));
 sg13g2_o21ai_1 _13678_ (.B1(_04635_),
    .Y(_00457_),
    .A1(net7701),
    .A2(net6598));
 sg13g2_nand3_1 _13679_ (.B(net7103),
    .C(net7099),
    .A(net7394),
    .Y(_04636_));
 sg13g2_nand2_1 _13680_ (.Y(_04637_),
    .A(net2876),
    .B(net6597));
 sg13g2_o21ai_1 _13681_ (.B1(_04637_),
    .Y(_00458_),
    .A1(net7341),
    .A2(net6597));
 sg13g2_nand2_1 _13682_ (.Y(_04638_),
    .A(net3334),
    .B(net6596));
 sg13g2_o21ai_1 _13683_ (.B1(_04638_),
    .Y(_00459_),
    .A1(net7539),
    .A2(net6596));
 sg13g2_nand2_1 _13684_ (.Y(_04639_),
    .A(net3847),
    .B(net6597));
 sg13g2_o21ai_1 _13685_ (.B1(_04639_),
    .Y(_00460_),
    .A1(net7701),
    .A2(net6596));
 sg13g2_nand3_1 _13686_ (.B(net7392),
    .C(_04234_),
    .A(net7114),
    .Y(_04640_));
 sg13g2_nand2_1 _13687_ (.Y(_04641_),
    .A(net3833),
    .B(net6595));
 sg13g2_o21ai_1 _13688_ (.B1(_04641_),
    .Y(_00461_),
    .A1(net7342),
    .A2(net6595));
 sg13g2_nand2_1 _13689_ (.Y(_04642_),
    .A(net2818),
    .B(net6594));
 sg13g2_o21ai_1 _13690_ (.B1(_04642_),
    .Y(_00462_),
    .A1(net7540),
    .A2(net6594));
 sg13g2_nand2_1 _13691_ (.Y(_04643_),
    .A(net2674),
    .B(net6594));
 sg13g2_o21ai_1 _13692_ (.B1(_04643_),
    .Y(_00463_),
    .A1(net7700),
    .A2(net6594));
 sg13g2_nand3_1 _13693_ (.B(net7099),
    .C(net7084),
    .A(net7390),
    .Y(_04644_));
 sg13g2_nand2_1 _13694_ (.Y(_04645_),
    .A(net2816),
    .B(net6593));
 sg13g2_o21ai_1 _13695_ (.B1(_04645_),
    .Y(_00464_),
    .A1(net7341),
    .A2(net6593));
 sg13g2_nand2_1 _13696_ (.Y(_04646_),
    .A(net3148),
    .B(net6592));
 sg13g2_o21ai_1 _13697_ (.B1(_04646_),
    .Y(_00465_),
    .A1(net7539),
    .A2(net6592));
 sg13g2_nand2_1 _13698_ (.Y(_04647_),
    .A(net2895),
    .B(net6592));
 sg13g2_o21ai_1 _13699_ (.B1(_04647_),
    .Y(_00466_),
    .A1(net7701),
    .A2(net6592));
 sg13g2_nor3_2 _13700_ (.A(net7374),
    .B(net7097),
    .C(net7234),
    .Y(_04648_));
 sg13g2_nor2_1 _13701_ (.A(net3632),
    .B(net6590),
    .Y(_04649_));
 sg13g2_a21oi_1 _13702_ (.A1(net7341),
    .A2(net6590),
    .Y(_00467_),
    .B1(_04649_));
 sg13g2_nor2_1 _13703_ (.A(net4006),
    .B(net6591),
    .Y(_04650_));
 sg13g2_a21oi_1 _13704_ (.A1(net7539),
    .A2(net6591),
    .Y(_00468_),
    .B1(_04650_));
 sg13g2_nor2_1 _13705_ (.A(net4601),
    .B(net6590),
    .Y(_04651_));
 sg13g2_a21oi_1 _13706_ (.A1(net7700),
    .A2(net6590),
    .Y(_00469_),
    .B1(_04651_));
 sg13g2_nand3_1 _13707_ (.B(net7391),
    .C(net7067),
    .A(net7114),
    .Y(_04652_));
 sg13g2_nand2_1 _13708_ (.Y(_04653_),
    .A(net3764),
    .B(net6588));
 sg13g2_o21ai_1 _13709_ (.B1(_04653_),
    .Y(_00470_),
    .A1(net7344),
    .A2(net6588));
 sg13g2_nand2_1 _13710_ (.Y(_04654_),
    .A(net2649),
    .B(net6588));
 sg13g2_o21ai_1 _13711_ (.B1(_04654_),
    .Y(_00471_),
    .A1(net7541),
    .A2(net6588));
 sg13g2_nand2_1 _13712_ (.Y(_04655_),
    .A(net3955),
    .B(net6589));
 sg13g2_o21ai_1 _13713_ (.B1(_04655_),
    .Y(_00472_),
    .A1(net7702),
    .A2(net6589));
 sg13g2_nand3_1 _13714_ (.B(net7390),
    .C(net7099),
    .A(net7408),
    .Y(_04656_));
 sg13g2_nand2_1 _13715_ (.Y(_04657_),
    .A(net2996),
    .B(net6586));
 sg13g2_o21ai_1 _13716_ (.B1(_04657_),
    .Y(_00473_),
    .A1(net7328),
    .A2(net6586));
 sg13g2_nand2_1 _13717_ (.Y(_04658_),
    .A(net2524),
    .B(net6586));
 sg13g2_o21ai_1 _13718_ (.B1(_04658_),
    .Y(_00474_),
    .A1(net7527),
    .A2(net6586));
 sg13g2_nand2_1 _13719_ (.Y(_04659_),
    .A(net3183),
    .B(net6587));
 sg13g2_o21ai_1 _13720_ (.B1(_04659_),
    .Y(_00475_),
    .A1(net7685),
    .A2(net6586));
 sg13g2_nand3_1 _13721_ (.B(net7282),
    .C(net7099),
    .A(net7390),
    .Y(_04660_));
 sg13g2_nand2_1 _13722_ (.Y(_04661_),
    .A(net2871),
    .B(net6584));
 sg13g2_o21ai_1 _13723_ (.B1(_04661_),
    .Y(_00476_),
    .A1(net7328),
    .A2(net6584));
 sg13g2_nand2_1 _13724_ (.Y(_04662_),
    .A(net3878),
    .B(net6584));
 sg13g2_o21ai_1 _13725_ (.B1(_04662_),
    .Y(_00477_),
    .A1(net7527),
    .A2(net6584));
 sg13g2_nand2_1 _13726_ (.Y(_04663_),
    .A(net3722),
    .B(net6584));
 sg13g2_o21ai_1 _13727_ (.B1(_04663_),
    .Y(_00478_),
    .A1(net7685),
    .A2(net6584));
 sg13g2_nand3_1 _13728_ (.B(net7362),
    .C(net7099),
    .A(net7390),
    .Y(_04664_));
 sg13g2_nand2_1 _13729_ (.Y(_04665_),
    .A(net2850),
    .B(net6582));
 sg13g2_o21ai_1 _13730_ (.B1(_04665_),
    .Y(_00479_),
    .A1(net7328),
    .A2(net6582));
 sg13g2_nand2_1 _13731_ (.Y(_04666_),
    .A(net3487),
    .B(net6582));
 sg13g2_o21ai_1 _13732_ (.B1(_04666_),
    .Y(_00480_),
    .A1(net7527),
    .A2(net6582));
 sg13g2_nand2_1 _13733_ (.Y(_04667_),
    .A(net3506),
    .B(net6582));
 sg13g2_o21ai_1 _13734_ (.B1(_04667_),
    .Y(_00481_),
    .A1(net7685),
    .A2(net6582));
 sg13g2_nor3_2 _13735_ (.A(net7366),
    .B(net7271),
    .C(net7251),
    .Y(_04668_));
 sg13g2_nor2_1 _13736_ (.A(net4094),
    .B(net6956),
    .Y(_04669_));
 sg13g2_a21oi_1 _13737_ (.A1(net7298),
    .A2(net6956),
    .Y(_00482_),
    .B1(_04669_));
 sg13g2_nor2_1 _13738_ (.A(net4582),
    .B(net6956),
    .Y(_04670_));
 sg13g2_a21oi_1 _13739_ (.A1(net7497),
    .A2(net6956),
    .Y(_00483_),
    .B1(_04670_));
 sg13g2_nor2_1 _13740_ (.A(net4559),
    .B(net6957),
    .Y(_04671_));
 sg13g2_a21oi_1 _13741_ (.A1(net7657),
    .A2(net6957),
    .Y(_00484_),
    .B1(_04671_));
 sg13g2_nor3_2 _13742_ (.A(net7374),
    .B(net7107),
    .C(net7097),
    .Y(_04672_));
 sg13g2_nor2_1 _13743_ (.A(net4511),
    .B(net6580),
    .Y(_04673_));
 sg13g2_a21oi_1 _13744_ (.A1(net7328),
    .A2(net6580),
    .Y(_00485_),
    .B1(_04673_));
 sg13g2_nor2_1 _13745_ (.A(net4488),
    .B(net6581),
    .Y(_04674_));
 sg13g2_a21oi_1 _13746_ (.A1(net7527),
    .A2(net6581),
    .Y(_00486_),
    .B1(_04674_));
 sg13g2_nor2_1 _13747_ (.A(net4327),
    .B(net6581),
    .Y(_04675_));
 sg13g2_a21oi_1 _13748_ (.A1(net7685),
    .A2(net6581),
    .Y(_00487_),
    .B1(_04675_));
 sg13g2_nor3_2 _13749_ (.A(net7372),
    .B(net7269),
    .C(net7246),
    .Y(_04676_));
 sg13g2_nor2_1 _13750_ (.A(net4712),
    .B(net6954),
    .Y(_04677_));
 sg13g2_a21oi_1 _13751_ (.A1(net7319),
    .A2(net6954),
    .Y(_00488_),
    .B1(_04677_));
 sg13g2_nor2_1 _13752_ (.A(net4458),
    .B(net6955),
    .Y(_04678_));
 sg13g2_a21oi_1 _13753_ (.A1(net7519),
    .A2(net6955),
    .Y(_00489_),
    .B1(_04678_));
 sg13g2_nor2_1 _13754_ (.A(net3390),
    .B(net6954),
    .Y(_04679_));
 sg13g2_a21oi_1 _13755_ (.A1(net7676),
    .A2(net6954),
    .Y(_00490_),
    .B1(_04679_));
 sg13g2_nor3_2 _13756_ (.A(net7366),
    .B(net7284),
    .C(net7251),
    .Y(_04680_));
 sg13g2_nor2_1 _13757_ (.A(net4038),
    .B(net6952),
    .Y(_04681_));
 sg13g2_a21oi_1 _13758_ (.A1(net7298),
    .A2(net6952),
    .Y(_00491_),
    .B1(_04681_));
 sg13g2_nor2_1 _13759_ (.A(net4577),
    .B(net6952),
    .Y(_04682_));
 sg13g2_a21oi_1 _13760_ (.A1(net7497),
    .A2(net6952),
    .Y(_00492_),
    .B1(_04682_));
 sg13g2_nor2_1 _13761_ (.A(net4744),
    .B(net6953),
    .Y(_04683_));
 sg13g2_a21oi_1 _13762_ (.A1(net7657),
    .A2(net6953),
    .Y(_00493_),
    .B1(_04683_));
 sg13g2_nor3_1 _13763_ (.A(net7374),
    .B(net7097),
    .C(net7272),
    .Y(_04684_));
 sg13g2_nor2_1 _13764_ (.A(net4364),
    .B(net6578),
    .Y(_04685_));
 sg13g2_a21oi_1 _13765_ (.A1(net7327),
    .A2(net6578),
    .Y(_00494_),
    .B1(_04685_));
 sg13g2_nor2_1 _13766_ (.A(net4730),
    .B(net6578),
    .Y(_04686_));
 sg13g2_a21oi_1 _13767_ (.A1(net7526),
    .A2(net6578),
    .Y(_00495_),
    .B1(_04686_));
 sg13g2_nor2_1 _13768_ (.A(net4107),
    .B(net6579),
    .Y(_04687_));
 sg13g2_a21oi_1 _13769_ (.A1(net7684),
    .A2(net6578),
    .Y(_00496_),
    .B1(_04687_));
 sg13g2_nor3_1 _13770_ (.A(net7365),
    .B(net7107),
    .C(net7052),
    .Y(_04688_));
 sg13g2_nor2_1 _13771_ (.A(net4720),
    .B(net6576),
    .Y(_04689_));
 sg13g2_a21oi_1 _13772_ (.A1(net7294),
    .A2(net6576),
    .Y(_00497_),
    .B1(_04689_));
 sg13g2_nor2_1 _13773_ (.A(net3989),
    .B(net6576),
    .Y(_04690_));
 sg13g2_a21oi_1 _13774_ (.A1(net7492),
    .A2(net6577),
    .Y(_00498_),
    .B1(_04690_));
 sg13g2_nor2_1 _13775_ (.A(net4204),
    .B(net6576),
    .Y(_04691_));
 sg13g2_a21oi_1 _13776_ (.A1(net7649),
    .A2(net6576),
    .Y(_00499_),
    .B1(_04691_));
 sg13g2_nor3_1 _13777_ (.A(net7364),
    .B(net7284),
    .C(net7049),
    .Y(_04692_));
 sg13g2_nor2_1 _13778_ (.A(net3865),
    .B(net6575),
    .Y(_04693_));
 sg13g2_a21oi_1 _13779_ (.A1(net7288),
    .A2(net6575),
    .Y(_00500_),
    .B1(_04693_));
 sg13g2_nor2_1 _13780_ (.A(net4383),
    .B(net6574),
    .Y(_04694_));
 sg13g2_a21oi_1 _13781_ (.A1(net7489),
    .A2(net6574),
    .Y(_00501_),
    .B1(_04694_));
 sg13g2_nor2_1 _13782_ (.A(net4512),
    .B(net6575),
    .Y(_04695_));
 sg13g2_a21oi_1 _13783_ (.A1(net7645),
    .A2(net6575),
    .Y(_00502_),
    .B1(_04695_));
 sg13g2_nand3_1 _13784_ (.B(net7094),
    .C(net7237),
    .A(net7375),
    .Y(_04696_));
 sg13g2_nand2_1 _13785_ (.Y(_04697_),
    .A(net3665),
    .B(net6572));
 sg13g2_o21ai_1 _13786_ (.B1(_04697_),
    .Y(_00503_),
    .A1(net7292),
    .A2(net6572));
 sg13g2_nand2_1 _13787_ (.Y(_04698_),
    .A(net3456),
    .B(net6573));
 sg13g2_o21ai_1 _13788_ (.B1(_04698_),
    .Y(_00504_),
    .A1(net7504),
    .A2(net6573));
 sg13g2_nand2_1 _13789_ (.Y(_04699_),
    .A(net3192),
    .B(net6573));
 sg13g2_o21ai_1 _13790_ (.B1(_04699_),
    .Y(_00505_),
    .A1(net7649),
    .A2(net6573));
 sg13g2_nor3_1 _13791_ (.A(net7364),
    .B(net7271),
    .C(net7049),
    .Y(_04700_));
 sg13g2_nor2_1 _13792_ (.A(net4404),
    .B(net6571),
    .Y(_04701_));
 sg13g2_a21oi_1 _13793_ (.A1(net7288),
    .A2(net6571),
    .Y(_00506_),
    .B1(_04701_));
 sg13g2_nor2_1 _13794_ (.A(net4341),
    .B(net6570),
    .Y(_04702_));
 sg13g2_a21oi_1 _13795_ (.A1(net7488),
    .A2(net6570),
    .Y(_00507_),
    .B1(_04702_));
 sg13g2_nor2_1 _13796_ (.A(net4817),
    .B(net6571),
    .Y(_04703_));
 sg13g2_a21oi_1 _13797_ (.A1(net7645),
    .A2(net6571),
    .Y(_00508_),
    .B1(_04703_));
 sg13g2_nor3_1 _13798_ (.A(net7364),
    .B(net7275),
    .C(net7049),
    .Y(_04704_));
 sg13g2_nor2_1 _13799_ (.A(net4703),
    .B(net6569),
    .Y(_04705_));
 sg13g2_a21oi_1 _13800_ (.A1(net7288),
    .A2(net6569),
    .Y(_00509_),
    .B1(_04705_));
 sg13g2_nor2_1 _13801_ (.A(net4770),
    .B(net6568),
    .Y(_04706_));
 sg13g2_a21oi_1 _13802_ (.A1(net7488),
    .A2(net6568),
    .Y(_00510_),
    .B1(_04706_));
 sg13g2_nor2_1 _13803_ (.A(net4422),
    .B(net6569),
    .Y(_04707_));
 sg13g2_a21oi_1 _13804_ (.A1(net7645),
    .A2(net6569),
    .Y(_00511_),
    .B1(_04707_));
 sg13g2_nand3_1 _13805_ (.B(net7094),
    .C(net7264),
    .A(net7375),
    .Y(_04708_));
 sg13g2_nand2_1 _13806_ (.Y(_04709_),
    .A(net2611),
    .B(net6566));
 sg13g2_o21ai_1 _13807_ (.B1(_04709_),
    .Y(_00512_),
    .A1(net7292),
    .A2(net6566));
 sg13g2_nand2_1 _13808_ (.Y(_04710_),
    .A(net2829),
    .B(net6566));
 sg13g2_o21ai_1 _13809_ (.B1(_04710_),
    .Y(_00513_),
    .A1(net7504),
    .A2(net6566));
 sg13g2_nand2_1 _13810_ (.Y(_04711_),
    .A(net3086),
    .B(net6566));
 sg13g2_o21ai_1 _13811_ (.B1(_04711_),
    .Y(_00514_),
    .A1(net7649),
    .A2(net6566));
 sg13g2_nor3_1 _13812_ (.A(net7364),
    .B(net7245),
    .C(net7048),
    .Y(_04712_));
 sg13g2_nor2_1 _13813_ (.A(net4090),
    .B(net6565),
    .Y(_04713_));
 sg13g2_a21oi_1 _13814_ (.A1(net7288),
    .A2(net6565),
    .Y(_00515_),
    .B1(_04713_));
 sg13g2_nor2_1 _13815_ (.A(net4768),
    .B(net6564),
    .Y(_04714_));
 sg13g2_a21oi_1 _13816_ (.A1(net7488),
    .A2(net6564),
    .Y(_00516_),
    .B1(_04714_));
 sg13g2_nor2_1 _13817_ (.A(net4665),
    .B(net6565),
    .Y(_04715_));
 sg13g2_a21oi_1 _13818_ (.A1(net7645),
    .A2(net6565),
    .Y(_00517_),
    .B1(_04715_));
 sg13g2_nor3_2 _13819_ (.A(net7562),
    .B(net7561),
    .C(_04049_),
    .Y(_04716_));
 sg13g2_nand3_1 _13820_ (.B(net7398),
    .C(net7229),
    .A(net7405),
    .Y(_04717_));
 sg13g2_nand2_1 _13821_ (.Y(_04718_),
    .A(net3530),
    .B(net6950));
 sg13g2_o21ai_1 _13822_ (.B1(_04718_),
    .Y(_00518_),
    .A1(net7357),
    .A2(net6950));
 sg13g2_nand2_1 _13823_ (.Y(_04719_),
    .A(net2997),
    .B(net6950));
 sg13g2_o21ai_1 _13824_ (.B1(_04719_),
    .Y(_00519_),
    .A1(net7554),
    .A2(net6950));
 sg13g2_nand2_1 _13825_ (.Y(_04720_),
    .A(net3870),
    .B(net6951));
 sg13g2_o21ai_1 _13826_ (.B1(_04720_),
    .Y(_00520_),
    .A1(net7714),
    .A2(net6951));
 sg13g2_nand3_1 _13827_ (.B(net7094),
    .C(net7236),
    .A(net7375),
    .Y(_04721_));
 sg13g2_nand2_1 _13828_ (.Y(_04722_),
    .A(net3787),
    .B(net6562));
 sg13g2_o21ai_1 _13829_ (.B1(_04722_),
    .Y(_00521_),
    .A1(net7292),
    .A2(net6562));
 sg13g2_nand2_1 _13830_ (.Y(_04723_),
    .A(net2686),
    .B(net6562));
 sg13g2_o21ai_1 _13831_ (.B1(_04723_),
    .Y(_00522_),
    .A1(net7491),
    .A2(net6562));
 sg13g2_nand2_1 _13832_ (.Y(_04724_),
    .A(net2557),
    .B(net6562));
 sg13g2_o21ai_1 _13833_ (.B1(_04724_),
    .Y(_00523_),
    .A1(net7649),
    .A2(net6562));
 sg13g2_nand3_1 _13834_ (.B(net7238),
    .C(net7229),
    .A(net7398),
    .Y(_04725_));
 sg13g2_nand2_1 _13835_ (.Y(_04726_),
    .A(net3239),
    .B(net6948));
 sg13g2_o21ai_1 _13836_ (.B1(_04726_),
    .Y(_00524_),
    .A1(net7351),
    .A2(net6948));
 sg13g2_nand2_1 _13837_ (.Y(_04727_),
    .A(net3331),
    .B(net6948));
 sg13g2_o21ai_1 _13838_ (.B1(_04727_),
    .Y(_00525_),
    .A1(net7554),
    .A2(net6948));
 sg13g2_nand2_1 _13839_ (.Y(_04728_),
    .A(net3621),
    .B(net6949));
 sg13g2_o21ai_1 _13840_ (.B1(_04728_),
    .Y(_00526_),
    .A1(net7714),
    .A2(net6949));
 sg13g2_nand3_1 _13841_ (.B(net7265),
    .C(net7229),
    .A(net7398),
    .Y(_04729_));
 sg13g2_nand2_1 _13842_ (.Y(_04730_),
    .A(net2969),
    .B(net6946));
 sg13g2_o21ai_1 _13843_ (.B1(_04730_),
    .Y(_00527_),
    .A1(net7351),
    .A2(net6946));
 sg13g2_nand2_1 _13844_ (.Y(_04731_),
    .A(net2470),
    .B(net6946));
 sg13g2_o21ai_1 _13845_ (.B1(_04731_),
    .Y(_00528_),
    .A1(net7554),
    .A2(net6946));
 sg13g2_nand2_1 _13846_ (.Y(_04732_),
    .A(net2787),
    .B(net6947));
 sg13g2_o21ai_1 _13847_ (.B1(_04732_),
    .Y(_00529_),
    .A1(net7714),
    .A2(net6947));
 sg13g2_nand3_1 _13848_ (.B(net7094),
    .C(net7065),
    .A(net7375),
    .Y(_04733_));
 sg13g2_nand2_1 _13849_ (.Y(_04734_),
    .A(net2469),
    .B(net6560));
 sg13g2_o21ai_1 _13850_ (.B1(_04734_),
    .Y(_00530_),
    .A1(net7293),
    .A2(net6560));
 sg13g2_nand2_1 _13851_ (.Y(_04735_),
    .A(net3898),
    .B(net6560));
 sg13g2_o21ai_1 _13852_ (.B1(_04735_),
    .Y(_00531_),
    .A1(net7491),
    .A2(net6560));
 sg13g2_nand2_1 _13853_ (.Y(_04736_),
    .A(net3041),
    .B(net6561));
 sg13g2_o21ai_1 _13854_ (.B1(_04736_),
    .Y(_00532_),
    .A1(net7651),
    .A2(net6561));
 sg13g2_nand3_1 _13855_ (.B(net7235),
    .C(net7228),
    .A(net7398),
    .Y(_04737_));
 sg13g2_nand2_1 _13856_ (.Y(_04738_),
    .A(net3097),
    .B(net6944));
 sg13g2_o21ai_1 _13857_ (.B1(_04738_),
    .Y(_00533_),
    .A1(net7351),
    .A2(net6944));
 sg13g2_nand2_1 _13858_ (.Y(_04739_),
    .A(net2857),
    .B(net6944));
 sg13g2_o21ai_1 _13859_ (.B1(_04739_),
    .Y(_00534_),
    .A1(net7554),
    .A2(net6944));
 sg13g2_nand2_1 _13860_ (.Y(_04740_),
    .A(net2761),
    .B(net6945));
 sg13g2_o21ai_1 _13861_ (.B1(_04740_),
    .Y(_00535_),
    .A1(net7711),
    .A2(net6945));
 sg13g2_nor3_1 _13862_ (.A(net7373),
    .B(_04065_),
    .C(net7269),
    .Y(_04741_));
 sg13g2_nor2_1 _13863_ (.A(net4607),
    .B(net6559),
    .Y(_04742_));
 sg13g2_a21oi_1 _13864_ (.A1(net7320),
    .A2(net6559),
    .Y(_00536_),
    .B1(_04742_));
 sg13g2_nor2_1 _13865_ (.A(net4363),
    .B(net6559),
    .Y(_04743_));
 sg13g2_a21oi_1 _13866_ (.A1(net7519),
    .A2(net6559),
    .Y(_00537_),
    .B1(_04743_));
 sg13g2_nor2_1 _13867_ (.A(net4604),
    .B(net6558),
    .Y(_04744_));
 sg13g2_a21oi_1 _13868_ (.A1(net7675),
    .A2(net6558),
    .Y(_00538_),
    .B1(_04744_));
 sg13g2_nand3_1 _13869_ (.B(net7104),
    .C(net7094),
    .A(net7375),
    .Y(_04745_));
 sg13g2_nand2_1 _13870_ (.Y(_04746_),
    .A(net4048),
    .B(net6557));
 sg13g2_o21ai_1 _13871_ (.B1(_04746_),
    .Y(_00539_),
    .A1(net7293),
    .A2(net6557));
 sg13g2_nand2_1 _13872_ (.Y(_04747_),
    .A(net2721),
    .B(net6556));
 sg13g2_o21ai_1 _13873_ (.B1(_04747_),
    .Y(_00540_),
    .A1(net7491),
    .A2(net6556));
 sg13g2_nand2_1 _13874_ (.Y(_04748_),
    .A(net3640),
    .B(net6557));
 sg13g2_o21ai_1 _13875_ (.B1(_04748_),
    .Y(_00541_),
    .A1(net7651),
    .A2(net6557));
 sg13g2_nand3_1 _13876_ (.B(net7103),
    .C(net7230),
    .A(net7399),
    .Y(_04749_));
 sg13g2_nand2_1 _13877_ (.Y(_04750_),
    .A(net4787),
    .B(net6555));
 sg13g2_o21ai_1 _13878_ (.B1(_04750_),
    .Y(_00542_),
    .A1(net7354),
    .A2(net6555));
 sg13g2_nand2_1 _13879_ (.Y(_04751_),
    .A(net4302),
    .B(net6555));
 sg13g2_o21ai_1 _13880_ (.B1(_04751_),
    .Y(_00543_),
    .A1(net7551),
    .A2(net6555));
 sg13g2_nand2_1 _13881_ (.Y(_04752_),
    .A(net3255),
    .B(net6554));
 sg13g2_o21ai_1 _13882_ (.B1(_04752_),
    .Y(_00544_),
    .A1(net7710),
    .A2(net6554));
 sg13g2_nand3_1 _13883_ (.B(net7084),
    .C(net7230),
    .A(net7399),
    .Y(_04753_));
 sg13g2_nand2_1 _13884_ (.Y(_04754_),
    .A(net3537),
    .B(net6553));
 sg13g2_o21ai_1 _13885_ (.B1(_04754_),
    .Y(_00545_),
    .A1(net7354),
    .A2(net6553));
 sg13g2_nand2_1 _13886_ (.Y(_04755_),
    .A(net3735),
    .B(net6553));
 sg13g2_o21ai_1 _13887_ (.B1(_04755_),
    .Y(_00546_),
    .A1(net7551),
    .A2(net6553));
 sg13g2_nand2_1 _13888_ (.Y(_04756_),
    .A(net2794),
    .B(net6552));
 sg13g2_o21ai_1 _13889_ (.B1(_04756_),
    .Y(_00547_),
    .A1(net7710),
    .A2(net6552));
 sg13g2_nor3_2 _13890_ (.A(net7373),
    .B(net7269),
    .C(net7234),
    .Y(_04757_));
 sg13g2_nor2_1 _13891_ (.A(net4792),
    .B(net6942),
    .Y(_04758_));
 sg13g2_a21oi_1 _13892_ (.A1(net7319),
    .A2(net6942),
    .Y(_00548_),
    .B1(_04758_));
 sg13g2_nor2_1 _13893_ (.A(net4850),
    .B(net6942),
    .Y(_04759_));
 sg13g2_a21oi_1 _13894_ (.A1(net7514),
    .A2(net6942),
    .Y(_00549_),
    .B1(_04759_));
 sg13g2_nor2_1 _13895_ (.A(net4522),
    .B(net6943),
    .Y(_04760_));
 sg13g2_a21oi_1 _13896_ (.A1(net7675),
    .A2(net6943),
    .Y(_00550_),
    .B1(_04760_));
 sg13g2_nand3_1 _13897_ (.B(net7042),
    .C(net7230),
    .A(net7399),
    .Y(_04761_));
 sg13g2_nand2_1 _13898_ (.Y(_04762_),
    .A(net2783),
    .B(net6551));
 sg13g2_o21ai_1 _13899_ (.B1(_04762_),
    .Y(_00551_),
    .A1(net7354),
    .A2(net6551));
 sg13g2_nand2_1 _13900_ (.Y(_04763_),
    .A(net2706),
    .B(net6551));
 sg13g2_o21ai_1 _13901_ (.B1(_04763_),
    .Y(_00552_),
    .A1(net7551),
    .A2(net6551));
 sg13g2_nand2_1 _13902_ (.Y(_04764_),
    .A(net2801),
    .B(net6550));
 sg13g2_o21ai_1 _13903_ (.B1(_04764_),
    .Y(_00553_),
    .A1(net7710),
    .A2(net6550));
 sg13g2_nand3_1 _13904_ (.B(net7397),
    .C(net7228),
    .A(net7409),
    .Y(_04765_));
 sg13g2_nand2_1 _13905_ (.Y(_04766_),
    .A(net3727),
    .B(net6941));
 sg13g2_o21ai_1 _13906_ (.B1(_04766_),
    .Y(_00554_),
    .A1(net7351),
    .A2(net6941));
 sg13g2_nand2_1 _13907_ (.Y(_04767_),
    .A(net3539),
    .B(net6941));
 sg13g2_o21ai_1 _13908_ (.B1(_04767_),
    .Y(_00555_),
    .A1(net7549),
    .A2(net6941));
 sg13g2_nand2_1 _13909_ (.Y(_04768_),
    .A(net2740),
    .B(net6940));
 sg13g2_o21ai_1 _13910_ (.B1(_04768_),
    .Y(_00556_),
    .A1(net7711),
    .A2(net6940));
 sg13g2_nor3_1 _13911_ (.A(net7369),
    .B(net7092),
    .C(net7234),
    .Y(_04769_));
 sg13g2_nor2_1 _13912_ (.A(net4350),
    .B(net6549),
    .Y(_04770_));
 sg13g2_a21oi_1 _13913_ (.A1(net7293),
    .A2(net6548),
    .Y(_00557_),
    .B1(_04770_));
 sg13g2_nor2_1 _13914_ (.A(net4669),
    .B(net6548),
    .Y(_04771_));
 sg13g2_a21oi_1 _13915_ (.A1(net7491),
    .A2(net6548),
    .Y(_00558_),
    .B1(_04771_));
 sg13g2_nor2_1 _13916_ (.A(net4325),
    .B(net6549),
    .Y(_04772_));
 sg13g2_a21oi_1 _13917_ (.A1(net7651),
    .A2(net6549),
    .Y(_00559_),
    .B1(_04772_));
 sg13g2_nand3_1 _13918_ (.B(net7283),
    .C(net7228),
    .A(net7397),
    .Y(_04773_));
 sg13g2_nand2_1 _13919_ (.Y(_04774_),
    .A(net3071),
    .B(net6939));
 sg13g2_o21ai_1 _13920_ (.B1(_04774_),
    .Y(_00560_),
    .A1(net7351),
    .A2(net6939));
 sg13g2_nand2_1 _13921_ (.Y(_04775_),
    .A(net2679),
    .B(net6939));
 sg13g2_o21ai_1 _13922_ (.B1(_04775_),
    .Y(_00561_),
    .A1(net7549),
    .A2(net6939));
 sg13g2_nand2_1 _13923_ (.Y(_04776_),
    .A(net4470),
    .B(net6938));
 sg13g2_o21ai_1 _13924_ (.B1(_04776_),
    .Y(_00562_),
    .A1(net7711),
    .A2(net6938));
 sg13g2_nand3_1 _13925_ (.B(net7363),
    .C(net7228),
    .A(net7397),
    .Y(_04777_));
 sg13g2_nand2_1 _13926_ (.Y(_04778_),
    .A(net2510),
    .B(net6937));
 sg13g2_o21ai_1 _13927_ (.B1(_04778_),
    .Y(_00563_),
    .A1(net7351),
    .A2(net6937));
 sg13g2_nand2_1 _13928_ (.Y(_04779_),
    .A(net3197),
    .B(net6937));
 sg13g2_o21ai_1 _13929_ (.B1(_04779_),
    .Y(_00564_),
    .A1(net7549),
    .A2(net6937));
 sg13g2_nand2_1 _13930_ (.Y(_04780_),
    .A(net3234),
    .B(net6936));
 sg13g2_o21ai_1 _13931_ (.B1(_04780_),
    .Y(_00565_),
    .A1(net7711),
    .A2(net6936));
 sg13g2_nand3_1 _13932_ (.B(net7376),
    .C(net7095),
    .A(net7406),
    .Y(_04781_));
 sg13g2_nand2_1 _13933_ (.Y(_04782_),
    .A(net3679),
    .B(net6547));
 sg13g2_o21ai_1 _13934_ (.B1(_04782_),
    .Y(_00566_),
    .A1(net7296),
    .A2(net6546));
 sg13g2_nand2_1 _13935_ (.Y(_04783_),
    .A(net3741),
    .B(net6547));
 sg13g2_o21ai_1 _13936_ (.B1(_04783_),
    .Y(_00567_),
    .A1(net7507),
    .A2(net6547));
 sg13g2_nand2_1 _13937_ (.Y(_04784_),
    .A(net2779),
    .B(net6546));
 sg13g2_o21ai_1 _13938_ (.B1(_04784_),
    .Y(_00568_),
    .A1(net7651),
    .A2(net6546));
 sg13g2_nand3_1 _13939_ (.B(net7279),
    .C(net7228),
    .A(net7397),
    .Y(_04785_));
 sg13g2_nand2_1 _13940_ (.Y(_04786_),
    .A(net2638),
    .B(net6935));
 sg13g2_o21ai_1 _13941_ (.B1(_04786_),
    .Y(_00569_),
    .A1(net7351),
    .A2(net6935));
 sg13g2_nand2_1 _13942_ (.Y(_04787_),
    .A(net3437),
    .B(net6934));
 sg13g2_o21ai_1 _13943_ (.B1(_04787_),
    .Y(_00570_),
    .A1(net7549),
    .A2(net6935));
 sg13g2_nand2_1 _13944_ (.Y(_04788_),
    .A(net4102),
    .B(net6934));
 sg13g2_o21ai_1 _13945_ (.B1(_04788_),
    .Y(_00571_),
    .A1(net7711),
    .A2(net6935));
 sg13g2_nand3_1 _13946_ (.B(net7286),
    .C(net7229),
    .A(net7397),
    .Y(_04789_));
 sg13g2_nand2_1 _13947_ (.Y(_04790_),
    .A(net4054),
    .B(net6933));
 sg13g2_o21ai_1 _13948_ (.B1(_04790_),
    .Y(_00572_),
    .A1(net7353),
    .A2(net6933));
 sg13g2_nand2_1 _13949_ (.Y(_04791_),
    .A(net2805),
    .B(net6932));
 sg13g2_o21ai_1 _13950_ (.B1(_04791_),
    .Y(_00573_),
    .A1(net7557),
    .A2(net6932));
 sg13g2_nand2_1 _13951_ (.Y(_04792_),
    .A(net2562),
    .B(net6932));
 sg13g2_o21ai_1 _13952_ (.B1(_04792_),
    .Y(_00574_),
    .A1(net7712),
    .A2(net6932));
 sg13g2_nand3_1 _13953_ (.B(net7281),
    .C(net7095),
    .A(net7376),
    .Y(_04793_));
 sg13g2_nand2_1 _13954_ (.Y(_04794_),
    .A(net3782),
    .B(net6545));
 sg13g2_o21ai_1 _13955_ (.B1(_04794_),
    .Y(_00575_),
    .A1(net7296),
    .A2(net6544));
 sg13g2_nand2_1 _13956_ (.Y(_04795_),
    .A(net2815),
    .B(net6545));
 sg13g2_o21ai_1 _13957_ (.B1(_04795_),
    .Y(_00576_),
    .A1(net7507),
    .A2(net6545));
 sg13g2_nand2_1 _13958_ (.Y(_04796_),
    .A(net3203),
    .B(net6544));
 sg13g2_o21ai_1 _13959_ (.B1(_04796_),
    .Y(_00577_),
    .A1(net7651),
    .A2(net6544));
 sg13g2_nand3_1 _13960_ (.B(net7274),
    .C(net7228),
    .A(net7397),
    .Y(_04797_));
 sg13g2_nand2_1 _13961_ (.Y(_04798_),
    .A(net4389),
    .B(net6931));
 sg13g2_o21ai_1 _13962_ (.B1(_04798_),
    .Y(_00578_),
    .A1(net7353),
    .A2(net6931));
 sg13g2_nand2_1 _13963_ (.Y(_04799_),
    .A(net2955),
    .B(net6930));
 sg13g2_o21ai_1 _13964_ (.B1(_04799_),
    .Y(_00579_),
    .A1(net7550),
    .A2(net6930));
 sg13g2_nand2_1 _13965_ (.Y(_04800_),
    .A(net3411),
    .B(net6930));
 sg13g2_o21ai_1 _13966_ (.B1(_04800_),
    .Y(_00580_),
    .A1(net7711),
    .A2(net6930));
 sg13g2_nor3_2 _13967_ (.A(net7372),
    .B(_04093_),
    .C(net7270),
    .Y(_04801_));
 sg13g2_nor2_1 _13968_ (.A(net4523),
    .B(net6543),
    .Y(_04802_));
 sg13g2_a21oi_1 _13969_ (.A1(net7320),
    .A2(net6543),
    .Y(_00581_),
    .B1(_04802_));
 sg13g2_nor2_1 _13970_ (.A(net4521),
    .B(net6543),
    .Y(_04803_));
 sg13g2_a21oi_1 _13971_ (.A1(net7519),
    .A2(net6543),
    .Y(_00582_),
    .B1(_04803_));
 sg13g2_nor2_1 _13972_ (.A(net4189),
    .B(net6542),
    .Y(_04804_));
 sg13g2_a21oi_1 _13973_ (.A1(net7675),
    .A2(net6542),
    .Y(_00583_),
    .B1(_04804_));
 sg13g2_nand3_1 _13974_ (.B(net7361),
    .C(net7094),
    .A(net7375),
    .Y(_04805_));
 sg13g2_nand2_1 _13975_ (.Y(_04806_),
    .A(net2966),
    .B(net6541));
 sg13g2_o21ai_1 _13976_ (.B1(_04806_),
    .Y(_00584_),
    .A1(net7296),
    .A2(net6540));
 sg13g2_nand2_1 _13977_ (.Y(_04807_),
    .A(net3631),
    .B(net6541));
 sg13g2_o21ai_1 _13978_ (.B1(_04807_),
    .Y(_00585_),
    .A1(net7507),
    .A2(net6541));
 sg13g2_nand2_1 _13979_ (.Y(_04808_),
    .A(net3475),
    .B(net6540));
 sg13g2_o21ai_1 _13980_ (.B1(_04808_),
    .Y(_00586_),
    .A1(net7651),
    .A2(net6540));
 sg13g2_nand3_1 _13981_ (.B(net7072),
    .C(net7235),
    .A(net7395),
    .Y(_04809_));
 sg13g2_nand2_1 _13982_ (.Y(_04810_),
    .A(net2893),
    .B(net6539));
 sg13g2_o21ai_1 _13983_ (.B1(_04810_),
    .Y(_00587_),
    .A1(net7352),
    .A2(net6539));
 sg13g2_nand2_1 _13984_ (.Y(_04811_),
    .A(net2590),
    .B(net6539));
 sg13g2_o21ai_1 _13985_ (.B1(_04811_),
    .Y(_00588_),
    .A1(net7550),
    .A2(net6539));
 sg13g2_nand2_1 _13986_ (.Y(_04812_),
    .A(net3400),
    .B(net6538));
 sg13g2_o21ai_1 _13987_ (.B1(_04812_),
    .Y(_00589_),
    .A1(net7696),
    .A2(net6538));
 sg13g2_nand3_1 _13988_ (.B(net7077),
    .C(net7067),
    .A(net7396),
    .Y(_04813_));
 sg13g2_nand2_1 _13989_ (.Y(_04814_),
    .A(net3426),
    .B(net6537));
 sg13g2_o21ai_1 _13990_ (.B1(_04814_),
    .Y(_00590_),
    .A1(net7352),
    .A2(net6537));
 sg13g2_nand2_1 _13991_ (.Y(_04815_),
    .A(net4126),
    .B(net6536));
 sg13g2_o21ai_1 _13992_ (.B1(_04815_),
    .Y(_00591_),
    .A1(net7549),
    .A2(net6536));
 sg13g2_nand2_1 _13993_ (.Y(_04816_),
    .A(net2860),
    .B(net6536));
 sg13g2_o21ai_1 _13994_ (.B1(_04816_),
    .Y(_00592_),
    .A1(net7709),
    .A2(net6536));
 sg13g2_nand3_1 _13995_ (.B(net7072),
    .C(net7238),
    .A(net7395),
    .Y(_04817_));
 sg13g2_nand2_1 _13996_ (.Y(_04818_),
    .A(net3515),
    .B(net6535));
 sg13g2_o21ai_1 _13997_ (.B1(_04818_),
    .Y(_00593_),
    .A1(net7352),
    .A2(net6535));
 sg13g2_nand2_1 _13998_ (.Y(_04819_),
    .A(net3035),
    .B(net6535));
 sg13g2_o21ai_1 _13999_ (.B1(_04819_),
    .Y(_00594_),
    .A1(net7550),
    .A2(net6535));
 sg13g2_nand2_1 _14000_ (.Y(_04820_),
    .A(net3751),
    .B(net6534));
 sg13g2_o21ai_1 _14001_ (.B1(_04820_),
    .Y(_00595_),
    .A1(net7696),
    .A2(net6534));
 sg13g2_nand3_1 _14002_ (.B(net7103),
    .C(net7072),
    .A(net7396),
    .Y(_04821_));
 sg13g2_nand2_1 _14003_ (.Y(_04822_),
    .A(net2848),
    .B(net6533));
 sg13g2_o21ai_1 _14004_ (.B1(_04822_),
    .Y(_00596_),
    .A1(net7352),
    .A2(net6533));
 sg13g2_nand2_1 _14005_ (.Y(_04823_),
    .A(net3789),
    .B(net6532));
 sg13g2_o21ai_1 _14006_ (.B1(_04823_),
    .Y(_00597_),
    .A1(net7549),
    .A2(net6532));
 sg13g2_nand2_1 _14007_ (.Y(_04824_),
    .A(net2702),
    .B(net6532));
 sg13g2_o21ai_1 _14008_ (.B1(_04824_),
    .Y(_00598_),
    .A1(net7709),
    .A2(net6532));
 sg13g2_nand3_1 _14009_ (.B(net7282),
    .C(net7072),
    .A(net7387),
    .Y(_04825_));
 sg13g2_nand2_1 _14010_ (.Y(_04826_),
    .A(net2581),
    .B(net6530));
 sg13g2_o21ai_1 _14011_ (.B1(_04826_),
    .Y(_00599_),
    .A1(net7339),
    .A2(net6530));
 sg13g2_nand2_1 _14012_ (.Y(_04827_),
    .A(net2532),
    .B(net6531));
 sg13g2_o21ai_1 _14013_ (.B1(_04827_),
    .Y(_00600_),
    .A1(net7537),
    .A2(net6531));
 sg13g2_nand2_1 _14014_ (.Y(_04828_),
    .A(net3690),
    .B(net6530));
 sg13g2_o21ai_1 _14015_ (.B1(_04828_),
    .Y(_00601_),
    .A1(net7697),
    .A2(net6530));
 sg13g2_nand3_1 _14016_ (.B(net7073),
    .C(net7042),
    .A(net7396),
    .Y(_04829_));
 sg13g2_nand2_1 _14017_ (.Y(_04830_),
    .A(net3408),
    .B(net6529));
 sg13g2_o21ai_1 _14018_ (.B1(_04830_),
    .Y(_00602_),
    .A1(net7352),
    .A2(net6529));
 sg13g2_nand2_1 _14019_ (.Y(_04831_),
    .A(net4033),
    .B(net6528));
 sg13g2_o21ai_1 _14020_ (.B1(_04831_),
    .Y(_00603_),
    .A1(net7549),
    .A2(net6528));
 sg13g2_nand2_1 _14021_ (.Y(_04832_),
    .A(net2931),
    .B(net6528));
 sg13g2_o21ai_1 _14022_ (.B1(_04832_),
    .Y(_00604_),
    .A1(net7709),
    .A2(net6528));
 sg13g2_nor3_1 _14023_ (.A(net7365),
    .B(_04065_),
    .C(net7051),
    .Y(_04833_));
 sg13g2_nor2_1 _14024_ (.A(net3644),
    .B(net6526),
    .Y(_04834_));
 sg13g2_a21oi_1 _14025_ (.A1(net7294),
    .A2(net6526),
    .Y(_00605_),
    .B1(_04834_));
 sg13g2_nor2_1 _14026_ (.A(net4143),
    .B(net6526),
    .Y(_04835_));
 sg13g2_a21oi_1 _14027_ (.A1(net7493),
    .A2(net6526),
    .Y(_00606_),
    .B1(_04835_));
 sg13g2_nor2_1 _14028_ (.A(net4666),
    .B(net6526),
    .Y(_04836_));
 sg13g2_a21oi_1 _14029_ (.A1(net7649),
    .A2(net6526),
    .Y(_00607_),
    .B1(_04836_));
 sg13g2_nand3_1 _14030_ (.B(net7066),
    .C(net7230),
    .A(net7399),
    .Y(_04837_));
 sg13g2_nand2_1 _14031_ (.Y(_04838_),
    .A(net4182),
    .B(net6525));
 sg13g2_o21ai_1 _14032_ (.B1(_04838_),
    .Y(_00608_),
    .A1(net7354),
    .A2(net6525));
 sg13g2_nand2_1 _14033_ (.Y(_04839_),
    .A(net4269),
    .B(net6525));
 sg13g2_o21ai_1 _14034_ (.B1(_04839_),
    .Y(_00609_),
    .A1(net7551),
    .A2(net6525));
 sg13g2_nand2_1 _14035_ (.Y(_04840_),
    .A(net3604),
    .B(net6524));
 sg13g2_o21ai_1 _14036_ (.B1(_04840_),
    .Y(_00610_),
    .A1(net7710),
    .A2(net6524));
 sg13g2_nand3_1 _14037_ (.B(net7104),
    .C(net7244),
    .A(net7381),
    .Y(_04841_));
 sg13g2_nand2_1 _14038_ (.Y(_04842_),
    .A(net3128),
    .B(net6522));
 sg13g2_o21ai_1 _14039_ (.B1(_04842_),
    .Y(_00611_),
    .A1(net7334),
    .A2(net6522));
 sg13g2_nand2_1 _14040_ (.Y(_04843_),
    .A(net3221),
    .B(net6522));
 sg13g2_o21ai_1 _14041_ (.B1(_04843_),
    .Y(_00612_),
    .A1(net7531),
    .A2(net6522));
 sg13g2_nand2_1 _14042_ (.Y(_04844_),
    .A(net3965),
    .B(net6523));
 sg13g2_o21ai_1 _14043_ (.B1(_04844_),
    .Y(_00613_),
    .A1(net7692),
    .A2(net6523));
 sg13g2_nand3_1 _14044_ (.B(net7278),
    .C(net7228),
    .A(net7397),
    .Y(_04845_));
 sg13g2_nand2_1 _14045_ (.Y(_04846_),
    .A(net4095),
    .B(net6929));
 sg13g2_o21ai_1 _14046_ (.B1(_04846_),
    .Y(_00614_),
    .A1(net7353),
    .A2(net6929));
 sg13g2_nand2_1 _14047_ (.Y(_04847_),
    .A(net3969),
    .B(net6928));
 sg13g2_o21ai_1 _14048_ (.B1(_04847_),
    .Y(_00615_),
    .A1(net7550),
    .A2(net6928));
 sg13g2_nand2_1 _14049_ (.Y(_04848_),
    .A(net3461),
    .B(net6928));
 sg13g2_o21ai_1 _14050_ (.B1(_04848_),
    .Y(_00616_),
    .A1(net7711),
    .A2(net6928));
 sg13g2_nand3_1 _14051_ (.B(net7387),
    .C(net7072),
    .A(net7408),
    .Y(_04849_));
 sg13g2_nand2_1 _14052_ (.Y(_04850_),
    .A(net3410),
    .B(net6520));
 sg13g2_o21ai_1 _14053_ (.B1(_04850_),
    .Y(_00617_),
    .A1(net7339),
    .A2(net6520));
 sg13g2_nand2_1 _14054_ (.Y(_04851_),
    .A(net3370),
    .B(net6521));
 sg13g2_o21ai_1 _14055_ (.B1(_04851_),
    .Y(_00618_),
    .A1(net7537),
    .A2(net6521));
 sg13g2_nand2_1 _14056_ (.Y(_04852_),
    .A(net3852),
    .B(net6520));
 sg13g2_o21ai_1 _14057_ (.B1(_04852_),
    .Y(_00619_),
    .A1(net7697),
    .A2(net6520));
 sg13g2_nand3_1 _14058_ (.B(net7085),
    .C(net7244),
    .A(net7385),
    .Y(_04853_));
 sg13g2_nand2_1 _14059_ (.Y(_04854_),
    .A(net3934),
    .B(net6518));
 sg13g2_o21ai_1 _14060_ (.B1(_04854_),
    .Y(_00620_),
    .A1(net7334),
    .A2(net6518));
 sg13g2_nand2_1 _14061_ (.Y(_04855_),
    .A(net3810),
    .B(net6518));
 sg13g2_o21ai_1 _14062_ (.B1(_04855_),
    .Y(_00621_),
    .A1(net7530),
    .A2(net6518));
 sg13g2_nand2_1 _14063_ (.Y(_04856_),
    .A(net3129),
    .B(net6519));
 sg13g2_o21ai_1 _14064_ (.B1(_04856_),
    .Y(_00622_),
    .A1(net7691),
    .A2(net6519));
 sg13g2_nand3_1 _14065_ (.B(net7264),
    .C(net7243),
    .A(net7381),
    .Y(_04857_));
 sg13g2_nand2_1 _14066_ (.Y(_04858_),
    .A(net4425),
    .B(net6927));
 sg13g2_o21ai_1 _14067_ (.B1(_04858_),
    .Y(_00623_),
    .A1(net7334),
    .A2(net6927));
 sg13g2_nand2_1 _14068_ (.Y(_04859_),
    .A(net4515),
    .B(net6926));
 sg13g2_o21ai_1 _14069_ (.B1(_04859_),
    .Y(_00624_),
    .A1(net7531),
    .A2(net6926));
 sg13g2_nand2_1 _14070_ (.Y(_04860_),
    .A(net3120),
    .B(net6926));
 sg13g2_o21ai_1 _14071_ (.B1(_04860_),
    .Y(_00625_),
    .A1(net7676),
    .A2(net6926));
 sg13g2_nand3_1 _14072_ (.B(net7285),
    .C(net7244),
    .A(net7385),
    .Y(_04861_));
 sg13g2_nand2_1 _14073_ (.Y(_04862_),
    .A(net2613),
    .B(net6924));
 sg13g2_o21ai_1 _14074_ (.B1(_04862_),
    .Y(_00626_),
    .A1(net7335),
    .A2(net6924));
 sg13g2_nand2_1 _14075_ (.Y(_04863_),
    .A(net3899),
    .B(net6925));
 sg13g2_o21ai_1 _14076_ (.B1(_04863_),
    .Y(_00627_),
    .A1(net7532),
    .A2(net6925));
 sg13g2_nand2_1 _14077_ (.Y(_04864_),
    .A(net3985),
    .B(net6925));
 sg13g2_o21ai_1 _14078_ (.B1(_04864_),
    .Y(_00628_),
    .A1(net7693),
    .A2(net6925));
 sg13g2_nand3_1 _14079_ (.B(net7243),
    .C(net7043),
    .A(net7381),
    .Y(_04865_));
 sg13g2_nand2_1 _14080_ (.Y(_04866_),
    .A(net3767),
    .B(net6516));
 sg13g2_o21ai_1 _14081_ (.B1(_04866_),
    .Y(_00629_),
    .A1(net7334),
    .A2(net6516));
 sg13g2_nand2_1 _14082_ (.Y(_04867_),
    .A(net3822),
    .B(net6516));
 sg13g2_o21ai_1 _14083_ (.B1(_04867_),
    .Y(_00630_),
    .A1(net7531),
    .A2(net6516));
 sg13g2_nand2_1 _14084_ (.Y(_04868_),
    .A(net4494),
    .B(net6517));
 sg13g2_o21ai_1 _14085_ (.B1(_04868_),
    .Y(_00631_),
    .A1(net7692),
    .A2(net6517));
 sg13g2_nor2_2 _14086_ (.A(\top1.addr_in[8] ),
    .B(_04059_),
    .Y(_04869_));
 sg13g2_nand2b_2 _14087_ (.Y(_04870_),
    .B(_04058_),
    .A_N(\top1.addr_in[8] ));
 sg13g2_nor3_1 _14088_ (.A(net7267),
    .B(_04152_),
    .C(net7199),
    .Y(_04871_));
 sg13g2_nor2_1 _14089_ (.A(net4424),
    .B(net6923),
    .Y(_04872_));
 sg13g2_a21oi_1 _14090_ (.A1(net7309),
    .A2(net6923),
    .Y(_00632_),
    .B1(_04872_));
 sg13g2_nor2_1 _14091_ (.A(net4836),
    .B(net6922),
    .Y(_04873_));
 sg13g2_a21oi_1 _14092_ (.A1(net7511),
    .A2(net6922),
    .Y(_00633_),
    .B1(_04873_));
 sg13g2_nor2_1 _14093_ (.A(net3730),
    .B(net6922),
    .Y(_04874_));
 sg13g2_a21oi_1 _14094_ (.A1(net7666),
    .A2(net6922),
    .Y(_00634_),
    .B1(_04874_));
 sg13g2_nand3_1 _14095_ (.B(net7383),
    .C(net7243),
    .A(net7407),
    .Y(_04875_));
 sg13g2_nand2_1 _14096_ (.Y(_04876_),
    .A(net4608),
    .B(net6921));
 sg13g2_o21ai_1 _14097_ (.B1(_04876_),
    .Y(_00635_),
    .A1(net7333),
    .A2(net6921));
 sg13g2_nand2_1 _14098_ (.Y(_04877_),
    .A(net2873),
    .B(net6920));
 sg13g2_o21ai_1 _14099_ (.B1(_04877_),
    .Y(_00636_),
    .A1(net7530),
    .A2(net6920));
 sg13g2_nand2_1 _14100_ (.Y(_04878_),
    .A(net2778),
    .B(net6921));
 sg13g2_o21ai_1 _14101_ (.B1(_04878_),
    .Y(_00637_),
    .A1(net7692),
    .A2(net6921));
 sg13g2_nand3_1 _14102_ (.B(net7283),
    .C(net7243),
    .A(net7383),
    .Y(_04879_));
 sg13g2_nand2_1 _14103_ (.Y(_04880_),
    .A(net2708),
    .B(net6919));
 sg13g2_o21ai_1 _14104_ (.B1(_04880_),
    .Y(_00638_),
    .A1(net7333),
    .A2(net6919));
 sg13g2_nand2_1 _14105_ (.Y(_04881_),
    .A(net3891),
    .B(net6918));
 sg13g2_o21ai_1 _14106_ (.B1(_04881_),
    .Y(_00639_),
    .A1(net7530),
    .A2(net6918));
 sg13g2_nand2_1 _14107_ (.Y(_04882_),
    .A(net4276),
    .B(net6919));
 sg13g2_o21ai_1 _14108_ (.B1(_04882_),
    .Y(_00640_),
    .A1(net7692),
    .A2(net6919));
 sg13g2_nand3_1 _14109_ (.B(net7363),
    .C(net7243),
    .A(net7381),
    .Y(_04883_));
 sg13g2_nand2_1 _14110_ (.Y(_04884_),
    .A(net3580),
    .B(net6917));
 sg13g2_o21ai_1 _14111_ (.B1(_04884_),
    .Y(_00641_),
    .A1(net7333),
    .A2(net6917));
 sg13g2_nand2_1 _14112_ (.Y(_04885_),
    .A(net2883),
    .B(net6916));
 sg13g2_o21ai_1 _14113_ (.B1(_04885_),
    .Y(_00642_),
    .A1(net7530),
    .A2(net6916));
 sg13g2_nand2_1 _14114_ (.Y(_04886_),
    .A(net4042),
    .B(net6917));
 sg13g2_o21ai_1 _14115_ (.B1(_04886_),
    .Y(_00643_),
    .A1(net7692),
    .A2(net6917));
 sg13g2_nor3_2 _14116_ (.A(net7367),
    .B(_04087_),
    .C(net7252),
    .Y(_04887_));
 sg13g2_nor2_1 _14117_ (.A(net4469),
    .B(net6514),
    .Y(_04888_));
 sg13g2_a21oi_1 _14118_ (.A1(net7299),
    .A2(net6514),
    .Y(_00644_),
    .B1(_04888_));
 sg13g2_nor2_1 _14119_ (.A(net4127),
    .B(net6514),
    .Y(_04889_));
 sg13g2_a21oi_1 _14120_ (.A1(net7498),
    .A2(net6514),
    .Y(_00645_),
    .B1(_04889_));
 sg13g2_nor2_1 _14121_ (.A(net4346),
    .B(net6515),
    .Y(_04890_));
 sg13g2_a21oi_1 _14122_ (.A1(net7658),
    .A2(net6515),
    .Y(_00646_),
    .B1(_04890_));
 sg13g2_nor3_1 _14123_ (.A(net7368),
    .B(_04065_),
    .C(net7252),
    .Y(_04891_));
 sg13g2_nor2_1 _14124_ (.A(net3901),
    .B(net6512),
    .Y(_04892_));
 sg13g2_a21oi_1 _14125_ (.A1(net7299),
    .A2(net6512),
    .Y(_00647_),
    .B1(_04892_));
 sg13g2_nor2_1 _14126_ (.A(net3906),
    .B(net6512),
    .Y(_04893_));
 sg13g2_a21oi_1 _14127_ (.A1(net7498),
    .A2(net6512),
    .Y(_00648_),
    .B1(_04893_));
 sg13g2_nor2_1 _14128_ (.A(net4092),
    .B(net6512),
    .Y(_04894_));
 sg13g2_a21oi_1 _14129_ (.A1(net7658),
    .A2(net6512),
    .Y(_00649_),
    .B1(_04894_));
 sg13g2_nor3_2 _14130_ (.A(net7368),
    .B(net7107),
    .C(net7252),
    .Y(_04895_));
 sg13g2_nor2_1 _14131_ (.A(net4719),
    .B(net6510),
    .Y(_04896_));
 sg13g2_a21oi_1 _14132_ (.A1(net7298),
    .A2(net6510),
    .Y(_00650_),
    .B1(_04896_));
 sg13g2_nor2_1 _14133_ (.A(net4480),
    .B(net6510),
    .Y(_04897_));
 sg13g2_a21oi_1 _14134_ (.A1(net7498),
    .A2(net6510),
    .Y(_00651_),
    .B1(_04897_));
 sg13g2_nor2_1 _14135_ (.A(net4560),
    .B(net6511),
    .Y(_04898_));
 sg13g2_a21oi_1 _14136_ (.A1(net7658),
    .A2(net6511),
    .Y(_00652_),
    .B1(_04898_));
 sg13g2_nor3_1 _14137_ (.A(net7369),
    .B(net7107),
    .C(net7092),
    .Y(_04899_));
 sg13g2_nor2_1 _14138_ (.A(net4741),
    .B(net6509),
    .Y(_04900_));
 sg13g2_a21oi_1 _14139_ (.A1(net7295),
    .A2(net6508),
    .Y(_00653_),
    .B1(_04900_));
 sg13g2_nor2_1 _14140_ (.A(net4534),
    .B(net6509),
    .Y(_04901_));
 sg13g2_a21oi_1 _14141_ (.A1(net7507),
    .A2(net6509),
    .Y(_00654_),
    .B1(_04901_));
 sg13g2_nor2_1 _14142_ (.A(net4618),
    .B(net6508),
    .Y(_04902_));
 sg13g2_a21oi_1 _14143_ (.A1(net7651),
    .A2(net6508),
    .Y(_00655_),
    .B1(_04902_));
 sg13g2_nor3_1 _14144_ (.A(net7369),
    .B(net7284),
    .C(net7092),
    .Y(_04903_));
 sg13g2_nor2_1 _14145_ (.A(net4845),
    .B(net6506),
    .Y(_04904_));
 sg13g2_a21oi_1 _14146_ (.A1(net7292),
    .A2(net6506),
    .Y(_00656_),
    .B1(_04904_));
 sg13g2_nor2_1 _14147_ (.A(net4001),
    .B(net6506),
    .Y(_04905_));
 sg13g2_a21oi_1 _14148_ (.A1(net7491),
    .A2(net6506),
    .Y(_00657_),
    .B1(_04905_));
 sg13g2_nor2_1 _14149_ (.A(net4495),
    .B(net6507),
    .Y(_04906_));
 sg13g2_a21oi_1 _14150_ (.A1(net7650),
    .A2(net6507),
    .Y(_00658_),
    .B1(_04906_));
 sg13g2_nand3_1 _14151_ (.B(net7396),
    .C(net7077),
    .A(net7405),
    .Y(_04907_));
 sg13g2_nand2_1 _14152_ (.Y(_04908_),
    .A(net2849),
    .B(net6505));
 sg13g2_o21ai_1 _14153_ (.B1(_04908_),
    .Y(_00659_),
    .A1(net7352),
    .A2(net6505));
 sg13g2_nand2_1 _14154_ (.Y(_04909_),
    .A(net3815),
    .B(net6505));
 sg13g2_o21ai_1 _14155_ (.B1(_04909_),
    .Y(_00660_),
    .A1(net7550),
    .A2(net6505));
 sg13g2_nand2_1 _14156_ (.Y(_04910_),
    .A(net3199),
    .B(net6504));
 sg13g2_o21ai_1 _14157_ (.B1(_04910_),
    .Y(_00661_),
    .A1(net7696),
    .A2(net6504));
 sg13g2_nand3_1 _14158_ (.B(net7084),
    .C(net7072),
    .A(net7395),
    .Y(_04911_));
 sg13g2_nand2_1 _14159_ (.Y(_04912_),
    .A(net3821),
    .B(net6503));
 sg13g2_o21ai_1 _14160_ (.B1(_04912_),
    .Y(_00662_),
    .A1(net7352),
    .A2(net6503));
 sg13g2_nand2_1 _14161_ (.Y(_04913_),
    .A(net4565),
    .B(net6502));
 sg13g2_o21ai_1 _14162_ (.B1(_04913_),
    .Y(_00663_),
    .A1(net7549),
    .A2(net6502));
 sg13g2_nand2_1 _14163_ (.Y(_04914_),
    .A(net3474),
    .B(net6502));
 sg13g2_o21ai_1 _14164_ (.B1(_04914_),
    .Y(_00664_),
    .A1(net7709),
    .A2(net6502));
 sg13g2_nand3_1 _14165_ (.B(net7248),
    .C(net7228),
    .A(net7397),
    .Y(_04915_));
 sg13g2_nand2_1 _14166_ (.Y(_04916_),
    .A(net3142),
    .B(net6915));
 sg13g2_o21ai_1 _14167_ (.B1(_04916_),
    .Y(_00665_),
    .A1(net7351),
    .A2(net6915));
 sg13g2_nand2_1 _14168_ (.Y(_04917_),
    .A(net4011),
    .B(net6914));
 sg13g2_o21ai_1 _14169_ (.B1(_04917_),
    .Y(_00666_),
    .A1(net7550),
    .A2(net6914));
 sg13g2_nand2_1 _14170_ (.Y(_04918_),
    .A(net3508),
    .B(net6914));
 sg13g2_o21ai_1 _14171_ (.B1(_04918_),
    .Y(_00667_),
    .A1(net7711),
    .A2(net6914));
 sg13g2_nand3_1 _14172_ (.B(net7280),
    .C(net7243),
    .A(net7381),
    .Y(_04919_));
 sg13g2_nand2_1 _14173_ (.Y(_04920_),
    .A(net3176),
    .B(net6913));
 sg13g2_o21ai_1 _14174_ (.B1(_04920_),
    .Y(_00668_),
    .A1(net7333),
    .A2(net6913));
 sg13g2_nand2_1 _14175_ (.Y(_04921_),
    .A(net2958),
    .B(net6912));
 sg13g2_o21ai_1 _14176_ (.B1(_04921_),
    .Y(_00669_),
    .A1(net7530),
    .A2(net6912));
 sg13g2_nand2_1 _14177_ (.Y(_04922_),
    .A(net3907),
    .B(net6913));
 sg13g2_o21ai_1 _14178_ (.B1(_04922_),
    .Y(_00670_),
    .A1(net7692),
    .A2(net6913));
 sg13g2_nand3_1 _14179_ (.B(net7362),
    .C(net7072),
    .A(net7387),
    .Y(_04923_));
 sg13g2_nand2_1 _14180_ (.Y(_04924_),
    .A(net4137),
    .B(net6500));
 sg13g2_o21ai_1 _14181_ (.B1(_04924_),
    .Y(_00671_),
    .A1(net7339),
    .A2(net6500));
 sg13g2_nand2_1 _14182_ (.Y(_04925_),
    .A(net4050),
    .B(net6501));
 sg13g2_o21ai_1 _14183_ (.B1(_04925_),
    .Y(_00672_),
    .A1(net7537),
    .A2(net6501));
 sg13g2_nand2_1 _14184_ (.Y(_04926_),
    .A(net2974),
    .B(net6500));
 sg13g2_o21ai_1 _14185_ (.B1(_04926_),
    .Y(_00673_),
    .A1(net7697),
    .A2(net6500));
 sg13g2_nand3_1 _14186_ (.B(net7236),
    .C(net7203),
    .A(net7096),
    .Y(_04927_));
 sg13g2_nand2_1 _14187_ (.Y(_04928_),
    .A(net2549),
    .B(net6499));
 sg13g2_o21ai_1 _14188_ (.B1(_04928_),
    .Y(_00674_),
    .A1(net7306),
    .A2(net6499));
 sg13g2_nand2_1 _14189_ (.Y(_04929_),
    .A(net3705),
    .B(net6498));
 sg13g2_o21ai_1 _14190_ (.B1(_04929_),
    .Y(_00675_),
    .A1(net7505),
    .A2(net6498));
 sg13g2_nand2_1 _14191_ (.Y(_04930_),
    .A(net3238),
    .B(net6498));
 sg13g2_o21ai_1 _14192_ (.B1(_04930_),
    .Y(_00676_),
    .A1(net7664),
    .A2(net6498));
 sg13g2_nand3_1 _14193_ (.B(net7264),
    .C(net7203),
    .A(net7096),
    .Y(_04931_));
 sg13g2_nand2_1 _14194_ (.Y(_04932_),
    .A(net2479),
    .B(net6497));
 sg13g2_o21ai_1 _14195_ (.B1(_04932_),
    .Y(_00677_),
    .A1(net7306),
    .A2(net6497));
 sg13g2_nand2_1 _14196_ (.Y(_04933_),
    .A(net2535),
    .B(net6496));
 sg13g2_o21ai_1 _14197_ (.B1(_04933_),
    .Y(_00678_),
    .A1(net7505),
    .A2(net6496));
 sg13g2_nand2_1 _14198_ (.Y(_04934_),
    .A(net3646),
    .B(net6496));
 sg13g2_o21ai_1 _14199_ (.B1(_04934_),
    .Y(_00679_),
    .A1(net7664),
    .A2(net6496));
 sg13g2_nand3_1 _14200_ (.B(net7237),
    .C(net7203),
    .A(net7096),
    .Y(_04935_));
 sg13g2_nand2_1 _14201_ (.Y(_04936_),
    .A(net2797),
    .B(net6495));
 sg13g2_o21ai_1 _14202_ (.B1(_04936_),
    .Y(_00680_),
    .A1(net7306),
    .A2(net6495));
 sg13g2_nand2_1 _14203_ (.Y(_04937_),
    .A(net3846),
    .B(net6494));
 sg13g2_o21ai_1 _14204_ (.B1(_04937_),
    .Y(_00681_),
    .A1(net7505),
    .A2(net6494));
 sg13g2_nand2_1 _14205_ (.Y(_04938_),
    .A(net3425),
    .B(net6494));
 sg13g2_o21ai_1 _14206_ (.B1(_04938_),
    .Y(_00682_),
    .A1(net7664),
    .A2(net6494));
 sg13g2_nand3_1 _14207_ (.B(net7096),
    .C(net7203),
    .A(net7403),
    .Y(_04939_));
 sg13g2_nand2_1 _14208_ (.Y(_04940_),
    .A(net2991),
    .B(net6493));
 sg13g2_o21ai_1 _14209_ (.B1(_04940_),
    .Y(_00683_),
    .A1(net7306),
    .A2(net6493));
 sg13g2_nand2_1 _14210_ (.Y(_04941_),
    .A(net3025),
    .B(net6492));
 sg13g2_o21ai_1 _14211_ (.B1(_04941_),
    .Y(_00684_),
    .A1(net7505),
    .A2(net6492));
 sg13g2_nand2_1 _14212_ (.Y(_04942_),
    .A(net2770),
    .B(net6492));
 sg13g2_o21ai_1 _14213_ (.B1(_04942_),
    .Y(_00685_),
    .A1(net7664),
    .A2(net6492));
 sg13g2_nand3_1 _14214_ (.B(net7080),
    .C(net7208),
    .A(net7083),
    .Y(_04943_));
 sg13g2_nand2_1 _14215_ (.Y(_04944_),
    .A(net2983),
    .B(net6490));
 sg13g2_o21ai_1 _14216_ (.B1(_04944_),
    .Y(_00686_),
    .A1(net7324),
    .A2(net6490));
 sg13g2_nand2_1 _14217_ (.Y(_04945_),
    .A(net2986),
    .B(net6490));
 sg13g2_o21ai_1 _14218_ (.B1(_04945_),
    .Y(_00687_),
    .A1(net7523),
    .A2(net6490));
 sg13g2_nand2_1 _14219_ (.Y(_04946_),
    .A(net4026),
    .B(net6490));
 sg13g2_o21ai_1 _14220_ (.B1(_04946_),
    .Y(_00688_),
    .A1(net7680),
    .A2(net6490));
 sg13g2_nand3_1 _14221_ (.B(net7065),
    .C(net7203),
    .A(_04118_),
    .Y(_04947_));
 sg13g2_nand2_1 _14222_ (.Y(_04948_),
    .A(net3186),
    .B(net6489));
 sg13g2_o21ai_1 _14223_ (.B1(_04948_),
    .Y(_00689_),
    .A1(net7307),
    .A2(net6489));
 sg13g2_nand2_1 _14224_ (.Y(_04949_),
    .A(net2457),
    .B(net6488));
 sg13g2_o21ai_1 _14225_ (.B1(_04949_),
    .Y(_00690_),
    .A1(net7505),
    .A2(net6488));
 sg13g2_nand2_1 _14226_ (.Y(_04950_),
    .A(net2530),
    .B(net6488));
 sg13g2_o21ai_1 _14227_ (.B1(_04950_),
    .Y(_00691_),
    .A1(net7664),
    .A2(net6488));
 sg13g2_nand3_1 _14228_ (.B(net7096),
    .C(net7203),
    .A(net7104),
    .Y(_04951_));
 sg13g2_nand2_1 _14229_ (.Y(_04952_),
    .A(net3045),
    .B(net6487));
 sg13g2_o21ai_1 _14230_ (.B1(_04952_),
    .Y(_00692_),
    .A1(net7307),
    .A2(net6487));
 sg13g2_nand2_1 _14231_ (.Y(_04953_),
    .A(net3528),
    .B(net6486));
 sg13g2_o21ai_1 _14232_ (.B1(_04953_),
    .Y(_00693_),
    .A1(net7505),
    .A2(net6486));
 sg13g2_nand2_1 _14233_ (.Y(_04954_),
    .A(net2550),
    .B(net6487));
 sg13g2_o21ai_1 _14234_ (.B1(_04954_),
    .Y(_00694_),
    .A1(net7665),
    .A2(net6486));
 sg13g2_nand3_1 _14235_ (.B(net7257),
    .C(net7205),
    .A(net7361),
    .Y(_04955_));
 sg13g2_nand2_1 _14236_ (.Y(_04956_),
    .A(net3494),
    .B(net6910));
 sg13g2_o21ai_1 _14237_ (.B1(_04956_),
    .Y(_00695_),
    .A1(net7295),
    .A2(net6910));
 sg13g2_nand2_1 _14238_ (.Y(_04957_),
    .A(net2972),
    .B(net6910));
 sg13g2_o21ai_1 _14239_ (.B1(_04957_),
    .Y(_00696_),
    .A1(net7493),
    .A2(net6910));
 sg13g2_nand2_1 _14240_ (.Y(_04958_),
    .A(net3189),
    .B(net6911));
 sg13g2_o21ai_1 _14241_ (.B1(_04958_),
    .Y(_00697_),
    .A1(net7652),
    .A2(net6911));
 sg13g2_nor3_1 _14242_ (.A(net7271),
    .B(net7093),
    .C(net7198),
    .Y(_04959_));
 sg13g2_nor2_1 _14243_ (.A(net4661),
    .B(net6484),
    .Y(_04960_));
 sg13g2_a21oi_1 _14244_ (.A1(net7306),
    .A2(net6484),
    .Y(_00698_),
    .B1(_04960_));
 sg13g2_nor2_1 _14245_ (.A(net4816),
    .B(net6485),
    .Y(_04961_));
 sg13g2_a21oi_1 _14246_ (.A1(net7504),
    .A2(net6485),
    .Y(_00699_),
    .B1(_04961_));
 sg13g2_nor2_1 _14247_ (.A(net4518),
    .B(net6484),
    .Y(_04962_));
 sg13g2_a21oi_1 _14248_ (.A1(net7663),
    .A2(net6484),
    .Y(_00700_),
    .B1(_04962_));
 sg13g2_nor3_1 _14249_ (.A(net7284),
    .B(net7093),
    .C(net7198),
    .Y(_04963_));
 sg13g2_nor2_1 _14250_ (.A(net4593),
    .B(net6482),
    .Y(_04964_));
 sg13g2_a21oi_1 _14251_ (.A1(net7306),
    .A2(net6482),
    .Y(_00701_),
    .B1(_04964_));
 sg13g2_nor2_1 _14252_ (.A(net4409),
    .B(net6483),
    .Y(_04965_));
 sg13g2_a21oi_1 _14253_ (.A1(net7504),
    .A2(net6483),
    .Y(_00702_),
    .B1(_04965_));
 sg13g2_nor2_1 _14254_ (.A(net4497),
    .B(net6482),
    .Y(_04966_));
 sg13g2_a21oi_1 _14255_ (.A1(net7663),
    .A2(net6482),
    .Y(_00703_),
    .B1(_04966_));
 sg13g2_nand3_1 _14256_ (.B(net7254),
    .C(net7207),
    .A(net7403),
    .Y(_04967_));
 sg13g2_nand2_1 _14257_ (.Y(_04968_),
    .A(net2488),
    .B(net6908));
 sg13g2_o21ai_1 _14258_ (.B1(_04968_),
    .Y(_00704_),
    .A1(net7304),
    .A2(net6908));
 sg13g2_nand2_1 _14259_ (.Y(_04969_),
    .A(net3414),
    .B(net6908));
 sg13g2_o21ai_1 _14260_ (.B1(_04969_),
    .Y(_00705_),
    .A1(net7502),
    .A2(net6908));
 sg13g2_nand2_1 _14261_ (.Y(_04970_),
    .A(net4075),
    .B(net6909));
 sg13g2_o21ai_1 _14262_ (.B1(_04970_),
    .Y(_00706_),
    .A1(net7661),
    .A2(net6909));
 sg13g2_nor3_1 _14263_ (.A(net7107),
    .B(net7093),
    .C(net7198),
    .Y(_04971_));
 sg13g2_nor2_1 _14264_ (.A(net4530),
    .B(net6480),
    .Y(_04972_));
 sg13g2_a21oi_1 _14265_ (.A1(net7314),
    .A2(net6480),
    .Y(_00707_),
    .B1(_04972_));
 sg13g2_nor2_1 _14266_ (.A(net4017),
    .B(net6481),
    .Y(_04973_));
 sg13g2_a21oi_1 _14267_ (.A1(net7506),
    .A2(net6481),
    .Y(_00708_),
    .B1(_04973_));
 sg13g2_nor2_1 _14268_ (.A(net4563),
    .B(net6480),
    .Y(_04974_));
 sg13g2_a21oi_1 _14269_ (.A1(net7664),
    .A2(net6480),
    .Y(_00709_),
    .B1(_04974_));
 sg13g2_nand3_1 _14270_ (.B(net7095),
    .C(net7205),
    .A(net7361),
    .Y(_04975_));
 sg13g2_nand2_1 _14271_ (.Y(_04976_),
    .A(net4440),
    .B(net6478));
 sg13g2_o21ai_1 _14272_ (.B1(_04976_),
    .Y(_00710_),
    .A1(net7308),
    .A2(net6478));
 sg13g2_nand2_1 _14273_ (.Y(_04977_),
    .A(net2898),
    .B(net6479));
 sg13g2_o21ai_1 _14274_ (.B1(_04977_),
    .Y(_00711_),
    .A1(net7507),
    .A2(net6479));
 sg13g2_nand2_1 _14275_ (.Y(_04978_),
    .A(net3381),
    .B(net6478));
 sg13g2_o21ai_1 _14276_ (.B1(_04978_),
    .Y(_00712_),
    .A1(net7663),
    .A2(net6478));
 sg13g2_nand3_1 _14277_ (.B(net7096),
    .C(net7205),
    .A(net7281),
    .Y(_04979_));
 sg13g2_nand2_1 _14278_ (.Y(_04980_),
    .A(net3538),
    .B(net6476));
 sg13g2_o21ai_1 _14279_ (.B1(_04980_),
    .Y(_00713_),
    .A1(net7308),
    .A2(net6476));
 sg13g2_nand2_1 _14280_ (.Y(_04981_),
    .A(net3268),
    .B(net6476));
 sg13g2_o21ai_1 _14281_ (.B1(_04981_),
    .Y(_00714_),
    .A1(net7506),
    .A2(net6476));
 sg13g2_nand2_1 _14282_ (.Y(_04982_),
    .A(net3190),
    .B(net6476));
 sg13g2_o21ai_1 _14283_ (.B1(_04982_),
    .Y(_00715_),
    .A1(net7663),
    .A2(net6476));
 sg13g2_nand3_1 _14284_ (.B(net7096),
    .C(net7203),
    .A(net7406),
    .Y(_04983_));
 sg13g2_nand2_1 _14285_ (.Y(_04984_),
    .A(net2792),
    .B(net6474));
 sg13g2_o21ai_1 _14286_ (.B1(_04984_),
    .Y(_00716_),
    .A1(net7308),
    .A2(net6474));
 sg13g2_nand2_1 _14287_ (.Y(_04985_),
    .A(net2930),
    .B(net6475));
 sg13g2_o21ai_1 _14288_ (.B1(_04985_),
    .Y(_00717_),
    .A1(net7506),
    .A2(net6475));
 sg13g2_nand2_1 _14289_ (.Y(_04986_),
    .A(net2807),
    .B(net6474));
 sg13g2_o21ai_1 _14290_ (.B1(_04986_),
    .Y(_00718_),
    .A1(net7663),
    .A2(net6474));
 sg13g2_nor3_1 _14291_ (.A(net7093),
    .B(net7234),
    .C(net7199),
    .Y(_04987_));
 sg13g2_nor2_1 _14292_ (.A(net3779),
    .B(net6472),
    .Y(_04988_));
 sg13g2_a21oi_1 _14293_ (.A1(net7307),
    .A2(net6472),
    .Y(_00719_),
    .B1(_04988_));
 sg13g2_nor2_1 _14294_ (.A(net3555),
    .B(net6472),
    .Y(_04989_));
 sg13g2_a21oi_1 _14295_ (.A1(net7505),
    .A2(net6472),
    .Y(_00720_),
    .B1(_04989_));
 sg13g2_nor2_1 _14296_ (.A(net4573),
    .B(net6473),
    .Y(_04990_));
 sg13g2_a21oi_1 _14297_ (.A1(net7663),
    .A2(net6473),
    .Y(_00721_),
    .B1(_04990_));
 sg13g2_nor3_1 _14298_ (.A(net7268),
    .B(_04291_),
    .C(net7201),
    .Y(_04991_));
 sg13g2_nor2_1 _14299_ (.A(net4446),
    .B(net6907),
    .Y(_04992_));
 sg13g2_a21oi_1 _14300_ (.A1(net7309),
    .A2(net6907),
    .Y(_00722_),
    .B1(_04992_));
 sg13g2_nor2_1 _14301_ (.A(net4776),
    .B(net6906),
    .Y(_04993_));
 sg13g2_a21oi_1 _14302_ (.A1(net7511),
    .A2(net6906),
    .Y(_00723_),
    .B1(_04993_));
 sg13g2_nor2_1 _14303_ (.A(net4600),
    .B(net6906),
    .Y(_04994_));
 sg13g2_a21oi_1 _14304_ (.A1(net7666),
    .A2(net6906),
    .Y(_00724_),
    .B1(_04994_));
 sg13g2_nand3_1 _14305_ (.B(net7117),
    .C(net7217),
    .A(net7409),
    .Y(_04995_));
 sg13g2_nand2_1 _14306_ (.Y(_04996_),
    .A(net3112),
    .B(net6470));
 sg13g2_o21ai_1 _14307_ (.B1(_04996_),
    .Y(_00725_),
    .A1(net7347),
    .A2(net6470));
 sg13g2_nand2_1 _14308_ (.Y(_04997_),
    .A(net4340),
    .B(net6471));
 sg13g2_o21ai_1 _14309_ (.B1(_04997_),
    .Y(_00726_),
    .A1(net7545),
    .A2(net6471));
 sg13g2_nand2_1 _14310_ (.Y(_04998_),
    .A(net3849),
    .B(net6470));
 sg13g2_o21ai_1 _14311_ (.B1(_04998_),
    .Y(_00727_),
    .A1(net7704),
    .A2(net6470));
 sg13g2_nor3_1 _14312_ (.A(net7275),
    .B(net7249),
    .C(net7194),
    .Y(_04999_));
 sg13g2_nor2_1 _14313_ (.A(net4735),
    .B(net6904),
    .Y(_05000_));
 sg13g2_a21oi_1 _14314_ (.A1(net7289),
    .A2(net6904),
    .Y(_00728_),
    .B1(_05000_));
 sg13g2_nor2_1 _14315_ (.A(net3592),
    .B(net6905),
    .Y(_05001_));
 sg13g2_a21oi_1 _14316_ (.A1(net7495),
    .A2(net6905),
    .Y(_00729_),
    .B1(_05001_));
 sg13g2_nor2_1 _14317_ (.A(net4214),
    .B(net6905),
    .Y(_05002_));
 sg13g2_a21oi_1 _14318_ (.A1(net7647),
    .A2(net6905),
    .Y(_00730_),
    .B1(_05002_));
 sg13g2_nor3_1 _14319_ (.A(net7250),
    .B(_04184_),
    .C(net7195),
    .Y(_05003_));
 sg13g2_nor2_1 _14320_ (.A(net4438),
    .B(net6903),
    .Y(_05004_));
 sg13g2_a21oi_1 _14321_ (.A1(net7297),
    .A2(net6903),
    .Y(_00731_),
    .B1(_05004_));
 sg13g2_nor2_1 _14322_ (.A(net4198),
    .B(net6903),
    .Y(_05005_));
 sg13g2_a21oi_1 _14323_ (.A1(net7496),
    .A2(net6903),
    .Y(_00732_),
    .B1(_05005_));
 sg13g2_nor2_1 _14324_ (.A(net3850),
    .B(net6902),
    .Y(_05006_));
 sg13g2_a21oi_1 _14325_ (.A1(net7655),
    .A2(net6902),
    .Y(_00733_),
    .B1(_05006_));
 sg13g2_nor3_1 _14326_ (.A(_04235_),
    .B(net7052),
    .C(net7192),
    .Y(_05007_));
 sg13g2_nor2_1 _14327_ (.A(net4673),
    .B(net6468),
    .Y(_05008_));
 sg13g2_a21oi_1 _14328_ (.A1(net7289),
    .A2(net6468),
    .Y(_00734_),
    .B1(_05008_));
 sg13g2_nor2_1 _14329_ (.A(net4284),
    .B(net6468),
    .Y(_05009_));
 sg13g2_a21oi_1 _14330_ (.A1(net7490),
    .A2(net6468),
    .Y(_00735_),
    .B1(_05009_));
 sg13g2_nor2_1 _14331_ (.A(net4386),
    .B(net6469),
    .Y(_05010_));
 sg13g2_a21oi_1 _14332_ (.A1(net7647),
    .A2(net6469),
    .Y(_00736_),
    .B1(_05010_));
 sg13g2_nor3_1 _14333_ (.A(_04141_),
    .B(net7050),
    .C(net7192),
    .Y(_05011_));
 sg13g2_nor2_1 _14334_ (.A(net4799),
    .B(net6466),
    .Y(_05012_));
 sg13g2_a21oi_1 _14335_ (.A1(net7289),
    .A2(net6466),
    .Y(_00737_),
    .B1(_05012_));
 sg13g2_nor2_1 _14336_ (.A(net4245),
    .B(net6466),
    .Y(_05013_));
 sg13g2_a21oi_1 _14337_ (.A1(net7490),
    .A2(net6466),
    .Y(_00738_),
    .B1(_05013_));
 sg13g2_nor2_1 _14338_ (.A(net3859),
    .B(net6467),
    .Y(_05014_));
 sg13g2_a21oi_1 _14339_ (.A1(net7647),
    .A2(net6467),
    .Y(_00739_),
    .B1(_05014_));
 sg13g2_nor3_1 _14340_ (.A(_04217_),
    .B(net7050),
    .C(net7192),
    .Y(_05015_));
 sg13g2_nor2_1 _14341_ (.A(net4658),
    .B(net6464),
    .Y(_05016_));
 sg13g2_a21oi_1 _14342_ (.A1(net7289),
    .A2(net6464),
    .Y(_00740_),
    .B1(_05016_));
 sg13g2_nor2_1 _14343_ (.A(net4857),
    .B(net6464),
    .Y(_05017_));
 sg13g2_a21oi_1 _14344_ (.A1(net7490),
    .A2(net6464),
    .Y(_00741_),
    .B1(_05017_));
 sg13g2_nor2_1 _14345_ (.A(net4270),
    .B(net6465),
    .Y(_05018_));
 sg13g2_a21oi_1 _14346_ (.A1(net7647),
    .A2(net6465),
    .Y(_00742_),
    .B1(_05018_));
 sg13g2_nand3_1 _14347_ (.B(_04129_),
    .C(net7211),
    .A(net7407),
    .Y(_05019_));
 sg13g2_nand2_1 _14348_ (.Y(_05020_),
    .A(net3108),
    .B(net6901));
 sg13g2_o21ai_1 _14349_ (.B1(_05020_),
    .Y(_00743_),
    .A1(net7312),
    .A2(net6901));
 sg13g2_nand2_1 _14350_ (.Y(_05021_),
    .A(net2603),
    .B(net6901));
 sg13g2_o21ai_1 _14351_ (.B1(_05021_),
    .Y(_00744_),
    .A1(net7510),
    .A2(net6900));
 sg13g2_nand2_1 _14352_ (.Y(_05022_),
    .A(net4141),
    .B(net6900));
 sg13g2_o21ai_1 _14353_ (.B1(_05022_),
    .Y(_00745_),
    .A1(net7669),
    .A2(net6900));
 sg13g2_nor3_1 _14354_ (.A(net7092),
    .B(net7245),
    .C(net7198),
    .Y(_05023_));
 sg13g2_nor2_1 _14355_ (.A(net4760),
    .B(net6462),
    .Y(_05024_));
 sg13g2_a21oi_1 _14356_ (.A1(net7306),
    .A2(net6462),
    .Y(_00746_),
    .B1(_05024_));
 sg13g2_nor2_1 _14357_ (.A(net4683),
    .B(net6463),
    .Y(_05025_));
 sg13g2_a21oi_1 _14358_ (.A1(net7504),
    .A2(net6462),
    .Y(_00747_),
    .B1(_05025_));
 sg13g2_nor2_1 _14359_ (.A(net4321),
    .B(net6462),
    .Y(_05026_));
 sg13g2_a21oi_1 _14360_ (.A1(net7663),
    .A2(net6463),
    .Y(_00748_),
    .B1(_05026_));
 sg13g2_nor3_1 _14361_ (.A(net7275),
    .B(net7092),
    .C(net7198),
    .Y(_05027_));
 sg13g2_nor2_1 _14362_ (.A(net3957),
    .B(net6460),
    .Y(_05028_));
 sg13g2_a21oi_1 _14363_ (.A1(net7306),
    .A2(net6460),
    .Y(_00749_),
    .B1(_05028_));
 sg13g2_nor2_1 _14364_ (.A(net3937),
    .B(net6461),
    .Y(_05029_));
 sg13g2_a21oi_1 _14365_ (.A1(net7504),
    .A2(net6461),
    .Y(_00750_),
    .B1(_05029_));
 sg13g2_nor2_1 _14366_ (.A(net4849),
    .B(net6460),
    .Y(_05030_));
 sg13g2_a21oi_1 _14367_ (.A1(net7663),
    .A2(net6460),
    .Y(_00751_),
    .B1(_05030_));
 sg13g2_nand3_1 _14368_ (.B(net7242),
    .C(net7210),
    .A(net7266),
    .Y(_05031_));
 sg13g2_nand2_1 _14369_ (.Y(_05032_),
    .A(net3740),
    .B(net6898));
 sg13g2_o21ai_1 _14370_ (.B1(_05032_),
    .Y(_00752_),
    .A1(net7332),
    .A2(net6898));
 sg13g2_nand2_1 _14371_ (.Y(_05033_),
    .A(net4093),
    .B(net6898));
 sg13g2_o21ai_1 _14372_ (.B1(_05033_),
    .Y(_00753_),
    .A1(net7529),
    .A2(net6898));
 sg13g2_nand2_1 _14373_ (.Y(_05034_),
    .A(net3451),
    .B(net6898));
 sg13g2_o21ai_1 _14374_ (.B1(_05034_),
    .Y(_00754_),
    .A1(net7682),
    .A2(net6898));
 sg13g2_nand3_1 _14375_ (.B(\top1.event_time[22] ),
    .C(\top1.event_time[24] ),
    .A(\top1.event_time[23] ),
    .Y(_05035_));
 sg13g2_nand4_1 _14376_ (.B(\top1.event_time[22] ),
    .C(\top1.event_time[24] ),
    .A(\top1.event_time[23] ),
    .Y(_05036_),
    .D(\top1.event_time[26] ));
 sg13g2_and4_1 _14377_ (.A(\top1.event_time[19] ),
    .B(_03840_),
    .C(\top1.event_time[20] ),
    .D(\top1.event_time[21] ),
    .X(_05037_));
 sg13g2_nand4_1 _14378_ (.B(\top1.event_time[13] ),
    .C(\top1.event_time[14] ),
    .A(_03837_),
    .Y(_05038_),
    .D(\top1.event_time[15] ));
 sg13g2_nand3_1 _14379_ (.B(\top1.event_time[10] ),
    .C(_04003_),
    .A(\top1.event_time[11] ),
    .Y(_05039_));
 sg13g2_nor4_2 _14380_ (.A(_03835_),
    .B(_03836_),
    .C(_04004_),
    .Y(_05040_),
    .D(_05038_));
 sg13g2_nand3_1 _14381_ (.B(\top1.event_time[16] ),
    .C(_05040_),
    .A(\top1.event_time[17] ),
    .Y(_05041_));
 sg13g2_and4_1 _14382_ (.A(\top1.event_time[17] ),
    .B(\top1.event_time[16] ),
    .C(_05037_),
    .D(_05040_),
    .X(_05042_));
 sg13g2_nand4_1 _14383_ (.B(\top1.event_time[16] ),
    .C(_05037_),
    .A(\top1.event_time[17] ),
    .Y(_05043_),
    .D(_05040_));
 sg13g2_nor2_1 _14384_ (.A(_05036_),
    .B(net6897),
    .Y(_05044_));
 sg13g2_nor3_1 _14385_ (.A(\top1.event_time[25] ),
    .B(_05036_),
    .C(net6897),
    .Y(_05045_));
 sg13g2_nor2_1 _14386_ (.A(\top1.event_time[27] ),
    .B(_05045_),
    .Y(_05046_));
 sg13g2_nand3_1 _14387_ (.B(\top1.event_time[30] ),
    .C(\top1.event_time[31] ),
    .A(\top1.event_time[29] ),
    .Y(_05047_));
 sg13g2_nor3_1 _14388_ (.A(_03842_),
    .B(\top1.event_time[27] ),
    .C(_05047_),
    .Y(_05048_));
 sg13g2_nor4_2 _14389_ (.A(\top1.event_time[25] ),
    .B(_03843_),
    .C(_05036_),
    .Y(_05049_),
    .D(net6897));
 sg13g2_nor3_1 _14390_ (.A(_05046_),
    .B(_05048_),
    .C(_05049_),
    .Y(_00755_));
 sg13g2_nand2_2 _14391_ (.Y(_05050_),
    .A(_05045_),
    .B(_05048_));
 sg13g2_o21ai_1 _14392_ (.B1(_05050_),
    .Y(_05051_),
    .A1(\top1.event_time[28] ),
    .A2(_05049_));
 sg13g2_a21oi_1 _14393_ (.A1(\top1.event_time[28] ),
    .A2(_05049_),
    .Y(_00756_),
    .B1(_05051_));
 sg13g2_a21oi_1 _14394_ (.A1(\top1.event_time[28] ),
    .A2(_05049_),
    .Y(_05052_),
    .B1(\top1.event_time[29] ));
 sg13g2_nand3_1 _14395_ (.B(\top1.event_time[29] ),
    .C(_05049_),
    .A(\top1.event_time[28] ),
    .Y(_05053_));
 sg13g2_nand2_1 _14396_ (.Y(_05054_),
    .A(_05050_),
    .B(_05053_));
 sg13g2_nor2_1 _14397_ (.A(_05052_),
    .B(_05054_),
    .Y(_00757_));
 sg13g2_nand4_1 _14398_ (.B(\top1.event_time[29] ),
    .C(\top1.event_time[30] ),
    .A(\top1.event_time[28] ),
    .Y(_05055_),
    .D(_05049_));
 sg13g2_nand3_1 _14399_ (.B(_05050_),
    .C(_05053_),
    .A(\top1.event_time[30] ),
    .Y(_05056_));
 sg13g2_o21ai_1 _14400_ (.B1(_05056_),
    .Y(_00758_),
    .A1(\top1.event_time[30] ),
    .A2(_05053_));
 sg13g2_o21ai_1 _14401_ (.B1(_05050_),
    .Y(_05057_),
    .A1(_03844_),
    .A2(_05055_));
 sg13g2_a21oi_1 _14402_ (.A1(_03844_),
    .A2(_05055_),
    .Y(_00759_),
    .B1(_05057_));
 sg13g2_nand3_1 _14403_ (.B(net7074),
    .C(net7223),
    .A(net7408),
    .Y(_05058_));
 sg13g2_nand2_1 _14404_ (.Y(_05059_),
    .A(net3169),
    .B(net6459));
 sg13g2_o21ai_1 _14405_ (.B1(_05059_),
    .Y(_00760_),
    .A1(net7358),
    .A2(net6459));
 sg13g2_nand2_1 _14406_ (.Y(_05060_),
    .A(net3038),
    .B(net6458));
 sg13g2_o21ai_1 _14407_ (.B1(_05060_),
    .Y(_00761_),
    .A1(net7555),
    .A2(net6458));
 sg13g2_nand2_1 _14408_ (.Y(_05061_),
    .A(net3841),
    .B(net6458));
 sg13g2_o21ai_1 _14409_ (.B1(_05061_),
    .Y(_00762_),
    .A1(net7715),
    .A2(net6458));
 sg13g2_nand3_1 _14410_ (.B(net7074),
    .C(net7223),
    .A(net7282),
    .Y(_05062_));
 sg13g2_nand2_1 _14411_ (.Y(_05063_),
    .A(net3588),
    .B(net6457));
 sg13g2_o21ai_1 _14412_ (.B1(_05063_),
    .Y(_00763_),
    .A1(net7358),
    .A2(net6456));
 sg13g2_nand2_1 _14413_ (.Y(_05064_),
    .A(net3459),
    .B(net6456));
 sg13g2_o21ai_1 _14414_ (.B1(_05064_),
    .Y(_00764_),
    .A1(net7555),
    .A2(net6456));
 sg13g2_nand2_1 _14415_ (.Y(_05065_),
    .A(net3336),
    .B(net6457));
 sg13g2_o21ai_1 _14416_ (.B1(_05065_),
    .Y(_00765_),
    .A1(net7715),
    .A2(net6456));
 sg13g2_nor3_1 _14417_ (.A(net7284),
    .B(net7267),
    .C(net7200),
    .Y(_05066_));
 sg13g2_nor2_1 _14418_ (.A(net4697),
    .B(net6896),
    .Y(_05067_));
 sg13g2_a21oi_1 _14419_ (.A1(net7310),
    .A2(net6896),
    .Y(_00766_),
    .B1(_05067_));
 sg13g2_nor2_1 _14420_ (.A(net4802),
    .B(net6896),
    .Y(_05068_));
 sg13g2_a21oi_1 _14421_ (.A1(net7509),
    .A2(net6896),
    .Y(_00767_),
    .B1(_05068_));
 sg13g2_nor2_1 _14422_ (.A(net3968),
    .B(net6895),
    .Y(_05069_));
 sg13g2_a21oi_1 _14423_ (.A1(net7666),
    .A2(net6895),
    .Y(_00768_),
    .B1(_05069_));
 sg13g2_nand3_1 _14424_ (.B(net7042),
    .C(net7224),
    .A(net7074),
    .Y(_05070_));
 sg13g2_nand2_1 _14425_ (.Y(_05071_),
    .A(net3922),
    .B(net6455));
 sg13g2_o21ai_1 _14426_ (.B1(_05071_),
    .Y(_00769_),
    .A1(net7357),
    .A2(net6455));
 sg13g2_nand2_1 _14427_ (.Y(_05072_),
    .A(net3049),
    .B(net6454));
 sg13g2_o21ai_1 _14428_ (.B1(_05072_),
    .Y(_00770_),
    .A1(net7552),
    .A2(net6454));
 sg13g2_nand2_1 _14429_ (.Y(_05073_),
    .A(net3416),
    .B(net6454));
 sg13g2_o21ai_1 _14430_ (.B1(_05073_),
    .Y(_00771_),
    .A1(net7713),
    .A2(net6454));
 sg13g2_nand3_1 _14431_ (.B(net7074),
    .C(net7224),
    .A(net7083),
    .Y(_05074_));
 sg13g2_nand2_1 _14432_ (.Y(_05075_),
    .A(net4308),
    .B(net6453));
 sg13g2_o21ai_1 _14433_ (.B1(_05075_),
    .Y(_00772_),
    .A1(net7357),
    .A2(net6453));
 sg13g2_nand2_1 _14434_ (.Y(_05076_),
    .A(net2880),
    .B(net6452));
 sg13g2_o21ai_1 _14435_ (.B1(_05076_),
    .Y(_00773_),
    .A1(net7552),
    .A2(net6452));
 sg13g2_nand2_1 _14436_ (.Y(_05077_),
    .A(net2672),
    .B(net6452));
 sg13g2_o21ai_1 _14437_ (.B1(_05077_),
    .Y(_00774_),
    .A1(net7714),
    .A2(net6452));
 sg13g2_nand3_1 _14438_ (.B(net7074),
    .C(net7224),
    .A(net7102),
    .Y(_05078_));
 sg13g2_nand2_1 _14439_ (.Y(_05079_),
    .A(net4105),
    .B(net6451));
 sg13g2_o21ai_1 _14440_ (.B1(_05079_),
    .Y(_00775_),
    .A1(net7357),
    .A2(net6451));
 sg13g2_nand2_1 _14441_ (.Y(_05080_),
    .A(net3709),
    .B(net6450));
 sg13g2_o21ai_1 _14442_ (.B1(_05080_),
    .Y(_00776_),
    .A1(net7552),
    .A2(net6450));
 sg13g2_nand2_1 _14443_ (.Y(_05081_),
    .A(net4119),
    .B(net6450));
 sg13g2_o21ai_1 _14444_ (.B1(_05081_),
    .Y(_00777_),
    .A1(net7714),
    .A2(net6450));
 sg13g2_nand3_1 _14445_ (.B(net7066),
    .C(net7224),
    .A(net7074),
    .Y(_05082_));
 sg13g2_nand2_1 _14446_ (.Y(_05083_),
    .A(net4070),
    .B(net6449));
 sg13g2_o21ai_1 _14447_ (.B1(_05083_),
    .Y(_00778_),
    .A1(net7357),
    .A2(net6449));
 sg13g2_nand2_1 _14448_ (.Y(_05084_),
    .A(net4148),
    .B(net6448));
 sg13g2_o21ai_1 _14449_ (.B1(_05084_),
    .Y(_00779_),
    .A1(net7552),
    .A2(net6448));
 sg13g2_nand2_1 _14450_ (.Y(_05085_),
    .A(net2891),
    .B(net6448));
 sg13g2_o21ai_1 _14451_ (.B1(_05085_),
    .Y(_00780_),
    .A1(net7714),
    .A2(net6448));
 sg13g2_nand3_1 _14452_ (.B(net7235),
    .C(net7222),
    .A(net7076),
    .Y(_05086_));
 sg13g2_nand2_1 _14453_ (.Y(_05087_),
    .A(net2464),
    .B(net6447));
 sg13g2_o21ai_1 _14454_ (.B1(_05087_),
    .Y(_00781_),
    .A1(net7359),
    .A2(net6447));
 sg13g2_nand2_1 _14455_ (.Y(_05088_),
    .A(net2700),
    .B(net6446));
 sg13g2_o21ai_1 _14456_ (.B1(_05088_),
    .Y(_00782_),
    .A1(net7553),
    .A2(net6446));
 sg13g2_nand2_1 _14457_ (.Y(_05089_),
    .A(net2633),
    .B(net6446));
 sg13g2_o21ai_1 _14458_ (.B1(_05089_),
    .Y(_00783_),
    .A1(net7713),
    .A2(net6446));
 sg13g2_nand3_1 _14459_ (.B(net7076),
    .C(net7222),
    .A(net7265),
    .Y(_05090_));
 sg13g2_nand2_1 _14460_ (.Y(_05091_),
    .A(net3420),
    .B(net6445));
 sg13g2_o21ai_1 _14461_ (.B1(_05091_),
    .Y(_00784_),
    .A1(net7355),
    .A2(net6445));
 sg13g2_nand2_1 _14462_ (.Y(_05092_),
    .A(net3605),
    .B(net6444));
 sg13g2_o21ai_1 _14463_ (.B1(_05092_),
    .Y(_00785_),
    .A1(net7553),
    .A2(net6444));
 sg13g2_nand2_1 _14464_ (.Y(_05093_),
    .A(net3623),
    .B(net6444));
 sg13g2_o21ai_1 _14465_ (.B1(_05093_),
    .Y(_00786_),
    .A1(net7713),
    .A2(net6444));
 sg13g2_nand3_1 _14466_ (.B(net7238),
    .C(net7222),
    .A(net7076),
    .Y(_05094_));
 sg13g2_nand2_1 _14467_ (.Y(_05095_),
    .A(net4128),
    .B(net6443));
 sg13g2_o21ai_1 _14468_ (.B1(_05095_),
    .Y(_00787_),
    .A1(net7355),
    .A2(net6443));
 sg13g2_nand2_1 _14469_ (.Y(_05096_),
    .A(net3266),
    .B(net6442));
 sg13g2_o21ai_1 _14470_ (.B1(_05096_),
    .Y(_00788_),
    .A1(net7553),
    .A2(net6442));
 sg13g2_nand2_1 _14471_ (.Y(_05097_),
    .A(net2835),
    .B(net6442));
 sg13g2_o21ai_1 _14472_ (.B1(_05097_),
    .Y(_00789_),
    .A1(net7713),
    .A2(net6442));
 sg13g2_nand3_1 _14473_ (.B(net7076),
    .C(net7222),
    .A(net7404),
    .Y(_05098_));
 sg13g2_nand2_1 _14474_ (.Y(_05099_),
    .A(net3469),
    .B(net6441));
 sg13g2_o21ai_1 _14475_ (.B1(_05099_),
    .Y(_00790_),
    .A1(net7355),
    .A2(net6440));
 sg13g2_nand2_1 _14476_ (.Y(_05100_),
    .A(net2806),
    .B(net6440));
 sg13g2_o21ai_1 _14477_ (.B1(_05100_),
    .Y(_00791_),
    .A1(net7553),
    .A2(net6440));
 sg13g2_nand2_1 _14478_ (.Y(_05101_),
    .A(net3434),
    .B(net6441));
 sg13g2_o21ai_1 _14479_ (.B1(_05101_),
    .Y(_00792_),
    .A1(net7713),
    .A2(net6440));
 sg13g2_nand3_1 _14480_ (.B(net7231),
    .C(net7221),
    .A(net7248),
    .Y(_05102_));
 sg13g2_nand2_1 _14481_ (.Y(_05103_),
    .A(net3372),
    .B(net6893));
 sg13g2_o21ai_1 _14482_ (.B1(_05103_),
    .Y(_00793_),
    .A1(net7355),
    .A2(net6893));
 sg13g2_nand2_1 _14483_ (.Y(_05104_),
    .A(net2637),
    .B(net6893));
 sg13g2_o21ai_1 _14484_ (.B1(_05104_),
    .Y(_00794_),
    .A1(net7553),
    .A2(net6893));
 sg13g2_nand2_1 _14485_ (.Y(_05105_),
    .A(net2942),
    .B(net6893));
 sg13g2_o21ai_1 _14486_ (.B1(_05105_),
    .Y(_00795_),
    .A1(net7716),
    .A2(net6893));
 sg13g2_nor3_1 _14487_ (.A(_04093_),
    .B(net7268),
    .C(net7201),
    .Y(_05106_));
 sg13g2_nor2_1 _14488_ (.A(net4758),
    .B(net6439),
    .Y(_05107_));
 sg13g2_a21oi_1 _14489_ (.A1(net7313),
    .A2(net6439),
    .Y(_00796_),
    .B1(_05107_));
 sg13g2_nor2_1 _14490_ (.A(net4032),
    .B(net6439),
    .Y(_05108_));
 sg13g2_a21oi_1 _14491_ (.A1(net7510),
    .A2(net6438),
    .Y(_00797_),
    .B1(_05108_));
 sg13g2_nor2_1 _14492_ (.A(net3917),
    .B(net6438),
    .Y(_05109_));
 sg13g2_a21oi_1 _14493_ (.A1(net7669),
    .A2(net6438),
    .Y(_00798_),
    .B1(_05109_));
 sg13g2_nand3_1 _14494_ (.B(net7231),
    .C(net7221),
    .A(net7274),
    .Y(_05110_));
 sg13g2_nand2_1 _14495_ (.Y(_05111_),
    .A(net3244),
    .B(net6891));
 sg13g2_o21ai_1 _14496_ (.B1(_05111_),
    .Y(_00799_),
    .A1(net7355),
    .A2(net6891));
 sg13g2_nand2_1 _14497_ (.Y(_05112_),
    .A(net2856),
    .B(net6891));
 sg13g2_o21ai_1 _14498_ (.B1(_05112_),
    .Y(_00800_),
    .A1(net7553),
    .A2(net6891));
 sg13g2_nand2_1 _14499_ (.Y(_05113_),
    .A(net4309),
    .B(net6891));
 sg13g2_o21ai_1 _14500_ (.B1(_05113_),
    .Y(_00801_),
    .A1(net7713),
    .A2(net6891));
 sg13g2_nand3_1 _14501_ (.B(net7232),
    .C(net7221),
    .A(net7286),
    .Y(_05114_));
 sg13g2_nand2_1 _14502_ (.Y(_05115_),
    .A(net3986),
    .B(net6889));
 sg13g2_o21ai_1 _14503_ (.B1(_05115_),
    .Y(_00802_),
    .A1(net7355),
    .A2(net6889));
 sg13g2_nand2_1 _14504_ (.Y(_05116_),
    .A(net3424),
    .B(net6889));
 sg13g2_o21ai_1 _14505_ (.B1(_05116_),
    .Y(_00803_),
    .A1(net7553),
    .A2(net6889));
 sg13g2_nand2_1 _14506_ (.Y(_05117_),
    .A(net2467),
    .B(net6889));
 sg13g2_o21ai_1 _14507_ (.B1(_05117_),
    .Y(_00804_),
    .A1(net7713),
    .A2(net6889));
 sg13g2_nand3_1 _14508_ (.B(net7233),
    .C(net7219),
    .A(net7279),
    .Y(_05118_));
 sg13g2_nand2_1 _14509_ (.Y(_05119_),
    .A(net3219),
    .B(net6888));
 sg13g2_o21ai_1 _14510_ (.B1(_05119_),
    .Y(_00805_),
    .A1(net7356),
    .A2(net6888));
 sg13g2_nand2_1 _14511_ (.Y(_05120_),
    .A(net3365),
    .B(net6888));
 sg13g2_o21ai_1 _14512_ (.B1(_05120_),
    .Y(_00806_),
    .A1(net7546),
    .A2(net6887));
 sg13g2_nand2_1 _14513_ (.Y(_05121_),
    .A(net3771),
    .B(net6887));
 sg13g2_o21ai_1 _14514_ (.B1(_05121_),
    .Y(_00807_),
    .A1(net7707),
    .A2(net6887));
 sg13g2_nand3_1 _14515_ (.B(net7231),
    .C(net7225),
    .A(net7363),
    .Y(_05122_));
 sg13g2_nand2_1 _14516_ (.Y(_05123_),
    .A(net4066),
    .B(net6886));
 sg13g2_o21ai_1 _14517_ (.B1(_05123_),
    .Y(_00808_),
    .A1(net7356),
    .A2(net6886));
 sg13g2_nand2_1 _14518_ (.Y(_05124_),
    .A(net3979),
    .B(net6886));
 sg13g2_o21ai_1 _14519_ (.B1(_05124_),
    .Y(_00809_),
    .A1(net7546),
    .A2(net6886));
 sg13g2_nand2_1 _14520_ (.Y(_05125_),
    .A(net3776),
    .B(net6885));
 sg13g2_o21ai_1 _14521_ (.B1(_05125_),
    .Y(_00810_),
    .A1(net7706),
    .A2(net6885));
 sg13g2_nand3_1 _14522_ (.B(net7231),
    .C(net7225),
    .A(net7282),
    .Y(_05126_));
 sg13g2_nand2_1 _14523_ (.Y(_05127_),
    .A(net3991),
    .B(net6884));
 sg13g2_o21ai_1 _14524_ (.B1(_05127_),
    .Y(_00811_),
    .A1(net7356),
    .A2(net6884));
 sg13g2_nand2_1 _14525_ (.Y(_05128_),
    .A(net3295),
    .B(net6884));
 sg13g2_o21ai_1 _14526_ (.B1(_05128_),
    .Y(_00812_),
    .A1(net7546),
    .A2(net6884));
 sg13g2_nand2_1 _14527_ (.Y(_05129_),
    .A(net3245),
    .B(net6883));
 sg13g2_o21ai_1 _14528_ (.B1(_05129_),
    .Y(_00813_),
    .A1(net7706),
    .A2(net6883));
 sg13g2_nand3_1 _14529_ (.B(net7231),
    .C(net7225),
    .A(net7408),
    .Y(_05130_));
 sg13g2_nand2_1 _14530_ (.Y(_05131_),
    .A(net3628),
    .B(net6882));
 sg13g2_o21ai_1 _14531_ (.B1(_05131_),
    .Y(_00814_),
    .A1(net7355),
    .A2(net6882));
 sg13g2_nand2_1 _14532_ (.Y(_05132_),
    .A(net3951),
    .B(net6882));
 sg13g2_o21ai_1 _14533_ (.B1(_05132_),
    .Y(_00815_),
    .A1(net7546),
    .A2(net6882));
 sg13g2_nand2_1 _14534_ (.Y(_05133_),
    .A(net3600),
    .B(net6881));
 sg13g2_o21ai_1 _14535_ (.B1(_05133_),
    .Y(_00816_),
    .A1(net7706),
    .A2(net6881));
 sg13g2_nand3_1 _14536_ (.B(net7233),
    .C(net7221),
    .A(net7042),
    .Y(_05134_));
 sg13g2_nand2_1 _14537_ (.Y(_05135_),
    .A(net2719),
    .B(net6437));
 sg13g2_o21ai_1 _14538_ (.B1(_05135_),
    .Y(_00817_),
    .A1(net7356),
    .A2(net6437));
 sg13g2_nand2_1 _14539_ (.Y(_05136_),
    .A(net4262),
    .B(net6437));
 sg13g2_o21ai_1 _14540_ (.B1(_05136_),
    .Y(_00818_),
    .A1(net7552),
    .A2(net6437));
 sg13g2_nand2_1 _14541_ (.Y(_05137_),
    .A(net2697),
    .B(net6436));
 sg13g2_o21ai_1 _14542_ (.B1(_05137_),
    .Y(_00819_),
    .A1(net7710),
    .A2(net6436));
 sg13g2_nand3_1 _14543_ (.B(net7233),
    .C(net7221),
    .A(net7083),
    .Y(_05138_));
 sg13g2_nand2_1 _14544_ (.Y(_05139_),
    .A(net3675),
    .B(net6435));
 sg13g2_o21ai_1 _14545_ (.B1(_05139_),
    .Y(_00820_),
    .A1(net7356),
    .A2(net6435));
 sg13g2_nand2_1 _14546_ (.Y(_05140_),
    .A(net3667),
    .B(net6435));
 sg13g2_o21ai_1 _14547_ (.B1(_05140_),
    .Y(_00821_),
    .A1(net7552),
    .A2(net6435));
 sg13g2_nand2_1 _14548_ (.Y(_05141_),
    .A(net2666),
    .B(net6434));
 sg13g2_o21ai_1 _14549_ (.B1(_05141_),
    .Y(_00822_),
    .A1(net7710),
    .A2(net6434));
 sg13g2_nand3_1 _14550_ (.B(net7233),
    .C(net7221),
    .A(net7102),
    .Y(_05142_));
 sg13g2_nand2_1 _14551_ (.Y(_05143_),
    .A(net3497),
    .B(net6433));
 sg13g2_o21ai_1 _14552_ (.B1(_05143_),
    .Y(_00823_),
    .A1(net7356),
    .A2(net6433));
 sg13g2_nand2_1 _14553_ (.Y(_05144_),
    .A(net3486),
    .B(net6433));
 sg13g2_o21ai_1 _14554_ (.B1(_05144_),
    .Y(_00824_),
    .A1(net7552),
    .A2(net6433));
 sg13g2_nand2_1 _14555_ (.Y(_05145_),
    .A(net2804),
    .B(net6432));
 sg13g2_o21ai_1 _14556_ (.B1(_05145_),
    .Y(_00825_),
    .A1(net7710),
    .A2(net6432));
 sg13g2_nor3_1 _14557_ (.A(_04065_),
    .B(net7268),
    .C(net7200),
    .Y(_05146_));
 sg13g2_nor2_1 _14558_ (.A(net4315),
    .B(net6431),
    .Y(_05147_));
 sg13g2_a21oi_1 _14559_ (.A1(net7313),
    .A2(net6431),
    .Y(_00826_),
    .B1(_05147_));
 sg13g2_nor2_1 _14560_ (.A(net4558),
    .B(net6430),
    .Y(_05148_));
 sg13g2_a21oi_1 _14561_ (.A1(net7510),
    .A2(net6431),
    .Y(_00827_),
    .B1(_05148_));
 sg13g2_nor2_1 _14562_ (.A(net4147),
    .B(net6430),
    .Y(_05149_));
 sg13g2_a21oi_1 _14563_ (.A1(net7669),
    .A2(net6430),
    .Y(_00828_),
    .B1(_05149_));
 sg13g2_nand3_1 _14564_ (.B(net7232),
    .C(net7218),
    .A(net7235),
    .Y(_05150_));
 sg13g2_nand2_1 _14565_ (.Y(_05151_),
    .A(net3725),
    .B(net6879));
 sg13g2_o21ai_1 _14566_ (.B1(_05151_),
    .Y(_00829_),
    .A1(net7349),
    .A2(net6879));
 sg13g2_nand2_1 _14567_ (.Y(_05152_),
    .A(net2890),
    .B(net6879));
 sg13g2_o21ai_1 _14568_ (.B1(_05152_),
    .Y(_00830_),
    .A1(net7547),
    .A2(net6879));
 sg13g2_nand2_1 _14569_ (.Y(_05153_),
    .A(net3584),
    .B(net6880));
 sg13g2_o21ai_1 _14570_ (.B1(_05153_),
    .Y(_00831_),
    .A1(net7706),
    .A2(net6879));
 sg13g2_nand3_1 _14571_ (.B(net7232),
    .C(net7218),
    .A(net7265),
    .Y(_05154_));
 sg13g2_nand2_1 _14572_ (.Y(_05155_),
    .A(net2963),
    .B(net6877));
 sg13g2_o21ai_1 _14573_ (.B1(_05155_),
    .Y(_00832_),
    .A1(net7349),
    .A2(net6877));
 sg13g2_nand2_1 _14574_ (.Y(_05156_),
    .A(net4024),
    .B(net6877));
 sg13g2_o21ai_1 _14575_ (.B1(_05156_),
    .Y(_00833_),
    .A1(net7547),
    .A2(net6877));
 sg13g2_nand2_1 _14576_ (.Y(_05157_),
    .A(net3560),
    .B(net6877));
 sg13g2_o21ai_1 _14577_ (.B1(_05157_),
    .Y(_00834_),
    .A1(net7706),
    .A2(net6877));
 sg13g2_nand3_1 _14578_ (.B(net7231),
    .C(net7218),
    .A(net7238),
    .Y(_05158_));
 sg13g2_nand2_1 _14579_ (.Y(_05159_),
    .A(net2830),
    .B(net6875));
 sg13g2_o21ai_1 _14580_ (.B1(_05159_),
    .Y(_00835_),
    .A1(net7349),
    .A2(net6875));
 sg13g2_nand2_1 _14581_ (.Y(_05160_),
    .A(net2594),
    .B(net6875));
 sg13g2_o21ai_1 _14582_ (.B1(_05160_),
    .Y(_00836_),
    .A1(net7547),
    .A2(net6875));
 sg13g2_nand2_1 _14583_ (.Y(_05161_),
    .A(net3524),
    .B(net6875));
 sg13g2_o21ai_1 _14584_ (.B1(_05161_),
    .Y(_00837_),
    .A1(net7706),
    .A2(net6875));
 sg13g2_nand3_1 _14585_ (.B(net7231),
    .C(net7221),
    .A(net7278),
    .Y(_05162_));
 sg13g2_nand2_1 _14586_ (.Y(_05163_),
    .A(net2586),
    .B(net6873));
 sg13g2_o21ai_1 _14587_ (.B1(_05163_),
    .Y(_00838_),
    .A1(net7355),
    .A2(net6873));
 sg13g2_nand2_1 _14588_ (.Y(_05164_),
    .A(net3383),
    .B(net6873));
 sg13g2_o21ai_1 _14589_ (.B1(_05164_),
    .Y(_00839_),
    .A1(net7553),
    .A2(net6873));
 sg13g2_nand2_1 _14590_ (.Y(_05165_),
    .A(net3101),
    .B(net6873));
 sg13g2_o21ai_1 _14591_ (.B1(_05165_),
    .Y(_00840_),
    .A1(net7713),
    .A2(net6873));
 sg13g2_nand3_1 _14592_ (.B(net7281),
    .C(net7204),
    .A(net7410),
    .Y(_05166_));
 sg13g2_nand2_1 _14593_ (.Y(_05167_),
    .A(net3251),
    .B(net6871));
 sg13g2_o21ai_1 _14594_ (.B1(_05167_),
    .Y(_00841_),
    .A1(net7308),
    .A2(net6871));
 sg13g2_nand2_1 _14595_ (.Y(_05168_),
    .A(net2691),
    .B(net6872));
 sg13g2_o21ai_1 _14596_ (.B1(_05168_),
    .Y(_00842_),
    .A1(net7506),
    .A2(net6872));
 sg13g2_nand2_1 _14597_ (.Y(_05169_),
    .A(net3975),
    .B(net6871));
 sg13g2_o21ai_1 _14598_ (.B1(_05169_),
    .Y(_00843_),
    .A1(net7665),
    .A2(net6871));
 sg13g2_nand3_1 _14599_ (.B(net7361),
    .C(net7205),
    .A(net7412),
    .Y(_05170_));
 sg13g2_nand2_1 _14600_ (.Y(_05171_),
    .A(net4252),
    .B(net6869));
 sg13g2_o21ai_1 _14601_ (.B1(_05171_),
    .Y(_00844_),
    .A1(net7308),
    .A2(net6869));
 sg13g2_nand2_1 _14602_ (.Y(_05172_),
    .A(net4224),
    .B(net6870));
 sg13g2_o21ai_1 _14603_ (.B1(_05172_),
    .Y(_00845_),
    .A1(net7507),
    .A2(net6870));
 sg13g2_nand2_1 _14604_ (.Y(_05173_),
    .A(net3067),
    .B(net6869));
 sg13g2_o21ai_1 _14605_ (.B1(_05173_),
    .Y(_00846_),
    .A1(net7665),
    .A2(net6869));
 sg13g2_nand3_1 _14606_ (.B(net7231),
    .C(net7218),
    .A(net7404),
    .Y(_05174_));
 sg13g2_nand2_1 _14607_ (.Y(_05175_),
    .A(net3638),
    .B(net6867));
 sg13g2_o21ai_1 _14608_ (.B1(_05175_),
    .Y(_00847_),
    .A1(net7349),
    .A2(net6867));
 sg13g2_nand2_1 _14609_ (.Y(_05176_),
    .A(net4199),
    .B(net6867));
 sg13g2_o21ai_1 _14610_ (.B1(_05176_),
    .Y(_00848_),
    .A1(net7547),
    .A2(net6867));
 sg13g2_nand2_1 _14611_ (.Y(_05177_),
    .A(net2777),
    .B(net6867));
 sg13g2_o21ai_1 _14612_ (.B1(_05177_),
    .Y(_00849_),
    .A1(net7706),
    .A2(net6867));
 sg13g2_nor3_1 _14613_ (.A(net7245),
    .B(net7048),
    .C(net7192),
    .Y(_05178_));
 sg13g2_nor2_1 _14614_ (.A(net3647),
    .B(net6429),
    .Y(_05179_));
 sg13g2_a21oi_1 _14615_ (.A1(net7287),
    .A2(net6429),
    .Y(_00850_),
    .B1(_05179_));
 sg13g2_nor2_1 _14616_ (.A(net4500),
    .B(net6429),
    .Y(_05180_));
 sg13g2_a21oi_1 _14617_ (.A1(net7489),
    .A2(net6428),
    .Y(_00851_),
    .B1(_05180_));
 sg13g2_nor2_1 _14618_ (.A(net4786),
    .B(net6428),
    .Y(_05181_));
 sg13g2_a21oi_1 _14619_ (.A1(net7646),
    .A2(net6429),
    .Y(_00852_),
    .B1(_05181_));
 sg13g2_nor3_1 _14620_ (.A(net7275),
    .B(net7048),
    .C(net7193),
    .Y(_05182_));
 sg13g2_nor2_1 _14621_ (.A(net4021),
    .B(net6427),
    .Y(_05183_));
 sg13g2_a21oi_1 _14622_ (.A1(net7287),
    .A2(net6427),
    .Y(_00853_),
    .B1(_05183_));
 sg13g2_nor2_1 _14623_ (.A(net4261),
    .B(net6427),
    .Y(_05184_));
 sg13g2_a21oi_1 _14624_ (.A1(net7489),
    .A2(net6426),
    .Y(_00854_),
    .B1(_05184_));
 sg13g2_nor2_1 _14625_ (.A(net4005),
    .B(net6426),
    .Y(_05185_));
 sg13g2_a21oi_1 _14626_ (.A1(net7646),
    .A2(net6427),
    .Y(_00855_),
    .B1(_05185_));
 sg13g2_nand3_1 _14627_ (.B(net7280),
    .C(net7204),
    .A(net7410),
    .Y(_05186_));
 sg13g2_nand2_1 _14628_ (.Y(_05187_),
    .A(net3576),
    .B(net6865));
 sg13g2_o21ai_1 _14629_ (.B1(_05187_),
    .Y(_00856_),
    .A1(net7308),
    .A2(net6865));
 sg13g2_nand2_1 _14630_ (.Y(_05188_),
    .A(net3146),
    .B(net6866));
 sg13g2_o21ai_1 _14631_ (.B1(_05188_),
    .Y(_00857_),
    .A1(net7508),
    .A2(net6866));
 sg13g2_nand2_1 _14632_ (.Y(_05189_),
    .A(net3910),
    .B(net6865));
 sg13g2_o21ai_1 _14633_ (.B1(_05189_),
    .Y(_00858_),
    .A1(net7665),
    .A2(net6865));
 sg13g2_nand3_1 _14634_ (.B(net7233),
    .C(net7221),
    .A(net7066),
    .Y(_05190_));
 sg13g2_nand2_1 _14635_ (.Y(_05191_),
    .A(net3473),
    .B(net6425));
 sg13g2_o21ai_1 _14636_ (.B1(_05191_),
    .Y(_00859_),
    .A1(net7356),
    .A2(net6425));
 sg13g2_nand2_1 _14637_ (.Y(_05192_),
    .A(net3232),
    .B(net6425));
 sg13g2_o21ai_1 _14638_ (.B1(_05192_),
    .Y(_00860_),
    .A1(net7552),
    .A2(net6425));
 sg13g2_nand2_1 _14639_ (.Y(_05193_),
    .A(net2774),
    .B(net6424));
 sg13g2_o21ai_1 _14640_ (.B1(_05193_),
    .Y(_00861_),
    .A1(net7710),
    .A2(net6424));
 sg13g2_nor3_1 _14641_ (.A(net7271),
    .B(net7048),
    .C(net7193),
    .Y(_05194_));
 sg13g2_nor2_1 _14642_ (.A(net4380),
    .B(net6423),
    .Y(_05195_));
 sg13g2_a21oi_1 _14643_ (.A1(net7287),
    .A2(net6423),
    .Y(_00862_),
    .B1(_05195_));
 sg13g2_nor2_1 _14644_ (.A(net4477),
    .B(net6423),
    .Y(_05196_));
 sg13g2_a21oi_1 _14645_ (.A1(net7489),
    .A2(net6422),
    .Y(_00863_),
    .B1(_05196_));
 sg13g2_nor2_1 _14646_ (.A(net4710),
    .B(net6422),
    .Y(_05197_));
 sg13g2_a21oi_1 _14647_ (.A1(net7646),
    .A2(net6423),
    .Y(_00864_),
    .B1(_05197_));
 sg13g2_nand3_1 _14648_ (.B(net7285),
    .C(net7204),
    .A(net7410),
    .Y(_05198_));
 sg13g2_nand2_1 _14649_ (.Y(_05199_),
    .A(net3792),
    .B(net6864));
 sg13g2_o21ai_1 _14650_ (.B1(_05199_),
    .Y(_00865_),
    .A1(net7312),
    .A2(net6864));
 sg13g2_nand2_1 _14651_ (.Y(_05200_),
    .A(net4111),
    .B(net6864));
 sg13g2_o21ai_1 _14652_ (.B1(_05200_),
    .Y(_00866_),
    .A1(net7506),
    .A2(net6863));
 sg13g2_nand2_1 _14653_ (.Y(_05201_),
    .A(net2644),
    .B(net6863));
 sg13g2_o21ai_1 _14654_ (.B1(_05201_),
    .Y(_00867_),
    .A1(net7665),
    .A2(net6863));
 sg13g2_nor3_1 _14655_ (.A(net7284),
    .B(net7049),
    .C(net7193),
    .Y(_05202_));
 sg13g2_nor2_1 _14656_ (.A(net4187),
    .B(net6421),
    .Y(_05203_));
 sg13g2_a21oi_1 _14657_ (.A1(net7287),
    .A2(net6421),
    .Y(_00868_),
    .B1(_05203_));
 sg13g2_nor2_1 _14658_ (.A(net4447),
    .B(net6421),
    .Y(_05204_));
 sg13g2_a21oi_1 _14659_ (.A1(net7488),
    .A2(net6420),
    .Y(_00869_),
    .B1(_05204_));
 sg13g2_nor2_1 _14660_ (.A(net4682),
    .B(net6420),
    .Y(_05205_));
 sg13g2_a21oi_1 _14661_ (.A1(net7645),
    .A2(net6421),
    .Y(_00870_),
    .B1(_05205_));
 sg13g2_nor3_1 _14662_ (.A(net7107),
    .B(net7051),
    .C(net7199),
    .Y(_05206_));
 sg13g2_nor2_1 _14663_ (.A(net4431),
    .B(net6418),
    .Y(_05207_));
 sg13g2_a21oi_1 _14664_ (.A1(net7290),
    .A2(net6418),
    .Y(_00871_),
    .B1(_05207_));
 sg13g2_nor2_1 _14665_ (.A(net4660),
    .B(net6419),
    .Y(_05208_));
 sg13g2_a21oi_1 _14666_ (.A1(net7493),
    .A2(net6419),
    .Y(_00872_),
    .B1(_05208_));
 sg13g2_nor2_1 _14667_ (.A(net4183),
    .B(net6418),
    .Y(_05209_));
 sg13g2_a21oi_1 _14668_ (.A1(net7648),
    .A2(net6418),
    .Y(_00873_),
    .B1(_05209_));
 sg13g2_nand3_1 _14669_ (.B(net7273),
    .C(net7204),
    .A(net7410),
    .Y(_05210_));
 sg13g2_nand2_1 _14670_ (.Y(_05211_),
    .A(net3565),
    .B(net6862));
 sg13g2_o21ai_1 _14671_ (.B1(_05211_),
    .Y(_00874_),
    .A1(net7312),
    .A2(net6862));
 sg13g2_nand2_1 _14672_ (.Y(_05212_),
    .A(net3431),
    .B(net6861));
 sg13g2_o21ai_1 _14673_ (.B1(_05212_),
    .Y(_00875_),
    .A1(net7506),
    .A2(net6861));
 sg13g2_nand2_1 _14674_ (.Y(_05213_),
    .A(net3468),
    .B(net6862));
 sg13g2_o21ai_1 _14675_ (.B1(_05213_),
    .Y(_00876_),
    .A1(net7665),
    .A2(net6862));
 sg13g2_nor3_1 _14676_ (.A(_04065_),
    .B(net7052),
    .C(net7197),
    .Y(_05214_));
 sg13g2_nor2_1 _14677_ (.A(net3884),
    .B(net6417),
    .Y(_05215_));
 sg13g2_a21oi_1 _14678_ (.A1(net7290),
    .A2(net6416),
    .Y(_00877_),
    .B1(_05215_));
 sg13g2_nor2_1 _14679_ (.A(net4213),
    .B(net6417),
    .Y(_05216_));
 sg13g2_a21oi_1 _14680_ (.A1(net7493),
    .A2(net6417),
    .Y(_00878_),
    .B1(_05216_));
 sg13g2_nor2_1 _14681_ (.A(net3944),
    .B(net6416),
    .Y(_05217_));
 sg13g2_a21oi_1 _14682_ (.A1(net7648),
    .A2(net6416),
    .Y(_00879_),
    .B1(_05217_));
 sg13g2_nor3_1 _14683_ (.A(_04087_),
    .B(net7268),
    .C(net7200),
    .Y(_05218_));
 sg13g2_nor2_1 _14684_ (.A(net4698),
    .B(net6415),
    .Y(_05219_));
 sg13g2_a21oi_1 _14685_ (.A1(net7313),
    .A2(net6415),
    .Y(_00880_),
    .B1(_05219_));
 sg13g2_nor2_1 _14686_ (.A(net4649),
    .B(net6414),
    .Y(_05220_));
 sg13g2_a21oi_1 _14687_ (.A1(net7510),
    .A2(net6415),
    .Y(_00881_),
    .B1(_05220_));
 sg13g2_nor2_1 _14688_ (.A(net4200),
    .B(net6414),
    .Y(_05221_));
 sg13g2_a21oi_1 _14689_ (.A1(net7669),
    .A2(net6414),
    .Y(_00882_),
    .B1(_05221_));
 sg13g2_nand3_1 _14690_ (.B(net7277),
    .C(net7204),
    .A(net7410),
    .Y(_05222_));
 sg13g2_nand2_1 _14691_ (.Y(_05223_),
    .A(net3033),
    .B(net6860));
 sg13g2_o21ai_1 _14692_ (.B1(_05223_),
    .Y(_00883_),
    .A1(net7312),
    .A2(net6860));
 sg13g2_nand2_1 _14693_ (.Y(_05224_),
    .A(net2571),
    .B(net6859));
 sg13g2_o21ai_1 _14694_ (.B1(_05224_),
    .Y(_00884_),
    .A1(net7506),
    .A2(net6859));
 sg13g2_nand2_1 _14695_ (.Y(_05225_),
    .A(net2589),
    .B(net6860));
 sg13g2_o21ai_1 _14696_ (.B1(_05225_),
    .Y(_00885_),
    .A1(net7679),
    .A2(net6860));
 sg13g2_nor3_1 _14697_ (.A(_04087_),
    .B(net7051),
    .C(net7197),
    .Y(_05226_));
 sg13g2_nor2_1 _14698_ (.A(net4065),
    .B(net6412),
    .Y(_05227_));
 sg13g2_a21oi_1 _14699_ (.A1(net7290),
    .A2(net6412),
    .Y(_00886_),
    .B1(_05227_));
 sg13g2_nor2_1 _14700_ (.A(net4588),
    .B(net6413),
    .Y(_05228_));
 sg13g2_a21oi_1 _14701_ (.A1(net7494),
    .A2(net6413),
    .Y(_00887_),
    .B1(_05228_));
 sg13g2_nor2_1 _14702_ (.A(net3941),
    .B(net6412),
    .Y(_05229_));
 sg13g2_a21oi_1 _14703_ (.A1(net7648),
    .A2(net6412),
    .Y(_00888_),
    .B1(_05229_));
 sg13g2_nand3_1 _14704_ (.B(_04240_),
    .C(net7205),
    .A(net7406),
    .Y(_05230_));
 sg13g2_nand2_1 _14705_ (.Y(_05231_),
    .A(net3396),
    .B(net6410));
 sg13g2_o21ai_1 _14706_ (.B1(_05231_),
    .Y(_00889_),
    .A1(net7290),
    .A2(net6410));
 sg13g2_nand2_1 _14707_ (.Y(_05232_),
    .A(net2583),
    .B(net6411));
 sg13g2_o21ai_1 _14708_ (.B1(_05232_),
    .Y(_00890_),
    .A1(net7493),
    .A2(net6411));
 sg13g2_nand2_1 _14709_ (.Y(_05233_),
    .A(net2948),
    .B(net6410));
 sg13g2_o21ai_1 _14710_ (.B1(_05233_),
    .Y(_00891_),
    .A1(net7648),
    .A2(net6410));
 sg13g2_nor3_1 _14711_ (.A(net7050),
    .B(net7234),
    .C(net7193),
    .Y(_05234_));
 sg13g2_nor2_1 _14712_ (.A(net4061),
    .B(net6409),
    .Y(_05235_));
 sg13g2_a21oi_1 _14713_ (.A1(net7290),
    .A2(net6409),
    .Y(_00892_),
    .B1(_05235_));
 sg13g2_nor2_1 _14714_ (.A(net4155),
    .B(net6408),
    .Y(_05236_));
 sg13g2_a21oi_1 _14715_ (.A1(net7494),
    .A2(net6408),
    .Y(_00893_),
    .B1(_05236_));
 sg13g2_nor2_1 _14716_ (.A(net4745),
    .B(net6409),
    .Y(_05237_));
 sg13g2_a21oi_1 _14717_ (.A1(net7648),
    .A2(net6409),
    .Y(_00894_),
    .B1(_05237_));
 sg13g2_nand3_1 _14718_ (.B(net7247),
    .C(net7204),
    .A(net7410),
    .Y(_05238_));
 sg13g2_nand2_1 _14719_ (.Y(_05239_),
    .A(net3684),
    .B(net6858));
 sg13g2_o21ai_1 _14720_ (.B1(_05239_),
    .Y(_00895_),
    .A1(net7312),
    .A2(net6858));
 sg13g2_nand2_1 _14721_ (.Y(_05240_),
    .A(net2964),
    .B(net6857));
 sg13g2_o21ai_1 _14722_ (.B1(_05240_),
    .Y(_00896_),
    .A1(net7506),
    .A2(net6857));
 sg13g2_nand2_1 _14723_ (.Y(_05241_),
    .A(net2940),
    .B(net6858));
 sg13g2_o21ai_1 _14724_ (.B1(_05241_),
    .Y(_00897_),
    .A1(net7665),
    .A2(net6858));
 sg13g2_nand3_1 _14725_ (.B(net7258),
    .C(net7214),
    .A(net7404),
    .Y(_05242_));
 sg13g2_nand2_1 _14726_ (.Y(_05243_),
    .A(net3178),
    .B(net6855));
 sg13g2_o21ai_1 _14727_ (.B1(_05243_),
    .Y(_00898_),
    .A1(net7329),
    .A2(net6855));
 sg13g2_nand2_1 _14728_ (.Y(_05244_),
    .A(net4462),
    .B(net6855));
 sg13g2_o21ai_1 _14729_ (.B1(_05244_),
    .Y(_00899_),
    .A1(net7528),
    .A2(net6855));
 sg13g2_nand2_1 _14730_ (.Y(_05245_),
    .A(net3007),
    .B(net6856));
 sg13g2_o21ai_1 _14731_ (.B1(_05245_),
    .Y(_00900_),
    .A1(net7687),
    .A2(net6856));
 sg13g2_nand3_1 _14732_ (.B(net7238),
    .C(net7214),
    .A(net7258),
    .Y(_05246_));
 sg13g2_nand2_1 _14733_ (.Y(_05247_),
    .A(net2710),
    .B(net6853));
 sg13g2_o21ai_1 _14734_ (.B1(_05247_),
    .Y(_00901_),
    .A1(net7329),
    .A2(net6853));
 sg13g2_nand2_1 _14735_ (.Y(_05248_),
    .A(net4403),
    .B(net6853));
 sg13g2_o21ai_1 _14736_ (.B1(_05248_),
    .Y(_00902_),
    .A1(net7528),
    .A2(net6853));
 sg13g2_nand2_1 _14737_ (.Y(_05249_),
    .A(net3201),
    .B(net6854));
 sg13g2_o21ai_1 _14738_ (.B1(_05249_),
    .Y(_00903_),
    .A1(net7687),
    .A2(net6854));
 sg13g2_nand3_1 _14739_ (.B(net7241),
    .C(net7212),
    .A(net7273),
    .Y(_05250_));
 sg13g2_nand2_1 _14740_ (.Y(_05251_),
    .A(net3495),
    .B(net6852));
 sg13g2_o21ai_1 _14741_ (.B1(_05251_),
    .Y(_00904_),
    .A1(net7333),
    .A2(net6851));
 sg13g2_nand2_1 _14742_ (.Y(_05252_),
    .A(net2825),
    .B(net6852));
 sg13g2_o21ai_1 _14743_ (.B1(_05252_),
    .Y(_00905_),
    .A1(net7533),
    .A2(net6851));
 sg13g2_nand2_1 _14744_ (.Y(_05253_),
    .A(net2539),
    .B(net6852));
 sg13g2_o21ai_1 _14745_ (.B1(_05253_),
    .Y(_00906_),
    .A1(net7689),
    .A2(net6852));
 sg13g2_nor3_1 _14746_ (.A(net7402),
    .B(net7052),
    .C(net7192),
    .Y(_05254_));
 sg13g2_nor2_1 _14747_ (.A(net4398),
    .B(net6406),
    .Y(_05255_));
 sg13g2_a21oi_1 _14748_ (.A1(net7289),
    .A2(net6406),
    .Y(_00907_),
    .B1(_05255_));
 sg13g2_nor2_1 _14749_ (.A(net4217),
    .B(net6406),
    .Y(_05256_));
 sg13g2_a21oi_1 _14750_ (.A1(net7490),
    .A2(net6406),
    .Y(_00908_),
    .B1(_05256_));
 sg13g2_nor2_1 _14751_ (.A(net4687),
    .B(net6407),
    .Y(_05257_));
 sg13g2_a21oi_1 _14752_ (.A1(net7647),
    .A2(net6407),
    .Y(_00909_),
    .B1(_05257_));
 sg13g2_nand3_1 _14753_ (.B(net7085),
    .C(net7203),
    .A(net7096),
    .Y(_05258_));
 sg13g2_nand2_1 _14754_ (.Y(_05259_),
    .A(net2493),
    .B(net6405));
 sg13g2_o21ai_1 _14755_ (.B1(_05259_),
    .Y(_00910_),
    .A1(net7307),
    .A2(net6405));
 sg13g2_nand2_1 _14756_ (.Y(_05260_),
    .A(net3800),
    .B(net6404));
 sg13g2_o21ai_1 _14757_ (.B1(_05260_),
    .Y(_00911_),
    .A1(net7504),
    .A2(net6404));
 sg13g2_nand2_1 _14758_ (.Y(_05261_),
    .A(net3187),
    .B(net6404));
 sg13g2_o21ai_1 _14759_ (.B1(_05261_),
    .Y(_00912_),
    .A1(net7664),
    .A2(net6404));
 sg13g2_nand3_1 _14760_ (.B(net7235),
    .C(net7214),
    .A(net7258),
    .Y(_05262_));
 sg13g2_nand2_1 _14761_ (.Y(_05263_),
    .A(net2839),
    .B(net6850));
 sg13g2_o21ai_1 _14762_ (.B1(_05263_),
    .Y(_00913_),
    .A1(net7329),
    .A2(net6850));
 sg13g2_nand2_1 _14763_ (.Y(_05264_),
    .A(net4109),
    .B(net6849));
 sg13g2_o21ai_1 _14764_ (.B1(_05264_),
    .Y(_00914_),
    .A1(net7528),
    .A2(net6849));
 sg13g2_nand2_1 _14765_ (.Y(_05265_),
    .A(net3432),
    .B(net6849));
 sg13g2_o21ai_1 _14766_ (.B1(_05265_),
    .Y(_00915_),
    .A1(net7687),
    .A2(net6849));
 sg13g2_nand3_1 _14767_ (.B(net7066),
    .C(net7215),
    .A(net7258),
    .Y(_05266_));
 sg13g2_nand2_1 _14768_ (.Y(_05267_),
    .A(net3689),
    .B(net6403));
 sg13g2_o21ai_1 _14769_ (.B1(_05267_),
    .Y(_00916_),
    .A1(net7327),
    .A2(net6403));
 sg13g2_nand2_1 _14770_ (.Y(_05268_),
    .A(net3088),
    .B(net6402));
 sg13g2_o21ai_1 _14771_ (.B1(_05268_),
    .Y(_00917_),
    .A1(net7524),
    .A2(net6402));
 sg13g2_nand2_1 _14772_ (.Y(_05269_),
    .A(net4058),
    .B(net6402));
 sg13g2_o21ai_1 _14773_ (.B1(_05269_),
    .Y(_00918_),
    .A1(net7681),
    .A2(net6402));
 sg13g2_nand3_1 _14774_ (.B(net7258),
    .C(net7215),
    .A(net7102),
    .Y(_05270_));
 sg13g2_nand2_1 _14775_ (.Y(_05271_),
    .A(net3276),
    .B(net6401));
 sg13g2_o21ai_1 _14776_ (.B1(_05271_),
    .Y(_00919_),
    .A1(net7327),
    .A2(net6400));
 sg13g2_nand2_1 _14777_ (.Y(_05272_),
    .A(net2762),
    .B(net6400));
 sg13g2_o21ai_1 _14778_ (.B1(_05272_),
    .Y(_00920_),
    .A1(net7524),
    .A2(net6400));
 sg13g2_nand2_1 _14779_ (.Y(_05273_),
    .A(net4651),
    .B(net6400));
 sg13g2_o21ai_1 _14780_ (.B1(_05273_),
    .Y(_00921_),
    .A1(net7681),
    .A2(net6400));
 sg13g2_nor3_1 _14781_ (.A(_04152_),
    .B(net7050),
    .C(net7192),
    .Y(_05274_));
 sg13g2_nor2_1 _14782_ (.A(net4246),
    .B(net6399),
    .Y(_05275_));
 sg13g2_a21oi_1 _14783_ (.A1(net7290),
    .A2(net6399),
    .Y(_00922_),
    .B1(_05275_));
 sg13g2_nor2_1 _14784_ (.A(net4250),
    .B(net6398),
    .Y(_05276_));
 sg13g2_a21oi_1 _14785_ (.A1(net7490),
    .A2(net6398),
    .Y(_00923_),
    .B1(_05276_));
 sg13g2_nor2_1 _14786_ (.A(net4100),
    .B(net6399),
    .Y(_05277_));
 sg13g2_a21oi_1 _14787_ (.A1(net7648),
    .A2(net6399),
    .Y(_00924_),
    .B1(_05277_));
 sg13g2_nand3_1 _14788_ (.B(net7083),
    .C(net7215),
    .A(net7258),
    .Y(_05278_));
 sg13g2_nand2_1 _14789_ (.Y(_05279_),
    .A(net2944),
    .B(net6397));
 sg13g2_o21ai_1 _14790_ (.B1(_05279_),
    .Y(_00925_),
    .A1(net7327),
    .A2(net6397));
 sg13g2_nand2_1 _14791_ (.Y(_05280_),
    .A(net2475),
    .B(net6396));
 sg13g2_o21ai_1 _14792_ (.B1(_05280_),
    .Y(_00926_),
    .A1(net7524),
    .A2(net6396));
 sg13g2_nand2_1 _14793_ (.Y(_05281_),
    .A(net3092),
    .B(net6396));
 sg13g2_o21ai_1 _14794_ (.B1(_05281_),
    .Y(_00927_),
    .A1(net7681),
    .A2(net6396));
 sg13g2_nor3_1 _14795_ (.A(_04101_),
    .B(net7050),
    .C(net7192),
    .Y(_05282_));
 sg13g2_nor2_1 _14796_ (.A(net4594),
    .B(net6395),
    .Y(_05283_));
 sg13g2_a21oi_1 _14797_ (.A1(net7290),
    .A2(net6395),
    .Y(_00928_),
    .B1(_05283_));
 sg13g2_nor2_1 _14798_ (.A(net4630),
    .B(net6394),
    .Y(_05284_));
 sg13g2_a21oi_1 _14799_ (.A1(net7494),
    .A2(net6394),
    .Y(_00929_),
    .B1(_05284_));
 sg13g2_nor2_1 _14800_ (.A(net4324),
    .B(net6395),
    .Y(_05285_));
 sg13g2_a21oi_1 _14801_ (.A1(net7648),
    .A2(net6395),
    .Y(_00930_),
    .B1(_05285_));
 sg13g2_nor3_1 _14802_ (.A(_04184_),
    .B(net7050),
    .C(net7192),
    .Y(_05286_));
 sg13g2_nor2_1 _14803_ (.A(net4116),
    .B(net6393),
    .Y(_05287_));
 sg13g2_a21oi_1 _14804_ (.A1(net7290),
    .A2(net6393),
    .Y(_00931_),
    .B1(_05287_));
 sg13g2_nor2_1 _14805_ (.A(net4619),
    .B(net6392),
    .Y(_05288_));
 sg13g2_a21oi_1 _14806_ (.A1(net7490),
    .A2(net6392),
    .Y(_00932_),
    .B1(_05288_));
 sg13g2_nor2_1 _14807_ (.A(net4501),
    .B(net6393),
    .Y(_05289_));
 sg13g2_a21oi_1 _14808_ (.A1(net7648),
    .A2(net6393),
    .Y(_00933_),
    .B1(_05289_));
 sg13g2_nand3_1 _14809_ (.B(net7042),
    .C(net7215),
    .A(net7258),
    .Y(_05290_));
 sg13g2_nand2_1 _14810_ (.Y(_05291_),
    .A(net2620),
    .B(net6391));
 sg13g2_o21ai_1 _14811_ (.B1(_05291_),
    .Y(_00934_),
    .A1(net7325),
    .A2(net6390));
 sg13g2_nand2_1 _14812_ (.Y(_05292_),
    .A(net2599),
    .B(net6390));
 sg13g2_o21ai_1 _14813_ (.B1(_05292_),
    .Y(_00935_),
    .A1(net7524),
    .A2(net6390));
 sg13g2_nand2_1 _14814_ (.Y(_05293_),
    .A(net3036),
    .B(net6390));
 sg13g2_o21ai_1 _14815_ (.B1(_05293_),
    .Y(_00936_),
    .A1(net7681),
    .A2(net6390));
 sg13g2_nand3_1 _14816_ (.B(net7259),
    .C(net7215),
    .A(net7408),
    .Y(_05294_));
 sg13g2_nand2_1 _14817_ (.Y(_05295_),
    .A(net3405),
    .B(net6847));
 sg13g2_o21ai_1 _14818_ (.B1(_05295_),
    .Y(_00937_),
    .A1(net7327),
    .A2(net6847));
 sg13g2_nand2_1 _14819_ (.Y(_05296_),
    .A(net3077),
    .B(net6847));
 sg13g2_o21ai_1 _14820_ (.B1(_05296_),
    .Y(_00938_),
    .A1(net7526),
    .A2(net6847));
 sg13g2_nand2_1 _14821_ (.Y(_05297_),
    .A(net2461),
    .B(net6848));
 sg13g2_o21ai_1 _14822_ (.B1(_05297_),
    .Y(_00939_),
    .A1(net7684),
    .A2(net6848));
 sg13g2_nand3_1 _14823_ (.B(net7259),
    .C(net7215),
    .A(net7282),
    .Y(_05298_));
 sg13g2_nand2_1 _14824_ (.Y(_05299_),
    .A(net2494),
    .B(net6845));
 sg13g2_o21ai_1 _14825_ (.B1(_05299_),
    .Y(_00940_),
    .A1(net7327),
    .A2(net6845));
 sg13g2_nand2_1 _14826_ (.Y(_05300_),
    .A(net4251),
    .B(net6845));
 sg13g2_o21ai_1 _14827_ (.B1(_05300_),
    .Y(_00941_),
    .A1(net7526),
    .A2(net6845));
 sg13g2_nand2_1 _14828_ (.Y(_05301_),
    .A(net3054),
    .B(net6846));
 sg13g2_o21ai_1 _14829_ (.B1(_05301_),
    .Y(_00942_),
    .A1(net7684),
    .A2(net6846));
 sg13g2_nand3_1 _14830_ (.B(net7259),
    .C(net7215),
    .A(net7362),
    .Y(_05302_));
 sg13g2_nand2_1 _14831_ (.Y(_05303_),
    .A(net3643),
    .B(net6843));
 sg13g2_o21ai_1 _14832_ (.B1(_05303_),
    .Y(_00943_),
    .A1(net7327),
    .A2(net6843));
 sg13g2_nand2_1 _14833_ (.Y(_05304_),
    .A(net4134),
    .B(net6843));
 sg13g2_o21ai_1 _14834_ (.B1(_05304_),
    .Y(_00944_),
    .A1(net7526),
    .A2(net6843));
 sg13g2_nand2_1 _14835_ (.Y(_05305_),
    .A(net3157),
    .B(net6843));
 sg13g2_o21ai_1 _14836_ (.B1(_05305_),
    .Y(_00945_),
    .A1(net7684),
    .A2(net6843));
 sg13g2_nand3_1 _14837_ (.B(net7259),
    .C(net7215),
    .A(net7279),
    .Y(_05306_));
 sg13g2_nand2_1 _14838_ (.Y(_05307_),
    .A(net3282),
    .B(net6841));
 sg13g2_o21ai_1 _14839_ (.B1(_05307_),
    .Y(_00946_),
    .A1(net7327),
    .A2(net6841));
 sg13g2_nand2_1 _14840_ (.Y(_05308_),
    .A(net3577),
    .B(net6841));
 sg13g2_o21ai_1 _14841_ (.B1(_05308_),
    .Y(_00947_),
    .A1(net7526),
    .A2(net6841));
 sg13g2_nand2_1 _14842_ (.Y(_05309_),
    .A(net2455),
    .B(net6841));
 sg13g2_o21ai_1 _14843_ (.B1(_05309_),
    .Y(_00948_),
    .A1(net7684),
    .A2(net6841));
 sg13g2_nand3_1 _14844_ (.B(net7241),
    .C(net7212),
    .A(net7277),
    .Y(_05310_));
 sg13g2_nand2_1 _14845_ (.Y(_05311_),
    .A(net2568),
    .B(net6839));
 sg13g2_o21ai_1 _14846_ (.B1(_05311_),
    .Y(_00949_),
    .A1(net7333),
    .A2(net6839));
 sg13g2_nand2_1 _14847_ (.Y(_05312_),
    .A(net3172),
    .B(net6840));
 sg13g2_o21ai_1 _14848_ (.B1(_05312_),
    .Y(_00950_),
    .A1(net7533),
    .A2(net6839));
 sg13g2_nand2_1 _14849_ (.Y(_05313_),
    .A(net3000),
    .B(net6840));
 sg13g2_o21ai_1 _14850_ (.B1(_05313_),
    .Y(_00951_),
    .A1(net7689),
    .A2(net6840));
 sg13g2_nor3_1 _14851_ (.A(_04079_),
    .B(net7098),
    .C(net7202),
    .Y(_05314_));
 sg13g2_nor2_1 _14852_ (.A(net4552),
    .B(net6388),
    .Y(_05315_));
 sg13g2_a21oi_1 _14853_ (.A1(net7330),
    .A2(net6389),
    .Y(_00952_),
    .B1(_05315_));
 sg13g2_nor2_1 _14854_ (.A(net4283),
    .B(net6388),
    .Y(_05316_));
 sg13g2_a21oi_1 _14855_ (.A1(net7535),
    .A2(net6388),
    .Y(_00953_),
    .B1(_05316_));
 sg13g2_nor2_1 _14856_ (.A(net4689),
    .B(net6388),
    .Y(_05317_));
 sg13g2_a21oi_1 _14857_ (.A1(net7688),
    .A2(net6388),
    .Y(_00954_),
    .B1(_05317_));
 sg13g2_nand3_1 _14858_ (.B(net7260),
    .C(net7213),
    .A(net7273),
    .Y(_05318_));
 sg13g2_nand2_1 _14859_ (.Y(_05319_),
    .A(net2928),
    .B(net6837));
 sg13g2_o21ai_1 _14860_ (.B1(_05319_),
    .Y(_00955_),
    .A1(net7329),
    .A2(net6837));
 sg13g2_nand2_1 _14861_ (.Y(_05320_),
    .A(net3206),
    .B(net6837));
 sg13g2_o21ai_1 _14862_ (.B1(_05320_),
    .Y(_00956_),
    .A1(net7529),
    .A2(net6837));
 sg13g2_nand2_1 _14863_ (.Y(_05321_),
    .A(net3845),
    .B(net6838));
 sg13g2_o21ai_1 _14864_ (.B1(_05321_),
    .Y(_00957_),
    .A1(net7687),
    .A2(net6838));
 sg13g2_nand3_1 _14865_ (.B(net7260),
    .C(net7213),
    .A(net7277),
    .Y(_05322_));
 sg13g2_nand2_1 _14866_ (.Y(_05323_),
    .A(net3694),
    .B(net6835));
 sg13g2_o21ai_1 _14867_ (.B1(_05323_),
    .Y(_00958_),
    .A1(net7329),
    .A2(net6835));
 sg13g2_nand2_1 _14868_ (.Y(_05324_),
    .A(net3686),
    .B(net6835));
 sg13g2_o21ai_1 _14869_ (.B1(_05324_),
    .Y(_00959_),
    .A1(net7529),
    .A2(net6835));
 sg13g2_nand2_1 _14870_ (.Y(_05325_),
    .A(net4318),
    .B(net6836));
 sg13g2_o21ai_1 _14871_ (.B1(_05325_),
    .Y(_00960_),
    .A1(net7687),
    .A2(net6836));
 sg13g2_nand3_1 _14872_ (.B(net7265),
    .C(net7220),
    .A(net7100),
    .Y(_05326_));
 sg13g2_nand2_1 _14873_ (.Y(_05327_),
    .A(net4349),
    .B(net6386));
 sg13g2_o21ai_1 _14874_ (.B1(_05327_),
    .Y(_00961_),
    .A1(net7343),
    .A2(net6386));
 sg13g2_nand2_1 _14875_ (.Y(_05328_),
    .A(net3563),
    .B(net6386));
 sg13g2_o21ai_1 _14876_ (.B1(_05328_),
    .Y(_00962_),
    .A1(net7541),
    .A2(net6386));
 sg13g2_nand2_1 _14877_ (.Y(_05329_),
    .A(net3721),
    .B(net6386));
 sg13g2_o21ai_1 _14878_ (.B1(_05329_),
    .Y(_00963_),
    .A1(net7702),
    .A2(net6386));
 sg13g2_nand3_1 _14879_ (.B(net7247),
    .C(net7214),
    .A(net7260),
    .Y(_05330_));
 sg13g2_nand2_1 _14880_ (.Y(_05331_),
    .A(net2600),
    .B(net6833));
 sg13g2_o21ai_1 _14881_ (.B1(_05331_),
    .Y(_00964_),
    .A1(net7329),
    .A2(net6833));
 sg13g2_nand2_1 _14882_ (.Y(_05332_),
    .A(net3057),
    .B(net6833));
 sg13g2_o21ai_1 _14883_ (.B1(_05332_),
    .Y(_00965_),
    .A1(net7528),
    .A2(net6833));
 sg13g2_nand2_1 _14884_ (.Y(_05333_),
    .A(net3053),
    .B(net6834));
 sg13g2_o21ai_1 _14885_ (.B1(_05333_),
    .Y(_00966_),
    .A1(net7687),
    .A2(net6834));
 sg13g2_nand3_1 _14886_ (.B(net7080),
    .C(net7208),
    .A(net7404),
    .Y(_05334_));
 sg13g2_nand2_1 _14887_ (.Y(_05335_),
    .A(net2654),
    .B(net6384));
 sg13g2_o21ai_1 _14888_ (.B1(_05335_),
    .Y(_00967_),
    .A1(net7324),
    .A2(net6384));
 sg13g2_nand2_1 _14889_ (.Y(_05336_),
    .A(net3269),
    .B(net6384));
 sg13g2_o21ai_1 _14890_ (.B1(_05336_),
    .Y(_00968_),
    .A1(net7523),
    .A2(net6384));
 sg13g2_nand2_1 _14891_ (.Y(_05337_),
    .A(net3892),
    .B(net6385));
 sg13g2_o21ai_1 _14892_ (.B1(_05337_),
    .Y(_00969_),
    .A1(net7680),
    .A2(net6385));
 sg13g2_nand3_1 _14893_ (.B(net7239),
    .C(net7208),
    .A(net7080),
    .Y(_05338_));
 sg13g2_nand2_1 _14894_ (.Y(_05339_),
    .A(net2858),
    .B(net6382));
 sg13g2_o21ai_1 _14895_ (.B1(_05339_),
    .Y(_00970_),
    .A1(net7324),
    .A2(net6382));
 sg13g2_nand2_1 _14896_ (.Y(_05340_),
    .A(net3406),
    .B(net6382));
 sg13g2_o21ai_1 _14897_ (.B1(_05340_),
    .Y(_00971_),
    .A1(net7523),
    .A2(net6382));
 sg13g2_nand2_1 _14898_ (.Y(_05341_),
    .A(net4074),
    .B(net6383));
 sg13g2_o21ai_1 _14899_ (.B1(_05341_),
    .Y(_00972_),
    .A1(net7680),
    .A2(net6383));
 sg13g2_nand3_1 _14900_ (.B(net7080),
    .C(net7208),
    .A(net7266),
    .Y(_05342_));
 sg13g2_nand2_1 _14901_ (.Y(_05343_),
    .A(net3466),
    .B(net6380));
 sg13g2_o21ai_1 _14902_ (.B1(_05343_),
    .Y(_00973_),
    .A1(net7324),
    .A2(net6380));
 sg13g2_nand2_1 _14903_ (.Y(_05344_),
    .A(net3554),
    .B(net6380));
 sg13g2_o21ai_1 _14904_ (.B1(_05344_),
    .Y(_00974_),
    .A1(net7523),
    .A2(net6380));
 sg13g2_nand2_1 _14905_ (.Y(_05345_),
    .A(net2692),
    .B(net6381));
 sg13g2_o21ai_1 _14906_ (.B1(_05345_),
    .Y(_00975_),
    .A1(net7680),
    .A2(net6381));
 sg13g2_nand3_1 _14907_ (.B(net7236),
    .C(net7208),
    .A(net7080),
    .Y(_05346_));
 sg13g2_nand2_1 _14908_ (.Y(_05347_),
    .A(net4159),
    .B(net6378));
 sg13g2_o21ai_1 _14909_ (.B1(_05347_),
    .Y(_00976_),
    .A1(net7324),
    .A2(net6378));
 sg13g2_nand2_1 _14910_ (.Y(_05348_),
    .A(net3573),
    .B(net6378));
 sg13g2_o21ai_1 _14911_ (.B1(_05348_),
    .Y(_00977_),
    .A1(net7523),
    .A2(net6378));
 sg13g2_nand2_1 _14912_ (.Y(_05349_),
    .A(net3490),
    .B(net6379));
 sg13g2_o21ai_1 _14913_ (.B1(_05349_),
    .Y(_00978_),
    .A1(net7680),
    .A2(net6379));
 sg13g2_nand3_1 _14914_ (.B(net7065),
    .C(net7208),
    .A(net7080),
    .Y(_05350_));
 sg13g2_nand2_1 _14915_ (.Y(_05351_),
    .A(net4241),
    .B(net6376));
 sg13g2_o21ai_1 _14916_ (.B1(_05351_),
    .Y(_00979_),
    .A1(net7324),
    .A2(net6376));
 sg13g2_nand2_1 _14917_ (.Y(_05352_),
    .A(net2614),
    .B(net6376));
 sg13g2_o21ai_1 _14918_ (.B1(_05352_),
    .Y(_00980_),
    .A1(net7523),
    .A2(net6376));
 sg13g2_nand2_1 _14919_ (.Y(_05353_),
    .A(net4077),
    .B(net6376));
 sg13g2_o21ai_1 _14920_ (.B1(_05353_),
    .Y(_00981_),
    .A1(net7680),
    .A2(net6376));
 sg13g2_nand3_1 _14921_ (.B(net7080),
    .C(net7208),
    .A(net7102),
    .Y(_05354_));
 sg13g2_nand2_1 _14922_ (.Y(_05355_),
    .A(net3200),
    .B(net6374));
 sg13g2_o21ai_1 _14923_ (.B1(_05355_),
    .Y(_00982_),
    .A1(net7324),
    .A2(net6374));
 sg13g2_nand2_1 _14924_ (.Y(_05356_),
    .A(net3371),
    .B(net6374));
 sg13g2_o21ai_1 _14925_ (.B1(_05356_),
    .Y(_00983_),
    .A1(net7523),
    .A2(net6374));
 sg13g2_nand2_1 _14926_ (.Y(_05357_),
    .A(net4209),
    .B(net6374));
 sg13g2_o21ai_1 _14927_ (.B1(_05357_),
    .Y(_00984_),
    .A1(net7680),
    .A2(net6374));
 sg13g2_nand3_1 _14928_ (.B(net7241),
    .C(net7212),
    .A(net7247),
    .Y(_05358_));
 sg13g2_nand2_1 _14929_ (.Y(_05359_),
    .A(net3877),
    .B(net6832));
 sg13g2_o21ai_1 _14930_ (.B1(_05359_),
    .Y(_00985_),
    .A1(net7333),
    .A2(net6831));
 sg13g2_nand2_1 _14931_ (.Y(_05360_),
    .A(net2977),
    .B(net6831));
 sg13g2_o21ai_1 _14932_ (.B1(_05360_),
    .Y(_00986_),
    .A1(net7533),
    .A2(net6831));
 sg13g2_nand2_1 _14933_ (.Y(_05361_),
    .A(net2498),
    .B(net6832));
 sg13g2_o21ai_1 _14934_ (.B1(_05361_),
    .Y(_00987_),
    .A1(net7689),
    .A2(net6832));
 sg13g2_nand3_1 _14935_ (.B(net7043),
    .C(net7209),
    .A(net7080),
    .Y(_05362_));
 sg13g2_nand2_1 _14936_ (.Y(_05363_),
    .A(net3662),
    .B(net6372));
 sg13g2_o21ai_1 _14937_ (.B1(_05363_),
    .Y(_00988_),
    .A1(net7324),
    .A2(net6372));
 sg13g2_nand2_1 _14938_ (.Y(_05364_),
    .A(net2903),
    .B(net6372));
 sg13g2_o21ai_1 _14939_ (.B1(_05364_),
    .Y(_00989_),
    .A1(net7523),
    .A2(net6372));
 sg13g2_nand2_1 _14940_ (.Y(_05365_),
    .A(net3294),
    .B(net6372));
 sg13g2_o21ai_1 _14941_ (.B1(_05365_),
    .Y(_00990_),
    .A1(net7680),
    .A2(net6372));
 sg13g2_nand3_1 _14942_ (.B(net7081),
    .C(net7209),
    .A(net7407),
    .Y(_05366_));
 sg13g2_nand2_1 _14943_ (.Y(_05367_),
    .A(net3648),
    .B(net6370));
 sg13g2_o21ai_1 _14944_ (.B1(_05367_),
    .Y(_00991_),
    .A1(net7325),
    .A2(net6370));
 sg13g2_nand2_1 _14945_ (.Y(_05368_),
    .A(net3175),
    .B(net6370));
 sg13g2_o21ai_1 _14946_ (.B1(_05368_),
    .Y(_00992_),
    .A1(net7524),
    .A2(net6370));
 sg13g2_nand2_1 _14947_ (.Y(_05369_),
    .A(net3457),
    .B(net6371));
 sg13g2_o21ai_1 _14948_ (.B1(_05369_),
    .Y(_00993_),
    .A1(net7681),
    .A2(net6370));
 sg13g2_nand3_1 _14949_ (.B(net7081),
    .C(net7209),
    .A(net7281),
    .Y(_05370_));
 sg13g2_nand2_1 _14950_ (.Y(_05371_),
    .A(net3685),
    .B(net6368));
 sg13g2_o21ai_1 _14951_ (.B1(_05371_),
    .Y(_00994_),
    .A1(net7325),
    .A2(net6368));
 sg13g2_nand2_1 _14952_ (.Y(_05372_),
    .A(net3162),
    .B(net6368));
 sg13g2_o21ai_1 _14953_ (.B1(_05372_),
    .Y(_00995_),
    .A1(net7524),
    .A2(net6368));
 sg13g2_nand2_1 _14954_ (.Y(_05373_),
    .A(net3788),
    .B(net6368));
 sg13g2_o21ai_1 _14955_ (.B1(_05373_),
    .Y(_00996_),
    .A1(net7681),
    .A2(net6368));
 sg13g2_nor3_1 _14956_ (.A(net7249),
    .B(net7245),
    .C(net7194),
    .Y(_05374_));
 sg13g2_nor2_1 _14957_ (.A(net4840),
    .B(net6829),
    .Y(_05375_));
 sg13g2_a21oi_1 _14958_ (.A1(net7289),
    .A2(net6829),
    .Y(_00997_),
    .B1(_05375_));
 sg13g2_nor2_1 _14959_ (.A(net4289),
    .B(net6830),
    .Y(_05376_));
 sg13g2_a21oi_1 _14960_ (.A1(net7495),
    .A2(net6830),
    .Y(_00998_),
    .B1(_05376_));
 sg13g2_nor2_1 _14961_ (.A(net3731),
    .B(net6830),
    .Y(_05377_));
 sg13g2_a21oi_1 _14962_ (.A1(net7647),
    .A2(net6830),
    .Y(_00999_),
    .B1(_05377_));
 sg13g2_nor2_2 _14963_ (.A(_04056_),
    .B(net7202),
    .Y(_05378_));
 sg13g2_nor2_1 _14964_ (.A(net4236),
    .B(net6366),
    .Y(_05379_));
 sg13g2_a21oi_1 _14965_ (.A1(net7348),
    .A2(net6367),
    .Y(_01000_),
    .B1(_05379_));
 sg13g2_nor2_1 _14966_ (.A(net4539),
    .B(net6366),
    .Y(_05380_));
 sg13g2_a21oi_1 _14967_ (.A1(net7547),
    .A2(net6366),
    .Y(_01001_),
    .B1(_05380_));
 sg13g2_nor2_1 _14968_ (.A(net4073),
    .B(net6367),
    .Y(_05381_));
 sg13g2_a21oi_1 _14969_ (.A1(net7705),
    .A2(net6367),
    .Y(_01002_),
    .B1(_05381_));
 sg13g2_nand3_1 _14970_ (.B(net7238),
    .C(net7219),
    .A(net7117),
    .Y(_05382_));
 sg13g2_nand2_1 _14971_ (.Y(_05383_),
    .A(net3546),
    .B(net6364));
 sg13g2_o21ai_1 _14972_ (.B1(_05383_),
    .Y(_01003_),
    .A1(net7348),
    .A2(net6364));
 sg13g2_nand2_1 _14973_ (.Y(_05384_),
    .A(net3616),
    .B(net6364));
 sg13g2_o21ai_1 _14974_ (.B1(_05384_),
    .Y(_01004_),
    .A1(net7547),
    .A2(net6364));
 sg13g2_nand2_1 _14975_ (.Y(_05385_),
    .A(net3784),
    .B(net6365));
 sg13g2_o21ai_1 _14976_ (.B1(_05385_),
    .Y(_01005_),
    .A1(net7705),
    .A2(net6365));
 sg13g2_nand3_1 _14977_ (.B(net7265),
    .C(net7219),
    .A(net7117),
    .Y(_05386_));
 sg13g2_nand2_1 _14978_ (.Y(_05387_),
    .A(net2665),
    .B(net6362));
 sg13g2_o21ai_1 _14979_ (.B1(_05387_),
    .Y(_01006_),
    .A1(net7348),
    .A2(net6362));
 sg13g2_nand2_1 _14980_ (.Y(_05388_),
    .A(net2908),
    .B(net6362));
 sg13g2_o21ai_1 _14981_ (.B1(_05388_),
    .Y(_01007_),
    .A1(net7547),
    .A2(net6362));
 sg13g2_nand2_1 _14982_ (.Y(_05389_),
    .A(net3267),
    .B(net6363));
 sg13g2_o21ai_1 _14983_ (.B1(_05389_),
    .Y(_01008_),
    .A1(net7705),
    .A2(net6363));
 sg13g2_nand3_1 _14984_ (.B(net7242),
    .C(net7210),
    .A(net7404),
    .Y(_05390_));
 sg13g2_nand2_1 _14985_ (.Y(_05391_),
    .A(net2877),
    .B(net6827));
 sg13g2_o21ai_1 _14986_ (.B1(_05391_),
    .Y(_01009_),
    .A1(net7326),
    .A2(net6827));
 sg13g2_nand2_1 _14987_ (.Y(_05392_),
    .A(net3205),
    .B(net6827));
 sg13g2_o21ai_1 _14988_ (.B1(_05392_),
    .Y(_01010_),
    .A1(net7529),
    .A2(net6827));
 sg13g2_nand2_1 _14989_ (.Y(_05393_),
    .A(net3422),
    .B(net6827));
 sg13g2_o21ai_1 _14990_ (.B1(_05393_),
    .Y(_01011_),
    .A1(net7682),
    .A2(net6827));
 sg13g2_xnor2_1 _14991_ (.Y(_01012_),
    .A(_03836_),
    .B(_04003_));
 sg13g2_o21ai_1 _14992_ (.B1(_03835_),
    .Y(_05394_),
    .A1(_03836_),
    .A2(_04004_));
 sg13g2_and2_1 _14993_ (.A(_05039_),
    .B(_05394_),
    .X(_01013_));
 sg13g2_or2_1 _14994_ (.X(_05395_),
    .B(_05039_),
    .A(_03837_));
 sg13g2_nand2_1 _14995_ (.Y(_05396_),
    .A(_05038_),
    .B(_05395_));
 sg13g2_a21oi_1 _14996_ (.A1(_03837_),
    .A2(_05039_),
    .Y(_01014_),
    .B1(_05396_));
 sg13g2_nand2b_1 _14997_ (.Y(_05397_),
    .B(\top1.event_time[13] ),
    .A_N(_05040_));
 sg13g2_nor2_1 _14998_ (.A(_03838_),
    .B(_05395_),
    .Y(_05398_));
 sg13g2_a21oi_1 _14999_ (.A1(_05395_),
    .A2(_05397_),
    .Y(_01015_),
    .B1(_05398_));
 sg13g2_nor2_1 _15000_ (.A(\top1.event_time[14] ),
    .B(_05398_),
    .Y(_05399_));
 sg13g2_a21o_1 _15001_ (.A2(_05398_),
    .A1(\top1.event_time[14] ),
    .B1(_05040_),
    .X(_05400_));
 sg13g2_nor2_1 _15002_ (.A(_05399_),
    .B(_05400_),
    .Y(_01016_));
 sg13g2_a21oi_1 _15003_ (.A1(\top1.event_time[14] ),
    .A2(_05398_),
    .Y(_05401_),
    .B1(\top1.event_time[15] ));
 sg13g2_a21oi_1 _15004_ (.A1(\top1.event_time[15] ),
    .A2(_05400_),
    .Y(_01017_),
    .B1(_05401_));
 sg13g2_nor2b_2 _15005_ (.A(net6127),
    .B_N(net6128),
    .Y(_05402_));
 sg13g2_nand2b_1 _15006_ (.Y(_05403_),
    .B(net6128),
    .A_N(net6127));
 sg13g2_nor2_1 _15007_ (.A(\top1.memory2.mem1[20][0] ),
    .B(net6045),
    .Y(_05404_));
 sg13g2_nor2b_2 _15008_ (.A(net6147),
    .B_N(net6212),
    .Y(_05405_));
 sg13g2_nand2b_1 _15009_ (.Y(_05406_),
    .B(net6202),
    .A_N(net6138));
 sg13g2_nor2_1 _15010_ (.A(\top1.memory2.mem1[21][0] ),
    .B(net5979),
    .Y(_05407_));
 sg13g2_and2_2 _15011_ (.A(net6212),
    .B(net6147),
    .X(_05408_));
 sg13g2_nand2_1 _15012_ (.Y(_05409_),
    .A(net6199),
    .B(net6135));
 sg13g2_nor2b_2 _15013_ (.A(net6212),
    .B_N(net6147),
    .Y(_05410_));
 sg13g2_nand2b_1 _15014_ (.Y(_05411_),
    .B(net6138),
    .A_N(net6202));
 sg13g2_nor2_1 _15015_ (.A(\top1.memory2.mem1[22][0] ),
    .B(net5899),
    .Y(_05412_));
 sg13g2_o21ai_1 _15016_ (.B1(net6026),
    .Y(_05413_),
    .A1(\top1.memory2.mem1[23][0] ),
    .A2(net5940));
 sg13g2_nor4_2 _15017_ (.A(_05404_),
    .B(_05407_),
    .C(_05412_),
    .Y(_05414_),
    .D(_05413_));
 sg13g2_a22oi_1 _15018_ (.Y(_05415_),
    .B1(net5959),
    .B2(\top1.memory2.mem1[27][0] ),
    .A2(net6064),
    .A1(\top1.memory2.mem1[24][0] ));
 sg13g2_a22oi_1 _15019_ (.Y(_05416_),
    .B1(net5919),
    .B2(\top1.memory2.mem1[26][0] ),
    .A2(net6000),
    .A1(\top1.memory2.mem1[25][0] ));
 sg13g2_a21oi_1 _15020_ (.A1(_05415_),
    .A2(_05416_),
    .Y(_05417_),
    .B1(net6081));
 sg13g2_nor2_2 _15021_ (.A(net6129),
    .B(net6127),
    .Y(_05418_));
 sg13g2_or2_1 _15022_ (.X(_05419_),
    .B(net6127),
    .A(net6128));
 sg13g2_mux4_1 _15023_ (.S0(net6229),
    .A0(\top1.memory2.mem1[16][0] ),
    .A1(\top1.memory2.mem1[17][0] ),
    .A2(\top1.memory2.mem1[18][0] ),
    .A3(\top1.memory2.mem1[19][0] ),
    .S1(net6164),
    .X(_05420_));
 sg13g2_and2_1 _15024_ (.A(net6128),
    .B(net6127),
    .X(_05421_));
 sg13g2_nand2_1 _15025_ (.Y(_05422_),
    .A(net6128),
    .B(net6127));
 sg13g2_a22oi_1 _15026_ (.Y(_05423_),
    .B1(net5959),
    .B2(\top1.memory2.mem1[31][0] ),
    .A2(net6000),
    .A1(\top1.memory2.mem1[29][0] ));
 sg13g2_a22oi_1 _15027_ (.Y(_05424_),
    .B1(net5919),
    .B2(\top1.memory2.mem1[30][0] ),
    .A2(net6064),
    .A1(\top1.memory2.mem1[28][0] ));
 sg13g2_a21oi_1 _15028_ (.A1(_05423_),
    .A2(_05424_),
    .Y(_05425_),
    .B1(net5847));
 sg13g2_a21o_1 _15029_ (.A2(_05420_),
    .A1(net5882),
    .B1(net6107),
    .X(_05426_));
 sg13g2_nor4_2 _15030_ (.A(_05414_),
    .B(_05417_),
    .C(_05425_),
    .Y(_05427_),
    .D(_05426_));
 sg13g2_mux4_1 _15031_ (.S0(net6211),
    .A0(\top1.memory2.mem1[0][0] ),
    .A1(\top1.memory2.mem1[1][0] ),
    .A2(\top1.memory2.mem1[2][0] ),
    .A3(\top1.memory2.mem1[3][0] ),
    .S1(net6146),
    .X(_05428_));
 sg13g2_a21o_1 _15032_ (.A2(_05428_),
    .A1(net5878),
    .B1(net6124),
    .X(_05429_));
 sg13g2_a22oi_1 _15033_ (.Y(_05430_),
    .B1(net5912),
    .B2(\top1.memory2.mem1[14][0] ),
    .A2(net5952),
    .A1(\top1.memory2.mem1[15][0] ));
 sg13g2_a22oi_1 _15034_ (.Y(_05431_),
    .B1(net5999),
    .B2(\top1.memory2.mem1[13][0] ),
    .A2(net6063),
    .A1(\top1.memory2.mem1[12][0] ));
 sg13g2_a21oi_1 _15035_ (.A1(_05430_),
    .A2(_05431_),
    .Y(_05432_),
    .B1(net5847));
 sg13g2_a22oi_1 _15036_ (.Y(_05433_),
    .B1(net5952),
    .B2(\top1.memory2.mem1[11][0] ),
    .A2(net5992),
    .A1(\top1.memory2.mem1[9][0] ));
 sg13g2_a22oi_1 _15037_ (.Y(_05434_),
    .B1(net5912),
    .B2(\top1.memory2.mem1[10][0] ),
    .A2(net6057),
    .A1(\top1.memory2.mem1[8][0] ));
 sg13g2_a21oi_1 _15038_ (.A1(_05433_),
    .A2(_05434_),
    .Y(_05435_),
    .B1(net6077));
 sg13g2_o21ai_1 _15039_ (.B1(net6022),
    .Y(_05436_),
    .A1(\top1.memory2.mem1[4][0] ),
    .A2(net6044));
 sg13g2_nor2_1 _15040_ (.A(\top1.memory2.mem1[7][0] ),
    .B(net5938),
    .Y(_05437_));
 sg13g2_nor2_1 _15041_ (.A(\top1.memory2.mem1[6][0] ),
    .B(net5898),
    .Y(_05438_));
 sg13g2_nor2_1 _15042_ (.A(\top1.memory2.mem1[5][0] ),
    .B(net5977),
    .Y(_05439_));
 sg13g2_nor4_2 _15043_ (.A(_05436_),
    .B(_05437_),
    .C(_05438_),
    .Y(_05440_),
    .D(_05439_));
 sg13g2_nor4_2 _15044_ (.A(_05429_),
    .B(_05432_),
    .C(_05435_),
    .Y(_05441_),
    .D(_05440_));
 sg13g2_or3_1 _15045_ (.A(net6118),
    .B(_05427_),
    .C(_05441_),
    .X(_05442_));
 sg13g2_nor2_2 _15046_ (.A(net6124),
    .B(_03829_),
    .Y(_05443_));
 sg13g2_nand2_2 _15047_ (.Y(_05444_),
    .A(net6106),
    .B(net6118));
 sg13g2_mux4_1 _15048_ (.S0(net6257),
    .A0(\top1.memory2.mem1[40][0] ),
    .A1(\top1.memory2.mem1[41][0] ),
    .A2(\top1.memory2.mem1[42][0] ),
    .A3(\top1.memory2.mem1[43][0] ),
    .S1(net6192),
    .X(_05445_));
 sg13g2_mux4_1 _15049_ (.S0(net6258),
    .A0(\top1.memory2.mem1[36][0] ),
    .A1(\top1.memory2.mem1[37][0] ),
    .A2(\top1.memory2.mem1[38][0] ),
    .A3(\top1.memory2.mem1[39][0] ),
    .S1(net6193),
    .X(_05446_));
 sg13g2_a22oi_1 _15050_ (.Y(_05447_),
    .B1(_05446_),
    .B2(net6035),
    .A2(_05445_),
    .A1(net6098));
 sg13g2_mux4_1 _15051_ (.S0(net6256),
    .A0(\top1.memory2.mem1[44][0] ),
    .A1(\top1.memory2.mem1[45][0] ),
    .A2(\top1.memory2.mem1[46][0] ),
    .A3(\top1.memory2.mem1[47][0] ),
    .S1(net6191),
    .X(_05448_));
 sg13g2_mux4_1 _15052_ (.S0(net6257),
    .A0(\top1.memory2.mem1[32][0] ),
    .A1(\top1.memory2.mem1[33][0] ),
    .A2(\top1.memory2.mem1[34][0] ),
    .A3(\top1.memory2.mem1[35][0] ),
    .S1(net6192),
    .X(_05449_));
 sg13g2_a22oi_1 _15053_ (.Y(_05450_),
    .B1(_05449_),
    .B2(net5887),
    .A2(_05448_),
    .A1(net5865));
 sg13g2_nand2_2 _15054_ (.Y(_05451_),
    .A(_05447_),
    .B(_05450_));
 sg13g2_nor2_2 _15055_ (.A(net6106),
    .B(net6103),
    .Y(_05452_));
 sg13g2_nand2_2 _15056_ (.Y(_05453_),
    .A(net6124),
    .B(net6118));
 sg13g2_mux4_1 _15057_ (.S0(net6240),
    .A0(\top1.memory2.mem1[52][0] ),
    .A1(\top1.memory2.mem1[53][0] ),
    .A2(\top1.memory2.mem1[54][0] ),
    .A3(\top1.memory2.mem1[55][0] ),
    .S1(net6175),
    .X(_05454_));
 sg13g2_mux4_1 _15058_ (.S0(net6250),
    .A0(\top1.memory2.mem1[56][0] ),
    .A1(\top1.memory2.mem1[57][0] ),
    .A2(\top1.memory2.mem1[58][0] ),
    .A3(\top1.memory2.mem1[59][0] ),
    .S1(net6185),
    .X(_05455_));
 sg13g2_a22oi_1 _15059_ (.Y(_05456_),
    .B1(_05455_),
    .B2(net6095),
    .A2(_05454_),
    .A1(net6033));
 sg13g2_mux4_1 _15060_ (.S0(net6255),
    .A0(\top1.memory2.mem1[48][0] ),
    .A1(\top1.memory2.mem1[49][0] ),
    .A2(\top1.memory2.mem1[50][0] ),
    .A3(\top1.memory2.mem1[51][0] ),
    .S1(net6190),
    .X(_05457_));
 sg13g2_mux4_1 _15061_ (.S0(net6247),
    .A0(\top1.memory2.mem1[60][0] ),
    .A1(\top1.memory2.mem1[61][0] ),
    .A2(\top1.memory2.mem1[62][0] ),
    .A3(\top1.memory2.mem1[63][0] ),
    .S1(net6182),
    .X(_05458_));
 sg13g2_a22oi_1 _15062_ (.Y(_05459_),
    .B1(_05458_),
    .B2(net5864),
    .A2(_05457_),
    .A1(net5886));
 sg13g2_nand2_2 _15063_ (.Y(_05460_),
    .A(_05456_),
    .B(_05459_));
 sg13g2_a22oi_1 _15064_ (.Y(_05461_),
    .B1(_05452_),
    .B2(_05460_),
    .A2(_05451_),
    .A1(_05443_));
 sg13g2_a21oi_2 _15065_ (.B1(net6115),
    .Y(_05462_),
    .A2(_05461_),
    .A1(_05442_));
 sg13g2_a22oi_1 _15066_ (.Y(_05463_),
    .B1(net5911),
    .B2(\top1.memory2.mem1[82][0] ),
    .A2(net5951),
    .A1(\top1.memory2.mem1[83][0] ));
 sg13g2_a22oi_1 _15067_ (.Y(_05464_),
    .B1(net5993),
    .B2(\top1.memory2.mem1[81][0] ),
    .A2(net6056),
    .A1(\top1.memory2.mem1[80][0] ));
 sg13g2_nand2_1 _15068_ (.Y(_05465_),
    .A(_05463_),
    .B(_05464_));
 sg13g2_a21oi_1 _15069_ (.A1(net5877),
    .A2(_05465_),
    .Y(_05466_),
    .B1(net6105));
 sg13g2_a22oi_1 _15070_ (.Y(_05467_),
    .B1(net5912),
    .B2(\top1.memory2.mem1[90][0] ),
    .A2(net6057),
    .A1(\top1.memory2.mem1[88][0] ));
 sg13g2_a22oi_1 _15071_ (.Y(_05468_),
    .B1(net5952),
    .B2(\top1.memory2.mem1[91][0] ),
    .A2(net5992),
    .A1(\top1.memory2.mem1[89][0] ));
 sg13g2_a21oi_1 _15072_ (.A1(_05467_),
    .A2(_05468_),
    .Y(_05469_),
    .B1(net6077));
 sg13g2_nor2_1 _15073_ (.A(\top1.memory2.mem1[85][0] ),
    .B(net5973),
    .Y(_05470_));
 sg13g2_nor2_1 _15074_ (.A(\top1.memory2.mem1[87][0] ),
    .B(net5937),
    .Y(_05471_));
 sg13g2_nor2_1 _15075_ (.A(\top1.memory2.mem1[86][0] ),
    .B(net5894),
    .Y(_05472_));
 sg13g2_o21ai_1 _15076_ (.B1(net6021),
    .Y(_05473_),
    .A1(\top1.memory2.mem1[84][0] ),
    .A2(net6039));
 sg13g2_nor4_2 _15077_ (.A(_05470_),
    .B(_05471_),
    .C(_05472_),
    .Y(_05474_),
    .D(_05473_));
 sg13g2_a22oi_1 _15078_ (.Y(_05475_),
    .B1(net5912),
    .B2(\top1.memory2.mem1[94][0] ),
    .A2(net6057),
    .A1(\top1.memory2.mem1[92][0] ));
 sg13g2_a22oi_1 _15079_ (.Y(_05476_),
    .B1(net5952),
    .B2(\top1.memory2.mem1[95][0] ),
    .A2(net5992),
    .A1(\top1.memory2.mem1[93][0] ));
 sg13g2_a21oi_1 _15080_ (.A1(_05475_),
    .A2(_05476_),
    .Y(_05477_),
    .B1(net5845));
 sg13g2_nor3_1 _15081_ (.A(_05469_),
    .B(_05474_),
    .C(_05477_),
    .Y(_05478_));
 sg13g2_nand2_2 _15082_ (.Y(_05479_),
    .A(net6103),
    .B(net6113));
 sg13g2_a22oi_1 _15083_ (.Y(_05480_),
    .B1(net5943),
    .B2(\top1.memory2.mem1[79][0] ),
    .A2(net5985),
    .A1(\top1.memory2.mem1[77][0] ));
 sg13g2_a22oi_1 _15084_ (.Y(_05481_),
    .B1(net5902),
    .B2(\top1.memory2.mem1[78][0] ),
    .A2(net6047),
    .A1(\top1.memory2.mem1[76][0] ));
 sg13g2_a21oi_1 _15085_ (.A1(_05480_),
    .A2(_05481_),
    .Y(_05482_),
    .B1(net5844));
 sg13g2_a22oi_1 _15086_ (.Y(_05483_),
    .B1(net5901),
    .B2(\top1.memory2.mem1[66][0] ),
    .A2(net6046),
    .A1(\top1.memory2.mem1[64][0] ));
 sg13g2_a22oi_1 _15087_ (.Y(_05484_),
    .B1(net5943),
    .B2(\top1.memory2.mem1[67][0] ),
    .A2(net5981),
    .A1(\top1.memory2.mem1[65][0] ));
 sg13g2_nand2_1 _15088_ (.Y(_05485_),
    .A(_05483_),
    .B(_05484_));
 sg13g2_a22oi_1 _15089_ (.Y(_05486_),
    .B1(net5902),
    .B2(\top1.memory2.mem1[74][0] ),
    .A2(net6049),
    .A1(\top1.memory2.mem1[72][0] ));
 sg13g2_a22oi_1 _15090_ (.Y(_05487_),
    .B1(net5943),
    .B2(\top1.memory2.mem1[75][0] ),
    .A2(net5982),
    .A1(\top1.memory2.mem1[73][0] ));
 sg13g2_a21oi_1 _15091_ (.A1(_05486_),
    .A2(_05487_),
    .Y(_05488_),
    .B1(net6075));
 sg13g2_o21ai_1 _15092_ (.B1(net6018),
    .Y(_05489_),
    .A1(\top1.memory2.mem1[70][0] ),
    .A2(net5890));
 sg13g2_nor2_1 _15093_ (.A(\top1.memory2.mem1[68][0] ),
    .B(net6036),
    .Y(_05490_));
 sg13g2_nor2_1 _15094_ (.A(\top1.memory2.mem1[69][0] ),
    .B(net5970),
    .Y(_05491_));
 sg13g2_nor2_1 _15095_ (.A(\top1.memory2.mem1[71][0] ),
    .B(net5932),
    .Y(_05492_));
 sg13g2_nor4_1 _15096_ (.A(_05489_),
    .B(_05490_),
    .C(_05491_),
    .D(_05492_),
    .Y(_05493_));
 sg13g2_a21o_1 _15097_ (.A2(_05485_),
    .A1(net5874),
    .B1(net6120),
    .X(_05494_));
 sg13g2_nor4_2 _15098_ (.A(_05482_),
    .B(_05488_),
    .C(_05493_),
    .Y(_05495_),
    .D(_05494_));
 sg13g2_a21o_1 _15099_ (.A2(_05478_),
    .A1(_05466_),
    .B1(_05479_),
    .X(_05496_));
 sg13g2_mux4_1 _15100_ (.S0(net6243),
    .A0(\top1.memory2.mem1[124][0] ),
    .A1(\top1.memory2.mem1[125][0] ),
    .A2(\top1.memory2.mem1[126][0] ),
    .A3(\top1.memory2.mem1[127][0] ),
    .S1(net6178),
    .X(_05497_));
 sg13g2_mux4_1 _15101_ (.S0(net6241),
    .A0(\top1.memory2.mem1[120][0] ),
    .A1(\top1.memory2.mem1[121][0] ),
    .A2(\top1.memory2.mem1[122][0] ),
    .A3(\top1.memory2.mem1[123][0] ),
    .S1(net6176),
    .X(_05498_));
 sg13g2_mux4_1 _15102_ (.S0(net6243),
    .A0(\top1.memory2.mem1[116][0] ),
    .A1(\top1.memory2.mem1[117][0] ),
    .A2(\top1.memory2.mem1[118][0] ),
    .A3(\top1.memory2.mem1[119][0] ),
    .S1(net6178),
    .X(_05499_));
 sg13g2_mux4_1 _15103_ (.S0(net6243),
    .A0(\top1.memory2.mem1[112][0] ),
    .A1(\top1.memory2.mem1[113][0] ),
    .A2(\top1.memory2.mem1[114][0] ),
    .A3(\top1.memory2.mem1[115][0] ),
    .S1(net6178),
    .X(_05500_));
 sg13g2_a22oi_1 _15104_ (.Y(_05501_),
    .B1(_05499_),
    .B2(net6030),
    .A2(_05497_),
    .A1(net5861));
 sg13g2_a22oi_1 _15105_ (.Y(_05502_),
    .B1(_05500_),
    .B2(net5884),
    .A2(_05498_),
    .A1(net6095));
 sg13g2_a21oi_2 _15106_ (.B1(net5839),
    .Y(_05503_),
    .A2(_05502_),
    .A1(_05501_));
 sg13g2_mux4_1 _15107_ (.S0(net6249),
    .A0(\top1.memory2.mem1[104][0] ),
    .A1(\top1.memory2.mem1[105][0] ),
    .A2(\top1.memory2.mem1[106][0] ),
    .A3(\top1.memory2.mem1[107][0] ),
    .S1(net6184),
    .X(_05504_));
 sg13g2_mux4_1 _15108_ (.S0(net6226),
    .A0(\top1.memory2.mem1[96][0] ),
    .A1(\top1.memory2.mem1[97][0] ),
    .A2(\top1.memory2.mem1[98][0] ),
    .A3(\top1.memory2.mem1[99][0] ),
    .S1(net6161),
    .X(_05505_));
 sg13g2_mux4_1 _15109_ (.S0(net6240),
    .A0(\top1.memory2.mem1[108][0] ),
    .A1(\top1.memory2.mem1[109][0] ),
    .A2(\top1.memory2.mem1[110][0] ),
    .A3(\top1.memory2.mem1[111][0] ),
    .S1(net6175),
    .X(_05506_));
 sg13g2_mux4_1 _15110_ (.S0(net6226),
    .A0(\top1.memory2.mem1[100][0] ),
    .A1(\top1.memory2.mem1[101][0] ),
    .A2(\top1.memory2.mem1[102][0] ),
    .A3(\top1.memory2.mem1[103][0] ),
    .S1(net6161),
    .X(_05507_));
 sg13g2_a22oi_1 _15111_ (.Y(_05508_),
    .B1(_05506_),
    .B2(net5863),
    .A2(_05504_),
    .A1(net6093));
 sg13g2_a22oi_1 _15112_ (.Y(_05509_),
    .B1(_05507_),
    .B2(net6025),
    .A2(_05505_),
    .A1(net5881));
 sg13g2_a21oi_1 _15113_ (.A1(_05508_),
    .A2(_05509_),
    .Y(_05510_),
    .B1(net5833));
 sg13g2_o21ai_1 _15114_ (.B1(net6116),
    .Y(_05511_),
    .A1(_05503_),
    .A2(_05510_));
 sg13g2_and2_1 _15115_ (.A(_03831_),
    .B(_05511_),
    .X(_05512_));
 sg13g2_o21ai_1 _15116_ (.B1(_05512_),
    .Y(_05513_),
    .A1(_05495_),
    .A2(_05496_));
 sg13g2_nor2_2 _15117_ (.A(net6113),
    .B(_03831_),
    .Y(_05514_));
 sg13g2_nand2_1 _15118_ (.Y(_05515_),
    .A(net6102),
    .B(net6112));
 sg13g2_nor2_2 _15119_ (.A(net6106),
    .B(net6118),
    .Y(_05516_));
 sg13g2_nand2_1 _15120_ (.Y(_05517_),
    .A(net6124),
    .B(net6103));
 sg13g2_a22oi_1 _15121_ (.Y(_05518_),
    .B1(net5949),
    .B2(\top1.memory2.mem1[155][0] ),
    .A2(net6053),
    .A1(\top1.memory2.mem1[152][0] ));
 sg13g2_a22oi_1 _15122_ (.Y(_05519_),
    .B1(net5908),
    .B2(\top1.memory2.mem1[154][0] ),
    .A2(net5989),
    .A1(\top1.memory2.mem1[153][0] ));
 sg13g2_a21oi_1 _15123_ (.A1(_05518_),
    .A2(_05519_),
    .Y(_05520_),
    .B1(net6076));
 sg13g2_o21ai_1 _15124_ (.B1(net6020),
    .Y(_05521_),
    .A1(\top1.memory2.mem1[149][0] ),
    .A2(net5974));
 sg13g2_nor2_1 _15125_ (.A(\top1.memory2.mem1[150][0] ),
    .B(net5895),
    .Y(_05522_));
 sg13g2_nor2_1 _15126_ (.A(\top1.memory2.mem1[148][0] ),
    .B(net6040),
    .Y(_05523_));
 sg13g2_nor2_1 _15127_ (.A(\top1.memory2.mem1[151][0] ),
    .B(net5934),
    .Y(_05524_));
 sg13g2_nor4_1 _15128_ (.A(_05521_),
    .B(_05522_),
    .C(_05523_),
    .D(_05524_),
    .Y(_05525_));
 sg13g2_a22oi_1 _15129_ (.Y(_05526_),
    .B1(net5908),
    .B2(\top1.memory2.mem1[146][0] ),
    .A2(net6053),
    .A1(\top1.memory2.mem1[144][0] ));
 sg13g2_a22oi_1 _15130_ (.Y(_05527_),
    .B1(net5949),
    .B2(\top1.memory2.mem1[147][0] ),
    .A2(net5989),
    .A1(\top1.memory2.mem1[145][0] ));
 sg13g2_a21oi_1 _15131_ (.A1(_05526_),
    .A2(_05527_),
    .Y(_05528_),
    .B1(net5869));
 sg13g2_a22oi_1 _15132_ (.Y(_05529_),
    .B1(net5909),
    .B2(\top1.memory2.mem1[158][0] ),
    .A2(net5948),
    .A1(\top1.memory2.mem1[159][0] ));
 sg13g2_a22oi_1 _15133_ (.Y(_05530_),
    .B1(net5990),
    .B2(\top1.memory2.mem1[157][0] ),
    .A2(net6054),
    .A1(\top1.memory2.mem1[156][0] ));
 sg13g2_a21oi_2 _15134_ (.B1(net5843),
    .Y(_05531_),
    .A2(_05530_),
    .A1(_05529_));
 sg13g2_or4_1 _15135_ (.A(_05520_),
    .B(_05525_),
    .C(_05528_),
    .D(_05531_),
    .X(_05532_));
 sg13g2_a22oi_1 _15136_ (.Y(_05533_),
    .B1(net5907),
    .B2(\top1.memory2.mem1[142][0] ),
    .A2(net5947),
    .A1(\top1.memory2.mem1[143][0] ));
 sg13g2_a22oi_1 _15137_ (.Y(_05534_),
    .B1(net5988),
    .B2(\top1.memory2.mem1[141][0] ),
    .A2(net6052),
    .A1(\top1.memory2.mem1[140][0] ));
 sg13g2_a21oi_1 _15138_ (.A1(_05533_),
    .A2(_05534_),
    .Y(_05535_),
    .B1(net5842));
 sg13g2_nor2_1 _15139_ (.A(\top1.memory2.mem1[135][0] ),
    .B(net5930),
    .Y(_05536_));
 sg13g2_nor2_1 _15140_ (.A(\top1.memory2.mem1[133][0] ),
    .B(net5971),
    .Y(_05537_));
 sg13g2_nor2_1 _15141_ (.A(\top1.memory2.mem1[132][0] ),
    .B(net6036),
    .Y(_05538_));
 sg13g2_o21ai_1 _15142_ (.B1(net6019),
    .Y(_05539_),
    .A1(\top1.memory2.mem1[134][0] ),
    .A2(net5891));
 sg13g2_nor4_1 _15143_ (.A(_05536_),
    .B(_05537_),
    .C(_05538_),
    .D(_05539_),
    .Y(_05540_));
 sg13g2_a22oi_1 _15144_ (.Y(_05541_),
    .B1(net5907),
    .B2(\top1.memory2.mem1[138][0] ),
    .A2(net5947),
    .A1(\top1.memory2.mem1[139][0] ));
 sg13g2_a22oi_1 _15145_ (.Y(_05542_),
    .B1(net5985),
    .B2(\top1.memory2.mem1[137][0] ),
    .A2(net6052),
    .A1(\top1.memory2.mem1[136][0] ));
 sg13g2_a21oi_1 _15146_ (.A1(_05541_),
    .A2(_05542_),
    .Y(_05543_),
    .B1(net6079));
 sg13g2_a22oi_1 _15147_ (.Y(_05544_),
    .B1(net5902),
    .B2(\top1.memory2.mem1[130][0] ),
    .A2(net5982),
    .A1(\top1.memory2.mem1[129][0] ));
 sg13g2_a22oi_1 _15148_ (.Y(_05545_),
    .B1(net5943),
    .B2(\top1.memory2.mem1[131][0] ),
    .A2(net6047),
    .A1(\top1.memory2.mem1[128][0] ));
 sg13g2_a21oi_1 _15149_ (.A1(_05544_),
    .A2(_05545_),
    .Y(_05546_),
    .B1(net5868));
 sg13g2_or4_2 _15150_ (.A(_05535_),
    .B(_05540_),
    .C(_05543_),
    .D(_05546_),
    .X(_05547_));
 sg13g2_a22oi_1 _15151_ (.Y(_05548_),
    .B1(net5926),
    .B2(\top1.memory2.mem1[190][0] ),
    .A2(net5966),
    .A1(\top1.memory2.mem1[191][0] ));
 sg13g2_a22oi_1 _15152_ (.Y(_05549_),
    .B1(net6006),
    .B2(\top1.memory2.mem1[189][0] ),
    .A2(net6070),
    .A1(\top1.memory2.mem1[188][0] ));
 sg13g2_a21oi_1 _15153_ (.A1(_05548_),
    .A2(_05549_),
    .Y(_05550_),
    .B1(net5848));
 sg13g2_a22oi_1 _15154_ (.Y(_05551_),
    .B1(net5919),
    .B2(\top1.memory2.mem1[186][0] ),
    .A2(net5959),
    .A1(\top1.memory2.mem1[187][0] ));
 sg13g2_a22oi_1 _15155_ (.Y(_05552_),
    .B1(net6000),
    .B2(\top1.memory2.mem1[185][0] ),
    .A2(net6069),
    .A1(\top1.memory2.mem1[184][0] ));
 sg13g2_a21oi_1 _15156_ (.A1(_05551_),
    .A2(_05552_),
    .Y(_05553_),
    .B1(net6081));
 sg13g2_a22oi_1 _15157_ (.Y(_05554_),
    .B1(net5926),
    .B2(\top1.memory2.mem1[182][0] ),
    .A2(net5966),
    .A1(\top1.memory2.mem1[183][0] ));
 sg13g2_a22oi_1 _15158_ (.Y(_05555_),
    .B1(net6006),
    .B2(\top1.memory2.mem1[181][0] ),
    .A2(net6070),
    .A1(\top1.memory2.mem1[180][0] ));
 sg13g2_a21oi_2 _15159_ (.B1(net6014),
    .Y(_05556_),
    .A2(_05555_),
    .A1(_05554_));
 sg13g2_a22oi_1 _15160_ (.Y(_05557_),
    .B1(net5926),
    .B2(\top1.memory2.mem1[178][0] ),
    .A2(net5966),
    .A1(\top1.memory2.mem1[179][0] ));
 sg13g2_a22oi_1 _15161_ (.Y(_05558_),
    .B1(net6006),
    .B2(\top1.memory2.mem1[177][0] ),
    .A2(net6070),
    .A1(\top1.memory2.mem1[176][0] ));
 sg13g2_a21oi_1 _15162_ (.A1(_05557_),
    .A2(_05558_),
    .Y(_05559_),
    .B1(net5871));
 sg13g2_or4_2 _15163_ (.A(_05550_),
    .B(_05553_),
    .C(_05556_),
    .D(_05559_),
    .X(_05560_));
 sg13g2_mux4_1 _15164_ (.S0(net6222),
    .A0(\top1.memory2.mem1[164][0] ),
    .A1(\top1.memory2.mem1[165][0] ),
    .A2(\top1.memory2.mem1[166][0] ),
    .A3(\top1.memory2.mem1[167][0] ),
    .S1(net6157),
    .X(_05561_));
 sg13g2_mux4_1 _15165_ (.S0(net6220),
    .A0(\top1.memory2.mem1[172][0] ),
    .A1(\top1.memory2.mem1[173][0] ),
    .A2(\top1.memory2.mem1[174][0] ),
    .A3(\top1.memory2.mem1[175][0] ),
    .S1(net6155),
    .X(_05562_));
 sg13g2_mux4_1 _15166_ (.S0(net6221),
    .A0(\top1.memory2.mem1[168][0] ),
    .A1(\top1.memory2.mem1[169][0] ),
    .A2(\top1.memory2.mem1[170][0] ),
    .A3(\top1.memory2.mem1[171][0] ),
    .S1(net6156),
    .X(_05563_));
 sg13g2_mux4_1 _15167_ (.S0(net6212),
    .A0(\top1.memory2.mem1[160][0] ),
    .A1(\top1.memory2.mem1[161][0] ),
    .A2(\top1.memory2.mem1[162][0] ),
    .A3(\top1.memory2.mem1[163][0] ),
    .S1(net6147),
    .X(_05564_));
 sg13g2_a22oi_1 _15168_ (.Y(_05565_),
    .B1(_05563_),
    .B2(net6089),
    .A2(_05561_),
    .A1(net6026));
 sg13g2_a22oi_1 _15169_ (.Y(_05566_),
    .B1(_05564_),
    .B2(net5877),
    .A2(_05562_),
    .A1(net5855));
 sg13g2_a21oi_2 _15170_ (.B1(net5836),
    .Y(_05567_),
    .A2(_05566_),
    .A1(_05565_));
 sg13g2_a21oi_1 _15171_ (.A1(_05452_),
    .A2(_05560_),
    .Y(_05568_),
    .B1(net5831));
 sg13g2_a221oi_1 _15172_ (.B2(_03976_),
    .C1(_05567_),
    .B1(_05547_),
    .A1(_05516_),
    .Y(_05569_),
    .A2(_05532_));
 sg13g2_nor2_1 _15173_ (.A(\top1.memory2.mem1[198][0] ),
    .B(net5896),
    .Y(_05570_));
 sg13g2_nor2_1 _15174_ (.A(\top1.memory2.mem1[197][0] ),
    .B(net5974),
    .Y(_05571_));
 sg13g2_o21ai_1 _15175_ (.B1(net6130),
    .Y(_05572_),
    .A1(\top1.memory2.mem1[199][0] ),
    .A2(net5933));
 sg13g2_nor3_1 _15176_ (.A(_05570_),
    .B(_05571_),
    .C(_05572_),
    .Y(_05573_));
 sg13g2_o21ai_1 _15177_ (.B1(_05573_),
    .Y(_05574_),
    .A1(\top1.memory2.mem1[196][0] ),
    .A2(net6041));
 sg13g2_nor2_1 _15178_ (.A(\top1.memory2.mem1[195][0] ),
    .B(net5937),
    .Y(_05575_));
 sg13g2_nor2_1 _15179_ (.A(\top1.memory2.mem1[192][0] ),
    .B(net6043),
    .Y(_05576_));
 sg13g2_nor2_1 _15180_ (.A(\top1.memory2.mem1[194][0] ),
    .B(net5897),
    .Y(_05577_));
 sg13g2_o21ai_1 _15181_ (.B1(_03827_),
    .Y(_05578_),
    .A1(\top1.memory2.mem1[193][0] ),
    .A2(net5977));
 sg13g2_nor4_2 _15182_ (.A(_05575_),
    .B(_05576_),
    .C(_05577_),
    .Y(_05579_),
    .D(_05578_));
 sg13g2_nor2_1 _15183_ (.A(_03979_),
    .B(_05579_),
    .Y(_05580_));
 sg13g2_a221oi_1 _15184_ (.B2(_05580_),
    .C1(net6108),
    .B1(_05574_),
    .A1(_05568_),
    .Y(_05581_),
    .A2(_05569_));
 sg13g2_o21ai_1 _15185_ (.B1(_05581_),
    .Y(_05582_),
    .A1(_05462_),
    .A2(_05513_));
 sg13g2_a22oi_1 _15186_ (.Y(_05583_),
    .B1(net5929),
    .B2(\top1.memory2.mem2[42][0] ),
    .A2(net5969),
    .A1(\top1.memory2.mem2[43][0] ));
 sg13g2_a22oi_1 _15187_ (.Y(_05584_),
    .B1(net6008),
    .B2(\top1.memory2.mem2[41][0] ),
    .A2(net6072),
    .A1(\top1.memory2.mem2[40][0] ));
 sg13g2_a21oi_1 _15188_ (.A1(_05583_),
    .A2(_05584_),
    .Y(_05585_),
    .B1(net6082));
 sg13g2_a22oi_1 _15189_ (.Y(_05586_),
    .B1(net5927),
    .B2(\top1.memory2.mem2[38][0] ),
    .A2(net5967),
    .A1(\top1.memory2.mem2[39][0] ));
 sg13g2_a22oi_1 _15190_ (.Y(_05587_),
    .B1(net6007),
    .B2(\top1.memory2.mem2[37][0] ),
    .A2(net6071),
    .A1(\top1.memory2.mem2[36][0] ));
 sg13g2_a21oi_1 _15191_ (.A1(_05586_),
    .A2(_05587_),
    .Y(_05588_),
    .B1(net6015));
 sg13g2_a22oi_1 _15192_ (.Y(_05589_),
    .B1(net5928),
    .B2(\top1.memory2.mem2[46][0] ),
    .A2(net5968),
    .A1(\top1.memory2.mem2[47][0] ));
 sg13g2_a22oi_1 _15193_ (.Y(_05590_),
    .B1(net6008),
    .B2(\top1.memory2.mem2[45][0] ),
    .A2(net6072),
    .A1(\top1.memory2.mem2[44][0] ));
 sg13g2_a21oi_1 _15194_ (.A1(_05589_),
    .A2(_05590_),
    .Y(_05591_),
    .B1(net5849));
 sg13g2_a22oi_1 _15195_ (.Y(_05592_),
    .B1(net5927),
    .B2(\top1.memory2.mem2[34][0] ),
    .A2(net5967),
    .A1(\top1.memory2.mem2[35][0] ));
 sg13g2_a22oi_1 _15196_ (.Y(_05593_),
    .B1(net6007),
    .B2(\top1.memory2.mem2[33][0] ),
    .A2(net6071),
    .A1(\top1.memory2.mem2[32][0] ));
 sg13g2_a21oi_1 _15197_ (.A1(_05592_),
    .A2(_05593_),
    .Y(_05594_),
    .B1(net5872));
 sg13g2_nor4_2 _15198_ (.A(_05585_),
    .B(_05588_),
    .C(_05591_),
    .Y(_05595_),
    .D(_05594_));
 sg13g2_nor2_1 _15199_ (.A(\top1.memory2.mem2[7][0] ),
    .B(net5939),
    .Y(_05596_));
 sg13g2_nor2_1 _15200_ (.A(\top1.memory2.mem2[4][0] ),
    .B(net6044),
    .Y(_05597_));
 sg13g2_nor2_1 _15201_ (.A(\top1.memory2.mem2[6][0] ),
    .B(net5899),
    .Y(_05598_));
 sg13g2_o21ai_1 _15202_ (.B1(net6024),
    .Y(_05599_),
    .A1(\top1.memory2.mem2[5][0] ),
    .A2(net5978));
 sg13g2_nor4_2 _15203_ (.A(_05596_),
    .B(_05597_),
    .C(_05598_),
    .Y(_05600_),
    .D(_05599_));
 sg13g2_a22oi_1 _15204_ (.Y(_05601_),
    .B1(net5916),
    .B2(\top1.memory2.mem2[14][0] ),
    .A2(net5956),
    .A1(\top1.memory2.mem2[15][0] ));
 sg13g2_a22oi_1 _15205_ (.Y(_05602_),
    .B1(net5996),
    .B2(\top1.memory2.mem2[13][0] ),
    .A2(net6061),
    .A1(\top1.memory2.mem2[12][0] ));
 sg13g2_a21oi_2 _15206_ (.B1(net5846),
    .Y(_05603_),
    .A2(_05602_),
    .A1(_05601_));
 sg13g2_a22oi_1 _15207_ (.Y(_05604_),
    .B1(net5921),
    .B2(\top1.memory2.mem2[2][0] ),
    .A2(net5961),
    .A1(\top1.memory2.mem2[3][0] ));
 sg13g2_a22oi_1 _15208_ (.Y(_05605_),
    .B1(net6002),
    .B2(\top1.memory2.mem2[1][0] ),
    .A2(net6068),
    .A1(\top1.memory2.mem2[0][0] ));
 sg13g2_a21oi_2 _15209_ (.B1(net5871),
    .Y(_05606_),
    .A2(_05605_),
    .A1(_05604_));
 sg13g2_a22oi_1 _15210_ (.Y(_05607_),
    .B1(net5915),
    .B2(\top1.memory2.mem2[10][0] ),
    .A2(net5955),
    .A1(\top1.memory2.mem2[11][0] ));
 sg13g2_a22oi_1 _15211_ (.Y(_05608_),
    .B1(net5996),
    .B2(\top1.memory2.mem2[9][0] ),
    .A2(net6061),
    .A1(\top1.memory2.mem2[8][0] ));
 sg13g2_a21oi_1 _15212_ (.A1(_05607_),
    .A2(_05608_),
    .Y(_05609_),
    .B1(net6078));
 sg13g2_nor4_2 _15213_ (.A(_05600_),
    .B(_05603_),
    .C(_05606_),
    .Y(_05610_),
    .D(_05609_));
 sg13g2_mux4_1 _15214_ (.S0(net6252),
    .A0(\top1.memory2.mem2[60][0] ),
    .A1(\top1.memory2.mem2[61][0] ),
    .A2(\top1.memory2.mem2[62][0] ),
    .A3(\top1.memory2.mem2[63][0] ),
    .S1(net6187),
    .X(_05611_));
 sg13g2_mux4_1 _15215_ (.S0(net6250),
    .A0(\top1.memory2.mem2[56][0] ),
    .A1(\top1.memory2.mem2[57][0] ),
    .A2(\top1.memory2.mem2[58][0] ),
    .A3(\top1.memory2.mem2[59][0] ),
    .S1(net6185),
    .X(_05612_));
 sg13g2_nand2_1 _15216_ (.Y(_05613_),
    .A(net6098),
    .B(_05612_));
 sg13g2_mux4_1 _15217_ (.S0(net6253),
    .A0(\top1.memory2.mem2[48][0] ),
    .A1(\top1.memory2.mem2[49][0] ),
    .A2(\top1.memory2.mem2[50][0] ),
    .A3(\top1.memory2.mem2[51][0] ),
    .S1(net6188),
    .X(_05614_));
 sg13g2_a22oi_1 _15218_ (.Y(_05615_),
    .B1(net5928),
    .B2(\top1.memory2.mem2[54][0] ),
    .A2(net5968),
    .A1(\top1.memory2.mem2[55][0] ));
 sg13g2_a22oi_1 _15219_ (.Y(_05616_),
    .B1(net6008),
    .B2(\top1.memory2.mem2[53][0] ),
    .A2(net6072),
    .A1(\top1.memory2.mem2[52][0] ));
 sg13g2_a21oi_1 _15220_ (.A1(_05615_),
    .A2(_05616_),
    .Y(_05617_),
    .B1(net6015));
 sg13g2_a22oi_1 _15221_ (.Y(_05618_),
    .B1(_05614_),
    .B2(net5888),
    .A2(_05611_),
    .A1(net5863));
 sg13g2_nand2_1 _15222_ (.Y(_05619_),
    .A(_05613_),
    .B(_05618_));
 sg13g2_nor2_2 _15223_ (.A(_05617_),
    .B(_05619_),
    .Y(_05620_));
 sg13g2_o21ai_1 _15224_ (.B1(net6027),
    .Y(_05621_),
    .A1(\top1.memory2.mem2[23][0] ),
    .A2(net5940));
 sg13g2_nor2_1 _15225_ (.A(\top1.memory2.mem2[21][0] ),
    .B(net5979),
    .Y(_05622_));
 sg13g2_nor2_1 _15226_ (.A(\top1.memory2.mem2[22][0] ),
    .B(net5899),
    .Y(_05623_));
 sg13g2_nor2_1 _15227_ (.A(\top1.memory2.mem2[20][0] ),
    .B(net6045),
    .Y(_05624_));
 sg13g2_nor4_2 _15228_ (.A(_05621_),
    .B(_05622_),
    .C(_05623_),
    .Y(_05625_),
    .D(_05624_));
 sg13g2_a22oi_1 _15229_ (.Y(_05626_),
    .B1(net5963),
    .B2(\top1.memory2.mem2[19][0] ),
    .A2(net6067),
    .A1(\top1.memory2.mem2[16][0] ));
 sg13g2_a22oi_1 _15230_ (.Y(_05627_),
    .B1(net5924),
    .B2(\top1.memory2.mem2[18][0] ),
    .A2(net6005),
    .A1(\top1.memory2.mem2[17][0] ));
 sg13g2_a21oi_2 _15231_ (.B1(net5870),
    .Y(_05628_),
    .A2(_05627_),
    .A1(_05626_));
 sg13g2_a22oi_1 _15232_ (.Y(_05629_),
    .B1(net5925),
    .B2(\top1.memory2.mem2[30][0] ),
    .A2(net5965),
    .A1(\top1.memory2.mem2[31][0] ));
 sg13g2_a22oi_1 _15233_ (.Y(_05630_),
    .B1(net6002),
    .B2(\top1.memory2.mem2[29][0] ),
    .A2(net6065),
    .A1(\top1.memory2.mem2[28][0] ));
 sg13g2_a21oi_1 _15234_ (.A1(_05629_),
    .A2(_05630_),
    .Y(_05631_),
    .B1(net5848));
 sg13g2_a22oi_1 _15235_ (.Y(_05632_),
    .B1(net5923),
    .B2(\top1.memory2.mem2[26][0] ),
    .A2(net5963),
    .A1(\top1.memory2.mem2[27][0] ));
 sg13g2_a22oi_1 _15236_ (.Y(_05633_),
    .B1(net6004),
    .B2(\top1.memory2.mem2[25][0] ),
    .A2(net6066),
    .A1(\top1.memory2.mem2[24][0] ));
 sg13g2_a21oi_1 _15237_ (.A1(_05632_),
    .A2(_05633_),
    .Y(_05634_),
    .B1(net6080));
 sg13g2_nor4_2 _15238_ (.A(_05625_),
    .B(_05628_),
    .C(_05631_),
    .Y(_05635_),
    .D(_05634_));
 sg13g2_mux4_1 _15239_ (.S0(net6103),
    .A0(_05595_),
    .A1(_05610_),
    .A2(_05620_),
    .A3(_05635_),
    .S1(net6125),
    .X(_05636_));
 sg13g2_mux4_1 _15240_ (.S0(net6236),
    .A0(\top1.memory2.mem2[108][0] ),
    .A1(\top1.memory2.mem2[109][0] ),
    .A2(\top1.memory2.mem2[110][0] ),
    .A3(\top1.memory2.mem2[111][0] ),
    .S1(net6171),
    .X(_05637_));
 sg13g2_mux4_1 _15241_ (.S0(net6223),
    .A0(\top1.memory2.mem2[96][0] ),
    .A1(\top1.memory2.mem2[97][0] ),
    .A2(\top1.memory2.mem2[98][0] ),
    .A3(\top1.memory2.mem2[99][0] ),
    .S1(net6158),
    .X(_05638_));
 sg13g2_mux4_1 _15242_ (.S0(net6223),
    .A0(\top1.memory2.mem2[100][0] ),
    .A1(\top1.memory2.mem2[101][0] ),
    .A2(\top1.memory2.mem2[102][0] ),
    .A3(\top1.memory2.mem2[103][0] ),
    .S1(net6158),
    .X(_05639_));
 sg13g2_mux4_1 _15243_ (.S0(net6238),
    .A0(\top1.memory2.mem2[104][0] ),
    .A1(\top1.memory2.mem2[105][0] ),
    .A2(\top1.memory2.mem2[106][0] ),
    .A3(\top1.memory2.mem2[107][0] ),
    .S1(net6173),
    .X(_05640_));
 sg13g2_a22oi_1 _15244_ (.Y(_05641_),
    .B1(_05639_),
    .B2(net6031),
    .A2(_05637_),
    .A1(net5857));
 sg13g2_a22oi_1 _15245_ (.Y(_05642_),
    .B1(_05640_),
    .B2(net6093),
    .A2(_05638_),
    .A1(net5885));
 sg13g2_a21oi_1 _15246_ (.A1(_05641_),
    .A2(_05642_),
    .Y(_05643_),
    .B1(net5832));
 sg13g2_mux4_1 _15247_ (.S0(net6242),
    .A0(\top1.memory2.mem2[112][0] ),
    .A1(\top1.memory2.mem2[113][0] ),
    .A2(\top1.memory2.mem2[114][0] ),
    .A3(\top1.memory2.mem2[115][0] ),
    .S1(net6177),
    .X(_05644_));
 sg13g2_mux4_1 _15248_ (.S0(net6238),
    .A0(\top1.memory2.mem2[120][0] ),
    .A1(\top1.memory2.mem2[121][0] ),
    .A2(\top1.memory2.mem2[122][0] ),
    .A3(\top1.memory2.mem2[123][0] ),
    .S1(net6173),
    .X(_05645_));
 sg13g2_mux4_1 _15249_ (.S0(net6241),
    .A0(\top1.memory2.mem2[116][0] ),
    .A1(\top1.memory2.mem2[117][0] ),
    .A2(\top1.memory2.mem2[118][0] ),
    .A3(\top1.memory2.mem2[119][0] ),
    .S1(net6176),
    .X(_05646_));
 sg13g2_mux4_1 _15250_ (.S0(net6238),
    .A0(\top1.memory2.mem2[124][0] ),
    .A1(\top1.memory2.mem2[125][0] ),
    .A2(\top1.memory2.mem2[126][0] ),
    .A3(\top1.memory2.mem2[127][0] ),
    .S1(net6173),
    .X(_05647_));
 sg13g2_a22oi_1 _15251_ (.Y(_05648_),
    .B1(_05646_),
    .B2(net6030),
    .A2(_05644_),
    .A1(net5884));
 sg13g2_a22oi_1 _15252_ (.Y(_05649_),
    .B1(_05647_),
    .B2(net5860),
    .A2(_05645_),
    .A1(net6094));
 sg13g2_a21oi_2 _15253_ (.B1(net5839),
    .Y(_05650_),
    .A2(_05649_),
    .A1(_05648_));
 sg13g2_or2_2 _15254_ (.X(_05651_),
    .B(_05650_),
    .A(_05643_));
 sg13g2_mux4_1 _15255_ (.S0(net6201),
    .A0(\top1.memory2.mem2[92][0] ),
    .A1(\top1.memory2.mem2[93][0] ),
    .A2(\top1.memory2.mem2[94][0] ),
    .A3(\top1.memory2.mem2[95][0] ),
    .S1(net6138),
    .X(_05652_));
 sg13g2_o21ai_1 _15256_ (.B1(net6017),
    .Y(_05653_),
    .A1(\top1.memory2.mem2[84][0] ),
    .A2(net6040));
 sg13g2_nor2_1 _15257_ (.A(\top1.memory2.mem2[87][0] ),
    .B(net5933),
    .Y(_05654_));
 sg13g2_nor2_1 _15258_ (.A(\top1.memory2.mem2[85][0] ),
    .B(net5974),
    .Y(_05655_));
 sg13g2_nor2_1 _15259_ (.A(\top1.memory2.mem2[86][0] ),
    .B(net5895),
    .Y(_05656_));
 sg13g2_or4_1 _15260_ (.A(_05653_),
    .B(_05654_),
    .C(_05655_),
    .D(_05656_),
    .X(_05657_));
 sg13g2_mux4_1 _15261_ (.S0(net6201),
    .A0(\top1.memory2.mem2[80][0] ),
    .A1(\top1.memory2.mem2[81][0] ),
    .A2(\top1.memory2.mem2[82][0] ),
    .A3(\top1.memory2.mem2[83][0] ),
    .S1(net6137),
    .X(_05658_));
 sg13g2_a22oi_1 _15262_ (.Y(_05659_),
    .B1(net5911),
    .B2(\top1.memory2.mem2[90][0] ),
    .A2(net6056),
    .A1(\top1.memory2.mem2[88][0] ));
 sg13g2_a22oi_1 _15263_ (.Y(_05660_),
    .B1(net5951),
    .B2(\top1.memory2.mem2[91][0] ),
    .A2(net5993),
    .A1(\top1.memory2.mem2[89][0] ));
 sg13g2_a21o_1 _15264_ (.A2(_05660_),
    .A1(_05659_),
    .B1(net6075),
    .X(_05661_));
 sg13g2_a221oi_1 _15265_ (.B2(net5874),
    .C1(net6104),
    .B1(_05658_),
    .A1(net5852),
    .Y(_05662_),
    .A2(_05652_));
 sg13g2_nand3_1 _15266_ (.B(_05661_),
    .C(_05662_),
    .A(_05657_),
    .Y(_05663_));
 sg13g2_mux4_1 _15267_ (.S0(net6197),
    .A0(\top1.memory2.mem2[64][0] ),
    .A1(\top1.memory2.mem2[65][0] ),
    .A2(\top1.memory2.mem2[66][0] ),
    .A3(\top1.memory2.mem2[67][0] ),
    .S1(net6133),
    .X(_05664_));
 sg13g2_mux4_1 _15268_ (.S0(net6200),
    .A0(\top1.memory2.mem2[72][0] ),
    .A1(\top1.memory2.mem2[73][0] ),
    .A2(\top1.memory2.mem2[74][0] ),
    .A3(\top1.memory2.mem2[75][0] ),
    .S1(net6136),
    .X(_05665_));
 sg13g2_a21oi_1 _15269_ (.A1(_03854_),
    .A2(net5983),
    .Y(_05666_),
    .B1(net6011));
 sg13g2_nor3_1 _15270_ (.A(net6201),
    .B(net6137),
    .C(\top1.memory2.mem2[68][0] ),
    .Y(_05667_));
 sg13g2_a221oi_1 _15271_ (.B2(_03855_),
    .C1(_05667_),
    .B1(net5903),
    .A1(_03856_),
    .Y(_05668_),
    .A2(net5944));
 sg13g2_mux4_1 _15272_ (.S0(net6197),
    .A0(\top1.memory2.mem2[76][0] ),
    .A1(\top1.memory2.mem2[77][0] ),
    .A2(\top1.memory2.mem2[78][0] ),
    .A3(\top1.memory2.mem2[79][0] ),
    .S1(net6133),
    .X(_05669_));
 sg13g2_a22oi_1 _15273_ (.Y(_05670_),
    .B1(_05666_),
    .B2(_05668_),
    .A2(_05665_),
    .A1(net6086));
 sg13g2_a221oi_1 _15274_ (.B2(net5850),
    .C1(net6120),
    .B1(_05669_),
    .A1(net5873),
    .Y(_05671_),
    .A2(_05664_));
 sg13g2_a21oi_2 _15275_ (.B1(_05479_),
    .Y(_05672_),
    .A2(_05671_),
    .A1(_05670_));
 sg13g2_a221oi_1 _15276_ (.B2(_05672_),
    .C1(net6111),
    .B1(_05663_),
    .A1(net6113),
    .Y(_05673_),
    .A2(_05651_));
 sg13g2_o21ai_1 _15277_ (.B1(_05673_),
    .Y(_05674_),
    .A1(net6114),
    .A2(_05636_));
 sg13g2_mux4_1 _15278_ (.S0(net6204),
    .A0(\top1.memory2.mem2[140][0] ),
    .A1(\top1.memory2.mem2[141][0] ),
    .A2(\top1.memory2.mem2[142][0] ),
    .A3(\top1.memory2.mem2[143][0] ),
    .S1(net6140),
    .X(_05675_));
 sg13g2_mux4_1 _15279_ (.S0(net6204),
    .A0(\top1.memory2.mem2[136][0] ),
    .A1(\top1.memory2.mem2[137][0] ),
    .A2(\top1.memory2.mem2[138][0] ),
    .A3(\top1.memory2.mem2[139][0] ),
    .S1(net6140),
    .X(_05676_));
 sg13g2_mux4_1 _15280_ (.S0(net6204),
    .A0(\top1.memory2.mem2[128][0] ),
    .A1(\top1.memory2.mem2[129][0] ),
    .A2(\top1.memory2.mem2[130][0] ),
    .A3(\top1.memory2.mem2[131][0] ),
    .S1(net6140),
    .X(_05677_));
 sg13g2_nor2_1 _15281_ (.A(\top1.memory2.mem2[134][0] ),
    .B(net5892),
    .Y(_05678_));
 sg13g2_nor2_1 _15282_ (.A(\top1.memory2.mem2[133][0] ),
    .B(net5976),
    .Y(_05679_));
 sg13g2_nor2_1 _15283_ (.A(\top1.memory2.mem2[135][0] ),
    .B(net5931),
    .Y(_05680_));
 sg13g2_o21ai_1 _15284_ (.B1(net6020),
    .Y(_05681_),
    .A1(\top1.memory2.mem2[132][0] ),
    .A2(net6038));
 sg13g2_or4_1 _15285_ (.A(_05678_),
    .B(_05679_),
    .C(_05680_),
    .D(_05681_),
    .X(_05682_));
 sg13g2_a21o_1 _15286_ (.A2(_05677_),
    .A1(net5875),
    .B1(net6122),
    .X(_05683_));
 sg13g2_a221oi_1 _15287_ (.B2(net6084),
    .C1(_05683_),
    .B1(_05676_),
    .A1(net5851),
    .Y(_05684_),
    .A2(_05675_));
 sg13g2_a22oi_1 _15288_ (.Y(_05685_),
    .B1(net5953),
    .B2(_03860_),
    .A2(net5994),
    .A1(_03858_));
 sg13g2_a221oi_1 _15289_ (.B2(_03859_),
    .C1(net6011),
    .B1(net5913),
    .A1(_03857_),
    .Y(_05686_),
    .A2(net6058));
 sg13g2_mux4_1 _15290_ (.S0(net6206),
    .A0(\top1.memory2.mem2[156][0] ),
    .A1(\top1.memory2.mem2[157][0] ),
    .A2(\top1.memory2.mem2[158][0] ),
    .A3(\top1.memory2.mem2[159][0] ),
    .S1(net6142),
    .X(_05687_));
 sg13g2_mux4_1 _15291_ (.S0(net6205),
    .A0(\top1.memory2.mem2[144][0] ),
    .A1(\top1.memory2.mem2[145][0] ),
    .A2(\top1.memory2.mem2[146][0] ),
    .A3(\top1.memory2.mem2[147][0] ),
    .S1(net6141),
    .X(_05688_));
 sg13g2_mux4_1 _15292_ (.S0(net6215),
    .A0(\top1.memory2.mem2[152][0] ),
    .A1(\top1.memory2.mem2[153][0] ),
    .A2(\top1.memory2.mem2[154][0] ),
    .A3(\top1.memory2.mem2[155][0] ),
    .S1(net6150),
    .X(_05689_));
 sg13g2_a22oi_1 _15293_ (.Y(_05690_),
    .B1(_05688_),
    .B2(net5875),
    .A2(_05687_),
    .A1(net5852));
 sg13g2_a221oi_1 _15294_ (.B2(net6084),
    .C1(net6107),
    .B1(_05689_),
    .A1(_05685_),
    .Y(_05691_),
    .A2(_05686_));
 sg13g2_a221oi_1 _15295_ (.B2(_05691_),
    .C1(net6119),
    .B1(_05690_),
    .A1(_05682_),
    .Y(_05692_),
    .A2(_05684_));
 sg13g2_mux4_1 _15296_ (.S0(net6214),
    .A0(\top1.memory2.mem2[172][0] ),
    .A1(\top1.memory2.mem2[173][0] ),
    .A2(\top1.memory2.mem2[174][0] ),
    .A3(\top1.memory2.mem2[175][0] ),
    .S1(net6149),
    .X(_05693_));
 sg13g2_mux4_1 _15297_ (.S0(net6217),
    .A0(\top1.memory2.mem2[164][0] ),
    .A1(\top1.memory2.mem2[165][0] ),
    .A2(\top1.memory2.mem2[166][0] ),
    .A3(\top1.memory2.mem2[167][0] ),
    .S1(net6152),
    .X(_05694_));
 sg13g2_mux4_1 _15298_ (.S0(net6229),
    .A0(\top1.memory2.mem2[168][0] ),
    .A1(\top1.memory2.mem2[169][0] ),
    .A2(\top1.memory2.mem2[170][0] ),
    .A3(\top1.memory2.mem2[171][0] ),
    .S1(net6164),
    .X(_05695_));
 sg13g2_mux4_1 _15299_ (.S0(net6217),
    .A0(\top1.memory2.mem2[160][0] ),
    .A1(\top1.memory2.mem2[161][0] ),
    .A2(\top1.memory2.mem2[162][0] ),
    .A3(\top1.memory2.mem2[163][0] ),
    .S1(net6152),
    .X(_05696_));
 sg13g2_a22oi_1 _15300_ (.Y(_05697_),
    .B1(_05695_),
    .B2(net6089),
    .A2(_05693_),
    .A1(net5854));
 sg13g2_a22oi_1 _15301_ (.Y(_05698_),
    .B1(_05696_),
    .B2(net5879),
    .A2(_05694_),
    .A1(net6023));
 sg13g2_a21oi_2 _15302_ (.B1(net5836),
    .Y(_05699_),
    .A2(_05698_),
    .A1(_05697_));
 sg13g2_mux4_1 _15303_ (.S0(net6232),
    .A0(\top1.memory2.mem2[180][0] ),
    .A1(\top1.memory2.mem2[181][0] ),
    .A2(\top1.memory2.mem2[182][0] ),
    .A3(\top1.memory2.mem2[183][0] ),
    .S1(net6167),
    .X(_05700_));
 sg13g2_a22oi_1 _15304_ (.Y(_05701_),
    .B1(net5923),
    .B2(\top1.memory2.mem2[186][0] ),
    .A2(net5964),
    .A1(\top1.memory2.mem2[187][0] ));
 sg13g2_a22oi_1 _15305_ (.Y(_05702_),
    .B1(net6005),
    .B2(\top1.memory2.mem2[185][0] ),
    .A2(net6066),
    .A1(\top1.memory2.mem2[184][0] ));
 sg13g2_a21o_1 _15306_ (.A2(_05702_),
    .A1(_05701_),
    .B1(net6080),
    .X(_05703_));
 sg13g2_mux4_1 _15307_ (.S0(net6234),
    .A0(\top1.memory2.mem2[176][0] ),
    .A1(\top1.memory2.mem2[177][0] ),
    .A2(\top1.memory2.mem2[178][0] ),
    .A3(\top1.memory2.mem2[179][0] ),
    .S1(net6169),
    .X(_05704_));
 sg13g2_mux4_1 _15308_ (.S0(net6234),
    .A0(\top1.memory2.mem2[188][0] ),
    .A1(\top1.memory2.mem2[189][0] ),
    .A2(\top1.memory2.mem2[190][0] ),
    .A3(\top1.memory2.mem2[191][0] ),
    .S1(net6169),
    .X(_05705_));
 sg13g2_and2_1 _15309_ (.A(net5858),
    .B(_05705_),
    .X(_05706_));
 sg13g2_a221oi_1 _15310_ (.B2(net5889),
    .C1(_05706_),
    .B1(_05704_),
    .A1(net6028),
    .Y(_05707_),
    .A2(_05700_));
 sg13g2_a21oi_2 _15311_ (.B1(_05453_),
    .Y(_05708_),
    .A2(_05707_),
    .A1(_05703_));
 sg13g2_nor4_1 _15312_ (.A(net5831),
    .B(_05692_),
    .C(_05699_),
    .D(_05708_),
    .Y(_05709_));
 sg13g2_a22oi_1 _15313_ (.Y(_05710_),
    .B1(net5995),
    .B2(\top1.memory2.mem2[197][0] ),
    .A2(net6060),
    .A1(\top1.memory2.mem2[196][0] ));
 sg13g2_a221oi_1 _15314_ (.B2(\top1.memory2.mem2[198][0] ),
    .C1(_03827_),
    .B1(net5914),
    .A1(\top1.memory2.mem2[199][0] ),
    .Y(_05711_),
    .A2(net5954));
 sg13g2_a22oi_1 _15315_ (.Y(_05712_),
    .B1(net5914),
    .B2(\top1.memory2.mem2[194][0] ),
    .A2(net5954),
    .A1(\top1.memory2.mem2[195][0] ));
 sg13g2_a221oi_1 _15316_ (.B2(\top1.memory2.mem2[193][0] ),
    .C1(net6131),
    .B1(net5995),
    .A1(\top1.memory2.mem2[192][0] ),
    .Y(_05713_),
    .A2(net6060));
 sg13g2_a22oi_1 _15317_ (.Y(_05714_),
    .B1(_05712_),
    .B2(_05713_),
    .A2(_05711_),
    .A1(_05710_));
 sg13g2_o21ai_1 _15318_ (.B1(net6109),
    .Y(_05715_),
    .A1(_03979_),
    .A2(_05714_));
 sg13g2_nor2_1 _15319_ (.A(_05709_),
    .B(_05715_),
    .Y(_05716_));
 sg13g2_a21oi_1 _15320_ (.A1(_05674_),
    .A2(_05716_),
    .Y(_05717_),
    .B1(_03832_));
 sg13g2_a22oi_1 _15321_ (.Y(_01018_),
    .B1(_05582_),
    .B2(_05717_),
    .A2(_03849_),
    .A1(net6101));
 sg13g2_mux4_1 _15322_ (.S0(net6235),
    .A0(\top1.memory2.mem2[36][1] ),
    .A1(\top1.memory2.mem2[37][1] ),
    .A2(\top1.memory2.mem2[38][1] ),
    .A3(\top1.memory2.mem2[39][1] ),
    .S1(net6170),
    .X(_05718_));
 sg13g2_mux4_1 _15323_ (.S0(net6251),
    .A0(\top1.memory2.mem2[40][1] ),
    .A1(\top1.memory2.mem2[41][1] ),
    .A2(\top1.memory2.mem2[42][1] ),
    .A3(\top1.memory2.mem2[43][1] ),
    .S1(net6186),
    .X(_05719_));
 sg13g2_mux4_1 _15324_ (.S0(net6233),
    .A0(\top1.memory2.mem2[32][1] ),
    .A1(\top1.memory2.mem2[33][1] ),
    .A2(\top1.memory2.mem2[34][1] ),
    .A3(\top1.memory2.mem2[35][1] ),
    .S1(net6168),
    .X(_05720_));
 sg13g2_mux4_1 _15325_ (.S0(net6253),
    .A0(\top1.memory2.mem2[44][1] ),
    .A1(\top1.memory2.mem2[45][1] ),
    .A2(\top1.memory2.mem2[46][1] ),
    .A3(\top1.memory2.mem2[47][1] ),
    .S1(net6188),
    .X(_05721_));
 sg13g2_a22oi_1 _15326_ (.Y(_05722_),
    .B1(_05720_),
    .B2(net5883),
    .A2(_05718_),
    .A1(net6028));
 sg13g2_a22oi_1 _15327_ (.Y(_05723_),
    .B1(_05721_),
    .B2(net5862),
    .A2(_05719_),
    .A1(net6099));
 sg13g2_a21oi_1 _15328_ (.A1(_05722_),
    .A2(_05723_),
    .Y(_05724_),
    .B1(net5834));
 sg13g2_mux4_1 _15329_ (.S0(net6231),
    .A0(\top1.memory2.mem2[16][1] ),
    .A1(\top1.memory2.mem2[17][1] ),
    .A2(\top1.memory2.mem2[18][1] ),
    .A3(\top1.memory2.mem2[19][1] ),
    .S1(net6166),
    .X(_05725_));
 sg13g2_mux4_1 _15330_ (.S0(net6216),
    .A0(\top1.memory2.mem2[28][1] ),
    .A1(\top1.memory2.mem2[29][1] ),
    .A2(\top1.memory2.mem2[30][1] ),
    .A3(\top1.memory2.mem2[31][1] ),
    .S1(net6151),
    .X(_05726_));
 sg13g2_a22oi_1 _15331_ (.Y(_05727_),
    .B1(net5921),
    .B2(_03870_),
    .A2(net6068),
    .A1(_03868_));
 sg13g2_a221oi_1 _15332_ (.B2(_03871_),
    .C1(net6012),
    .B1(net5961),
    .A1(_03869_),
    .Y(_05728_),
    .A2(net6003));
 sg13g2_mux4_1 _15333_ (.S0(net6230),
    .A0(\top1.memory2.mem2[24][1] ),
    .A1(\top1.memory2.mem2[25][1] ),
    .A2(\top1.memory2.mem2[26][1] ),
    .A3(\top1.memory2.mem2[27][1] ),
    .S1(net6165),
    .X(_05729_));
 sg13g2_mux4_1 _15334_ (.S0(net6250),
    .A0(\top1.memory2.mem2[56][1] ),
    .A1(\top1.memory2.mem2[57][1] ),
    .A2(\top1.memory2.mem2[58][1] ),
    .A3(\top1.memory2.mem2[59][1] ),
    .S1(net6185),
    .X(_05730_));
 sg13g2_mux4_1 _15335_ (.S0(net6252),
    .A0(\top1.memory2.mem2[60][1] ),
    .A1(\top1.memory2.mem2[61][1] ),
    .A2(\top1.memory2.mem2[62][1] ),
    .A3(\top1.memory2.mem2[63][1] ),
    .S1(net6187),
    .X(_05731_));
 sg13g2_mux4_1 _15336_ (.S0(net6249),
    .A0(\top1.memory2.mem2[52][1] ),
    .A1(\top1.memory2.mem2[53][1] ),
    .A2(\top1.memory2.mem2[54][1] ),
    .A3(\top1.memory2.mem2[55][1] ),
    .S1(net6184),
    .X(_05732_));
 sg13g2_mux4_1 _15337_ (.S0(net6252),
    .A0(\top1.memory2.mem2[48][1] ),
    .A1(\top1.memory2.mem2[49][1] ),
    .A2(\top1.memory2.mem2[50][1] ),
    .A3(\top1.memory2.mem2[51][1] ),
    .S1(net6187),
    .X(_05733_));
 sg13g2_a22oi_1 _15338_ (.Y(_05734_),
    .B1(_05732_),
    .B2(net6034),
    .A2(_05730_),
    .A1(net6099));
 sg13g2_a22oi_1 _15339_ (.Y(_05735_),
    .B1(_05733_),
    .B2(net5888),
    .A2(_05731_),
    .A1(net5862));
 sg13g2_a21oi_2 _15340_ (.B1(net5840),
    .Y(_05736_),
    .A2(_05735_),
    .A1(_05734_));
 sg13g2_mux4_1 _15341_ (.S0(net6216),
    .A0(\top1.memory2.mem2[0][1] ),
    .A1(\top1.memory2.mem2[1][1] ),
    .A2(\top1.memory2.mem2[2][1] ),
    .A3(\top1.memory2.mem2[3][1] ),
    .S1(net6151),
    .X(_05737_));
 sg13g2_and2_1 _15342_ (.A(net5879),
    .B(_05737_),
    .X(_05738_));
 sg13g2_mux4_1 _15343_ (.S0(net6215),
    .A0(\top1.memory2.mem2[12][1] ),
    .A1(\top1.memory2.mem2[13][1] ),
    .A2(\top1.memory2.mem2[14][1] ),
    .A3(\top1.memory2.mem2[15][1] ),
    .S1(net6150),
    .X(_05739_));
 sg13g2_mux4_1 _15344_ (.S0(net6216),
    .A0(\top1.memory2.mem2[8][1] ),
    .A1(\top1.memory2.mem2[9][1] ),
    .A2(\top1.memory2.mem2[10][1] ),
    .A3(\top1.memory2.mem2[11][1] ),
    .S1(net6151),
    .X(_05740_));
 sg13g2_nor3_1 _15345_ (.A(net6218),
    .B(net6153),
    .C(\top1.memory2.mem2[4][1] ),
    .Y(_05741_));
 sg13g2_a21oi_1 _15346_ (.A1(_03867_),
    .A2(net5961),
    .Y(_05742_),
    .B1(net6013));
 sg13g2_a221oi_1 _15347_ (.B2(_03866_),
    .C1(_05741_),
    .B1(net5921),
    .A1(_03865_),
    .Y(_05743_),
    .A2(net6002));
 sg13g2_a22oi_1 _15348_ (.Y(_05744_),
    .B1(_05727_),
    .B2(_05728_),
    .A2(_05726_),
    .A1(net5854));
 sg13g2_a221oi_1 _15349_ (.B2(net6091),
    .C1(net6106),
    .B1(_05729_),
    .A1(net5883),
    .Y(_05745_),
    .A2(_05725_));
 sg13g2_a21oi_1 _15350_ (.A1(net6087),
    .A2(_05740_),
    .Y(_05746_),
    .B1(net6125));
 sg13g2_a221oi_1 _15351_ (.B2(_05743_),
    .C1(_05738_),
    .B1(_05742_),
    .A1(net5854),
    .Y(_05747_),
    .A2(_05739_));
 sg13g2_a221oi_1 _15352_ (.B2(_05747_),
    .C1(net6119),
    .B1(_05746_),
    .A1(_05744_),
    .Y(_05748_),
    .A2(_05745_));
 sg13g2_or2_2 _15353_ (.X(_05749_),
    .B(_05736_),
    .A(_05724_));
 sg13g2_o21ai_1 _15354_ (.B1(net6102),
    .Y(_05750_),
    .A1(_05748_),
    .A2(_05749_));
 sg13g2_mux4_1 _15355_ (.S0(net6198),
    .A0(\top1.memory2.mem2[72][1] ),
    .A1(\top1.memory2.mem2[73][1] ),
    .A2(\top1.memory2.mem2[74][1] ),
    .A3(\top1.memory2.mem2[75][1] ),
    .S1(net6134),
    .X(_05751_));
 sg13g2_a21o_1 _15356_ (.A2(_05751_),
    .A1(net6083),
    .B1(net6120),
    .X(_05752_));
 sg13g2_o21ai_1 _15357_ (.B1(net6016),
    .Y(_05753_),
    .A1(\top1.memory2.mem2[71][1] ),
    .A2(net5932));
 sg13g2_or3_1 _15358_ (.A(net6202),
    .B(net6138),
    .C(\top1.memory2.mem2[68][1] ),
    .X(_05754_));
 sg13g2_o21ai_1 _15359_ (.B1(_05754_),
    .Y(_05755_),
    .A1(\top1.memory2.mem2[69][1] ),
    .A2(net5970));
 sg13g2_nor2_1 _15360_ (.A(\top1.memory2.mem2[70][1] ),
    .B(net5893),
    .Y(_05756_));
 sg13g2_nor3_2 _15361_ (.A(_05753_),
    .B(_05755_),
    .C(_05756_),
    .Y(_05757_));
 sg13g2_a22oi_1 _15362_ (.Y(_05758_),
    .B1(net5901),
    .B2(\top1.memory2.mem2[78][1] ),
    .A2(net5942),
    .A1(\top1.memory2.mem2[79][1] ));
 sg13g2_a22oi_1 _15363_ (.Y(_05759_),
    .B1(net5981),
    .B2(\top1.memory2.mem2[77][1] ),
    .A2(net6046),
    .A1(\top1.memory2.mem2[76][1] ));
 sg13g2_a21oi_2 _15364_ (.B1(net5844),
    .Y(_05760_),
    .A2(_05759_),
    .A1(_05758_));
 sg13g2_a22oi_1 _15365_ (.Y(_05761_),
    .B1(net5902),
    .B2(\top1.memory2.mem2[66][1] ),
    .A2(net5942),
    .A1(\top1.memory2.mem2[67][1] ));
 sg13g2_a22oi_1 _15366_ (.Y(_05762_),
    .B1(net5981),
    .B2(\top1.memory2.mem2[65][1] ),
    .A2(net6047),
    .A1(\top1.memory2.mem2[64][1] ));
 sg13g2_a21oi_1 _15367_ (.A1(_05761_),
    .A2(_05762_),
    .Y(_05763_),
    .B1(net5868));
 sg13g2_nor4_2 _15368_ (.A(_05752_),
    .B(_05757_),
    .C(_05760_),
    .Y(_05764_),
    .D(_05763_));
 sg13g2_a22oi_1 _15369_ (.Y(_05765_),
    .B1(net5903),
    .B2(\top1.memory2.mem2[94][1] ),
    .A2(net5944),
    .A1(\top1.memory2.mem2[95][1] ));
 sg13g2_a22oi_1 _15370_ (.Y(_05766_),
    .B1(net5983),
    .B2(\top1.memory2.mem2[93][1] ),
    .A2(net6048),
    .A1(\top1.memory2.mem2[92][1] ));
 sg13g2_a21oi_1 _15371_ (.A1(_05765_),
    .A2(_05766_),
    .Y(_05767_),
    .B1(net5845));
 sg13g2_mux4_1 _15372_ (.S0(net6200),
    .A0(\top1.memory2.mem2[80][1] ),
    .A1(\top1.memory2.mem2[81][1] ),
    .A2(\top1.memory2.mem2[82][1] ),
    .A3(\top1.memory2.mem2[83][1] ),
    .S1(net6136),
    .X(_05768_));
 sg13g2_a22oi_1 _15373_ (.Y(_05769_),
    .B1(net5904),
    .B2(\top1.memory2.mem2[90][1] ),
    .A2(net6048),
    .A1(\top1.memory2.mem2[88][1] ));
 sg13g2_a22oi_1 _15374_ (.Y(_05770_),
    .B1(net5944),
    .B2(\top1.memory2.mem2[91][1] ),
    .A2(net5983),
    .A1(\top1.memory2.mem2[89][1] ));
 sg13g2_a21oi_1 _15375_ (.A1(_05769_),
    .A2(_05770_),
    .Y(_05771_),
    .B1(net6076));
 sg13g2_nor2_1 _15376_ (.A(\top1.memory2.mem2[87][1] ),
    .B(net5934),
    .Y(_05772_));
 sg13g2_nor2_1 _15377_ (.A(\top1.memory2.mem2[85][1] ),
    .B(net5972),
    .Y(_05773_));
 sg13g2_nor2_1 _15378_ (.A(\top1.memory2.mem2[84][1] ),
    .B(net6040),
    .Y(_05774_));
 sg13g2_o21ai_1 _15379_ (.B1(net6017),
    .Y(_05775_),
    .A1(\top1.memory2.mem2[86][1] ),
    .A2(net5895));
 sg13g2_nor4_2 _15380_ (.A(_05772_),
    .B(_05773_),
    .C(_05774_),
    .Y(_05776_),
    .D(_05775_));
 sg13g2_a21o_1 _15381_ (.A2(_05768_),
    .A1(net5874),
    .B1(net6104),
    .X(_05777_));
 sg13g2_nor4_1 _15382_ (.A(_05767_),
    .B(_05771_),
    .C(_05776_),
    .D(_05777_),
    .Y(_05778_));
 sg13g2_or3_2 _15383_ (.A(_05479_),
    .B(_05764_),
    .C(_05778_),
    .X(_05779_));
 sg13g2_mux4_1 _15384_ (.S0(net6246),
    .A0(\top1.memory2.mem2[112][1] ),
    .A1(\top1.memory2.mem2[113][1] ),
    .A2(\top1.memory2.mem2[114][1] ),
    .A3(\top1.memory2.mem2[115][1] ),
    .S1(net6181),
    .X(_05780_));
 sg13g2_mux4_1 _15385_ (.S0(net6237),
    .A0(\top1.memory2.mem2[124][1] ),
    .A1(\top1.memory2.mem2[125][1] ),
    .A2(\top1.memory2.mem2[126][1] ),
    .A3(\top1.memory2.mem2[127][1] ),
    .S1(net6172),
    .X(_05781_));
 sg13g2_mux4_1 _15386_ (.S0(net6241),
    .A0(\top1.memory2.mem2[116][1] ),
    .A1(\top1.memory2.mem2[117][1] ),
    .A2(\top1.memory2.mem2[118][1] ),
    .A3(\top1.memory2.mem2[119][1] ),
    .S1(net6176),
    .X(_05782_));
 sg13g2_mux4_1 _15387_ (.S0(net6240),
    .A0(\top1.memory2.mem2[120][1] ),
    .A1(\top1.memory2.mem2[121][1] ),
    .A2(\top1.memory2.mem2[122][1] ),
    .A3(\top1.memory2.mem2[123][1] ),
    .S1(net6175),
    .X(_05783_));
 sg13g2_a22oi_1 _15388_ (.Y(_05784_),
    .B1(_05782_),
    .B2(net6032),
    .A2(_05780_),
    .A1(net5885));
 sg13g2_a22oi_1 _15389_ (.Y(_05785_),
    .B1(_05783_),
    .B2(net6094),
    .A2(_05781_),
    .A1(net5860));
 sg13g2_a21oi_2 _15390_ (.B1(net5838),
    .Y(_05786_),
    .A2(_05785_),
    .A1(_05784_));
 sg13g2_mux4_1 _15391_ (.S0(net6223),
    .A0(\top1.memory2.mem2[96][1] ),
    .A1(\top1.memory2.mem2[97][1] ),
    .A2(\top1.memory2.mem2[98][1] ),
    .A3(\top1.memory2.mem2[99][1] ),
    .S1(net6158),
    .X(_05787_));
 sg13g2_mux4_1 _15392_ (.S0(net6236),
    .A0(\top1.memory2.mem2[108][1] ),
    .A1(\top1.memory2.mem2[109][1] ),
    .A2(\top1.memory2.mem2[110][1] ),
    .A3(\top1.memory2.mem2[111][1] ),
    .S1(net6171),
    .X(_05788_));
 sg13g2_and2_1 _15393_ (.A(net5859),
    .B(_05788_),
    .X(_05789_));
 sg13g2_mux4_1 _15394_ (.S0(net6223),
    .A0(\top1.memory2.mem2[100][1] ),
    .A1(\top1.memory2.mem2[101][1] ),
    .A2(\top1.memory2.mem2[102][1] ),
    .A3(\top1.memory2.mem2[103][1] ),
    .S1(net6158),
    .X(_05790_));
 sg13g2_a22oi_1 _15395_ (.Y(_05791_),
    .B1(net5929),
    .B2(\top1.memory2.mem2[106][1] ),
    .A2(net5969),
    .A1(\top1.memory2.mem2[107][1] ));
 sg13g2_a22oi_1 _15396_ (.Y(_05792_),
    .B1(net6009),
    .B2(\top1.memory2.mem2[105][1] ),
    .A2(net6073),
    .A1(\top1.memory2.mem2[104][1] ));
 sg13g2_a21o_1 _15397_ (.A2(_05792_),
    .A1(_05791_),
    .B1(net6082),
    .X(_05793_));
 sg13g2_a221oi_1 _15398_ (.B2(net6031),
    .C1(_05789_),
    .B1(_05790_),
    .A1(net5885),
    .Y(_05794_),
    .A2(_05787_));
 sg13g2_a21oi_1 _15399_ (.A1(_05793_),
    .A2(_05794_),
    .Y(_05795_),
    .B1(net5832));
 sg13g2_o21ai_1 _15400_ (.B1(net6116),
    .Y(_05796_),
    .A1(_05786_),
    .A2(_05795_));
 sg13g2_nand4_1 _15401_ (.B(_05750_),
    .C(_05779_),
    .A(_03831_),
    .Y(_05797_),
    .D(_05796_));
 sg13g2_a22oi_1 _15402_ (.Y(_05798_),
    .B1(net5906),
    .B2(\top1.memory2.mem2[138][1] ),
    .A2(net5947),
    .A1(\top1.memory2.mem2[139][1] ));
 sg13g2_a22oi_1 _15403_ (.Y(_05799_),
    .B1(net5987),
    .B2(\top1.memory2.mem2[137][1] ),
    .A2(net6051),
    .A1(\top1.memory2.mem2[136][1] ));
 sg13g2_a21oi_1 _15404_ (.A1(_05798_),
    .A2(_05799_),
    .Y(_05800_),
    .B1(net6076));
 sg13g2_nor2_1 _15405_ (.A(\top1.memory2.mem2[133][1] ),
    .B(net5972),
    .Y(_05801_));
 sg13g2_nor2_1 _15406_ (.A(\top1.memory2.mem2[134][1] ),
    .B(net5892),
    .Y(_05802_));
 sg13g2_nor2_1 _15407_ (.A(\top1.memory2.mem2[132][1] ),
    .B(net6038),
    .Y(_05803_));
 sg13g2_o21ai_1 _15408_ (.B1(net6020),
    .Y(_05804_),
    .A1(\top1.memory2.mem2[135][1] ),
    .A2(net5930));
 sg13g2_nor4_1 _15409_ (.A(_05801_),
    .B(_05802_),
    .C(_05803_),
    .D(_05804_),
    .Y(_05805_));
 sg13g2_a22oi_1 _15410_ (.Y(_05806_),
    .B1(net5905),
    .B2(\top1.memory2.mem2[130][1] ),
    .A2(net5946),
    .A1(\top1.memory2.mem2[131][1] ));
 sg13g2_a22oi_1 _15411_ (.Y(_05807_),
    .B1(net5986),
    .B2(\top1.memory2.mem2[129][1] ),
    .A2(net6051),
    .A1(\top1.memory2.mem2[128][1] ));
 sg13g2_a21oi_1 _15412_ (.A1(_05806_),
    .A2(_05807_),
    .Y(_05808_),
    .B1(net5867));
 sg13g2_a22oi_1 _15413_ (.Y(_05809_),
    .B1(net5905),
    .B2(\top1.memory2.mem2[142][1] ),
    .A2(net5986),
    .A1(\top1.memory2.mem2[141][1] ));
 sg13g2_a22oi_1 _15414_ (.Y(_05810_),
    .B1(net5946),
    .B2(\top1.memory2.mem2[143][1] ),
    .A2(net6050),
    .A1(\top1.memory2.mem2[140][1] ));
 sg13g2_a21oi_1 _15415_ (.A1(_05809_),
    .A2(_05810_),
    .Y(_05811_),
    .B1(net5842));
 sg13g2_nor4_2 _15416_ (.A(_05800_),
    .B(_05805_),
    .C(_05808_),
    .Y(_05812_),
    .D(_05811_));
 sg13g2_o21ai_1 _15417_ (.B1(_05514_),
    .Y(_05813_),
    .A1(_03977_),
    .A2(_05812_));
 sg13g2_a22oi_1 _15418_ (.Y(_05814_),
    .B1(net5913),
    .B2(\top1.memory2.mem2[158][1] ),
    .A2(net5953),
    .A1(\top1.memory2.mem2[159][1] ));
 sg13g2_a22oi_1 _15419_ (.Y(_05815_),
    .B1(net5994),
    .B2(\top1.memory2.mem2[157][1] ),
    .A2(net6058),
    .A1(\top1.memory2.mem2[156][1] ));
 sg13g2_a21oi_1 _15420_ (.A1(_05814_),
    .A2(_05815_),
    .Y(_05816_),
    .B1(net5845));
 sg13g2_a22oi_1 _15421_ (.Y(_05817_),
    .B1(net5913),
    .B2(\top1.memory2.mem2[154][1] ),
    .A2(net5953),
    .A1(\top1.memory2.mem2[155][1] ));
 sg13g2_a22oi_1 _15422_ (.Y(_05818_),
    .B1(net5994),
    .B2(\top1.memory2.mem2[153][1] ),
    .A2(net6058),
    .A1(\top1.memory2.mem2[152][1] ));
 sg13g2_a21oi_1 _15423_ (.A1(_05817_),
    .A2(_05818_),
    .Y(_05819_),
    .B1(net6078));
 sg13g2_nor2_1 _15424_ (.A(\top1.memory2.mem2[148][1] ),
    .B(net6042),
    .Y(_05820_));
 sg13g2_nor2_1 _15425_ (.A(\top1.memory2.mem2[149][1] ),
    .B(net5975),
    .Y(_05821_));
 sg13g2_nor2_1 _15426_ (.A(\top1.memory2.mem2[151][1] ),
    .B(net5935),
    .Y(_05822_));
 sg13g2_o21ai_1 _15427_ (.B1(net6024),
    .Y(_05823_),
    .A1(\top1.memory2.mem2[150][1] ),
    .A2(net5896));
 sg13g2_nor4_2 _15428_ (.A(_05820_),
    .B(_05821_),
    .C(_05822_),
    .Y(_05824_),
    .D(_05823_));
 sg13g2_a22oi_1 _15429_ (.Y(_05825_),
    .B1(net5913),
    .B2(\top1.memory2.mem2[146][1] ),
    .A2(net5953),
    .A1(\top1.memory2.mem2[147][1] ));
 sg13g2_a22oi_1 _15430_ (.Y(_05826_),
    .B1(net5994),
    .B2(\top1.memory2.mem2[145][1] ),
    .A2(net6058),
    .A1(\top1.memory2.mem2[144][1] ));
 sg13g2_a21oi_1 _15431_ (.A1(_05825_),
    .A2(_05826_),
    .Y(_05827_),
    .B1(net5869));
 sg13g2_or4_2 _15432_ (.A(_05816_),
    .B(_05819_),
    .C(_05824_),
    .D(_05827_),
    .X(_05828_));
 sg13g2_a22oi_1 _15433_ (.Y(_05829_),
    .B1(net5922),
    .B2(\top1.memory2.mem2[162][1] ),
    .A2(net5962),
    .A1(\top1.memory2.mem2[163][1] ));
 sg13g2_a22oi_1 _15434_ (.Y(_05830_),
    .B1(net5996),
    .B2(\top1.memory2.mem2[161][1] ),
    .A2(net6061),
    .A1(\top1.memory2.mem2[160][1] ));
 sg13g2_a21oi_1 _15435_ (.A1(_05829_),
    .A2(_05830_),
    .Y(_05831_),
    .B1(net5870));
 sg13g2_a22oi_1 _15436_ (.Y(_05832_),
    .B1(net5922),
    .B2(\top1.memory2.mem2[166][1] ),
    .A2(net5962),
    .A1(\top1.memory2.mem2[167][1] ));
 sg13g2_a22oi_1 _15437_ (.Y(_05833_),
    .B1(net6003),
    .B2(\top1.memory2.mem2[165][1] ),
    .A2(net6065),
    .A1(\top1.memory2.mem2[164][1] ));
 sg13g2_a21oi_1 _15438_ (.A1(_05832_),
    .A2(_05833_),
    .Y(_05834_),
    .B1(net6013));
 sg13g2_a22oi_1 _15439_ (.Y(_05835_),
    .B1(net5922),
    .B2(\top1.memory2.mem2[170][1] ),
    .A2(net5962),
    .A1(\top1.memory2.mem2[171][1] ));
 sg13g2_a22oi_1 _15440_ (.Y(_05836_),
    .B1(net6003),
    .B2(\top1.memory2.mem2[169][1] ),
    .A2(net6065),
    .A1(\top1.memory2.mem2[168][1] ));
 sg13g2_a21oi_1 _15441_ (.A1(_05835_),
    .A2(_05836_),
    .Y(_05837_),
    .B1(net6080));
 sg13g2_a22oi_1 _15442_ (.Y(_05838_),
    .B1(net5918),
    .B2(\top1.memory2.mem2[174][1] ),
    .A2(net5958),
    .A1(\top1.memory2.mem2[175][1] ));
 sg13g2_a22oi_1 _15443_ (.Y(_05839_),
    .B1(net6001),
    .B2(\top1.memory2.mem2[173][1] ),
    .A2(net6064),
    .A1(\top1.memory2.mem2[172][1] ));
 sg13g2_a21oi_2 _15444_ (.B1(net5847),
    .Y(_05840_),
    .A2(_05839_),
    .A1(_05838_));
 sg13g2_or4_1 _15445_ (.A(_05831_),
    .B(_05834_),
    .C(_05837_),
    .D(_05840_),
    .X(_05841_));
 sg13g2_mux4_1 _15446_ (.S0(net6234),
    .A0(\top1.memory2.mem2[176][1] ),
    .A1(\top1.memory2.mem2[177][1] ),
    .A2(\top1.memory2.mem2[178][1] ),
    .A3(\top1.memory2.mem2[179][1] ),
    .S1(net6169),
    .X(_05842_));
 sg13g2_mux4_1 _15447_ (.S0(net6232),
    .A0(\top1.memory2.mem2[180][1] ),
    .A1(\top1.memory2.mem2[181][1] ),
    .A2(\top1.memory2.mem2[182][1] ),
    .A3(\top1.memory2.mem2[183][1] ),
    .S1(net6167),
    .X(_05843_));
 sg13g2_mux4_1 _15448_ (.S0(net6230),
    .A0(\top1.memory2.mem2[184][1] ),
    .A1(\top1.memory2.mem2[185][1] ),
    .A2(\top1.memory2.mem2[186][1] ),
    .A3(\top1.memory2.mem2[187][1] ),
    .S1(net6165),
    .X(_05844_));
 sg13g2_mux4_1 _15449_ (.S0(net6232),
    .A0(\top1.memory2.mem2[188][1] ),
    .A1(\top1.memory2.mem2[189][1] ),
    .A2(\top1.memory2.mem2[190][1] ),
    .A3(\top1.memory2.mem2[191][1] ),
    .S1(net6167),
    .X(_05845_));
 sg13g2_a22oi_1 _15450_ (.Y(_05846_),
    .B1(_05844_),
    .B2(net6092),
    .A2(_05842_),
    .A1(net5883));
 sg13g2_a22oi_1 _15451_ (.Y(_05847_),
    .B1(_05845_),
    .B2(net5858),
    .A2(_05843_),
    .A1(net6028));
 sg13g2_a21oi_2 _15452_ (.B1(net5837),
    .Y(_05848_),
    .A2(_05847_),
    .A1(_05846_));
 sg13g2_a221oi_1 _15453_ (.B2(_05443_),
    .C1(_05848_),
    .B1(_05841_),
    .A1(_05516_),
    .Y(_05849_),
    .A2(_05828_));
 sg13g2_nand2b_1 _15454_ (.Y(_05850_),
    .B(_05849_),
    .A_N(_05813_));
 sg13g2_nor2_1 _15455_ (.A(\top1.memory2.mem2[198][1] ),
    .B(net5898),
    .Y(_05851_));
 sg13g2_nor2_1 _15456_ (.A(\top1.memory2.mem2[197][1] ),
    .B(net5978),
    .Y(_05852_));
 sg13g2_nor2_1 _15457_ (.A(\top1.memory2.mem2[199][1] ),
    .B(net5937),
    .Y(_05853_));
 sg13g2_o21ai_1 _15458_ (.B1(net6132),
    .Y(_05854_),
    .A1(\top1.memory2.mem2[196][1] ),
    .A2(net6043));
 sg13g2_or4_1 _15459_ (.A(_05851_),
    .B(_05852_),
    .C(_05853_),
    .D(_05854_),
    .X(_05855_));
 sg13g2_nor2_1 _15460_ (.A(\top1.memory2.mem2[193][1] ),
    .B(net5975),
    .Y(_05856_));
 sg13g2_nor2_1 _15461_ (.A(\top1.memory2.mem2[195][1] ),
    .B(net5939),
    .Y(_05857_));
 sg13g2_o21ai_1 _15462_ (.B1(_03827_),
    .Y(_05858_),
    .A1(\top1.memory2.mem2[192][1] ),
    .A2(net6041));
 sg13g2_nor3_1 _15463_ (.A(_05856_),
    .B(_05857_),
    .C(_05858_),
    .Y(_05859_));
 sg13g2_o21ai_1 _15464_ (.B1(_05859_),
    .Y(_05860_),
    .A1(\top1.memory2.mem2[194][1] ),
    .A2(net5898));
 sg13g2_nand3_1 _15465_ (.B(_05855_),
    .C(_05860_),
    .A(_03978_),
    .Y(_05861_));
 sg13g2_nand4_1 _15466_ (.B(_05797_),
    .C(_05850_),
    .A(net6108),
    .Y(_05862_),
    .D(_05861_));
 sg13g2_mux4_1 _15467_ (.S0(net6245),
    .A0(\top1.memory2.mem1[60][1] ),
    .A1(\top1.memory2.mem1[61][1] ),
    .A2(\top1.memory2.mem1[62][1] ),
    .A3(\top1.memory2.mem1[63][1] ),
    .S1(net6180),
    .X(_05863_));
 sg13g2_mux4_1 _15468_ (.S0(net6255),
    .A0(\top1.memory2.mem1[48][1] ),
    .A1(\top1.memory2.mem1[49][1] ),
    .A2(\top1.memory2.mem1[50][1] ),
    .A3(\top1.memory2.mem1[51][1] ),
    .S1(net6190),
    .X(_05864_));
 sg13g2_a22oi_1 _15469_ (.Y(_05865_),
    .B1(_05864_),
    .B2(net5886),
    .A2(_05863_),
    .A1(net5864));
 sg13g2_mux4_1 _15470_ (.S0(net6250),
    .A0(\top1.memory2.mem1[56][1] ),
    .A1(\top1.memory2.mem1[57][1] ),
    .A2(\top1.memory2.mem1[58][1] ),
    .A3(\top1.memory2.mem1[59][1] ),
    .S1(net6185),
    .X(_05866_));
 sg13g2_mux4_1 _15471_ (.S0(net6254),
    .A0(\top1.memory2.mem1[52][1] ),
    .A1(\top1.memory2.mem1[53][1] ),
    .A2(\top1.memory2.mem1[54][1] ),
    .A3(\top1.memory2.mem1[55][1] ),
    .S1(net6189),
    .X(_05867_));
 sg13g2_a22oi_1 _15472_ (.Y(_05868_),
    .B1(_05867_),
    .B2(net6033),
    .A2(_05866_),
    .A1(net6097));
 sg13g2_a21oi_2 _15473_ (.B1(net5841),
    .Y(_05869_),
    .A2(_05868_),
    .A1(_05865_));
 sg13g2_mux4_1 _15474_ (.S0(net6214),
    .A0(\top1.memory2.mem1[8][1] ),
    .A1(\top1.memory2.mem1[9][1] ),
    .A2(\top1.memory2.mem1[10][1] ),
    .A3(\top1.memory2.mem1[11][1] ),
    .S1(net6149),
    .X(_05870_));
 sg13g2_mux4_1 _15475_ (.S0(net6211),
    .A0(\top1.memory2.mem1[0][1] ),
    .A1(\top1.memory2.mem1[1][1] ),
    .A2(\top1.memory2.mem1[2][1] ),
    .A3(\top1.memory2.mem1[3][1] ),
    .S1(net6146),
    .X(_05871_));
 sg13g2_nand2_1 _15476_ (.Y(_05872_),
    .A(net5878),
    .B(_05871_));
 sg13g2_mux4_1 _15477_ (.S0(net6213),
    .A0(\top1.memory2.mem1[12][1] ),
    .A1(\top1.memory2.mem1[13][1] ),
    .A2(\top1.memory2.mem1[14][1] ),
    .A3(\top1.memory2.mem1[15][1] ),
    .S1(net6148),
    .X(_05873_));
 sg13g2_o21ai_1 _15478_ (.B1(net6022),
    .Y(_05874_),
    .A1(\top1.memory2.mem1[6][1] ),
    .A2(net5897));
 sg13g2_nor2_1 _15479_ (.A(\top1.memory2.mem1[5][1] ),
    .B(net5978),
    .Y(_05875_));
 sg13g2_nor2_1 _15480_ (.A(\top1.memory2.mem1[4][1] ),
    .B(net6043),
    .Y(_05876_));
 sg13g2_nor2_1 _15481_ (.A(\top1.memory2.mem1[7][1] ),
    .B(net5938),
    .Y(_05877_));
 sg13g2_nor4_1 _15482_ (.A(_05874_),
    .B(_05875_),
    .C(_05876_),
    .D(_05877_),
    .Y(_05878_));
 sg13g2_a22oi_1 _15483_ (.Y(_05879_),
    .B1(_05873_),
    .B2(net5855),
    .A2(_05870_),
    .A1(net6087));
 sg13g2_nand2_2 _15484_ (.Y(_05880_),
    .A(_05872_),
    .B(_05879_));
 sg13g2_o21ai_1 _15485_ (.B1(_03976_),
    .Y(_05881_),
    .A1(_05878_),
    .A2(_05880_));
 sg13g2_mux4_1 _15486_ (.S0(net6258),
    .A0(\top1.memory2.mem1[36][1] ),
    .A1(\top1.memory2.mem1[37][1] ),
    .A2(\top1.memory2.mem1[38][1] ),
    .A3(\top1.memory2.mem1[39][1] ),
    .S1(net6193),
    .X(_05882_));
 sg13g2_mux4_1 _15487_ (.S0(net6259),
    .A0(\top1.memory2.mem1[44][1] ),
    .A1(\top1.memory2.mem1[45][1] ),
    .A2(\top1.memory2.mem1[46][1] ),
    .A3(\top1.memory2.mem1[47][1] ),
    .S1(net6194),
    .X(_05883_));
 sg13g2_a22oi_1 _15488_ (.Y(_05884_),
    .B1(_05883_),
    .B2(net5865),
    .A2(_05882_),
    .A1(net6034));
 sg13g2_mux4_1 _15489_ (.S0(net6257),
    .A0(\top1.memory2.mem1[40][1] ),
    .A1(\top1.memory2.mem1[41][1] ),
    .A2(\top1.memory2.mem1[42][1] ),
    .A3(\top1.memory2.mem1[43][1] ),
    .S1(net6192),
    .X(_05885_));
 sg13g2_mux4_1 _15490_ (.S0(net6258),
    .A0(\top1.memory2.mem1[32][1] ),
    .A1(\top1.memory2.mem1[33][1] ),
    .A2(\top1.memory2.mem1[34][1] ),
    .A3(\top1.memory2.mem1[35][1] ),
    .S1(net6193),
    .X(_05886_));
 sg13g2_a22oi_1 _15491_ (.Y(_05887_),
    .B1(_05886_),
    .B2(net5887),
    .A2(_05885_),
    .A1(net6098));
 sg13g2_a21oi_2 _15492_ (.B1(net5835),
    .Y(_05888_),
    .A2(_05887_),
    .A1(_05884_));
 sg13g2_mux4_1 _15493_ (.S0(net6232),
    .A0(\top1.memory2.mem1[24][1] ),
    .A1(\top1.memory2.mem1[25][1] ),
    .A2(\top1.memory2.mem1[26][1] ),
    .A3(\top1.memory2.mem1[27][1] ),
    .S1(net6167),
    .X(_05889_));
 sg13g2_a22oi_1 _15494_ (.Y(_05890_),
    .B1(net5959),
    .B2(_03864_),
    .A2(net6000),
    .A1(_03862_));
 sg13g2_a221oi_1 _15495_ (.B2(_03863_),
    .C1(net6012),
    .B1(net5919),
    .A1(_03861_),
    .Y(_05891_),
    .A2(net6064));
 sg13g2_mux4_1 _15496_ (.S0(net6229),
    .A0(\top1.memory2.mem1[16][1] ),
    .A1(\top1.memory2.mem1[17][1] ),
    .A2(\top1.memory2.mem1[18][1] ),
    .A3(\top1.memory2.mem1[19][1] ),
    .S1(net6164),
    .X(_05892_));
 sg13g2_and2_1 _15497_ (.A(net5882),
    .B(_05892_),
    .X(_05893_));
 sg13g2_a22oi_1 _15498_ (.Y(_05894_),
    .B1(net5959),
    .B2(\top1.memory2.mem1[31][1] ),
    .A2(net6000),
    .A1(\top1.memory2.mem1[29][1] ));
 sg13g2_a22oi_1 _15499_ (.Y(_05895_),
    .B1(net5919),
    .B2(\top1.memory2.mem1[30][1] ),
    .A2(net6064),
    .A1(\top1.memory2.mem1[28][1] ));
 sg13g2_a21o_1 _15500_ (.A2(_05895_),
    .A1(_05894_),
    .B1(net5847),
    .X(_05896_));
 sg13g2_a221oi_1 _15501_ (.B2(_05891_),
    .C1(_05893_),
    .B1(_05890_),
    .A1(net6091),
    .Y(_05897_),
    .A2(_05889_));
 sg13g2_a21o_1 _15502_ (.A2(_05897_),
    .A1(_05896_),
    .B1(_05517_),
    .X(_05898_));
 sg13g2_mux4_1 _15503_ (.S0(net6199),
    .A0(\top1.memory2.mem1[72][1] ),
    .A1(\top1.memory2.mem1[73][1] ),
    .A2(\top1.memory2.mem1[74][1] ),
    .A3(\top1.memory2.mem1[75][1] ),
    .S1(net6135),
    .X(_05899_));
 sg13g2_nor2_1 _15504_ (.A(\top1.memory2.mem1[69][1] ),
    .B(net5971),
    .Y(_05900_));
 sg13g2_nor2_1 _15505_ (.A(\top1.memory2.mem1[71][1] ),
    .B(net5932),
    .Y(_05901_));
 sg13g2_nor2_1 _15506_ (.A(\top1.memory2.mem1[70][1] ),
    .B(net5893),
    .Y(_05902_));
 sg13g2_o21ai_1 _15507_ (.B1(net6016),
    .Y(_05903_),
    .A1(\top1.memory2.mem1[68][1] ),
    .A2(net6037));
 sg13g2_nor4_2 _15508_ (.A(_05900_),
    .B(_05901_),
    .C(_05902_),
    .Y(_05904_),
    .D(_05903_));
 sg13g2_mux4_1 _15509_ (.S0(net6198),
    .A0(\top1.memory2.mem1[64][1] ),
    .A1(\top1.memory2.mem1[65][1] ),
    .A2(\top1.memory2.mem1[66][1] ),
    .A3(\top1.memory2.mem1[67][1] ),
    .S1(net6134),
    .X(_05905_));
 sg13g2_mux4_1 _15510_ (.S0(net6199),
    .A0(\top1.memory2.mem1[76][1] ),
    .A1(\top1.memory2.mem1[77][1] ),
    .A2(\top1.memory2.mem1[78][1] ),
    .A3(\top1.memory2.mem1[79][1] ),
    .S1(net6135),
    .X(_05906_));
 sg13g2_nand2_1 _15511_ (.Y(_05907_),
    .A(net5850),
    .B(_05906_));
 sg13g2_a22oi_1 _15512_ (.Y(_05908_),
    .B1(_05905_),
    .B2(net5873),
    .A2(_05899_),
    .A1(net6083));
 sg13g2_nand2_2 _15513_ (.Y(_05909_),
    .A(_05907_),
    .B(_05908_));
 sg13g2_o21ai_1 _15514_ (.B1(_03976_),
    .Y(_05910_),
    .A1(_05904_),
    .A2(_05909_));
 sg13g2_mux4_1 _15515_ (.S0(net6246),
    .A0(\top1.memory2.mem1[124][1] ),
    .A1(\top1.memory2.mem1[125][1] ),
    .A2(\top1.memory2.mem1[126][1] ),
    .A3(\top1.memory2.mem1[127][1] ),
    .S1(net6181),
    .X(_05911_));
 sg13g2_mux4_1 _15516_ (.S0(net6243),
    .A0(\top1.memory2.mem1[116][1] ),
    .A1(\top1.memory2.mem1[117][1] ),
    .A2(\top1.memory2.mem1[118][1] ),
    .A3(\top1.memory2.mem1[119][1] ),
    .S1(net6178),
    .X(_05912_));
 sg13g2_mux4_1 _15517_ (.S0(net6242),
    .A0(\top1.memory2.mem1[120][1] ),
    .A1(\top1.memory2.mem1[121][1] ),
    .A2(\top1.memory2.mem1[122][1] ),
    .A3(\top1.memory2.mem1[123][1] ),
    .S1(net6177),
    .X(_05913_));
 sg13g2_mux4_1 _15518_ (.S0(net6245),
    .A0(\top1.memory2.mem1[112][1] ),
    .A1(\top1.memory2.mem1[113][1] ),
    .A2(\top1.memory2.mem1[114][1] ),
    .A3(\top1.memory2.mem1[115][1] ),
    .S1(net6180),
    .X(_05914_));
 sg13g2_a22oi_1 _15519_ (.Y(_05915_),
    .B1(_05913_),
    .B2(net6095),
    .A2(_05911_),
    .A1(net5861));
 sg13g2_a22oi_1 _15520_ (.Y(_05916_),
    .B1(_05914_),
    .B2(net5884),
    .A2(_05912_),
    .A1(net6032));
 sg13g2_a21oi_2 _15521_ (.B1(net5839),
    .Y(_05917_),
    .A2(_05916_),
    .A1(_05915_));
 sg13g2_mux4_1 _15522_ (.S0(net6239),
    .A0(\top1.memory2.mem1[108][1] ),
    .A1(\top1.memory2.mem1[109][1] ),
    .A2(\top1.memory2.mem1[110][1] ),
    .A3(\top1.memory2.mem1[111][1] ),
    .S1(net6174),
    .X(_05918_));
 sg13g2_mux4_1 _15523_ (.S0(net6249),
    .A0(\top1.memory2.mem1[104][1] ),
    .A1(\top1.memory2.mem1[105][1] ),
    .A2(\top1.memory2.mem1[106][1] ),
    .A3(\top1.memory2.mem1[107][1] ),
    .S1(net6184),
    .X(_05919_));
 sg13g2_a22oi_1 _15524_ (.Y(_05920_),
    .B1(_05919_),
    .B2(net6096),
    .A2(_05918_),
    .A1(net5863));
 sg13g2_mux4_1 _15525_ (.S0(net6226),
    .A0(\top1.memory2.mem1[96][1] ),
    .A1(\top1.memory2.mem1[97][1] ),
    .A2(\top1.memory2.mem1[98][1] ),
    .A3(\top1.memory2.mem1[99][1] ),
    .S1(net6161),
    .X(_05921_));
 sg13g2_mux4_1 _15526_ (.S0(net6226),
    .A0(\top1.memory2.mem1[100][1] ),
    .A1(\top1.memory2.mem1[101][1] ),
    .A2(\top1.memory2.mem1[102][1] ),
    .A3(\top1.memory2.mem1[103][1] ),
    .S1(net6161),
    .X(_05922_));
 sg13g2_a22oi_1 _15527_ (.Y(_05923_),
    .B1(_05922_),
    .B2(net6025),
    .A2(_05921_),
    .A1(net5880));
 sg13g2_a21oi_1 _15528_ (.A1(_05920_),
    .A2(_05923_),
    .Y(_05924_),
    .B1(net5832));
 sg13g2_mux4_1 _15529_ (.S0(net6209),
    .A0(\top1.memory2.mem1[80][1] ),
    .A1(\top1.memory2.mem1[81][1] ),
    .A2(\top1.memory2.mem1[82][1] ),
    .A3(\top1.memory2.mem1[83][1] ),
    .S1(net6144),
    .X(_05925_));
 sg13g2_mux4_1 _15530_ (.S0(net6210),
    .A0(\top1.memory2.mem1[92][1] ),
    .A1(\top1.memory2.mem1[93][1] ),
    .A2(\top1.memory2.mem1[94][1] ),
    .A3(\top1.memory2.mem1[95][1] ),
    .S1(net6145),
    .X(_05926_));
 sg13g2_a22oi_1 _15531_ (.Y(_05927_),
    .B1(_05926_),
    .B2(net5853),
    .A2(_05925_),
    .A1(net5877));
 sg13g2_o21ai_1 _15532_ (.B1(net6021),
    .Y(_05928_),
    .A1(\top1.memory2.mem1[86][1] ),
    .A2(net5894));
 sg13g2_nor2_1 _15533_ (.A(\top1.memory2.mem1[87][1] ),
    .B(net5937),
    .Y(_05929_));
 sg13g2_nor2_1 _15534_ (.A(\top1.memory2.mem1[85][1] ),
    .B(net5973),
    .Y(_05930_));
 sg13g2_nor2_1 _15535_ (.A(\top1.memory2.mem1[84][1] ),
    .B(net6039),
    .Y(_05931_));
 sg13g2_nor4_2 _15536_ (.A(_05928_),
    .B(_05929_),
    .C(_05930_),
    .Y(_05932_),
    .D(_05931_));
 sg13g2_mux4_1 _15537_ (.S0(net6210),
    .A0(\top1.memory2.mem1[88][1] ),
    .A1(\top1.memory2.mem1[89][1] ),
    .A2(\top1.memory2.mem1[90][1] ),
    .A3(\top1.memory2.mem1[91][1] ),
    .S1(net6145),
    .X(_05933_));
 sg13g2_nand2_1 _15538_ (.Y(_05934_),
    .A(net6087),
    .B(_05933_));
 sg13g2_nand2_1 _15539_ (.Y(_05935_),
    .A(_05927_),
    .B(_05934_));
 sg13g2_o21ai_1 _15540_ (.B1(_05516_),
    .Y(_05936_),
    .A1(_05932_),
    .A2(_05935_));
 sg13g2_nor3_2 _15541_ (.A(net6116),
    .B(_05869_),
    .C(_05888_),
    .Y(_05937_));
 sg13g2_nand3_1 _15542_ (.B(_05898_),
    .C(_05937_),
    .A(_05881_),
    .Y(_05938_));
 sg13g2_nor3_2 _15543_ (.A(net6102),
    .B(_05917_),
    .C(_05924_),
    .Y(_05939_));
 sg13g2_nand3_1 _15544_ (.B(_05936_),
    .C(_05939_),
    .A(_05910_),
    .Y(_05940_));
 sg13g2_a21o_1 _15545_ (.A2(_05940_),
    .A1(_05938_),
    .B1(net6111),
    .X(_05941_));
 sg13g2_a22oi_1 _15546_ (.Y(_05942_),
    .B1(net5907),
    .B2(\top1.memory2.mem1[138][1] ),
    .A2(net5947),
    .A1(\top1.memory2.mem1[139][1] ));
 sg13g2_a22oi_1 _15547_ (.Y(_05943_),
    .B1(net5982),
    .B2(\top1.memory2.mem1[137][1] ),
    .A2(net6047),
    .A1(\top1.memory2.mem1[136][1] ));
 sg13g2_a21oi_1 _15548_ (.A1(_05942_),
    .A2(_05943_),
    .Y(_05944_),
    .B1(net6075));
 sg13g2_o21ai_1 _15549_ (.B1(net6019),
    .Y(_05945_),
    .A1(\top1.memory2.mem1[135][1] ),
    .A2(net5930));
 sg13g2_nor2_1 _15550_ (.A(\top1.memory2.mem1[132][1] ),
    .B(net6036),
    .Y(_05946_));
 sg13g2_nor2_1 _15551_ (.A(\top1.memory2.mem1[133][1] ),
    .B(net5970),
    .Y(_05947_));
 sg13g2_nor2_1 _15552_ (.A(\top1.memory2.mem1[134][1] ),
    .B(net5891),
    .Y(_05948_));
 sg13g2_nor4_1 _15553_ (.A(_05945_),
    .B(_05946_),
    .C(_05947_),
    .D(_05948_),
    .Y(_05949_));
 sg13g2_mux4_1 _15554_ (.S0(net6208),
    .A0(\top1.memory2.mem1[128][1] ),
    .A1(\top1.memory2.mem1[129][1] ),
    .A2(\top1.memory2.mem1[130][1] ),
    .A3(\top1.memory2.mem1[131][1] ),
    .S1(net6143),
    .X(_05950_));
 sg13g2_mux4_1 _15555_ (.S0(net6203),
    .A0(\top1.memory2.mem1[140][1] ),
    .A1(\top1.memory2.mem1[141][1] ),
    .A2(\top1.memory2.mem1[142][1] ),
    .A3(\top1.memory2.mem1[143][1] ),
    .S1(net6139),
    .X(_05951_));
 sg13g2_a22oi_1 _15556_ (.Y(_05952_),
    .B1(_05951_),
    .B2(net5851),
    .A2(_05950_),
    .A1(net5875));
 sg13g2_inv_1 _15557_ (.Y(_05953_),
    .A(_05952_));
 sg13g2_nor4_2 _15558_ (.A(net6122),
    .B(_05944_),
    .C(_05949_),
    .Y(_05954_),
    .D(_05953_));
 sg13g2_nor2_1 _15559_ (.A(\top1.memory2.mem1[148][1] ),
    .B(net6037),
    .Y(_05955_));
 sg13g2_nor2_1 _15560_ (.A(\top1.memory2.mem1[149][1] ),
    .B(net5971),
    .Y(_05956_));
 sg13g2_nor2_1 _15561_ (.A(\top1.memory2.mem1[151][1] ),
    .B(net5934),
    .Y(_05957_));
 sg13g2_o21ai_1 _15562_ (.B1(net6016),
    .Y(_05958_),
    .A1(\top1.memory2.mem1[150][1] ),
    .A2(net5890));
 sg13g2_nor4_2 _15563_ (.A(_05955_),
    .B(_05956_),
    .C(_05957_),
    .Y(_05959_),
    .D(_05958_));
 sg13g2_mux4_1 _15564_ (.S0(net6205),
    .A0(\top1.memory2.mem1[144][1] ),
    .A1(\top1.memory2.mem1[145][1] ),
    .A2(\top1.memory2.mem1[146][1] ),
    .A3(\top1.memory2.mem1[147][1] ),
    .S1(net6141),
    .X(_05960_));
 sg13g2_nand2_1 _15565_ (.Y(_05961_),
    .A(net5876),
    .B(_05960_));
 sg13g2_mux4_1 _15566_ (.S0(net6205),
    .A0(\top1.memory2.mem1[152][1] ),
    .A1(\top1.memory2.mem1[153][1] ),
    .A2(\top1.memory2.mem1[154][1] ),
    .A3(\top1.memory2.mem1[155][1] ),
    .S1(net6141),
    .X(_05962_));
 sg13g2_mux4_1 _15567_ (.S0(net6206),
    .A0(\top1.memory2.mem1[156][1] ),
    .A1(\top1.memory2.mem1[157][1] ),
    .A2(\top1.memory2.mem1[158][1] ),
    .A3(\top1.memory2.mem1[159][1] ),
    .S1(net6142),
    .X(_05963_));
 sg13g2_a22oi_1 _15568_ (.Y(_05964_),
    .B1(_05963_),
    .B2(net5852),
    .A2(_05962_),
    .A1(net6085));
 sg13g2_nand2_1 _15569_ (.Y(_05965_),
    .A(_05961_),
    .B(_05964_));
 sg13g2_nor3_1 _15570_ (.A(net6107),
    .B(_05959_),
    .C(_05965_),
    .Y(_05966_));
 sg13g2_or3_2 _15571_ (.A(net6117),
    .B(_05954_),
    .C(_05966_),
    .X(_05967_));
 sg13g2_mux4_1 _15572_ (.S0(net6224),
    .A0(\top1.memory2.mem1[176][1] ),
    .A1(\top1.memory2.mem1[177][1] ),
    .A2(\top1.memory2.mem1[178][1] ),
    .A3(\top1.memory2.mem1[179][1] ),
    .S1(net6159),
    .X(_05968_));
 sg13g2_mux4_1 _15573_ (.S0(net6224),
    .A0(\top1.memory2.mem1[184][1] ),
    .A1(\top1.memory2.mem1[185][1] ),
    .A2(\top1.memory2.mem1[186][1] ),
    .A3(\top1.memory2.mem1[187][1] ),
    .S1(net6159),
    .X(_05969_));
 sg13g2_and2_1 _15574_ (.A(net6090),
    .B(_05969_),
    .X(_05970_));
 sg13g2_mux4_1 _15575_ (.S0(net6224),
    .A0(\top1.memory2.mem1[180][1] ),
    .A1(\top1.memory2.mem1[181][1] ),
    .A2(\top1.memory2.mem1[182][1] ),
    .A3(\top1.memory2.mem1[183][1] ),
    .S1(net6159),
    .X(_05971_));
 sg13g2_a22oi_1 _15576_ (.Y(_05972_),
    .B1(net5926),
    .B2(\top1.memory2.mem1[190][1] ),
    .A2(net5966),
    .A1(\top1.memory2.mem1[191][1] ));
 sg13g2_a22oi_1 _15577_ (.Y(_05973_),
    .B1(net6006),
    .B2(\top1.memory2.mem1[189][1] ),
    .A2(net6070),
    .A1(\top1.memory2.mem1[188][1] ));
 sg13g2_a21o_1 _15578_ (.A2(_05973_),
    .A1(_05972_),
    .B1(net5848),
    .X(_05974_));
 sg13g2_a221oi_1 _15579_ (.B2(net6025),
    .C1(_05970_),
    .B1(_05971_),
    .A1(net5880),
    .Y(_05975_),
    .A2(_05968_));
 sg13g2_a21oi_2 _15580_ (.B1(net5837),
    .Y(_05976_),
    .A2(_05975_),
    .A1(_05974_));
 sg13g2_mux4_1 _15581_ (.S0(net6221),
    .A0(\top1.memory2.mem1[168][1] ),
    .A1(\top1.memory2.mem1[169][1] ),
    .A2(\top1.memory2.mem1[170][1] ),
    .A3(\top1.memory2.mem1[171][1] ),
    .S1(net6156),
    .X(_05977_));
 sg13g2_mux4_1 _15582_ (.S0(net6212),
    .A0(\top1.memory2.mem1[160][1] ),
    .A1(\top1.memory2.mem1[161][1] ),
    .A2(\top1.memory2.mem1[162][1] ),
    .A3(\top1.memory2.mem1[163][1] ),
    .S1(net6147),
    .X(_05978_));
 sg13g2_mux4_1 _15583_ (.S0(net6222),
    .A0(\top1.memory2.mem1[164][1] ),
    .A1(\top1.memory2.mem1[165][1] ),
    .A2(\top1.memory2.mem1[166][1] ),
    .A3(\top1.memory2.mem1[167][1] ),
    .S1(net6157),
    .X(_05979_));
 sg13g2_mux4_1 _15584_ (.S0(net6220),
    .A0(\top1.memory2.mem1[172][1] ),
    .A1(\top1.memory2.mem1[173][1] ),
    .A2(\top1.memory2.mem1[174][1] ),
    .A3(\top1.memory2.mem1[175][1] ),
    .S1(net6155),
    .X(_05980_));
 sg13g2_a22oi_1 _15585_ (.Y(_05981_),
    .B1(_05979_),
    .B2(net6026),
    .A2(_05977_),
    .A1(net6089));
 sg13g2_a22oi_1 _15586_ (.Y(_05982_),
    .B1(_05980_),
    .B2(net5856),
    .A2(_05978_),
    .A1(net5881));
 sg13g2_a21oi_2 _15587_ (.B1(net5836),
    .Y(_05983_),
    .A2(_05982_),
    .A1(_05981_));
 sg13g2_nor3_1 _15588_ (.A(_05515_),
    .B(_05976_),
    .C(_05983_),
    .Y(_05984_));
 sg13g2_a21oi_1 _15589_ (.A1(\top1.memory2.mem1[199][1] ),
    .A2(net5951),
    .Y(_05985_),
    .B1(_03827_));
 sg13g2_a22oi_1 _15590_ (.Y(_05986_),
    .B1(net5993),
    .B2(\top1.memory2.mem1[197][1] ),
    .A2(net6056),
    .A1(\top1.memory2.mem1[196][1] ));
 sg13g2_nand2_1 _15591_ (.Y(_05987_),
    .A(_05985_),
    .B(_05986_));
 sg13g2_a21oi_1 _15592_ (.A1(\top1.memory2.mem1[198][1] ),
    .A2(net5911),
    .Y(_05988_),
    .B1(_05987_));
 sg13g2_a22oi_1 _15593_ (.Y(_05989_),
    .B1(net5952),
    .B2(\top1.memory2.mem1[195][1] ),
    .A2(net5998),
    .A1(\top1.memory2.mem1[193][1] ));
 sg13g2_a221oi_1 _15594_ (.B2(\top1.memory2.mem1[194][1] ),
    .C1(net6131),
    .B1(net5912),
    .A1(\top1.memory2.mem1[192][1] ),
    .Y(_05990_),
    .A2(net6057));
 sg13g2_a21o_1 _15595_ (.A2(_05990_),
    .A1(_05989_),
    .B1(_05988_),
    .X(_05991_));
 sg13g2_a221oi_1 _15596_ (.B2(_03978_),
    .C1(net6108),
    .B1(_05991_),
    .A1(_05967_),
    .Y(_05992_),
    .A2(_05984_));
 sg13g2_a21oi_1 _15597_ (.A1(_05941_),
    .A2(_05992_),
    .Y(_05993_),
    .B1(net6101));
 sg13g2_a22oi_1 _15598_ (.Y(_01019_),
    .B1(_05862_),
    .B2(_05993_),
    .A2(_03850_),
    .A1(net6101));
 sg13g2_nand2_1 _15599_ (.Y(_05994_),
    .A(_03832_),
    .B(\top1.memory2.data_out[2] ));
 sg13g2_nor3_1 _15600_ (.A(net6222),
    .B(net6163),
    .C(\top1.memory2.mem1[20][2] ),
    .Y(_05995_));
 sg13g2_a21oi_1 _15601_ (.A1(_03873_),
    .A2(net5919),
    .Y(_05996_),
    .B1(net6012));
 sg13g2_a221oi_1 _15602_ (.B2(_03874_),
    .C1(_05995_),
    .B1(net5959),
    .A1(_03872_),
    .Y(_05997_),
    .A2(net6000));
 sg13g2_mux4_1 _15603_ (.S0(net6229),
    .A0(\top1.memory2.mem1[16][2] ),
    .A1(\top1.memory2.mem1[17][2] ),
    .A2(\top1.memory2.mem1[18][2] ),
    .A3(\top1.memory2.mem1[19][2] ),
    .S1(net6164),
    .X(_05998_));
 sg13g2_mux4_1 _15604_ (.S0(net6225),
    .A0(\top1.memory2.mem1[24][2] ),
    .A1(\top1.memory2.mem1[25][2] ),
    .A2(\top1.memory2.mem1[26][2] ),
    .A3(\top1.memory2.mem1[27][2] ),
    .S1(net6160),
    .X(_05999_));
 sg13g2_and2_1 _15605_ (.A(net6090),
    .B(_05999_),
    .X(_06000_));
 sg13g2_mux4_1 _15606_ (.S0(net6228),
    .A0(\top1.memory2.mem1[28][2] ),
    .A1(\top1.memory2.mem1[29][2] ),
    .A2(\top1.memory2.mem1[30][2] ),
    .A3(\top1.memory2.mem1[31][2] ),
    .S1(net6163),
    .X(_06001_));
 sg13g2_a21oi_2 _15607_ (.B1(net6107),
    .Y(_06002_),
    .A2(_05998_),
    .A1(net5882));
 sg13g2_a221oi_1 _15608_ (.B2(net5856),
    .C1(_06000_),
    .B1(_06001_),
    .A1(_05996_),
    .Y(_06003_),
    .A2(_05997_));
 sg13g2_mux4_1 _15609_ (.S0(net6213),
    .A0(\top1.memory2.mem1[8][2] ),
    .A1(\top1.memory2.mem1[9][2] ),
    .A2(\top1.memory2.mem1[10][2] ),
    .A3(\top1.memory2.mem1[11][2] ),
    .S1(net6148),
    .X(_06004_));
 sg13g2_mux4_1 _15610_ (.S0(net6213),
    .A0(\top1.memory2.mem1[12][2] ),
    .A1(\top1.memory2.mem1[13][2] ),
    .A2(\top1.memory2.mem1[14][2] ),
    .A3(\top1.memory2.mem1[15][2] ),
    .S1(net6148),
    .X(_06005_));
 sg13g2_o21ai_1 _15611_ (.B1(net6022),
    .Y(_06006_),
    .A1(\top1.memory2.mem1[7][2] ),
    .A2(net5938));
 sg13g2_nor2_1 _15612_ (.A(\top1.memory2.mem1[4][2] ),
    .B(net6043),
    .Y(_06007_));
 sg13g2_nor2_1 _15613_ (.A(\top1.memory2.mem1[6][2] ),
    .B(net5897),
    .Y(_06008_));
 sg13g2_nor2_1 _15614_ (.A(\top1.memory2.mem1[5][2] ),
    .B(net5977),
    .Y(_06009_));
 sg13g2_or4_2 _15615_ (.A(_06006_),
    .B(_06007_),
    .C(_06008_),
    .D(_06009_),
    .X(_06010_));
 sg13g2_mux4_1 _15616_ (.S0(net6211),
    .A0(\top1.memory2.mem1[0][2] ),
    .A1(\top1.memory2.mem1[1][2] ),
    .A2(\top1.memory2.mem1[2][2] ),
    .A3(\top1.memory2.mem1[3][2] ),
    .S1(net6146),
    .X(_06011_));
 sg13g2_a21o_1 _15617_ (.A2(_06005_),
    .A1(net5853),
    .B1(net6124),
    .X(_06012_));
 sg13g2_a221oi_1 _15618_ (.B2(net5877),
    .C1(_06012_),
    .B1(_06011_),
    .A1(net6087),
    .Y(_06013_),
    .A2(_06004_));
 sg13g2_a221oi_1 _15619_ (.B2(_06013_),
    .C1(net6118),
    .B1(_06010_),
    .A1(_06002_),
    .Y(_06014_),
    .A2(_06003_));
 sg13g2_mux4_1 _15620_ (.S0(net6258),
    .A0(\top1.memory2.mem1[36][2] ),
    .A1(\top1.memory2.mem1[37][2] ),
    .A2(\top1.memory2.mem1[38][2] ),
    .A3(\top1.memory2.mem1[39][2] ),
    .S1(net6193),
    .X(_06015_));
 sg13g2_mux4_1 _15621_ (.S0(net6256),
    .A0(\top1.memory2.mem1[40][2] ),
    .A1(\top1.memory2.mem1[41][2] ),
    .A2(\top1.memory2.mem1[42][2] ),
    .A3(\top1.memory2.mem1[43][2] ),
    .S1(net6191),
    .X(_06016_));
 sg13g2_mux4_1 _15622_ (.S0(net6257),
    .A0(\top1.memory2.mem1[32][2] ),
    .A1(\top1.memory2.mem1[33][2] ),
    .A2(\top1.memory2.mem1[34][2] ),
    .A3(\top1.memory2.mem1[35][2] ),
    .S1(net6192),
    .X(_06017_));
 sg13g2_mux4_1 _15623_ (.S0(net6255),
    .A0(\top1.memory2.mem1[44][2] ),
    .A1(\top1.memory2.mem1[45][2] ),
    .A2(\top1.memory2.mem1[46][2] ),
    .A3(\top1.memory2.mem1[47][2] ),
    .S1(net6190),
    .X(_06018_));
 sg13g2_a22oi_1 _15624_ (.Y(_06019_),
    .B1(_06017_),
    .B2(net5887),
    .A2(_06015_),
    .A1(net6034));
 sg13g2_a22oi_1 _15625_ (.Y(_06020_),
    .B1(_06018_),
    .B2(net5864),
    .A2(_06016_),
    .A1(net6097));
 sg13g2_a21oi_1 _15626_ (.A1(_06019_),
    .A2(_06020_),
    .Y(_06021_),
    .B1(net5835));
 sg13g2_mux4_1 _15627_ (.S0(net6255),
    .A0(\top1.memory2.mem1[48][2] ),
    .A1(\top1.memory2.mem1[49][2] ),
    .A2(\top1.memory2.mem1[50][2] ),
    .A3(\top1.memory2.mem1[51][2] ),
    .S1(net6190),
    .X(_06022_));
 sg13g2_mux4_1 _15628_ (.S0(net6254),
    .A0(\top1.memory2.mem1[56][2] ),
    .A1(\top1.memory2.mem1[57][2] ),
    .A2(\top1.memory2.mem1[58][2] ),
    .A3(\top1.memory2.mem1[59][2] ),
    .S1(net6189),
    .X(_06023_));
 sg13g2_mux4_1 _15629_ (.S0(net6255),
    .A0(\top1.memory2.mem1[60][2] ),
    .A1(\top1.memory2.mem1[61][2] ),
    .A2(\top1.memory2.mem1[62][2] ),
    .A3(\top1.memory2.mem1[63][2] ),
    .S1(net6190),
    .X(_06024_));
 sg13g2_mux4_1 _15630_ (.S0(net6254),
    .A0(\top1.memory2.mem1[52][2] ),
    .A1(\top1.memory2.mem1[53][2] ),
    .A2(\top1.memory2.mem1[54][2] ),
    .A3(\top1.memory2.mem1[55][2] ),
    .S1(net6189),
    .X(_06025_));
 sg13g2_a22oi_1 _15631_ (.Y(_06026_),
    .B1(_06024_),
    .B2(net5864),
    .A2(_06022_),
    .A1(net5886));
 sg13g2_a22oi_1 _15632_ (.Y(_06027_),
    .B1(_06025_),
    .B2(net6033),
    .A2(_06023_),
    .A1(net6097));
 sg13g2_a21oi_1 _15633_ (.A1(_06026_),
    .A2(_06027_),
    .Y(_06028_),
    .B1(net5840));
 sg13g2_or2_2 _15634_ (.X(_06029_),
    .B(_06028_),
    .A(_06021_));
 sg13g2_o21ai_1 _15635_ (.B1(net6102),
    .Y(_06030_),
    .A1(_06014_),
    .A2(_06029_));
 sg13g2_mux4_1 _15636_ (.S0(net6209),
    .A0(\top1.memory2.mem1[80][2] ),
    .A1(\top1.memory2.mem1[81][2] ),
    .A2(\top1.memory2.mem1[82][2] ),
    .A3(\top1.memory2.mem1[83][2] ),
    .S1(net6144),
    .X(_06031_));
 sg13g2_a21o_1 _15637_ (.A2(_06031_),
    .A1(net5877),
    .B1(net6105),
    .X(_06032_));
 sg13g2_a22oi_1 _15638_ (.Y(_06033_),
    .B1(net5911),
    .B2(\top1.memory2.mem1[90][2] ),
    .A2(net6056),
    .A1(\top1.memory2.mem1[88][2] ));
 sg13g2_a22oi_1 _15639_ (.Y(_06034_),
    .B1(net5952),
    .B2(\top1.memory2.mem1[91][2] ),
    .A2(net5992),
    .A1(\top1.memory2.mem1[89][2] ));
 sg13g2_a21oi_1 _15640_ (.A1(_06033_),
    .A2(_06034_),
    .Y(_06035_),
    .B1(net6077));
 sg13g2_nor2_1 _15641_ (.A(\top1.memory2.mem1[87][2] ),
    .B(net5933),
    .Y(_06036_));
 sg13g2_nor2_1 _15642_ (.A(\top1.memory2.mem1[85][2] ),
    .B(net5973),
    .Y(_06037_));
 sg13g2_nor2_1 _15643_ (.A(\top1.memory2.mem1[84][2] ),
    .B(net6039),
    .Y(_06038_));
 sg13g2_o21ai_1 _15644_ (.B1(net6021),
    .Y(_06039_),
    .A1(\top1.memory2.mem1[86][2] ),
    .A2(net5894));
 sg13g2_nor4_2 _15645_ (.A(_06036_),
    .B(_06037_),
    .C(_06038_),
    .Y(_06040_),
    .D(_06039_));
 sg13g2_a22oi_1 _15646_ (.Y(_06041_),
    .B1(net5912),
    .B2(\top1.memory2.mem1[94][2] ),
    .A2(net5952),
    .A1(\top1.memory2.mem1[95][2] ));
 sg13g2_a22oi_1 _15647_ (.Y(_06042_),
    .B1(net5992),
    .B2(\top1.memory2.mem1[93][2] ),
    .A2(net6057),
    .A1(\top1.memory2.mem1[92][2] ));
 sg13g2_a21oi_1 _15648_ (.A1(_06041_),
    .A2(_06042_),
    .Y(_06043_),
    .B1(net5845));
 sg13g2_nor4_2 _15649_ (.A(_06032_),
    .B(_06035_),
    .C(_06040_),
    .Y(_06044_),
    .D(_06043_));
 sg13g2_mux4_1 _15650_ (.S0(net6198),
    .A0(\top1.memory2.mem1[64][2] ),
    .A1(\top1.memory2.mem1[65][2] ),
    .A2(\top1.memory2.mem1[66][2] ),
    .A3(\top1.memory2.mem1[67][2] ),
    .S1(net6134),
    .X(_06045_));
 sg13g2_a21o_1 _15651_ (.A2(_06045_),
    .A1(net5873),
    .B1(net6120),
    .X(_06046_));
 sg13g2_a22oi_1 _15652_ (.Y(_06047_),
    .B1(net5901),
    .B2(\top1.memory2.mem1[78][2] ),
    .A2(net5942),
    .A1(\top1.memory2.mem1[79][2] ));
 sg13g2_a22oi_1 _15653_ (.Y(_06048_),
    .B1(net5981),
    .B2(\top1.memory2.mem1[77][2] ),
    .A2(net6046),
    .A1(\top1.memory2.mem1[76][2] ));
 sg13g2_a21oi_1 _15654_ (.A1(_06047_),
    .A2(_06048_),
    .Y(_06049_),
    .B1(net5844));
 sg13g2_nor2_1 _15655_ (.A(\top1.memory2.mem1[68][2] ),
    .B(net6036),
    .Y(_06050_));
 sg13g2_nor2_1 _15656_ (.A(\top1.memory2.mem1[70][2] ),
    .B(net5890),
    .Y(_06051_));
 sg13g2_nor2_1 _15657_ (.A(\top1.memory2.mem1[69][2] ),
    .B(net5970),
    .Y(_06052_));
 sg13g2_o21ai_1 _15658_ (.B1(net6018),
    .Y(_06053_),
    .A1(\top1.memory2.mem1[71][2] ),
    .A2(net5932));
 sg13g2_nor4_2 _15659_ (.A(_06050_),
    .B(_06051_),
    .C(_06052_),
    .Y(_06054_),
    .D(_06053_));
 sg13g2_a22oi_1 _15660_ (.Y(_06055_),
    .B1(net5901),
    .B2(\top1.memory2.mem1[74][2] ),
    .A2(net6046),
    .A1(\top1.memory2.mem1[72][2] ));
 sg13g2_a22oi_1 _15661_ (.Y(_06056_),
    .B1(net5942),
    .B2(\top1.memory2.mem1[75][2] ),
    .A2(net5981),
    .A1(\top1.memory2.mem1[73][2] ));
 sg13g2_a21oi_1 _15662_ (.A1(_06055_),
    .A2(_06056_),
    .Y(_06057_),
    .B1(net6075));
 sg13g2_nor4_2 _15663_ (.A(_06046_),
    .B(_06049_),
    .C(_06054_),
    .Y(_06058_),
    .D(_06057_));
 sg13g2_or3_2 _15664_ (.A(_05479_),
    .B(_06044_),
    .C(_06058_),
    .X(_06059_));
 sg13g2_mux4_1 _15665_ (.S0(net6243),
    .A0(\top1.memory2.mem1[116][2] ),
    .A1(\top1.memory2.mem1[117][2] ),
    .A2(\top1.memory2.mem1[118][2] ),
    .A3(\top1.memory2.mem1[119][2] ),
    .S1(net6178),
    .X(_06060_));
 sg13g2_mux4_1 _15666_ (.S0(net6242),
    .A0(\top1.memory2.mem1[120][2] ),
    .A1(\top1.memory2.mem1[121][2] ),
    .A2(\top1.memory2.mem1[122][2] ),
    .A3(\top1.memory2.mem1[123][2] ),
    .S1(net6177),
    .X(_06061_));
 sg13g2_mux4_1 _15667_ (.S0(net6244),
    .A0(\top1.memory2.mem1[112][2] ),
    .A1(\top1.memory2.mem1[113][2] ),
    .A2(\top1.memory2.mem1[114][2] ),
    .A3(\top1.memory2.mem1[115][2] ),
    .S1(net6179),
    .X(_06062_));
 sg13g2_mux4_1 _15668_ (.S0(net6246),
    .A0(\top1.memory2.mem1[124][2] ),
    .A1(\top1.memory2.mem1[125][2] ),
    .A2(\top1.memory2.mem1[126][2] ),
    .A3(\top1.memory2.mem1[127][2] ),
    .S1(net6181),
    .X(_06063_));
 sg13g2_a22oi_1 _15669_ (.Y(_06064_),
    .B1(_06062_),
    .B2(net5884),
    .A2(_06060_),
    .A1(net6030));
 sg13g2_a22oi_1 _15670_ (.Y(_06065_),
    .B1(_06063_),
    .B2(net5861),
    .A2(_06061_),
    .A1(net6094));
 sg13g2_a21oi_2 _15671_ (.B1(net5839),
    .Y(_06066_),
    .A2(_06065_),
    .A1(_06064_));
 sg13g2_mux4_1 _15672_ (.S0(net6249),
    .A0(\top1.memory2.mem1[104][2] ),
    .A1(\top1.memory2.mem1[105][2] ),
    .A2(\top1.memory2.mem1[106][2] ),
    .A3(\top1.memory2.mem1[107][2] ),
    .S1(net6184),
    .X(_06067_));
 sg13g2_mux4_1 _15673_ (.S0(net6233),
    .A0(\top1.memory2.mem1[96][2] ),
    .A1(\top1.memory2.mem1[97][2] ),
    .A2(\top1.memory2.mem1[98][2] ),
    .A3(\top1.memory2.mem1[99][2] ),
    .S1(net6168),
    .X(_06068_));
 sg13g2_mux4_1 _15674_ (.S0(net6239),
    .A0(\top1.memory2.mem1[100][2] ),
    .A1(\top1.memory2.mem1[101][2] ),
    .A2(\top1.memory2.mem1[102][2] ),
    .A3(\top1.memory2.mem1[103][2] ),
    .S1(net6174),
    .X(_06069_));
 sg13g2_mux4_1 _15675_ (.S0(net6239),
    .A0(\top1.memory2.mem1[108][2] ),
    .A1(\top1.memory2.mem1[109][2] ),
    .A2(\top1.memory2.mem1[110][2] ),
    .A3(\top1.memory2.mem1[111][2] ),
    .S1(net6174),
    .X(_06070_));
 sg13g2_a22oi_1 _15676_ (.Y(_06071_),
    .B1(_06069_),
    .B2(net6031),
    .A2(_06067_),
    .A1(net6096));
 sg13g2_a22oi_1 _15677_ (.Y(_06072_),
    .B1(_06070_),
    .B2(net5860),
    .A2(_06068_),
    .A1(net5885));
 sg13g2_a21oi_1 _15678_ (.A1(_06071_),
    .A2(_06072_),
    .Y(_06073_),
    .B1(net5833));
 sg13g2_o21ai_1 _15679_ (.B1(net6116),
    .Y(_06074_),
    .A1(_06066_),
    .A2(_06073_));
 sg13g2_nand4_1 _15680_ (.B(_06030_),
    .C(_06059_),
    .A(_03831_),
    .Y(_06075_),
    .D(_06074_));
 sg13g2_mux4_1 _15681_ (.S0(net6203),
    .A0(\top1.memory2.mem1[136][2] ),
    .A1(\top1.memory2.mem1[137][2] ),
    .A2(\top1.memory2.mem1[138][2] ),
    .A3(\top1.memory2.mem1[139][2] ),
    .S1(net6139),
    .X(_06076_));
 sg13g2_a21oi_1 _15682_ (.A1(net6084),
    .A2(_06076_),
    .Y(_06077_),
    .B1(net6122));
 sg13g2_nor2_1 _15683_ (.A(\top1.memory2.mem1[135][2] ),
    .B(net5930),
    .Y(_06078_));
 sg13g2_nor2_1 _15684_ (.A(\top1.memory2.mem1[133][2] ),
    .B(net5976),
    .Y(_06079_));
 sg13g2_nor2_1 _15685_ (.A(\top1.memory2.mem1[134][2] ),
    .B(net5891),
    .Y(_06080_));
 sg13g2_o21ai_1 _15686_ (.B1(net6019),
    .Y(_06081_),
    .A1(\top1.memory2.mem1[132][2] ),
    .A2(net6042));
 sg13g2_or4_1 _15687_ (.A(_06078_),
    .B(_06079_),
    .C(_06080_),
    .D(_06081_),
    .X(_06082_));
 sg13g2_mux4_1 _15688_ (.S0(net6203),
    .A0(\top1.memory2.mem1[128][2] ),
    .A1(\top1.memory2.mem1[129][2] ),
    .A2(\top1.memory2.mem1[130][2] ),
    .A3(\top1.memory2.mem1[131][2] ),
    .S1(net6139),
    .X(_06083_));
 sg13g2_mux4_1 _15689_ (.S0(net6203),
    .A0(\top1.memory2.mem1[140][2] ),
    .A1(\top1.memory2.mem1[141][2] ),
    .A2(\top1.memory2.mem1[142][2] ),
    .A3(\top1.memory2.mem1[143][2] ),
    .S1(net6139),
    .X(_06084_));
 sg13g2_a22oi_1 _15690_ (.Y(_06085_),
    .B1(_06084_),
    .B2(net5851),
    .A2(_06083_),
    .A1(net5875));
 sg13g2_nand3_1 _15691_ (.B(_06082_),
    .C(_06085_),
    .A(_06077_),
    .Y(_06086_));
 sg13g2_mux4_1 _15692_ (.S0(net6205),
    .A0(\top1.memory2.mem1[152][2] ),
    .A1(\top1.memory2.mem1[153][2] ),
    .A2(\top1.memory2.mem1[154][2] ),
    .A3(\top1.memory2.mem1[155][2] ),
    .S1(net6141),
    .X(_06087_));
 sg13g2_a22oi_1 _15693_ (.Y(_06088_),
    .B1(net5908),
    .B2(\top1.memory2.mem1[146][2] ),
    .A2(net5949),
    .A1(\top1.memory2.mem1[147][2] ));
 sg13g2_a22oi_1 _15694_ (.Y(_06089_),
    .B1(net5989),
    .B2(\top1.memory2.mem1[145][2] ),
    .A2(net6053),
    .A1(\top1.memory2.mem1[144][2] ));
 sg13g2_a21o_1 _15695_ (.A2(_06089_),
    .A1(_06088_),
    .B1(net5867),
    .X(_06090_));
 sg13g2_o21ai_1 _15696_ (.B1(net6016),
    .Y(_06091_),
    .A1(\top1.memory2.mem1[150][2] ),
    .A2(net5890));
 sg13g2_nor2_1 _15697_ (.A(\top1.memory2.mem1[149][2] ),
    .B(net5971),
    .Y(_06092_));
 sg13g2_nor2_1 _15698_ (.A(\top1.memory2.mem1[151][2] ),
    .B(net5934),
    .Y(_06093_));
 sg13g2_nor2_1 _15699_ (.A(\top1.memory2.mem1[148][2] ),
    .B(net6037),
    .Y(_06094_));
 sg13g2_or4_1 _15700_ (.A(_06091_),
    .B(_06092_),
    .C(_06093_),
    .D(_06094_),
    .X(_06095_));
 sg13g2_mux4_1 _15701_ (.S0(net6206),
    .A0(\top1.memory2.mem1[156][2] ),
    .A1(\top1.memory2.mem1[157][2] ),
    .A2(\top1.memory2.mem1[158][2] ),
    .A3(\top1.memory2.mem1[159][2] ),
    .S1(net6142),
    .X(_06096_));
 sg13g2_a22oi_1 _15702_ (.Y(_06097_),
    .B1(_06096_),
    .B2(net5852),
    .A2(_06087_),
    .A1(net6085));
 sg13g2_nand4_1 _15703_ (.B(_06090_),
    .C(_06095_),
    .A(net6122),
    .Y(_06098_),
    .D(_06097_));
 sg13g2_nand3_1 _15704_ (.B(_06086_),
    .C(_06098_),
    .A(net6103),
    .Y(_06099_));
 sg13g2_mux4_1 _15705_ (.S0(net6220),
    .A0(\top1.memory2.mem1[168][2] ),
    .A1(\top1.memory2.mem1[169][2] ),
    .A2(\top1.memory2.mem1[170][2] ),
    .A3(\top1.memory2.mem1[171][2] ),
    .S1(net6155),
    .X(_06100_));
 sg13g2_mux4_1 _15706_ (.S0(net6212),
    .A0(\top1.memory2.mem1[160][2] ),
    .A1(\top1.memory2.mem1[161][2] ),
    .A2(\top1.memory2.mem1[162][2] ),
    .A3(\top1.memory2.mem1[163][2] ),
    .S1(net6147),
    .X(_06101_));
 sg13g2_mux4_1 _15707_ (.S0(net6221),
    .A0(\top1.memory2.mem1[164][2] ),
    .A1(\top1.memory2.mem1[165][2] ),
    .A2(\top1.memory2.mem1[166][2] ),
    .A3(\top1.memory2.mem1[167][2] ),
    .S1(net6156),
    .X(_06102_));
 sg13g2_mux4_1 _15708_ (.S0(net6220),
    .A0(\top1.memory2.mem1[172][2] ),
    .A1(\top1.memory2.mem1[173][2] ),
    .A2(\top1.memory2.mem1[174][2] ),
    .A3(\top1.memory2.mem1[175][2] ),
    .S1(net6155),
    .X(_06103_));
 sg13g2_a22oi_1 _15709_ (.Y(_06104_),
    .B1(_06102_),
    .B2(net6026),
    .A2(_06100_),
    .A1(net6089));
 sg13g2_a22oi_1 _15710_ (.Y(_06105_),
    .B1(_06103_),
    .B2(net5856),
    .A2(_06101_),
    .A1(net5881));
 sg13g2_a21oi_2 _15711_ (.B1(net5836),
    .Y(_06106_),
    .A2(_06105_),
    .A1(_06104_));
 sg13g2_mux4_1 _15712_ (.S0(net6225),
    .A0(\top1.memory2.mem1[188][2] ),
    .A1(\top1.memory2.mem1[189][2] ),
    .A2(\top1.memory2.mem1[190][2] ),
    .A3(\top1.memory2.mem1[191][2] ),
    .S1(net6160),
    .X(_06107_));
 sg13g2_mux4_1 _15713_ (.S0(net6225),
    .A0(\top1.memory2.mem1[176][2] ),
    .A1(\top1.memory2.mem1[177][2] ),
    .A2(\top1.memory2.mem1[178][2] ),
    .A3(\top1.memory2.mem1[179][2] ),
    .S1(net6160),
    .X(_06108_));
 sg13g2_mux4_1 _15714_ (.S0(net6224),
    .A0(\top1.memory2.mem1[180][2] ),
    .A1(\top1.memory2.mem1[181][2] ),
    .A2(\top1.memory2.mem1[182][2] ),
    .A3(\top1.memory2.mem1[183][2] ),
    .S1(net6159),
    .X(_06109_));
 sg13g2_mux4_1 _15715_ (.S0(net6224),
    .A0(\top1.memory2.mem1[184][2] ),
    .A1(\top1.memory2.mem1[185][2] ),
    .A2(\top1.memory2.mem1[186][2] ),
    .A3(\top1.memory2.mem1[187][2] ),
    .S1(net6159),
    .X(_06110_));
 sg13g2_a22oi_1 _15716_ (.Y(_06111_),
    .B1(_06109_),
    .B2(net6025),
    .A2(_06107_),
    .A1(net5857));
 sg13g2_a22oi_1 _15717_ (.Y(_06112_),
    .B1(_06110_),
    .B2(net6090),
    .A2(_06108_),
    .A1(net5880));
 sg13g2_a21oi_2 _15718_ (.B1(net5837),
    .Y(_06113_),
    .A2(_06112_),
    .A1(_06111_));
 sg13g2_nor3_2 _15719_ (.A(net5831),
    .B(_06106_),
    .C(_06113_),
    .Y(_06114_));
 sg13g2_o21ai_1 _15720_ (.B1(_03827_),
    .Y(_06115_),
    .A1(\top1.memory2.mem1[195][2] ),
    .A2(net5937));
 sg13g2_nor2_1 _15721_ (.A(\top1.memory2.mem1[194][2] ),
    .B(net5897),
    .Y(_06116_));
 sg13g2_nor2_1 _15722_ (.A(\top1.memory2.mem1[192][2] ),
    .B(net6043),
    .Y(_06117_));
 sg13g2_nor2_1 _15723_ (.A(\top1.memory2.mem1[193][2] ),
    .B(net5977),
    .Y(_06118_));
 sg13g2_nor4_1 _15724_ (.A(_06115_),
    .B(_06116_),
    .C(_06117_),
    .D(_06118_),
    .Y(_06119_));
 sg13g2_o21ai_1 _15725_ (.B1(net6130),
    .Y(_06120_),
    .A1(\top1.memory2.mem1[199][2] ),
    .A2(net5938));
 sg13g2_nor2_1 _15726_ (.A(\top1.memory2.mem1[198][2] ),
    .B(net5896),
    .Y(_06121_));
 sg13g2_nor2_1 _15727_ (.A(\top1.memory2.mem1[196][2] ),
    .B(net6039),
    .Y(_06122_));
 sg13g2_nor2_1 _15728_ (.A(\top1.memory2.mem1[197][2] ),
    .B(net5973),
    .Y(_06123_));
 sg13g2_nor4_2 _15729_ (.A(_06120_),
    .B(_06121_),
    .C(_06122_),
    .Y(_06124_),
    .D(_06123_));
 sg13g2_nor3_1 _15730_ (.A(_03979_),
    .B(_06119_),
    .C(_06124_),
    .Y(_06125_));
 sg13g2_a21oi_1 _15731_ (.A1(_06099_),
    .A2(_06114_),
    .Y(_06126_),
    .B1(_06125_));
 sg13g2_a21oi_1 _15732_ (.A1(_06075_),
    .A2(_06126_),
    .Y(_06127_),
    .B1(net6108));
 sg13g2_a22oi_1 _15733_ (.Y(_06128_),
    .B1(net5955),
    .B2(\top1.memory2.mem2[3][2] ),
    .A2(net5996),
    .A1(\top1.memory2.mem2[1][2] ));
 sg13g2_a22oi_1 _15734_ (.Y(_06129_),
    .B1(net5916),
    .B2(\top1.memory2.mem2[2][2] ),
    .A2(net6061),
    .A1(\top1.memory2.mem2[0][2] ));
 sg13g2_a21oi_1 _15735_ (.A1(_06128_),
    .A2(_06129_),
    .Y(_06130_),
    .B1(net5869));
 sg13g2_o21ai_1 _15736_ (.B1(net6023),
    .Y(_06131_),
    .A1(\top1.memory2.mem2[6][2] ),
    .A2(net5898));
 sg13g2_nor2_1 _15737_ (.A(\top1.memory2.mem2[4][2] ),
    .B(net6044),
    .Y(_06132_));
 sg13g2_nor2_1 _15738_ (.A(\top1.memory2.mem2[5][2] ),
    .B(net5978),
    .Y(_06133_));
 sg13g2_nor2_1 _15739_ (.A(\top1.memory2.mem2[7][2] ),
    .B(net5939),
    .Y(_06134_));
 sg13g2_nor4_2 _15740_ (.A(_06131_),
    .B(_06132_),
    .C(_06133_),
    .Y(_06135_),
    .D(_06134_));
 sg13g2_a22oi_1 _15741_ (.Y(_06136_),
    .B1(net5915),
    .B2(\top1.memory2.mem2[10][2] ),
    .A2(net5955),
    .A1(\top1.memory2.mem2[11][2] ));
 sg13g2_a22oi_1 _15742_ (.Y(_06137_),
    .B1(net5996),
    .B2(\top1.memory2.mem2[9][2] ),
    .A2(net6061),
    .A1(\top1.memory2.mem2[8][2] ));
 sg13g2_a21oi_1 _15743_ (.A1(_06136_),
    .A2(_06137_),
    .Y(_06138_),
    .B1(net6077));
 sg13g2_a22oi_1 _15744_ (.Y(_06139_),
    .B1(net5916),
    .B2(\top1.memory2.mem2[14][2] ),
    .A2(net5956),
    .A1(\top1.memory2.mem2[15][2] ));
 sg13g2_a22oi_1 _15745_ (.Y(_06140_),
    .B1(net5996),
    .B2(\top1.memory2.mem2[13][2] ),
    .A2(net6061),
    .A1(\top1.memory2.mem2[12][2] ));
 sg13g2_a21oi_1 _15746_ (.A1(_06139_),
    .A2(_06140_),
    .Y(_06141_),
    .B1(net5846));
 sg13g2_or4_2 _15747_ (.A(_06130_),
    .B(_06135_),
    .C(_06138_),
    .D(_06141_),
    .X(_06142_));
 sg13g2_a22oi_1 _15748_ (.Y(_06143_),
    .B1(net5924),
    .B2(\top1.memory2.mem2[18][2] ),
    .A2(net5964),
    .A1(\top1.memory2.mem2[19][2] ));
 sg13g2_a22oi_1 _15749_ (.Y(_06144_),
    .B1(net6004),
    .B2(\top1.memory2.mem2[17][2] ),
    .A2(net6066),
    .A1(\top1.memory2.mem2[16][2] ));
 sg13g2_a21oi_1 _15750_ (.A1(_06143_),
    .A2(_06144_),
    .Y(_06145_),
    .B1(net5870));
 sg13g2_a22oi_1 _15751_ (.Y(_06146_),
    .B1(net5921),
    .B2(\top1.memory2.mem2[30][2] ),
    .A2(net5961),
    .A1(\top1.memory2.mem2[31][2] ));
 sg13g2_a22oi_1 _15752_ (.Y(_06147_),
    .B1(net6002),
    .B2(\top1.memory2.mem2[29][2] ),
    .A2(net6065),
    .A1(\top1.memory2.mem2[28][2] ));
 sg13g2_a21oi_2 _15753_ (.B1(net5848),
    .Y(_06148_),
    .A2(_06147_),
    .A1(_06146_));
 sg13g2_a22oi_1 _15754_ (.Y(_06149_),
    .B1(net5923),
    .B2(\top1.memory2.mem2[26][2] ),
    .A2(net5963),
    .A1(\top1.memory2.mem2[27][2] ));
 sg13g2_a22oi_1 _15755_ (.Y(_06150_),
    .B1(net6004),
    .B2(\top1.memory2.mem2[25][2] ),
    .A2(net6066),
    .A1(\top1.memory2.mem2[24][2] ));
 sg13g2_a21oi_1 _15756_ (.A1(_06149_),
    .A2(_06150_),
    .Y(_06151_),
    .B1(net6080));
 sg13g2_nor2_1 _15757_ (.A(\top1.memory2.mem2[22][2] ),
    .B(net5899),
    .Y(_06152_));
 sg13g2_nor2_1 _15758_ (.A(\top1.memory2.mem2[21][2] ),
    .B(net5979),
    .Y(_06153_));
 sg13g2_nor2_1 _15759_ (.A(\top1.memory2.mem2[23][2] ),
    .B(net5940),
    .Y(_06154_));
 sg13g2_o21ai_1 _15760_ (.B1(net6027),
    .Y(_06155_),
    .A1(\top1.memory2.mem2[20][2] ),
    .A2(net6045));
 sg13g2_nor4_1 _15761_ (.A(_06152_),
    .B(_06153_),
    .C(_06154_),
    .D(_06155_),
    .Y(_06156_));
 sg13g2_or4_1 _15762_ (.A(_06145_),
    .B(_06148_),
    .C(_06151_),
    .D(_06156_),
    .X(_06157_));
 sg13g2_a22oi_1 _15763_ (.Y(_06158_),
    .B1(net5927),
    .B2(\top1.memory2.mem2[34][2] ),
    .A2(net5967),
    .A1(\top1.memory2.mem2[35][2] ));
 sg13g2_a22oi_1 _15764_ (.Y(_06159_),
    .B1(net6007),
    .B2(\top1.memory2.mem2[33][2] ),
    .A2(net6071),
    .A1(\top1.memory2.mem2[32][2] ));
 sg13g2_a21oi_1 _15765_ (.A1(_06158_),
    .A2(_06159_),
    .Y(_06160_),
    .B1(net5872));
 sg13g2_a22oi_1 _15766_ (.Y(_06161_),
    .B1(net5927),
    .B2(\top1.memory2.mem2[38][2] ),
    .A2(net5967),
    .A1(\top1.memory2.mem2[39][2] ));
 sg13g2_a22oi_1 _15767_ (.Y(_06162_),
    .B1(net6007),
    .B2(\top1.memory2.mem2[37][2] ),
    .A2(net6071),
    .A1(\top1.memory2.mem2[36][2] ));
 sg13g2_a21oi_1 _15768_ (.A1(_06161_),
    .A2(_06162_),
    .Y(_06163_),
    .B1(net6014));
 sg13g2_a22oi_1 _15769_ (.Y(_06164_),
    .B1(net5928),
    .B2(\top1.memory2.mem2[46][2] ),
    .A2(net5968),
    .A1(\top1.memory2.mem2[47][2] ));
 sg13g2_a22oi_1 _15770_ (.Y(_06165_),
    .B1(net6008),
    .B2(\top1.memory2.mem2[45][2] ),
    .A2(net6072),
    .A1(\top1.memory2.mem2[44][2] ));
 sg13g2_a21oi_2 _15771_ (.B1(net5849),
    .Y(_06166_),
    .A2(_06165_),
    .A1(_06164_));
 sg13g2_a22oi_1 _15772_ (.Y(_06167_),
    .B1(net5929),
    .B2(\top1.memory2.mem2[42][2] ),
    .A2(net5969),
    .A1(\top1.memory2.mem2[43][2] ));
 sg13g2_a22oi_1 _15773_ (.Y(_06168_),
    .B1(net6008),
    .B2(\top1.memory2.mem2[41][2] ),
    .A2(net6072),
    .A1(\top1.memory2.mem2[40][2] ));
 sg13g2_a21oi_1 _15774_ (.A1(_06167_),
    .A2(_06168_),
    .Y(_06169_),
    .B1(net6082));
 sg13g2_or4_2 _15775_ (.A(_06160_),
    .B(_06163_),
    .C(_06166_),
    .D(_06169_),
    .X(_06170_));
 sg13g2_a22oi_1 _15776_ (.Y(_06171_),
    .B1(_06170_),
    .B2(_05443_),
    .A2(_06157_),
    .A1(_05516_));
 sg13g2_mux4_1 _15777_ (.S0(net6252),
    .A0(\top1.memory2.mem2[60][2] ),
    .A1(\top1.memory2.mem2[61][2] ),
    .A2(\top1.memory2.mem2[62][2] ),
    .A3(\top1.memory2.mem2[63][2] ),
    .S1(net6187),
    .X(_06172_));
 sg13g2_a22oi_1 _15778_ (.Y(_06173_),
    .B1(net5928),
    .B2(\top1.memory2.mem2[50][2] ),
    .A2(net5968),
    .A1(\top1.memory2.mem2[51][2] ));
 sg13g2_a22oi_1 _15779_ (.Y(_06174_),
    .B1(net6008),
    .B2(\top1.memory2.mem2[49][2] ),
    .A2(net6072),
    .A1(\top1.memory2.mem2[48][2] ));
 sg13g2_a21o_1 _15780_ (.A2(_06174_),
    .A1(_06173_),
    .B1(net5872),
    .X(_06175_));
 sg13g2_mux4_1 _15781_ (.S0(net6251),
    .A0(\top1.memory2.mem2[52][2] ),
    .A1(\top1.memory2.mem2[53][2] ),
    .A2(\top1.memory2.mem2[54][2] ),
    .A3(\top1.memory2.mem2[55][2] ),
    .S1(net6186),
    .X(_06176_));
 sg13g2_a22oi_1 _15782_ (.Y(_06177_),
    .B1(net5928),
    .B2(\top1.memory2.mem2[58][2] ),
    .A2(net5968),
    .A1(\top1.memory2.mem2[59][2] ));
 sg13g2_a22oi_1 _15783_ (.Y(_06178_),
    .B1(net6008),
    .B2(\top1.memory2.mem2[57][2] ),
    .A2(net6072),
    .A1(\top1.memory2.mem2[56][2] ));
 sg13g2_a21o_1 _15784_ (.A2(_06178_),
    .A1(_06177_),
    .B1(net6082),
    .X(_06179_));
 sg13g2_a22oi_1 _15785_ (.Y(_06180_),
    .B1(_06176_),
    .B2(net6034),
    .A2(_06172_),
    .A1(net5862));
 sg13g2_nand3_1 _15786_ (.B(_06179_),
    .C(_06180_),
    .A(_06175_),
    .Y(_06181_));
 sg13g2_a221oi_1 _15787_ (.B2(_05452_),
    .C1(net6114),
    .B1(_06181_),
    .A1(_03976_),
    .Y(_06182_),
    .A2(_06142_));
 sg13g2_mux4_1 _15788_ (.S0(net6236),
    .A0(\top1.memory2.mem2[108][2] ),
    .A1(\top1.memory2.mem2[109][2] ),
    .A2(\top1.memory2.mem2[110][2] ),
    .A3(\top1.memory2.mem2[111][2] ),
    .S1(net6171),
    .X(_06183_));
 sg13g2_mux4_1 _15789_ (.S0(net6223),
    .A0(\top1.memory2.mem2[96][2] ),
    .A1(\top1.memory2.mem2[97][2] ),
    .A2(\top1.memory2.mem2[98][2] ),
    .A3(\top1.memory2.mem2[99][2] ),
    .S1(net6158),
    .X(_06184_));
 sg13g2_mux4_1 _15790_ (.S0(net6223),
    .A0(\top1.memory2.mem2[100][2] ),
    .A1(\top1.memory2.mem2[101][2] ),
    .A2(\top1.memory2.mem2[102][2] ),
    .A3(\top1.memory2.mem2[103][2] ),
    .S1(net6158),
    .X(_06185_));
 sg13g2_mux4_1 _15791_ (.S0(net6238),
    .A0(\top1.memory2.mem2[104][2] ),
    .A1(\top1.memory2.mem2[105][2] ),
    .A2(\top1.memory2.mem2[106][2] ),
    .A3(\top1.memory2.mem2[107][2] ),
    .S1(net6173),
    .X(_06186_));
 sg13g2_a22oi_1 _15792_ (.Y(_06187_),
    .B1(_06185_),
    .B2(net6031),
    .A2(_06183_),
    .A1(net5857));
 sg13g2_a22oi_1 _15793_ (.Y(_06188_),
    .B1(_06186_),
    .B2(net6093),
    .A2(_06184_),
    .A1(net5880));
 sg13g2_a21oi_1 _15794_ (.A1(_06187_),
    .A2(_06188_),
    .Y(_06189_),
    .B1(net5832));
 sg13g2_o21ai_1 _15795_ (.B1(net6016),
    .Y(_06190_),
    .A1(\top1.memory2.mem2[85][2] ),
    .A2(net5971));
 sg13g2_nor2_1 _15796_ (.A(\top1.memory2.mem2[87][2] ),
    .B(net5934),
    .Y(_06191_));
 sg13g2_nor2_1 _15797_ (.A(\top1.memory2.mem2[84][2] ),
    .B(net6040),
    .Y(_06192_));
 sg13g2_nor2_1 _15798_ (.A(\top1.memory2.mem2[86][2] ),
    .B(net5895),
    .Y(_06193_));
 sg13g2_nor4_2 _15799_ (.A(_06190_),
    .B(_06191_),
    .C(_06192_),
    .Y(_06194_),
    .D(_06193_));
 sg13g2_a22oi_1 _15800_ (.Y(_06195_),
    .B1(net5903),
    .B2(\top1.memory2.mem2[90][2] ),
    .A2(net5944),
    .A1(\top1.memory2.mem2[91][2] ));
 sg13g2_a22oi_1 _15801_ (.Y(_06196_),
    .B1(net5983),
    .B2(\top1.memory2.mem2[89][2] ),
    .A2(net6048),
    .A1(\top1.memory2.mem2[88][2] ));
 sg13g2_a21oi_1 _15802_ (.A1(_06195_),
    .A2(_06196_),
    .Y(_06197_),
    .B1(net6075));
 sg13g2_mux4_1 _15803_ (.S0(net6200),
    .A0(\top1.memory2.mem2[80][2] ),
    .A1(\top1.memory2.mem2[81][2] ),
    .A2(\top1.memory2.mem2[82][2] ),
    .A3(\top1.memory2.mem2[83][2] ),
    .S1(net6136),
    .X(_06198_));
 sg13g2_a22oi_1 _15804_ (.Y(_06199_),
    .B1(net5903),
    .B2(\top1.memory2.mem2[94][2] ),
    .A2(net6048),
    .A1(\top1.memory2.mem2[92][2] ));
 sg13g2_a22oi_1 _15805_ (.Y(_06200_),
    .B1(net5951),
    .B2(\top1.memory2.mem2[95][2] ),
    .A2(net5993),
    .A1(\top1.memory2.mem2[93][2] ));
 sg13g2_a21oi_1 _15806_ (.A1(_06199_),
    .A2(_06200_),
    .Y(_06201_),
    .B1(net5845));
 sg13g2_mux4_1 _15807_ (.S0(net6240),
    .A0(\top1.memory2.mem2[120][2] ),
    .A1(\top1.memory2.mem2[121][2] ),
    .A2(\top1.memory2.mem2[122][2] ),
    .A3(\top1.memory2.mem2[123][2] ),
    .S1(net6175),
    .X(_06202_));
 sg13g2_mux4_1 _15808_ (.S0(net6237),
    .A0(\top1.memory2.mem2[116][2] ),
    .A1(\top1.memory2.mem2[117][2] ),
    .A2(\top1.memory2.mem2[118][2] ),
    .A3(\top1.memory2.mem2[119][2] ),
    .S1(net6172),
    .X(_06203_));
 sg13g2_mux4_1 _15809_ (.S0(net6246),
    .A0(\top1.memory2.mem2[112][2] ),
    .A1(\top1.memory2.mem2[113][2] ),
    .A2(\top1.memory2.mem2[114][2] ),
    .A3(\top1.memory2.mem2[115][2] ),
    .S1(net6181),
    .X(_06204_));
 sg13g2_mux4_1 _15810_ (.S0(net6237),
    .A0(\top1.memory2.mem2[124][2] ),
    .A1(\top1.memory2.mem2[125][2] ),
    .A2(\top1.memory2.mem2[126][2] ),
    .A3(\top1.memory2.mem2[127][2] ),
    .S1(net6172),
    .X(_06205_));
 sg13g2_a22oi_1 _15811_ (.Y(_06206_),
    .B1(_06204_),
    .B2(net5885),
    .A2(_06202_),
    .A1(net6095));
 sg13g2_a22oi_1 _15812_ (.Y(_06207_),
    .B1(_06205_),
    .B2(net5859),
    .A2(_06203_),
    .A1(net6031));
 sg13g2_a21oi_2 _15813_ (.B1(net5838),
    .Y(_06208_),
    .A2(_06207_),
    .A1(_06206_));
 sg13g2_mux4_1 _15814_ (.S0(net6197),
    .A0(\top1.memory2.mem2[64][2] ),
    .A1(\top1.memory2.mem2[65][2] ),
    .A2(\top1.memory2.mem2[66][2] ),
    .A3(\top1.memory2.mem2[67][2] ),
    .S1(net6133),
    .X(_06209_));
 sg13g2_mux4_1 _15815_ (.S0(net6197),
    .A0(\top1.memory2.mem2[76][2] ),
    .A1(\top1.memory2.mem2[77][2] ),
    .A2(\top1.memory2.mem2[78][2] ),
    .A3(\top1.memory2.mem2[79][2] ),
    .S1(net6133),
    .X(_06210_));
 sg13g2_a22oi_1 _15816_ (.Y(_06211_),
    .B1(_06210_),
    .B2(net5850),
    .A2(_06209_),
    .A1(net5873));
 sg13g2_mux4_1 _15817_ (.S0(net6200),
    .A0(\top1.memory2.mem2[72][2] ),
    .A1(\top1.memory2.mem2[73][2] ),
    .A2(\top1.memory2.mem2[74][2] ),
    .A3(\top1.memory2.mem2[75][2] ),
    .S1(net6136),
    .X(_06212_));
 sg13g2_nor2_1 _15818_ (.A(\top1.memory2.mem2[70][2] ),
    .B(net5893),
    .Y(_06213_));
 sg13g2_nor2_1 _15819_ (.A(\top1.memory2.mem2[69][2] ),
    .B(net5972),
    .Y(_06214_));
 sg13g2_nor2_1 _15820_ (.A(\top1.memory2.mem2[71][2] ),
    .B(net5934),
    .Y(_06215_));
 sg13g2_o21ai_1 _15821_ (.B1(net6016),
    .Y(_06216_),
    .A1(\top1.memory2.mem2[68][2] ),
    .A2(net6037));
 sg13g2_nor4_1 _15822_ (.A(_06213_),
    .B(_06214_),
    .C(_06215_),
    .D(_06216_),
    .Y(_06217_));
 sg13g2_a21oi_1 _15823_ (.A1(net6083),
    .A2(_06212_),
    .Y(_06218_),
    .B1(net6120));
 sg13g2_nand2_2 _15824_ (.Y(_06219_),
    .A(_06211_),
    .B(_06218_));
 sg13g2_a21o_1 _15825_ (.A2(_06198_),
    .A1(net5874),
    .B1(net6104),
    .X(_06220_));
 sg13g2_nor4_1 _15826_ (.A(_06194_),
    .B(_06197_),
    .C(_06201_),
    .D(_06220_),
    .Y(_06221_));
 sg13g2_o21ai_1 _15827_ (.B1(net6103),
    .Y(_06222_),
    .A1(_06217_),
    .A2(_06219_));
 sg13g2_or2_2 _15828_ (.X(_06223_),
    .B(_06222_),
    .A(_06221_));
 sg13g2_nor3_2 _15829_ (.A(_03830_),
    .B(_06189_),
    .C(_06208_),
    .Y(_06224_));
 sg13g2_a221oi_1 _15830_ (.B2(_06224_),
    .C1(net6112),
    .B1(_06223_),
    .A1(_06171_),
    .Y(_06225_),
    .A2(_06182_));
 sg13g2_nor2_1 _15831_ (.A(\top1.memory2.mem2[149][2] ),
    .B(net5975),
    .Y(_06226_));
 sg13g2_nor2_1 _15832_ (.A(\top1.memory2.mem2[148][2] ),
    .B(net6042),
    .Y(_06227_));
 sg13g2_nor2_1 _15833_ (.A(\top1.memory2.mem2[150][2] ),
    .B(net5896),
    .Y(_06228_));
 sg13g2_o21ai_1 _15834_ (.B1(net6020),
    .Y(_06229_),
    .A1(\top1.memory2.mem2[151][2] ),
    .A2(net5935));
 sg13g2_or4_1 _15835_ (.A(_06226_),
    .B(_06227_),
    .C(_06228_),
    .D(_06229_),
    .X(_06230_));
 sg13g2_mux4_1 _15836_ (.S0(net6205),
    .A0(\top1.memory2.mem2[144][2] ),
    .A1(\top1.memory2.mem2[145][2] ),
    .A2(\top1.memory2.mem2[146][2] ),
    .A3(\top1.memory2.mem2[147][2] ),
    .S1(net6141),
    .X(_06231_));
 sg13g2_mux4_1 _15837_ (.S0(net6215),
    .A0(\top1.memory2.mem2[152][2] ),
    .A1(\top1.memory2.mem2[153][2] ),
    .A2(\top1.memory2.mem2[154][2] ),
    .A3(\top1.memory2.mem2[155][2] ),
    .S1(net6150),
    .X(_06232_));
 sg13g2_mux4_1 _15838_ (.S0(net6206),
    .A0(\top1.memory2.mem2[156][2] ),
    .A1(\top1.memory2.mem2[157][2] ),
    .A2(\top1.memory2.mem2[158][2] ),
    .A3(\top1.memory2.mem2[159][2] ),
    .S1(net6141),
    .X(_06233_));
 sg13g2_a21o_1 _15839_ (.A2(_06231_),
    .A1(net5875),
    .B1(net6105),
    .X(_06234_));
 sg13g2_a221oi_1 _15840_ (.B2(net5851),
    .C1(_06234_),
    .B1(_06233_),
    .A1(net6085),
    .Y(_06235_),
    .A2(_06232_));
 sg13g2_nor3_1 _15841_ (.A(net6204),
    .B(net6140),
    .C(\top1.memory2.mem2[132][2] ),
    .Y(_06236_));
 sg13g2_a21oi_1 _15842_ (.A1(_03877_),
    .A2(net5950),
    .Y(_06237_),
    .B1(net6011));
 sg13g2_a221oi_1 _15843_ (.B2(_03876_),
    .C1(_06236_),
    .B1(net5906),
    .A1(_03875_),
    .Y(_06238_),
    .A2(net5987));
 sg13g2_mux4_1 _15844_ (.S0(net6204),
    .A0(\top1.memory2.mem2[128][2] ),
    .A1(\top1.memory2.mem2[129][2] ),
    .A2(\top1.memory2.mem2[130][2] ),
    .A3(\top1.memory2.mem2[131][2] ),
    .S1(net6140),
    .X(_06239_));
 sg13g2_mux4_1 _15845_ (.S0(net6204),
    .A0(\top1.memory2.mem2[140][2] ),
    .A1(\top1.memory2.mem2[141][2] ),
    .A2(\top1.memory2.mem2[142][2] ),
    .A3(\top1.memory2.mem2[143][2] ),
    .S1(net6140),
    .X(_06240_));
 sg13g2_mux4_1 _15846_ (.S0(net6203),
    .A0(\top1.memory2.mem2[136][2] ),
    .A1(\top1.memory2.mem2[137][2] ),
    .A2(\top1.memory2.mem2[138][2] ),
    .A3(\top1.memory2.mem2[139][2] ),
    .S1(net6139),
    .X(_06241_));
 sg13g2_and2_1 _15847_ (.A(net6084),
    .B(_06241_),
    .X(_06242_));
 sg13g2_a21oi_1 _15848_ (.A1(net5851),
    .A2(_06240_),
    .Y(_06243_),
    .B1(net6123));
 sg13g2_a221oi_1 _15849_ (.B2(net5875),
    .C1(_06242_),
    .B1(_06239_),
    .A1(_06237_),
    .Y(_06244_),
    .A2(_06238_));
 sg13g2_a22oi_1 _15850_ (.Y(_06245_),
    .B1(_06243_),
    .B2(_06244_),
    .A2(_06235_),
    .A1(_06230_));
 sg13g2_mux4_1 _15851_ (.S0(net6214),
    .A0(\top1.memory2.mem2[172][2] ),
    .A1(\top1.memory2.mem2[173][2] ),
    .A2(\top1.memory2.mem2[174][2] ),
    .A3(\top1.memory2.mem2[175][2] ),
    .S1(net6149),
    .X(_06246_));
 sg13g2_mux4_1 _15852_ (.S0(net6217),
    .A0(\top1.memory2.mem2[160][2] ),
    .A1(\top1.memory2.mem2[161][2] ),
    .A2(\top1.memory2.mem2[162][2] ),
    .A3(\top1.memory2.mem2[163][2] ),
    .S1(net6152),
    .X(_06247_));
 sg13g2_a22oi_1 _15853_ (.Y(_06248_),
    .B1(_06247_),
    .B2(net5879),
    .A2(_06246_),
    .A1(net5855));
 sg13g2_mux4_1 _15854_ (.S0(net6217),
    .A0(\top1.memory2.mem2[168][2] ),
    .A1(\top1.memory2.mem2[169][2] ),
    .A2(\top1.memory2.mem2[170][2] ),
    .A3(\top1.memory2.mem2[171][2] ),
    .S1(net6152),
    .X(_06249_));
 sg13g2_mux4_1 _15855_ (.S0(net6217),
    .A0(\top1.memory2.mem2[164][2] ),
    .A1(\top1.memory2.mem2[165][2] ),
    .A2(\top1.memory2.mem2[166][2] ),
    .A3(\top1.memory2.mem2[167][2] ),
    .S1(net6152),
    .X(_06250_));
 sg13g2_a22oi_1 _15856_ (.Y(_06251_),
    .B1(_06250_),
    .B2(net6023),
    .A2(_06249_),
    .A1(net6087));
 sg13g2_nand2_2 _15857_ (.Y(_06252_),
    .A(_06248_),
    .B(_06251_));
 sg13g2_mux4_1 _15858_ (.S0(net6234),
    .A0(\top1.memory2.mem2[188][2] ),
    .A1(\top1.memory2.mem2[189][2] ),
    .A2(\top1.memory2.mem2[190][2] ),
    .A3(\top1.memory2.mem2[191][2] ),
    .S1(net6169),
    .X(_06253_));
 sg13g2_mux4_1 _15859_ (.S0(net6234),
    .A0(\top1.memory2.mem2[176][2] ),
    .A1(\top1.memory2.mem2[177][2] ),
    .A2(\top1.memory2.mem2[178][2] ),
    .A3(\top1.memory2.mem2[179][2] ),
    .S1(net6169),
    .X(_06254_));
 sg13g2_mux4_1 _15860_ (.S0(net6230),
    .A0(\top1.memory2.mem2[184][2] ),
    .A1(\top1.memory2.mem2[185][2] ),
    .A2(\top1.memory2.mem2[186][2] ),
    .A3(\top1.memory2.mem2[187][2] ),
    .S1(net6165),
    .X(_06255_));
 sg13g2_mux4_1 _15861_ (.S0(net6229),
    .A0(\top1.memory2.mem2[180][2] ),
    .A1(\top1.memory2.mem2[181][2] ),
    .A2(\top1.memory2.mem2[182][2] ),
    .A3(\top1.memory2.mem2[183][2] ),
    .S1(net6164),
    .X(_06256_));
 sg13g2_a22oi_1 _15862_ (.Y(_06257_),
    .B1(_06255_),
    .B2(net6092),
    .A2(_06253_),
    .A1(net5858));
 sg13g2_a22oi_1 _15863_ (.Y(_06258_),
    .B1(_06256_),
    .B2(net6028),
    .A2(_06254_),
    .A1(net5883));
 sg13g2_a21oi_2 _15864_ (.B1(net5837),
    .Y(_06259_),
    .A2(_06258_),
    .A1(_06257_));
 sg13g2_a221oi_1 _15865_ (.B2(_05443_),
    .C1(_06259_),
    .B1(_06252_),
    .A1(net6103),
    .Y(_06260_),
    .A2(_06245_));
 sg13g2_a21oi_1 _15866_ (.A1(\top1.memory2.mem2[195][2] ),
    .A2(net5954),
    .Y(_06261_),
    .B1(net6129));
 sg13g2_and2_1 _15867_ (.A(\top1.memory2.mem2[193][2] ),
    .B(net5995),
    .X(_06262_));
 sg13g2_a221oi_1 _15868_ (.B2(\top1.memory2.mem2[194][2] ),
    .C1(_06262_),
    .B1(net5915),
    .A1(\top1.memory2.mem2[192][2] ),
    .Y(_06263_),
    .A2(net6060));
 sg13g2_a22oi_1 _15869_ (.Y(_06264_),
    .B1(net5955),
    .B2(\top1.memory2.mem2[199][2] ),
    .A2(net5995),
    .A1(\top1.memory2.mem2[197][2] ));
 sg13g2_a221oi_1 _15870_ (.B2(\top1.memory2.mem2[198][2] ),
    .C1(_03827_),
    .B1(net5915),
    .A1(\top1.memory2.mem2[196][2] ),
    .Y(_06265_),
    .A2(net6060));
 sg13g2_a221oi_1 _15871_ (.B2(_06265_),
    .C1(_03979_),
    .B1(_06264_),
    .A1(_06261_),
    .Y(_06266_),
    .A2(_06263_));
 sg13g2_nor2b_1 _15872_ (.A(_06266_),
    .B_N(net6109),
    .Y(_06267_));
 sg13g2_o21ai_1 _15873_ (.B1(_06267_),
    .Y(_06268_),
    .A1(net5831),
    .A2(_06260_));
 sg13g2_o21ai_1 _15874_ (.B1(\top1.fsm.re ),
    .Y(_06269_),
    .A1(_06225_),
    .A2(_06268_));
 sg13g2_o21ai_1 _15875_ (.B1(_05994_),
    .Y(_01020_),
    .A1(_06127_),
    .A2(_06269_));
 sg13g2_xor2_1 _15876_ (.B(_05040_),
    .A(\top1.event_time[16] ),
    .X(_01021_));
 sg13g2_a21o_1 _15877_ (.A2(_05040_),
    .A1(\top1.event_time[16] ),
    .B1(\top1.event_time[17] ),
    .X(_06270_));
 sg13g2_and2_1 _15878_ (.A(_05041_),
    .B(_06270_),
    .X(_01022_));
 sg13g2_nand4_1 _15879_ (.B(\top1.event_time[16] ),
    .C(\top1.event_time[18] ),
    .A(\top1.event_time[17] ),
    .Y(_06271_),
    .D(_05040_));
 sg13g2_nand2_1 _15880_ (.Y(_06272_),
    .A(net6897),
    .B(_06271_));
 sg13g2_a21oi_1 _15881_ (.A1(_03840_),
    .A2(_05041_),
    .Y(_01023_),
    .B1(_06272_));
 sg13g2_nor2_1 _15882_ (.A(_03839_),
    .B(_06271_),
    .Y(_06273_));
 sg13g2_nand2_1 _15883_ (.Y(_06274_),
    .A(\top1.event_time[19] ),
    .B(net6897));
 sg13g2_a21oi_1 _15884_ (.A1(_06271_),
    .A2(_06274_),
    .Y(_01024_),
    .B1(_06273_));
 sg13g2_nor2_1 _15885_ (.A(\top1.event_time[20] ),
    .B(_06273_),
    .Y(_06275_));
 sg13g2_nand2_1 _15886_ (.Y(_06276_),
    .A(\top1.event_time[20] ),
    .B(_06273_));
 sg13g2_nand2_1 _15887_ (.Y(_06277_),
    .A(_05043_),
    .B(_06276_));
 sg13g2_nor2_1 _15888_ (.A(_06275_),
    .B(_06277_),
    .Y(_01025_));
 sg13g2_nand3_1 _15889_ (.B(_05043_),
    .C(_06276_),
    .A(\top1.event_time[21] ),
    .Y(_06278_));
 sg13g2_o21ai_1 _15890_ (.B1(_06278_),
    .Y(_01026_),
    .A1(\top1.event_time[21] ),
    .A2(_06276_));
 sg13g2_nand3_1 _15891_ (.B(net7260),
    .C(net7214),
    .A(net7265),
    .Y(_06279_));
 sg13g2_nand2_1 _15892_ (.Y(_06280_),
    .A(net3703),
    .B(net6826));
 sg13g2_o21ai_1 _15893_ (.B1(_06280_),
    .Y(_01027_),
    .A1(net7329),
    .A2(net6826));
 sg13g2_nand2_1 _15894_ (.Y(_06281_),
    .A(net4338),
    .B(net6825));
 sg13g2_o21ai_1 _15895_ (.B1(_06281_),
    .Y(_01028_),
    .A1(net7528),
    .A2(net6825));
 sg13g2_nand2_1 _15896_ (.Y(_06282_),
    .A(net3561),
    .B(net6825));
 sg13g2_o21ai_1 _15897_ (.B1(_06282_),
    .Y(_01029_),
    .A1(net7687),
    .A2(net6825));
 sg13g2_nand3_1 _15898_ (.B(net7075),
    .C(net7222),
    .A(net7277),
    .Y(_06283_));
 sg13g2_nand2_1 _15899_ (.Y(_06284_),
    .A(net3060),
    .B(net6360));
 sg13g2_o21ai_1 _15900_ (.B1(_06284_),
    .Y(_01030_),
    .A1(net7358),
    .A2(net6360));
 sg13g2_nand2_1 _15901_ (.Y(_06285_),
    .A(net2509),
    .B(net6361));
 sg13g2_o21ai_1 _15902_ (.B1(_06285_),
    .Y(_01031_),
    .A1(net7554),
    .A2(net6361));
 sg13g2_nand2_1 _15903_ (.Y(_06286_),
    .A(net3382),
    .B(net6360));
 sg13g2_o21ai_1 _15904_ (.B1(_06286_),
    .Y(_01032_),
    .A1(net7715),
    .A2(net6360));
 sg13g2_nand3_1 _15905_ (.B(net7075),
    .C(net7222),
    .A(net7273),
    .Y(_06287_));
 sg13g2_nand2_1 _15906_ (.Y(_06288_),
    .A(net3249),
    .B(net6358));
 sg13g2_o21ai_1 _15907_ (.B1(_06288_),
    .Y(_01033_),
    .A1(net7357),
    .A2(net6358));
 sg13g2_nand2_1 _15908_ (.Y(_06289_),
    .A(net3872),
    .B(net6359));
 sg13g2_o21ai_1 _15909_ (.B1(_06289_),
    .Y(_01034_),
    .A1(net7554),
    .A2(net6359));
 sg13g2_nand2_1 _15910_ (.Y(_06290_),
    .A(net3839),
    .B(net6358));
 sg13g2_o21ai_1 _15911_ (.B1(_06290_),
    .Y(_01035_),
    .A1(net7715),
    .A2(net6358));
 sg13g2_nand3_1 _15912_ (.B(net7241),
    .C(net7212),
    .A(net7285),
    .Y(_06291_));
 sg13g2_nand2_1 _15913_ (.Y(_06292_),
    .A(net3430),
    .B(net6824));
 sg13g2_o21ai_1 _15914_ (.B1(_06292_),
    .Y(_01036_),
    .A1(net7333),
    .A2(net6823));
 sg13g2_nand2_1 _15915_ (.Y(_06293_),
    .A(net3830),
    .B(net6824));
 sg13g2_o21ai_1 _15916_ (.B1(_06293_),
    .Y(_01037_),
    .A1(net7533),
    .A2(net6823));
 sg13g2_nand2_1 _15917_ (.Y(_06294_),
    .A(net2989),
    .B(net6824));
 sg13g2_o21ai_1 _15918_ (.B1(_06294_),
    .Y(_01038_),
    .A1(net7689),
    .A2(net6824));
 sg13g2_nor3_1 _15919_ (.A(net7098),
    .B(net7272),
    .C(net7202),
    .Y(_06295_));
 sg13g2_nor2_1 _15920_ (.A(net4280),
    .B(net6356),
    .Y(_06296_));
 sg13g2_a21oi_1 _15921_ (.A1(net7330),
    .A2(net6357),
    .Y(_01039_),
    .B1(_06296_));
 sg13g2_nor2_1 _15922_ (.A(net4838),
    .B(net6356),
    .Y(_06297_));
 sg13g2_a21oi_1 _15923_ (.A1(net7535),
    .A2(net6356),
    .Y(_01040_),
    .B1(_06297_));
 sg13g2_nor2_1 _15924_ (.A(net4264),
    .B(net6356),
    .Y(_06298_));
 sg13g2_a21oi_1 _15925_ (.A1(net7686),
    .A2(net6356),
    .Y(_01041_),
    .B1(_06298_));
 sg13g2_nor3_2 _15926_ (.A(net7272),
    .B(net7267),
    .C(net7200),
    .Y(_06299_));
 sg13g2_nor2_1 _15927_ (.A(net4348),
    .B(net6822),
    .Y(_06300_));
 sg13g2_a21oi_1 _15928_ (.A1(net7311),
    .A2(net6822),
    .Y(_01042_),
    .B1(_06300_));
 sg13g2_nor2_1 _15929_ (.A(net4361),
    .B(net6822),
    .Y(_06301_));
 sg13g2_a21oi_1 _15930_ (.A1(net7509),
    .A2(net6822),
    .Y(_01043_),
    .B1(_06301_));
 sg13g2_nor2_1 _15931_ (.A(net4253),
    .B(net6821),
    .Y(_06302_));
 sg13g2_a21oi_1 _15932_ (.A1(net7666),
    .A2(net6821),
    .Y(_01044_),
    .B1(_06302_));
 sg13g2_nor3_1 _15933_ (.A(net7276),
    .B(net7098),
    .C(net7202),
    .Y(_06303_));
 sg13g2_nor2_1 _15934_ (.A(net4019),
    .B(net6354),
    .Y(_06304_));
 sg13g2_a21oi_1 _15935_ (.A1(net7330),
    .A2(net6355),
    .Y(_01045_),
    .B1(_06304_));
 sg13g2_nor2_1 _15936_ (.A(net4587),
    .B(net6354),
    .Y(_06305_));
 sg13g2_a21oi_1 _15937_ (.A1(net7535),
    .A2(net6354),
    .Y(_01046_),
    .B1(_06305_));
 sg13g2_nor2_1 _15938_ (.A(net4700),
    .B(net6354),
    .Y(_06306_));
 sg13g2_a21oi_1 _15939_ (.A1(net7686),
    .A2(net6354),
    .Y(_01047_),
    .B1(_06306_));
 sg13g2_nor3_1 _15940_ (.A(net7097),
    .B(net7246),
    .C(net7202),
    .Y(_06307_));
 sg13g2_nor2_1 _15941_ (.A(net4220),
    .B(net6353),
    .Y(_06308_));
 sg13g2_a21oi_1 _15942_ (.A1(net7330),
    .A2(net6352),
    .Y(_01048_),
    .B1(_06308_));
 sg13g2_nor2_1 _15943_ (.A(net4813),
    .B(net6352),
    .Y(_06309_));
 sg13g2_a21oi_1 _15944_ (.A1(net7535),
    .A2(net6352),
    .Y(_01049_),
    .B1(_06309_));
 sg13g2_nor2_1 _15945_ (.A(net4103),
    .B(net6352),
    .Y(_06310_));
 sg13g2_a21oi_1 _15946_ (.A1(net7686),
    .A2(net6352),
    .Y(_01050_),
    .B1(_06310_));
 sg13g2_nand3_1 _15947_ (.B(net7236),
    .C(net7210),
    .A(net7242),
    .Y(_06311_));
 sg13g2_nand2_1 _15948_ (.Y(_06312_),
    .A(net2643),
    .B(net6819));
 sg13g2_o21ai_1 _15949_ (.B1(_06312_),
    .Y(_01051_),
    .A1(net7326),
    .A2(net6819));
 sg13g2_nand2_1 _15950_ (.Y(_06313_),
    .A(net2564),
    .B(net6819));
 sg13g2_o21ai_1 _15951_ (.B1(_06313_),
    .Y(_01052_),
    .A1(net7525),
    .A2(net6819));
 sg13g2_nand2_1 _15952_ (.Y(_06314_),
    .A(net3718),
    .B(net6819));
 sg13g2_o21ai_1 _15953_ (.B1(_06314_),
    .Y(_01053_),
    .A1(net7682),
    .A2(net6819));
 sg13g2_nor2_1 _15954_ (.A(\top1.memory1.mem1[85][0] ),
    .B(net5973),
    .Y(_06315_));
 sg13g2_nor2_1 _15955_ (.A(\top1.memory1.mem1[86][0] ),
    .B(net5894),
    .Y(_06316_));
 sg13g2_nor2_1 _15956_ (.A(\top1.memory1.mem1[87][0] ),
    .B(net5933),
    .Y(_06317_));
 sg13g2_o21ai_1 _15957_ (.B1(net6021),
    .Y(_06318_),
    .A1(\top1.memory1.mem1[84][0] ),
    .A2(net6039));
 sg13g2_nor4_1 _15958_ (.A(_06315_),
    .B(_06316_),
    .C(_06317_),
    .D(_06318_),
    .Y(_06319_));
 sg13g2_a22oi_1 _15959_ (.Y(_06320_),
    .B1(net5952),
    .B2(\top1.memory1.mem1[95][0] ),
    .A2(net6057),
    .A1(\top1.memory1.mem1[92][0] ));
 sg13g2_a22oi_1 _15960_ (.Y(_06321_),
    .B1(net5912),
    .B2(\top1.memory1.mem1[94][0] ),
    .A2(net5992),
    .A1(\top1.memory1.mem1[93][0] ));
 sg13g2_a21oi_1 _15961_ (.A1(_06320_),
    .A2(_06321_),
    .Y(_06322_),
    .B1(net5845));
 sg13g2_mux4_1 _15962_ (.S0(net6209),
    .A0(\top1.memory1.mem1[80][0] ),
    .A1(\top1.memory1.mem1[81][0] ),
    .A2(\top1.memory1.mem1[82][0] ),
    .A3(\top1.memory1.mem1[83][0] ),
    .S1(net6144),
    .X(_06323_));
 sg13g2_a22oi_1 _15963_ (.Y(_06324_),
    .B1(net5911),
    .B2(\top1.memory1.mem1[90][0] ),
    .A2(net6056),
    .A1(\top1.memory1.mem1[88][0] ));
 sg13g2_a22oi_1 _15964_ (.Y(_06325_),
    .B1(net5951),
    .B2(\top1.memory1.mem1[91][0] ),
    .A2(net5993),
    .A1(\top1.memory1.mem1[89][0] ));
 sg13g2_a21oi_1 _15965_ (.A1(_06324_),
    .A2(_06325_),
    .Y(_06326_),
    .B1(net6077));
 sg13g2_a21o_1 _15966_ (.A2(_06323_),
    .A1(net5877),
    .B1(net6104),
    .X(_06327_));
 sg13g2_nor4_1 _15967_ (.A(_06319_),
    .B(_06322_),
    .C(_06326_),
    .D(_06327_),
    .Y(_06328_));
 sg13g2_nor2_1 _15968_ (.A(\top1.memory1.mem1[70][0] ),
    .B(net5890),
    .Y(_06329_));
 sg13g2_nor2_1 _15969_ (.A(\top1.memory1.mem1[68][0] ),
    .B(net6036),
    .Y(_06330_));
 sg13g2_nor2_1 _15970_ (.A(\top1.memory1.mem1[69][0] ),
    .B(net5970),
    .Y(_06331_));
 sg13g2_o21ai_1 _15971_ (.B1(net6018),
    .Y(_06332_),
    .A1(\top1.memory1.mem1[71][0] ),
    .A2(net5932));
 sg13g2_nor4_2 _15972_ (.A(_06329_),
    .B(_06330_),
    .C(_06331_),
    .Y(_06333_),
    .D(_06332_));
 sg13g2_a22oi_1 _15973_ (.Y(_06334_),
    .B1(net5901),
    .B2(\top1.memory1.mem1[74][0] ),
    .A2(net5942),
    .A1(\top1.memory1.mem1[75][0] ));
 sg13g2_a22oi_1 _15974_ (.Y(_06335_),
    .B1(net5981),
    .B2(\top1.memory1.mem1[73][0] ),
    .A2(net6046),
    .A1(\top1.memory1.mem1[72][0] ));
 sg13g2_a21oi_1 _15975_ (.A1(_06334_),
    .A2(_06335_),
    .Y(_06336_),
    .B1(net6075));
 sg13g2_mux4_1 _15976_ (.S0(net6197),
    .A0(\top1.memory1.mem1[76][0] ),
    .A1(\top1.memory1.mem1[77][0] ),
    .A2(\top1.memory1.mem1[78][0] ),
    .A3(\top1.memory1.mem1[79][0] ),
    .S1(net6133),
    .X(_06337_));
 sg13g2_a22oi_1 _15977_ (.Y(_06338_),
    .B1(net5942),
    .B2(\top1.memory1.mem1[67][0] ),
    .A2(net6046),
    .A1(\top1.memory1.mem1[64][0] ));
 sg13g2_a22oi_1 _15978_ (.Y(_06339_),
    .B1(net5901),
    .B2(\top1.memory1.mem1[66][0] ),
    .A2(net5982),
    .A1(\top1.memory1.mem1[65][0] ));
 sg13g2_a21oi_1 _15979_ (.A1(_06338_),
    .A2(_06339_),
    .Y(_06340_),
    .B1(net5868));
 sg13g2_a21o_1 _15980_ (.A2(_06337_),
    .A1(net5850),
    .B1(net6120),
    .X(_06341_));
 sg13g2_nor4_2 _15981_ (.A(_06333_),
    .B(_06336_),
    .C(_06340_),
    .Y(_06342_),
    .D(_06341_));
 sg13g2_mux4_1 _15982_ (.S0(net6244),
    .A0(\top1.memory1.mem1[116][0] ),
    .A1(\top1.memory1.mem1[117][0] ),
    .A2(\top1.memory1.mem1[118][0] ),
    .A3(\top1.memory1.mem1[119][0] ),
    .S1(net6179),
    .X(_06343_));
 sg13g2_mux4_1 _15983_ (.S0(net6245),
    .A0(\top1.memory1.mem1[124][0] ),
    .A1(\top1.memory1.mem1[125][0] ),
    .A2(\top1.memory1.mem1[126][0] ),
    .A3(\top1.memory1.mem1[127][0] ),
    .S1(net6180),
    .X(_06344_));
 sg13g2_a22oi_1 _15984_ (.Y(_06345_),
    .B1(_06344_),
    .B2(net5861),
    .A2(_06343_),
    .A1(net6030));
 sg13g2_mux4_1 _15985_ (.S0(net6241),
    .A0(\top1.memory1.mem1[120][0] ),
    .A1(\top1.memory1.mem1[121][0] ),
    .A2(\top1.memory1.mem1[122][0] ),
    .A3(\top1.memory1.mem1[123][0] ),
    .S1(net6176),
    .X(_06346_));
 sg13g2_mux4_1 _15986_ (.S0(net6245),
    .A0(\top1.memory1.mem1[112][0] ),
    .A1(\top1.memory1.mem1[113][0] ),
    .A2(\top1.memory1.mem1[114][0] ),
    .A3(\top1.memory1.mem1[115][0] ),
    .S1(net6180),
    .X(_06347_));
 sg13g2_a22oi_1 _15987_ (.Y(_06348_),
    .B1(_06347_),
    .B2(net5889),
    .A2(_06346_),
    .A1(net6094));
 sg13g2_a21oi_2 _15988_ (.B1(net5838),
    .Y(_06349_),
    .A2(_06348_),
    .A1(_06345_));
 sg13g2_mux4_1 _15989_ (.S0(net6239),
    .A0(\top1.memory1.mem1[108][0] ),
    .A1(\top1.memory1.mem1[109][0] ),
    .A2(\top1.memory1.mem1[110][0] ),
    .A3(\top1.memory1.mem1[111][0] ),
    .S1(net6174),
    .X(_06350_));
 sg13g2_mux4_1 _15990_ (.S0(net6239),
    .A0(\top1.memory1.mem1[100][0] ),
    .A1(\top1.memory1.mem1[101][0] ),
    .A2(\top1.memory1.mem1[102][0] ),
    .A3(\top1.memory1.mem1[103][0] ),
    .S1(net6174),
    .X(_06351_));
 sg13g2_mux4_1 _15991_ (.S0(net6226),
    .A0(\top1.memory1.mem1[96][0] ),
    .A1(\top1.memory1.mem1[97][0] ),
    .A2(\top1.memory1.mem1[98][0] ),
    .A3(\top1.memory1.mem1[99][0] ),
    .S1(net6161),
    .X(_06352_));
 sg13g2_mux4_1 _15992_ (.S0(net6249),
    .A0(\top1.memory1.mem1[104][0] ),
    .A1(\top1.memory1.mem1[105][0] ),
    .A2(\top1.memory1.mem1[106][0] ),
    .A3(\top1.memory1.mem1[107][0] ),
    .S1(net6184),
    .X(_06353_));
 sg13g2_a22oi_1 _15993_ (.Y(_06354_),
    .B1(_06352_),
    .B2(net5885),
    .A2(_06350_),
    .A1(net5860));
 sg13g2_a22oi_1 _15994_ (.Y(_06355_),
    .B1(_06353_),
    .B2(net6093),
    .A2(_06351_),
    .A1(net6031));
 sg13g2_a21oi_1 _15995_ (.A1(_06354_),
    .A2(_06355_),
    .Y(_06356_),
    .B1(net5833));
 sg13g2_mux4_1 _15996_ (.S0(net6211),
    .A0(\top1.memory1.mem1[0][0] ),
    .A1(\top1.memory1.mem1[1][0] ),
    .A2(\top1.memory1.mem1[2][0] ),
    .A3(\top1.memory1.mem1[3][0] ),
    .S1(net6146),
    .X(_06357_));
 sg13g2_a21o_1 _15997_ (.A2(_06357_),
    .A1(net5878),
    .B1(net6124),
    .X(_06358_));
 sg13g2_o21ai_1 _15998_ (.B1(net6022),
    .Y(_06359_),
    .A1(\top1.memory1.mem1[4][0] ),
    .A2(net6043));
 sg13g2_nor2_1 _15999_ (.A(\top1.memory1.mem1[6][0] ),
    .B(net5897),
    .Y(_06360_));
 sg13g2_nor2_1 _16000_ (.A(\top1.memory1.mem1[7][0] ),
    .B(net5938),
    .Y(_06361_));
 sg13g2_nor2_1 _16001_ (.A(\top1.memory1.mem1[5][0] ),
    .B(net5977),
    .Y(_06362_));
 sg13g2_or4_1 _16002_ (.A(_06359_),
    .B(_06360_),
    .C(_06361_),
    .D(_06362_),
    .X(_06363_));
 sg13g2_mux4_1 _16003_ (.S0(net6212),
    .A0(\top1.memory1.mem1[8][0] ),
    .A1(\top1.memory1.mem1[9][0] ),
    .A2(\top1.memory1.mem1[10][0] ),
    .A3(\top1.memory1.mem1[11][0] ),
    .S1(net6147),
    .X(_06364_));
 sg13g2_mux4_1 _16004_ (.S0(net6213),
    .A0(\top1.memory1.mem1[12][0] ),
    .A1(\top1.memory1.mem1[13][0] ),
    .A2(\top1.memory1.mem1[14][0] ),
    .A3(\top1.memory1.mem1[15][0] ),
    .S1(net6148),
    .X(_06365_));
 sg13g2_a221oi_1 _16005_ (.B2(net5853),
    .C1(_06358_),
    .B1(_06365_),
    .A1(net6087),
    .Y(_06366_),
    .A2(_06364_));
 sg13g2_mux4_1 _16006_ (.S0(net6229),
    .A0(\top1.memory1.mem1[16][0] ),
    .A1(\top1.memory1.mem1[17][0] ),
    .A2(\top1.memory1.mem1[18][0] ),
    .A3(\top1.memory1.mem1[19][0] ),
    .S1(net6164),
    .X(_06367_));
 sg13g2_mux4_1 _16007_ (.S0(net6231),
    .A0(\top1.memory1.mem1[24][0] ),
    .A1(\top1.memory1.mem1[25][0] ),
    .A2(\top1.memory1.mem1[26][0] ),
    .A3(\top1.memory1.mem1[27][0] ),
    .S1(net6166),
    .X(_06368_));
 sg13g2_nor3_1 _16008_ (.A(net6228),
    .B(net6157),
    .C(\top1.memory1.mem1[20][0] ),
    .Y(_06369_));
 sg13g2_a21oi_1 _16009_ (.A1(_03880_),
    .A2(net5959),
    .Y(_06370_),
    .B1(net6012));
 sg13g2_a221oi_1 _16010_ (.B2(_03879_),
    .C1(_06369_),
    .B1(net5919),
    .A1(_03878_),
    .Y(_06371_),
    .A2(net6001));
 sg13g2_mux4_1 _16011_ (.S0(net6222),
    .A0(\top1.memory1.mem1[28][0] ),
    .A1(\top1.memory1.mem1[29][0] ),
    .A2(\top1.memory1.mem1[30][0] ),
    .A3(\top1.memory1.mem1[31][0] ),
    .S1(net6157),
    .X(_06372_));
 sg13g2_a22oi_1 _16012_ (.Y(_06373_),
    .B1(_06372_),
    .B2(net5856),
    .A2(_06371_),
    .A1(_06370_));
 sg13g2_a221oi_1 _16013_ (.B2(net6091),
    .C1(net6107),
    .B1(_06368_),
    .A1(net5882),
    .Y(_06374_),
    .A2(_06367_));
 sg13g2_a221oi_1 _16014_ (.B2(_06374_),
    .C1(net6118),
    .B1(_06373_),
    .A1(_06363_),
    .Y(_06375_),
    .A2(_06366_));
 sg13g2_mux4_1 _16015_ (.S0(net6245),
    .A0(\top1.memory1.mem1[60][0] ),
    .A1(\top1.memory1.mem1[61][0] ),
    .A2(\top1.memory1.mem1[62][0] ),
    .A3(\top1.memory1.mem1[63][0] ),
    .S1(net6180),
    .X(_06376_));
 sg13g2_mux4_1 _16016_ (.S0(net6255),
    .A0(\top1.memory1.mem1[48][0] ),
    .A1(\top1.memory1.mem1[49][0] ),
    .A2(\top1.memory1.mem1[50][0] ),
    .A3(\top1.memory1.mem1[51][0] ),
    .S1(net6190),
    .X(_06377_));
 sg13g2_mux4_1 _16017_ (.S0(net6254),
    .A0(\top1.memory1.mem1[56][0] ),
    .A1(\top1.memory1.mem1[57][0] ),
    .A2(\top1.memory1.mem1[58][0] ),
    .A3(\top1.memory1.mem1[59][0] ),
    .S1(net6189),
    .X(_06378_));
 sg13g2_mux4_1 _16018_ (.S0(net6254),
    .A0(\top1.memory1.mem1[52][0] ),
    .A1(\top1.memory1.mem1[53][0] ),
    .A2(\top1.memory1.mem1[54][0] ),
    .A3(\top1.memory1.mem1[55][0] ),
    .S1(net6189),
    .X(_06379_));
 sg13g2_a22oi_1 _16019_ (.Y(_06380_),
    .B1(_06378_),
    .B2(net6097),
    .A2(_06376_),
    .A1(net5864));
 sg13g2_a22oi_1 _16020_ (.Y(_06381_),
    .B1(_06379_),
    .B2(net6033),
    .A2(_06377_),
    .A1(net5886));
 sg13g2_a21oi_1 _16021_ (.A1(_06380_),
    .A2(_06381_),
    .Y(_06382_),
    .B1(net5840));
 sg13g2_mux4_1 _16022_ (.S0(net6255),
    .A0(\top1.memory1.mem1[44][0] ),
    .A1(\top1.memory1.mem1[45][0] ),
    .A2(\top1.memory1.mem1[46][0] ),
    .A3(\top1.memory1.mem1[47][0] ),
    .S1(net6190),
    .X(_06383_));
 sg13g2_mux4_1 _16023_ (.S0(net6257),
    .A0(\top1.memory1.mem1[32][0] ),
    .A1(\top1.memory1.mem1[33][0] ),
    .A2(\top1.memory1.mem1[34][0] ),
    .A3(\top1.memory1.mem1[35][0] ),
    .S1(net6192),
    .X(_06384_));
 sg13g2_mux4_1 _16024_ (.S0(net6258),
    .A0(\top1.memory1.mem1[36][0] ),
    .A1(\top1.memory1.mem1[37][0] ),
    .A2(\top1.memory1.mem1[38][0] ),
    .A3(\top1.memory1.mem1[39][0] ),
    .S1(net6193),
    .X(_06385_));
 sg13g2_mux4_1 _16025_ (.S0(net6257),
    .A0(\top1.memory1.mem1[40][0] ),
    .A1(\top1.memory1.mem1[41][0] ),
    .A2(\top1.memory1.mem1[42][0] ),
    .A3(\top1.memory1.mem1[43][0] ),
    .S1(net6192),
    .X(_06386_));
 sg13g2_a22oi_1 _16026_ (.Y(_06387_),
    .B1(_06385_),
    .B2(net6033),
    .A2(_06383_),
    .A1(net5865));
 sg13g2_a22oi_1 _16027_ (.Y(_06388_),
    .B1(_06386_),
    .B2(net6098),
    .A2(_06384_),
    .A1(net5886));
 sg13g2_a21oi_1 _16028_ (.A1(_06387_),
    .A2(_06388_),
    .Y(_06389_),
    .B1(net5835));
 sg13g2_or2_2 _16029_ (.X(_06390_),
    .B(_06389_),
    .A(_06382_));
 sg13g2_o21ai_1 _16030_ (.B1(net6102),
    .Y(_06391_),
    .A1(_06375_),
    .A2(_06390_));
 sg13g2_or3_2 _16031_ (.A(_05479_),
    .B(_06328_),
    .C(_06342_),
    .X(_06392_));
 sg13g2_o21ai_1 _16032_ (.B1(net6116),
    .Y(_06393_),
    .A1(_06349_),
    .A2(_06356_));
 sg13g2_nand4_1 _16033_ (.B(_06391_),
    .C(_06392_),
    .A(_03831_),
    .Y(_06394_),
    .D(_06393_));
 sg13g2_o21ai_1 _16034_ (.B1(net6016),
    .Y(_06395_),
    .A1(\top1.memory1.mem1[149][0] ),
    .A2(net5971));
 sg13g2_nor2_1 _16035_ (.A(\top1.memory1.mem1[148][0] ),
    .B(net6037),
    .Y(_06396_));
 sg13g2_nor2_1 _16036_ (.A(\top1.memory1.mem1[151][0] ),
    .B(net5934),
    .Y(_06397_));
 sg13g2_nor2_1 _16037_ (.A(\top1.memory1.mem1[150][0] ),
    .B(net5890),
    .Y(_06398_));
 sg13g2_nor4_2 _16038_ (.A(_06395_),
    .B(_06396_),
    .C(_06397_),
    .Y(_06399_),
    .D(_06398_));
 sg13g2_a22oi_1 _16039_ (.Y(_06400_),
    .B1(net5909),
    .B2(\top1.memory1.mem1[158][0] ),
    .A2(net5948),
    .A1(\top1.memory1.mem1[159][0] ));
 sg13g2_a22oi_1 _16040_ (.Y(_06401_),
    .B1(net5990),
    .B2(\top1.memory1.mem1[157][0] ),
    .A2(net6054),
    .A1(\top1.memory1.mem1[156][0] ));
 sg13g2_a21oi_2 _16041_ (.B1(net5843),
    .Y(_06402_),
    .A2(_06401_),
    .A1(_06400_));
 sg13g2_mux4_1 _16042_ (.S0(net6205),
    .A0(\top1.memory1.mem1[144][0] ),
    .A1(\top1.memory1.mem1[145][0] ),
    .A2(\top1.memory1.mem1[146][0] ),
    .A3(\top1.memory1.mem1[147][0] ),
    .S1(net6141),
    .X(_06403_));
 sg13g2_a22oi_1 _16043_ (.Y(_06404_),
    .B1(net5908),
    .B2(\top1.memory1.mem1[154][0] ),
    .A2(net6053),
    .A1(\top1.memory1.mem1[152][0] ));
 sg13g2_a22oi_1 _16044_ (.Y(_06405_),
    .B1(net5949),
    .B2(\top1.memory1.mem1[155][0] ),
    .A2(net5989),
    .A1(\top1.memory1.mem1[153][0] ));
 sg13g2_a21oi_1 _16045_ (.A1(_06404_),
    .A2(_06405_),
    .Y(_06406_),
    .B1(net6076));
 sg13g2_a21o_1 _16046_ (.A2(_06403_),
    .A1(net5876),
    .B1(net6105),
    .X(_06407_));
 sg13g2_nor4_1 _16047_ (.A(_06399_),
    .B(_06402_),
    .C(_06406_),
    .D(_06407_),
    .Y(_06408_));
 sg13g2_mux4_1 _16048_ (.S0(net6199),
    .A0(\top1.memory1.mem1[128][0] ),
    .A1(\top1.memory1.mem1[129][0] ),
    .A2(\top1.memory1.mem1[130][0] ),
    .A3(\top1.memory1.mem1[131][0] ),
    .S1(net6135),
    .X(_06409_));
 sg13g2_nand2_1 _16049_ (.Y(_06410_),
    .A(net5875),
    .B(_06409_));
 sg13g2_mux4_1 _16050_ (.S0(net6203),
    .A0(\top1.memory1.mem1[140][0] ),
    .A1(\top1.memory1.mem1[141][0] ),
    .A2(\top1.memory1.mem1[142][0] ),
    .A3(\top1.memory1.mem1[143][0] ),
    .S1(net6139),
    .X(_06411_));
 sg13g2_o21ai_1 _16051_ (.B1(net6019),
    .Y(_06412_),
    .A1(\top1.memory1.mem1[134][0] ),
    .A2(net5891));
 sg13g2_nor2_1 _16052_ (.A(\top1.memory1.mem1[135][0] ),
    .B(net5930),
    .Y(_06413_));
 sg13g2_nor2_1 _16053_ (.A(\top1.memory1.mem1[133][0] ),
    .B(net5970),
    .Y(_06414_));
 sg13g2_nor2_1 _16054_ (.A(\top1.memory1.mem1[132][0] ),
    .B(net6036),
    .Y(_06415_));
 sg13g2_nor4_1 _16055_ (.A(_06412_),
    .B(_06413_),
    .C(_06414_),
    .D(_06415_),
    .Y(_06416_));
 sg13g2_mux4_1 _16056_ (.S0(net6203),
    .A0(\top1.memory1.mem1[136][0] ),
    .A1(\top1.memory1.mem1[137][0] ),
    .A2(\top1.memory1.mem1[138][0] ),
    .A3(\top1.memory1.mem1[139][0] ),
    .S1(net6139),
    .X(_06417_));
 sg13g2_a22oi_1 _16057_ (.Y(_06418_),
    .B1(_06417_),
    .B2(net6084),
    .A2(_06411_),
    .A1(net5851));
 sg13g2_nand2_1 _16058_ (.Y(_06419_),
    .A(_06410_),
    .B(_06418_));
 sg13g2_nor3_1 _16059_ (.A(net6122),
    .B(_06416_),
    .C(_06419_),
    .Y(_06420_));
 sg13g2_or3_2 _16060_ (.A(net6117),
    .B(_06408_),
    .C(_06420_),
    .X(_06421_));
 sg13g2_mux4_1 _16061_ (.S0(net6220),
    .A0(\top1.memory1.mem1[164][0] ),
    .A1(\top1.memory1.mem1[165][0] ),
    .A2(\top1.memory1.mem1[166][0] ),
    .A3(\top1.memory1.mem1[167][0] ),
    .S1(net6155),
    .X(_06422_));
 sg13g2_a22oi_1 _16062_ (.Y(_06423_),
    .B1(net5918),
    .B2(\top1.memory1.mem1[162][0] ),
    .A2(net5958),
    .A1(\top1.memory1.mem1[163][0] ));
 sg13g2_a22oi_1 _16063_ (.Y(_06424_),
    .B1(net5999),
    .B2(\top1.memory1.mem1[161][0] ),
    .A2(net6063),
    .A1(\top1.memory1.mem1[160][0] ));
 sg13g2_a21o_1 _16064_ (.A2(_06424_),
    .A1(_06423_),
    .B1(net5870),
    .X(_06425_));
 sg13g2_mux4_1 _16065_ (.S0(net6220),
    .A0(\top1.memory1.mem1[172][0] ),
    .A1(\top1.memory1.mem1[173][0] ),
    .A2(\top1.memory1.mem1[174][0] ),
    .A3(\top1.memory1.mem1[175][0] ),
    .S1(net6155),
    .X(_06426_));
 sg13g2_mux4_1 _16066_ (.S0(net6221),
    .A0(\top1.memory1.mem1[168][0] ),
    .A1(\top1.memory1.mem1[169][0] ),
    .A2(\top1.memory1.mem1[170][0] ),
    .A3(\top1.memory1.mem1[171][0] ),
    .S1(net6156),
    .X(_06427_));
 sg13g2_and2_1 _16067_ (.A(net6089),
    .B(_06427_),
    .X(_06428_));
 sg13g2_a221oi_1 _16068_ (.B2(net5856),
    .C1(_06428_),
    .B1(_06426_),
    .A1(net6026),
    .Y(_06429_),
    .A2(_06422_));
 sg13g2_a21oi_1 _16069_ (.A1(_06425_),
    .A2(_06429_),
    .Y(_06430_),
    .B1(net5836));
 sg13g2_mux4_1 _16070_ (.S0(net6225),
    .A0(\top1.memory1.mem1[188][0] ),
    .A1(\top1.memory1.mem1[189][0] ),
    .A2(\top1.memory1.mem1[190][0] ),
    .A3(\top1.memory1.mem1[191][0] ),
    .S1(net6160),
    .X(_06431_));
 sg13g2_mux4_1 _16071_ (.S0(net6221),
    .A0(\top1.memory1.mem1[184][0] ),
    .A1(\top1.memory1.mem1[185][0] ),
    .A2(\top1.memory1.mem1[186][0] ),
    .A3(\top1.memory1.mem1[187][0] ),
    .S1(net6156),
    .X(_06432_));
 sg13g2_mux4_1 _16072_ (.S0(net6225),
    .A0(\top1.memory1.mem1[176][0] ),
    .A1(\top1.memory1.mem1[177][0] ),
    .A2(\top1.memory1.mem1[178][0] ),
    .A3(\top1.memory1.mem1[179][0] ),
    .S1(net6160),
    .X(_06433_));
 sg13g2_mux4_1 _16073_ (.S0(net6224),
    .A0(\top1.memory1.mem1[180][0] ),
    .A1(\top1.memory1.mem1[181][0] ),
    .A2(\top1.memory1.mem1[182][0] ),
    .A3(\top1.memory1.mem1[183][0] ),
    .S1(net6159),
    .X(_06434_));
 sg13g2_a22oi_1 _16074_ (.Y(_06435_),
    .B1(_06433_),
    .B2(net5881),
    .A2(_06431_),
    .A1(net5857));
 sg13g2_a22oi_1 _16075_ (.Y(_06436_),
    .B1(_06434_),
    .B2(net6025),
    .A2(_06432_),
    .A1(net6090));
 sg13g2_a21oi_2 _16076_ (.B1(net5837),
    .Y(_06437_),
    .A2(_06436_),
    .A1(_06435_));
 sg13g2_nor3_2 _16077_ (.A(net5831),
    .B(_06430_),
    .C(_06437_),
    .Y(_06438_));
 sg13g2_nor2_1 _16078_ (.A(\top1.memory1.mem1[193][0] ),
    .B(net5977),
    .Y(_06439_));
 sg13g2_nor2_1 _16079_ (.A(\top1.memory1.mem1[194][0] ),
    .B(net5897),
    .Y(_06440_));
 sg13g2_nor2_1 _16080_ (.A(\top1.memory1.mem1[192][0] ),
    .B(net6043),
    .Y(_06441_));
 sg13g2_nor4_1 _16081_ (.A(net6131),
    .B(_06439_),
    .C(_06440_),
    .D(_06441_),
    .Y(_06442_));
 sg13g2_o21ai_1 _16082_ (.B1(_06442_),
    .Y(_06443_),
    .A1(\top1.memory1.mem1[195][0] ),
    .A2(net5938));
 sg13g2_nor2_1 _16083_ (.A(\top1.memory1.mem1[199][0] ),
    .B(net5936),
    .Y(_06444_));
 sg13g2_nor2_1 _16084_ (.A(\top1.memory1.mem1[196][0] ),
    .B(net6041),
    .Y(_06445_));
 sg13g2_nor2_1 _16085_ (.A(\top1.memory1.mem1[197][0] ),
    .B(net5974),
    .Y(_06446_));
 sg13g2_o21ai_1 _16086_ (.B1(net6130),
    .Y(_06447_),
    .A1(\top1.memory1.mem1[198][0] ),
    .A2(net5894));
 sg13g2_nor4_2 _16087_ (.A(_06444_),
    .B(_06445_),
    .C(_06446_),
    .Y(_06448_),
    .D(_06447_));
 sg13g2_nor2_1 _16088_ (.A(_03979_),
    .B(_06448_),
    .Y(_06449_));
 sg13g2_a221oi_1 _16089_ (.B2(_06449_),
    .C1(net6108),
    .B1(_06443_),
    .A1(_06421_),
    .Y(_06450_),
    .A2(_06438_));
 sg13g2_nor2_1 _16090_ (.A(\top1.memory1.mem2[84][0] ),
    .B(net6040),
    .Y(_06451_));
 sg13g2_nor2_1 _16091_ (.A(\top1.memory1.mem2[85][0] ),
    .B(net5974),
    .Y(_06452_));
 sg13g2_nor2_1 _16092_ (.A(\top1.memory1.mem2[86][0] ),
    .B(net5895),
    .Y(_06453_));
 sg13g2_o21ai_1 _16093_ (.B1(net6016),
    .Y(_06454_),
    .A1(\top1.memory1.mem2[87][0] ),
    .A2(net5933));
 sg13g2_nor4_2 _16094_ (.A(_06451_),
    .B(_06452_),
    .C(_06453_),
    .Y(_06455_),
    .D(_06454_));
 sg13g2_mux4_1 _16095_ (.S0(net6201),
    .A0(\top1.memory1.mem2[92][0] ),
    .A1(\top1.memory1.mem2[93][0] ),
    .A2(\top1.memory1.mem2[94][0] ),
    .A3(\top1.memory1.mem2[95][0] ),
    .S1(net6137),
    .X(_06456_));
 sg13g2_a22oi_1 _16096_ (.Y(_06457_),
    .B1(net5904),
    .B2(\top1.memory1.mem2[82][0] ),
    .A2(net6048),
    .A1(\top1.memory1.mem2[80][0] ));
 sg13g2_a22oi_1 _16097_ (.Y(_06458_),
    .B1(net5945),
    .B2(\top1.memory1.mem2[83][0] ),
    .A2(net5984),
    .A1(\top1.memory1.mem2[81][0] ));
 sg13g2_a21oi_1 _16098_ (.A1(_06457_),
    .A2(_06458_),
    .Y(_06459_),
    .B1(net5868));
 sg13g2_a22oi_1 _16099_ (.Y(_06460_),
    .B1(net5903),
    .B2(\top1.memory1.mem2[90][0] ),
    .A2(net5944),
    .A1(\top1.memory1.mem2[91][0] ));
 sg13g2_a22oi_1 _16100_ (.Y(_06461_),
    .B1(net5983),
    .B2(\top1.memory1.mem2[89][0] ),
    .A2(net6048),
    .A1(\top1.memory1.mem2[88][0] ));
 sg13g2_a21oi_1 _16101_ (.A1(_06460_),
    .A2(_06461_),
    .Y(_06462_),
    .B1(net6075));
 sg13g2_a21o_1 _16102_ (.A2(_06456_),
    .A1(net5852),
    .B1(net6104),
    .X(_06463_));
 sg13g2_nor4_2 _16103_ (.A(_06455_),
    .B(_06459_),
    .C(_06462_),
    .Y(_06464_),
    .D(_06463_));
 sg13g2_mux4_1 _16104_ (.S0(net6198),
    .A0(\top1.memory1.mem2[76][0] ),
    .A1(\top1.memory1.mem2[77][0] ),
    .A2(\top1.memory1.mem2[78][0] ),
    .A3(\top1.memory1.mem2[79][0] ),
    .S1(net6134),
    .X(_06465_));
 sg13g2_and2_1 _16105_ (.A(net5850),
    .B(_06465_),
    .X(_06466_));
 sg13g2_mux4_1 _16106_ (.S0(net6198),
    .A0(\top1.memory1.mem2[64][0] ),
    .A1(\top1.memory1.mem2[65][0] ),
    .A2(\top1.memory1.mem2[66][0] ),
    .A3(\top1.memory1.mem2[67][0] ),
    .S1(net6134),
    .X(_06467_));
 sg13g2_mux4_1 _16107_ (.S0(net6200),
    .A0(\top1.memory1.mem2[72][0] ),
    .A1(\top1.memory1.mem2[73][0] ),
    .A2(\top1.memory1.mem2[74][0] ),
    .A3(\top1.memory1.mem2[75][0] ),
    .S1(net6136),
    .X(_06468_));
 sg13g2_a221oi_1 _16108_ (.B2(_03882_),
    .C1(net6011),
    .B1(net5983),
    .A1(_03881_),
    .Y(_06469_),
    .A2(net6048));
 sg13g2_a22oi_1 _16109_ (.Y(_06470_),
    .B1(net5903),
    .B2(_03883_),
    .A2(net5944),
    .A1(_03884_));
 sg13g2_a21oi_1 _16110_ (.A1(net6083),
    .A2(_06468_),
    .Y(_06471_),
    .B1(net6120));
 sg13g2_a221oi_1 _16111_ (.B2(_06470_),
    .C1(_06466_),
    .B1(_06469_),
    .A1(net5873),
    .Y(_06472_),
    .A2(_06467_));
 sg13g2_a21o_2 _16112_ (.A2(_06472_),
    .A1(_06471_),
    .B1(net6117),
    .X(_06473_));
 sg13g2_mux4_1 _16113_ (.S0(net6242),
    .A0(\top1.memory1.mem2[112][0] ),
    .A1(\top1.memory1.mem2[113][0] ),
    .A2(\top1.memory1.mem2[114][0] ),
    .A3(\top1.memory1.mem2[115][0] ),
    .S1(net6177),
    .X(_06474_));
 sg13g2_mux4_1 _16114_ (.S0(net6237),
    .A0(\top1.memory1.mem2[124][0] ),
    .A1(\top1.memory1.mem2[125][0] ),
    .A2(\top1.memory1.mem2[126][0] ),
    .A3(\top1.memory1.mem2[127][0] ),
    .S1(net6172),
    .X(_06475_));
 sg13g2_mux4_1 _16115_ (.S0(net6241),
    .A0(\top1.memory1.mem2[116][0] ),
    .A1(\top1.memory1.mem2[117][0] ),
    .A2(\top1.memory1.mem2[118][0] ),
    .A3(\top1.memory1.mem2[119][0] ),
    .S1(net6176),
    .X(_06476_));
 sg13g2_mux4_1 _16116_ (.S0(net6238),
    .A0(\top1.memory1.mem2[120][0] ),
    .A1(\top1.memory1.mem2[121][0] ),
    .A2(\top1.memory1.mem2[122][0] ),
    .A3(\top1.memory1.mem2[123][0] ),
    .S1(net6173),
    .X(_06477_));
 sg13g2_a22oi_1 _16117_ (.Y(_06478_),
    .B1(_06476_),
    .B2(net6030),
    .A2(_06474_),
    .A1(net5884));
 sg13g2_a22oi_1 _16118_ (.Y(_06479_),
    .B1(_06477_),
    .B2(net6094),
    .A2(_06475_),
    .A1(net5859));
 sg13g2_a21oi_2 _16119_ (.B1(net5838),
    .Y(_06480_),
    .A2(_06479_),
    .A1(_06478_));
 sg13g2_mux4_1 _16120_ (.S0(net6227),
    .A0(\top1.memory1.mem2[96][0] ),
    .A1(\top1.memory1.mem2[97][0] ),
    .A2(\top1.memory1.mem2[98][0] ),
    .A3(\top1.memory1.mem2[99][0] ),
    .S1(net6162),
    .X(_06481_));
 sg13g2_mux4_1 _16121_ (.S0(net6236),
    .A0(\top1.memory1.mem2[108][0] ),
    .A1(\top1.memory1.mem2[109][0] ),
    .A2(\top1.memory1.mem2[110][0] ),
    .A3(\top1.memory1.mem2[111][0] ),
    .S1(net6171),
    .X(_06482_));
 sg13g2_mux4_1 _16122_ (.S0(net6223),
    .A0(\top1.memory1.mem2[100][0] ),
    .A1(\top1.memory1.mem2[101][0] ),
    .A2(\top1.memory1.mem2[102][0] ),
    .A3(\top1.memory1.mem2[103][0] ),
    .S1(net6158),
    .X(_06483_));
 sg13g2_mux4_1 _16123_ (.S0(net6236),
    .A0(\top1.memory1.mem2[104][0] ),
    .A1(\top1.memory1.mem2[105][0] ),
    .A2(\top1.memory1.mem2[106][0] ),
    .A3(\top1.memory1.mem2[107][0] ),
    .S1(net6171),
    .X(_06484_));
 sg13g2_a22oi_1 _16124_ (.Y(_06485_),
    .B1(_06483_),
    .B2(net6025),
    .A2(_06481_),
    .A1(net5880));
 sg13g2_a22oi_1 _16125_ (.Y(_06486_),
    .B1(_06484_),
    .B2(net6093),
    .A2(_06482_),
    .A1(net5859));
 sg13g2_a21oi_1 _16126_ (.A1(_06485_),
    .A2(_06486_),
    .Y(_06487_),
    .B1(net5832));
 sg13g2_nor3_2 _16127_ (.A(_03830_),
    .B(_06480_),
    .C(_06487_),
    .Y(_06488_));
 sg13g2_o21ai_1 _16128_ (.B1(_06488_),
    .Y(_06489_),
    .A1(_06464_),
    .A2(_06473_));
 sg13g2_mux4_1 _16129_ (.S0(net6230),
    .A0(\top1.memory1.mem2[24][0] ),
    .A1(\top1.memory1.mem2[25][0] ),
    .A2(\top1.memory1.mem2[26][0] ),
    .A3(\top1.memory1.mem2[27][0] ),
    .S1(net6165),
    .X(_06490_));
 sg13g2_a21o_1 _16130_ (.A2(_06490_),
    .A1(net6091),
    .B1(net6106),
    .X(_06491_));
 sg13g2_a22oi_1 _16131_ (.Y(_06492_),
    .B1(net5923),
    .B2(\top1.memory1.mem2[18][0] ),
    .A2(net6066),
    .A1(\top1.memory1.mem2[16][0] ));
 sg13g2_a22oi_1 _16132_ (.Y(_06493_),
    .B1(net5963),
    .B2(\top1.memory1.mem2[19][0] ),
    .A2(net6004),
    .A1(\top1.memory1.mem2[17][0] ));
 sg13g2_a21oi_1 _16133_ (.A1(_06492_),
    .A2(_06493_),
    .Y(_06494_),
    .B1(net5870));
 sg13g2_a22oi_1 _16134_ (.Y(_06495_),
    .B1(net5921),
    .B2(\top1.memory1.mem2[30][0] ),
    .A2(net5961),
    .A1(\top1.memory1.mem2[31][0] ));
 sg13g2_a22oi_1 _16135_ (.Y(_06496_),
    .B1(net6002),
    .B2(\top1.memory1.mem2[29][0] ),
    .A2(net6068),
    .A1(\top1.memory1.mem2[28][0] ));
 sg13g2_a21oi_1 _16136_ (.A1(_06495_),
    .A2(_06496_),
    .Y(_06497_),
    .B1(net5848));
 sg13g2_o21ai_1 _16137_ (.B1(net6027),
    .Y(_06498_),
    .A1(\top1.memory1.mem2[20][0] ),
    .A2(net6045));
 sg13g2_nor2_1 _16138_ (.A(\top1.memory1.mem2[22][0] ),
    .B(net5899),
    .Y(_06499_));
 sg13g2_nor2_1 _16139_ (.A(\top1.memory1.mem2[23][0] ),
    .B(net5940),
    .Y(_06500_));
 sg13g2_nor2_1 _16140_ (.A(\top1.memory1.mem2[21][0] ),
    .B(net5979),
    .Y(_06501_));
 sg13g2_nor4_1 _16141_ (.A(_06498_),
    .B(_06499_),
    .C(_06500_),
    .D(_06501_),
    .Y(_06502_));
 sg13g2_nor4_1 _16142_ (.A(_06491_),
    .B(_06494_),
    .C(_06497_),
    .D(_06502_),
    .Y(_06503_));
 sg13g2_mux4_1 _16143_ (.S0(net6215),
    .A0(\top1.memory1.mem2[12][0] ),
    .A1(\top1.memory1.mem2[13][0] ),
    .A2(\top1.memory1.mem2[14][0] ),
    .A3(\top1.memory1.mem2[15][0] ),
    .S1(net6150),
    .X(_06504_));
 sg13g2_mux4_1 _16144_ (.S0(net6216),
    .A0(\top1.memory1.mem2[0][0] ),
    .A1(\top1.memory1.mem2[1][0] ),
    .A2(\top1.memory1.mem2[2][0] ),
    .A3(\top1.memory1.mem2[3][0] ),
    .S1(net6151),
    .X(_06505_));
 sg13g2_mux4_1 _16145_ (.S0(net6216),
    .A0(\top1.memory1.mem2[8][0] ),
    .A1(\top1.memory1.mem2[9][0] ),
    .A2(\top1.memory1.mem2[10][0] ),
    .A3(\top1.memory1.mem2[11][0] ),
    .S1(net6151),
    .X(_06506_));
 sg13g2_o21ai_1 _16146_ (.B1(net6023),
    .Y(_06507_),
    .A1(\top1.memory1.mem2[4][0] ),
    .A2(_03984_));
 sg13g2_nor2_1 _16147_ (.A(\top1.memory1.mem2[5][0] ),
    .B(net5980),
    .Y(_06508_));
 sg13g2_nor2_1 _16148_ (.A(\top1.memory1.mem2[7][0] ),
    .B(net5940),
    .Y(_06509_));
 sg13g2_nor2_1 _16149_ (.A(\top1.memory1.mem2[6][0] ),
    .B(net5900),
    .Y(_06510_));
 sg13g2_nor4_1 _16150_ (.A(_06507_),
    .B(_06508_),
    .C(_06509_),
    .D(_06510_),
    .Y(_06511_));
 sg13g2_a21oi_1 _16151_ (.A1(net5879),
    .A2(_06505_),
    .Y(_06512_),
    .B1(net6125));
 sg13g2_a22oi_1 _16152_ (.Y(_06513_),
    .B1(_06506_),
    .B2(net6088),
    .A2(_06504_),
    .A1(net5854));
 sg13g2_nand2_1 _16153_ (.Y(_06514_),
    .A(_06512_),
    .B(_06513_));
 sg13g2_o21ai_1 _16154_ (.B1(net6103),
    .Y(_06515_),
    .A1(_06511_),
    .A2(_06514_));
 sg13g2_mux4_1 _16155_ (.S0(net6251),
    .A0(\top1.memory1.mem2[44][0] ),
    .A1(\top1.memory1.mem2[45][0] ),
    .A2(\top1.memory1.mem2[46][0] ),
    .A3(\top1.memory1.mem2[47][0] ),
    .S1(net6186),
    .X(_06516_));
 sg13g2_mux4_1 _16156_ (.S0(net6235),
    .A0(\top1.memory1.mem2[36][0] ),
    .A1(\top1.memory1.mem2[37][0] ),
    .A2(\top1.memory1.mem2[38][0] ),
    .A3(\top1.memory1.mem2[39][0] ),
    .S1(net6170),
    .X(_06517_));
 sg13g2_mux4_1 _16157_ (.S0(net6251),
    .A0(\top1.memory1.mem2[40][0] ),
    .A1(\top1.memory1.mem2[41][0] ),
    .A2(\top1.memory1.mem2[42][0] ),
    .A3(\top1.memory1.mem2[43][0] ),
    .S1(net6186),
    .X(_06518_));
 sg13g2_mux4_1 _16158_ (.S0(net6233),
    .A0(\top1.memory1.mem2[32][0] ),
    .A1(\top1.memory1.mem2[33][0] ),
    .A2(\top1.memory1.mem2[34][0] ),
    .A3(\top1.memory1.mem2[35][0] ),
    .S1(net6168),
    .X(_06519_));
 sg13g2_a22oi_1 _16159_ (.Y(_06520_),
    .B1(_06518_),
    .B2(net6099),
    .A2(_06516_),
    .A1(net5862));
 sg13g2_a22oi_1 _16160_ (.Y(_06521_),
    .B1(_06519_),
    .B2(net5883),
    .A2(_06517_),
    .A1(net6028));
 sg13g2_a21oi_1 _16161_ (.A1(_06520_),
    .A2(_06521_),
    .Y(_06522_),
    .B1(net5834));
 sg13g2_mux4_1 _16162_ (.S0(net6252),
    .A0(\top1.memory1.mem2[60][0] ),
    .A1(\top1.memory1.mem2[61][0] ),
    .A2(\top1.memory1.mem2[62][0] ),
    .A3(\top1.memory1.mem2[63][0] ),
    .S1(net6187),
    .X(_06523_));
 sg13g2_mux4_1 _16163_ (.S0(net6253),
    .A0(\top1.memory1.mem2[48][0] ),
    .A1(\top1.memory1.mem2[49][0] ),
    .A2(\top1.memory1.mem2[50][0] ),
    .A3(\top1.memory1.mem2[51][0] ),
    .S1(net6188),
    .X(_06524_));
 sg13g2_mux4_1 _16164_ (.S0(net6250),
    .A0(\top1.memory1.mem2[56][0] ),
    .A1(\top1.memory1.mem2[57][0] ),
    .A2(\top1.memory1.mem2[58][0] ),
    .A3(\top1.memory1.mem2[59][0] ),
    .S1(net6185),
    .X(_06525_));
 sg13g2_mux4_1 _16165_ (.S0(net6252),
    .A0(\top1.memory1.mem2[52][0] ),
    .A1(\top1.memory1.mem2[53][0] ),
    .A2(\top1.memory1.mem2[54][0] ),
    .A3(\top1.memory1.mem2[55][0] ),
    .S1(net6187),
    .X(_06526_));
 sg13g2_a22oi_1 _16166_ (.Y(_06527_),
    .B1(_06525_),
    .B2(net6098),
    .A2(_06523_),
    .A1(net5862));
 sg13g2_a22oi_1 _16167_ (.Y(_06528_),
    .B1(_06526_),
    .B2(net6034),
    .A2(_06524_),
    .A1(net5888));
 sg13g2_a21oi_2 _16168_ (.B1(net5840),
    .Y(_06529_),
    .A2(_06528_),
    .A1(_06527_));
 sg13g2_nor3_2 _16169_ (.A(net6116),
    .B(_06522_),
    .C(_06529_),
    .Y(_06530_));
 sg13g2_o21ai_1 _16170_ (.B1(_06530_),
    .Y(_06531_),
    .A1(_06503_),
    .A2(_06515_));
 sg13g2_a21o_1 _16171_ (.A2(_06531_),
    .A1(_06489_),
    .B1(net6111),
    .X(_06532_));
 sg13g2_nor2_1 _16172_ (.A(\top1.memory1.mem2[151][0] ),
    .B(net5936),
    .Y(_06533_));
 sg13g2_nor2_1 _16173_ (.A(\top1.memory1.mem2[149][0] ),
    .B(net5975),
    .Y(_06534_));
 sg13g2_nor2_1 _16174_ (.A(\top1.memory1.mem2[148][0] ),
    .B(net6041),
    .Y(_06535_));
 sg13g2_o21ai_1 _16175_ (.B1(net6020),
    .Y(_06536_),
    .A1(\top1.memory1.mem2[150][0] ),
    .A2(net5896));
 sg13g2_nor4_1 _16176_ (.A(_06533_),
    .B(_06534_),
    .C(_06535_),
    .D(_06536_),
    .Y(_06537_));
 sg13g2_nor2_1 _16177_ (.A(net6105),
    .B(_06537_),
    .Y(_06538_));
 sg13g2_a22oi_1 _16178_ (.Y(_06539_),
    .B1(net5914),
    .B2(\top1.memory1.mem2[154][0] ),
    .A2(net5997),
    .A1(\top1.memory1.mem2[153][0] ));
 sg13g2_a22oi_1 _16179_ (.Y(_06540_),
    .B1(net5956),
    .B2(\top1.memory1.mem2[155][0] ),
    .A2(net6059),
    .A1(\top1.memory1.mem2[152][0] ));
 sg13g2_a21oi_2 _16180_ (.B1(net6078),
    .Y(_06541_),
    .A2(_06540_),
    .A1(_06539_));
 sg13g2_a22oi_1 _16181_ (.Y(_06542_),
    .B1(net5909),
    .B2(\top1.memory1.mem2[146][0] ),
    .A2(net5948),
    .A1(\top1.memory1.mem2[147][0] ));
 sg13g2_a22oi_1 _16182_ (.Y(_06543_),
    .B1(net5990),
    .B2(\top1.memory1.mem2[145][0] ),
    .A2(net6054),
    .A1(\top1.memory1.mem2[144][0] ));
 sg13g2_a21oi_1 _16183_ (.A1(_06542_),
    .A2(_06543_),
    .Y(_06544_),
    .B1(net5867));
 sg13g2_a22oi_1 _16184_ (.Y(_06545_),
    .B1(net5994),
    .B2(\top1.memory1.mem2[157][0] ),
    .A2(net6058),
    .A1(\top1.memory1.mem2[156][0] ));
 sg13g2_a22oi_1 _16185_ (.Y(_06546_),
    .B1(net5913),
    .B2(\top1.memory1.mem2[158][0] ),
    .A2(net5953),
    .A1(\top1.memory1.mem2[159][0] ));
 sg13g2_a21oi_1 _16186_ (.A1(_06545_),
    .A2(_06546_),
    .Y(_06547_),
    .B1(net5846));
 sg13g2_nor3_2 _16187_ (.A(_06541_),
    .B(_06544_),
    .C(_06547_),
    .Y(_06548_));
 sg13g2_a22oi_1 _16188_ (.Y(_06549_),
    .B1(net5905),
    .B2(\top1.memory1.mem2[142][0] ),
    .A2(net5946),
    .A1(\top1.memory1.mem2[143][0] ));
 sg13g2_a22oi_1 _16189_ (.Y(_06550_),
    .B1(net5986),
    .B2(\top1.memory1.mem2[141][0] ),
    .A2(net6050),
    .A1(\top1.memory1.mem2[140][0] ));
 sg13g2_a21oi_1 _16190_ (.A1(_06549_),
    .A2(_06550_),
    .Y(_06551_),
    .B1(net5842));
 sg13g2_a22oi_1 _16191_ (.Y(_06552_),
    .B1(net5909),
    .B2(\top1.memory1.mem2[138][0] ),
    .A2(net6054),
    .A1(\top1.memory1.mem2[136][0] ));
 sg13g2_a22oi_1 _16192_ (.Y(_06553_),
    .B1(net5948),
    .B2(\top1.memory1.mem2[139][0] ),
    .A2(net5990),
    .A1(\top1.memory1.mem2[137][0] ));
 sg13g2_a21o_2 _16193_ (.A2(_06553_),
    .A1(_06552_),
    .B1(net6076),
    .X(_06554_));
 sg13g2_a22oi_1 _16194_ (.Y(_06555_),
    .B1(net5905),
    .B2(\top1.memory1.mem2[130][0] ),
    .A2(net5946),
    .A1(\top1.memory1.mem2[131][0] ));
 sg13g2_a22oi_1 _16195_ (.Y(_06556_),
    .B1(net5986),
    .B2(\top1.memory1.mem2[129][0] ),
    .A2(net6050),
    .A1(\top1.memory1.mem2[128][0] ));
 sg13g2_a21oi_2 _16196_ (.B1(net5867),
    .Y(_06557_),
    .A2(_06556_),
    .A1(_06555_));
 sg13g2_nor2_1 _16197_ (.A(\top1.memory1.mem2[132][0] ),
    .B(net6038),
    .Y(_06558_));
 sg13g2_nor2_1 _16198_ (.A(\top1.memory1.mem2[133][0] ),
    .B(net5972),
    .Y(_06559_));
 sg13g2_nor2_1 _16199_ (.A(\top1.memory1.mem2[135][0] ),
    .B(net5930),
    .Y(_06560_));
 sg13g2_o21ai_1 _16200_ (.B1(net6019),
    .Y(_06561_),
    .A1(\top1.memory1.mem2[134][0] ),
    .A2(net5892));
 sg13g2_nor4_1 _16201_ (.A(_06558_),
    .B(_06559_),
    .C(_06560_),
    .D(_06561_),
    .Y(_06562_));
 sg13g2_nor4_2 _16202_ (.A(net6122),
    .B(_06551_),
    .C(_06557_),
    .Y(_06563_),
    .D(_06562_));
 sg13g2_a221oi_1 _16203_ (.B2(_06563_),
    .C1(net6117),
    .B1(_06554_),
    .A1(_06538_),
    .Y(_06564_),
    .A2(_06548_));
 sg13g2_a22oi_1 _16204_ (.Y(_06565_),
    .B1(net5928),
    .B2(\top1.memory1.mem2[178][0] ),
    .A2(net5968),
    .A1(\top1.memory1.mem2[179][0] ));
 sg13g2_a22oi_1 _16205_ (.Y(_06566_),
    .B1(net6007),
    .B2(\top1.memory1.mem2[177][0] ),
    .A2(net6071),
    .A1(\top1.memory1.mem2[176][0] ));
 sg13g2_a21oi_1 _16206_ (.A1(_06565_),
    .A2(_06566_),
    .Y(_06567_),
    .B1(net5871));
 sg13g2_a22oi_1 _16207_ (.Y(_06568_),
    .B1(net5928),
    .B2(\top1.memory1.mem2[190][0] ),
    .A2(net5968),
    .A1(\top1.memory1.mem2[191][0] ));
 sg13g2_a22oi_1 _16208_ (.Y(_06569_),
    .B1(net6007),
    .B2(\top1.memory1.mem2[189][0] ),
    .A2(net6071),
    .A1(\top1.memory1.mem2[188][0] ));
 sg13g2_a21oi_1 _16209_ (.A1(_06568_),
    .A2(_06569_),
    .Y(_06570_),
    .B1(net5849));
 sg13g2_a22oi_1 _16210_ (.Y(_06571_),
    .B1(net5927),
    .B2(\top1.memory1.mem2[182][0] ),
    .A2(net5967),
    .A1(\top1.memory1.mem2[183][0] ));
 sg13g2_a22oi_1 _16211_ (.Y(_06572_),
    .B1(net6005),
    .B2(\top1.memory1.mem2[181][0] ),
    .A2(net6067),
    .A1(\top1.memory1.mem2[180][0] ));
 sg13g2_a21oi_1 _16212_ (.A1(_06571_),
    .A2(_06572_),
    .Y(_06573_),
    .B1(net6014));
 sg13g2_a22oi_1 _16213_ (.Y(_06574_),
    .B1(net5923),
    .B2(\top1.memory1.mem2[186][0] ),
    .A2(net5963),
    .A1(\top1.memory1.mem2[187][0] ));
 sg13g2_a22oi_1 _16214_ (.Y(_06575_),
    .B1(net6004),
    .B2(\top1.memory1.mem2[185][0] ),
    .A2(net6066),
    .A1(\top1.memory1.mem2[184][0] ));
 sg13g2_a21oi_1 _16215_ (.A1(_06574_),
    .A2(_06575_),
    .Y(_06576_),
    .B1(net6080));
 sg13g2_or4_2 _16216_ (.A(_06567_),
    .B(_06570_),
    .C(_06573_),
    .D(_06576_),
    .X(_06577_));
 sg13g2_a22oi_1 _16217_ (.Y(_06578_),
    .B1(net5922),
    .B2(\top1.memory1.mem2[170][0] ),
    .A2(net5962),
    .A1(\top1.memory1.mem2[171][0] ));
 sg13g2_a22oi_1 _16218_ (.Y(_06579_),
    .B1(net5999),
    .B2(\top1.memory1.mem2[169][0] ),
    .A2(net6063),
    .A1(\top1.memory1.mem2[168][0] ));
 sg13g2_a21oi_1 _16219_ (.A1(_06578_),
    .A2(_06579_),
    .Y(_06580_),
    .B1(net6080));
 sg13g2_a22oi_1 _16220_ (.Y(_06581_),
    .B1(net5922),
    .B2(\top1.memory1.mem2[166][0] ),
    .A2(net5962),
    .A1(\top1.memory1.mem2[167][0] ));
 sg13g2_a22oi_1 _16221_ (.Y(_06582_),
    .B1(net6003),
    .B2(\top1.memory1.mem2[165][0] ),
    .A2(net6065),
    .A1(\top1.memory1.mem2[164][0] ));
 sg13g2_a21oi_2 _16222_ (.B1(net6013),
    .Y(_06583_),
    .A2(_06582_),
    .A1(_06581_));
 sg13g2_a22oi_1 _16223_ (.Y(_06584_),
    .B1(net5918),
    .B2(\top1.memory1.mem2[174][0] ),
    .A2(net5958),
    .A1(\top1.memory1.mem2[175][0] ));
 sg13g2_a22oi_1 _16224_ (.Y(_06585_),
    .B1(net5999),
    .B2(\top1.memory1.mem2[173][0] ),
    .A2(net6064),
    .A1(\top1.memory1.mem2[172][0] ));
 sg13g2_a21oi_2 _16225_ (.B1(net5847),
    .Y(_06586_),
    .A2(_06585_),
    .A1(_06584_));
 sg13g2_a22oi_1 _16226_ (.Y(_06587_),
    .B1(net5922),
    .B2(\top1.memory1.mem2[162][0] ),
    .A2(net5962),
    .A1(\top1.memory1.mem2[163][0] ));
 sg13g2_a22oi_1 _16227_ (.Y(_06588_),
    .B1(net5995),
    .B2(\top1.memory1.mem2[161][0] ),
    .A2(net6060),
    .A1(\top1.memory1.mem2[160][0] ));
 sg13g2_a21oi_1 _16228_ (.A1(_06587_),
    .A2(_06588_),
    .Y(_06589_),
    .B1(net5871));
 sg13g2_nor4_2 _16229_ (.A(_06580_),
    .B(_06583_),
    .C(_06586_),
    .Y(_06590_),
    .D(_06589_));
 sg13g2_nand2b_1 _16230_ (.Y(_06591_),
    .B(_05443_),
    .A_N(_06590_));
 sg13g2_a21oi_1 _16231_ (.A1(_05452_),
    .A2(_06577_),
    .Y(_06592_),
    .B1(net5831));
 sg13g2_nand3b_1 _16232_ (.B(_06591_),
    .C(_06592_),
    .Y(_06593_),
    .A_N(_06564_));
 sg13g2_nand2_1 _16233_ (.Y(_06594_),
    .A(\top1.memory1.mem2[199][0] ),
    .B(net5955));
 sg13g2_a22oi_1 _16234_ (.Y(_06595_),
    .B1(net5995),
    .B2(\top1.memory1.mem2[197][0] ),
    .A2(net6060),
    .A1(\top1.memory1.mem2[196][0] ));
 sg13g2_nand3_1 _16235_ (.B(_06594_),
    .C(_06595_),
    .A(net6132),
    .Y(_06596_));
 sg13g2_a21oi_1 _16236_ (.A1(\top1.memory1.mem2[198][0] ),
    .A2(net5915),
    .Y(_06597_),
    .B1(_06596_));
 sg13g2_a22oi_1 _16237_ (.Y(_06598_),
    .B1(net5995),
    .B2(\top1.memory1.mem2[193][0] ),
    .A2(net6060),
    .A1(\top1.memory1.mem2[192][0] ));
 sg13g2_a221oi_1 _16238_ (.B2(\top1.memory1.mem2[194][0] ),
    .C1(net6129),
    .B1(net5914),
    .A1(\top1.memory1.mem2[195][0] ),
    .Y(_06599_),
    .A2(net5954));
 sg13g2_and2_1 _16239_ (.A(_06598_),
    .B(_06599_),
    .X(_06600_));
 sg13g2_o21ai_1 _16240_ (.B1(_03978_),
    .Y(_06601_),
    .A1(_06597_),
    .A2(_06600_));
 sg13g2_nand4_1 _16241_ (.B(_06532_),
    .C(_06593_),
    .A(net6109),
    .Y(_06602_),
    .D(_06601_));
 sg13g2_a21oi_1 _16242_ (.A1(_06394_),
    .A2(_06450_),
    .Y(_06603_),
    .B1(net6101));
 sg13g2_a22oi_1 _16243_ (.Y(_01054_),
    .B1(_06602_),
    .B2(_06603_),
    .A2(_03851_),
    .A1(net6101));
 sg13g2_mux4_1 _16244_ (.S0(net6230),
    .A0(\top1.memory1.mem2[24][1] ),
    .A1(\top1.memory1.mem2[25][1] ),
    .A2(\top1.memory1.mem2[26][1] ),
    .A3(\top1.memory1.mem2[27][1] ),
    .S1(net6165),
    .X(_06604_));
 sg13g2_a21o_1 _16245_ (.A2(_06604_),
    .A1(net6091),
    .B1(net6106),
    .X(_06605_));
 sg13g2_a22oi_1 _16246_ (.Y(_06606_),
    .B1(net5963),
    .B2(\top1.memory1.mem2[19][1] ),
    .A2(net6066),
    .A1(\top1.memory1.mem2[16][1] ));
 sg13g2_a22oi_1 _16247_ (.Y(_06607_),
    .B1(net5923),
    .B2(\top1.memory1.mem2[18][1] ),
    .A2(net6004),
    .A1(\top1.memory1.mem2[17][1] ));
 sg13g2_a21oi_1 _16248_ (.A1(_06606_),
    .A2(_06607_),
    .Y(_06608_),
    .B1(net5870));
 sg13g2_o21ai_1 _16249_ (.B1(net6027),
    .Y(_06609_),
    .A1(\top1.memory1.mem2[21][1] ),
    .A2(net5979));
 sg13g2_nor2_1 _16250_ (.A(\top1.memory1.mem2[23][1] ),
    .B(net5940),
    .Y(_06610_));
 sg13g2_nor2_1 _16251_ (.A(\top1.memory1.mem2[20][1] ),
    .B(net6045),
    .Y(_06611_));
 sg13g2_nor2_1 _16252_ (.A(\top1.memory1.mem2[22][1] ),
    .B(net5899),
    .Y(_06612_));
 sg13g2_nor4_1 _16253_ (.A(_06609_),
    .B(_06610_),
    .C(_06611_),
    .D(_06612_),
    .Y(_06613_));
 sg13g2_a22oi_1 _16254_ (.Y(_06614_),
    .B1(net5921),
    .B2(\top1.memory1.mem2[30][1] ),
    .A2(net5961),
    .A1(\top1.memory1.mem2[31][1] ));
 sg13g2_a22oi_1 _16255_ (.Y(_06615_),
    .B1(net6002),
    .B2(\top1.memory1.mem2[29][1] ),
    .A2(net6065),
    .A1(\top1.memory1.mem2[28][1] ));
 sg13g2_a21oi_2 _16256_ (.B1(net5847),
    .Y(_06616_),
    .A2(_06615_),
    .A1(_06614_));
 sg13g2_nor4_2 _16257_ (.A(_06605_),
    .B(_06608_),
    .C(_06613_),
    .Y(_06617_),
    .D(_06616_));
 sg13g2_a21oi_1 _16258_ (.A1(_03898_),
    .A2(net5921),
    .Y(_06618_),
    .B1(net6013));
 sg13g2_nor3_1 _16259_ (.A(net6217),
    .B(net6152),
    .C(\top1.memory1.mem2[4][1] ),
    .Y(_06619_));
 sg13g2_a221oi_1 _16260_ (.B2(_03899_),
    .C1(_06619_),
    .B1(net5961),
    .A1(_03897_),
    .Y(_06620_),
    .A2(net6002));
 sg13g2_mux4_1 _16261_ (.S0(net6218),
    .A0(\top1.memory1.mem2[0][1] ),
    .A1(\top1.memory1.mem2[1][1] ),
    .A2(\top1.memory1.mem2[2][1] ),
    .A3(\top1.memory1.mem2[3][1] ),
    .S1(net6153),
    .X(_06621_));
 sg13g2_mux4_1 _16262_ (.S0(net6218),
    .A0(\top1.memory1.mem2[8][1] ),
    .A1(\top1.memory1.mem2[9][1] ),
    .A2(\top1.memory1.mem2[10][1] ),
    .A3(\top1.memory1.mem2[11][1] ),
    .S1(net6153),
    .X(_06622_));
 sg13g2_mux4_1 _16263_ (.S0(net6215),
    .A0(\top1.memory1.mem2[12][1] ),
    .A1(\top1.memory1.mem2[13][1] ),
    .A2(\top1.memory1.mem2[14][1] ),
    .A3(\top1.memory1.mem2[15][1] ),
    .S1(net6150),
    .X(_06623_));
 sg13g2_a22oi_1 _16264_ (.Y(_06624_),
    .B1(_06621_),
    .B2(net5879),
    .A2(_06620_),
    .A1(_06618_));
 sg13g2_a221oi_1 _16265_ (.B2(net5854),
    .C1(net6125),
    .B1(_06623_),
    .A1(net6087),
    .Y(_06625_),
    .A2(_06622_));
 sg13g2_a21o_1 _16266_ (.A2(_06625_),
    .A1(_06624_),
    .B1(net6119),
    .X(_06626_));
 sg13g2_mux4_1 _16267_ (.S0(net6253),
    .A0(\top1.memory1.mem2[48][1] ),
    .A1(\top1.memory1.mem2[49][1] ),
    .A2(\top1.memory1.mem2[50][1] ),
    .A3(\top1.memory1.mem2[51][1] ),
    .S1(net6188),
    .X(_06627_));
 sg13g2_mux4_1 _16268_ (.S0(net6250),
    .A0(\top1.memory1.mem2[56][1] ),
    .A1(\top1.memory1.mem2[57][1] ),
    .A2(\top1.memory1.mem2[58][1] ),
    .A3(\top1.memory1.mem2[59][1] ),
    .S1(net6185),
    .X(_06628_));
 sg13g2_mux4_1 _16269_ (.S0(net6251),
    .A0(\top1.memory1.mem2[52][1] ),
    .A1(\top1.memory1.mem2[53][1] ),
    .A2(\top1.memory1.mem2[54][1] ),
    .A3(\top1.memory1.mem2[55][1] ),
    .S1(net6186),
    .X(_06629_));
 sg13g2_mux4_1 _16270_ (.S0(net6252),
    .A0(\top1.memory1.mem2[60][1] ),
    .A1(\top1.memory1.mem2[61][1] ),
    .A2(\top1.memory1.mem2[62][1] ),
    .A3(\top1.memory1.mem2[63][1] ),
    .S1(net6187),
    .X(_06630_));
 sg13g2_a22oi_1 _16271_ (.Y(_06631_),
    .B1(_06629_),
    .B2(net6034),
    .A2(_06627_),
    .A1(net5888));
 sg13g2_a22oi_1 _16272_ (.Y(_06632_),
    .B1(_06630_),
    .B2(net5862),
    .A2(_06628_),
    .A1(net6098));
 sg13g2_a21oi_2 _16273_ (.B1(net5840),
    .Y(_06633_),
    .A2(_06632_),
    .A1(_06631_));
 sg13g2_mux4_1 _16274_ (.S0(net6235),
    .A0(\top1.memory1.mem2[36][1] ),
    .A1(\top1.memory1.mem2[37][1] ),
    .A2(\top1.memory1.mem2[38][1] ),
    .A3(\top1.memory1.mem2[39][1] ),
    .S1(net6170),
    .X(_06634_));
 sg13g2_mux4_1 _16275_ (.S0(net6251),
    .A0(\top1.memory1.mem2[40][1] ),
    .A1(\top1.memory1.mem2[41][1] ),
    .A2(\top1.memory1.mem2[42][1] ),
    .A3(\top1.memory1.mem2[43][1] ),
    .S1(net6186),
    .X(_06635_));
 sg13g2_mux4_1 _16276_ (.S0(net6233),
    .A0(\top1.memory1.mem2[32][1] ),
    .A1(\top1.memory1.mem2[33][1] ),
    .A2(\top1.memory1.mem2[34][1] ),
    .A3(\top1.memory1.mem2[35][1] ),
    .S1(net6168),
    .X(_06636_));
 sg13g2_mux4_1 _16277_ (.S0(net6251),
    .A0(\top1.memory1.mem2[44][1] ),
    .A1(\top1.memory1.mem2[45][1] ),
    .A2(\top1.memory1.mem2[46][1] ),
    .A3(\top1.memory1.mem2[47][1] ),
    .S1(net6186),
    .X(_06637_));
 sg13g2_a22oi_1 _16278_ (.Y(_06638_),
    .B1(_06636_),
    .B2(net5883),
    .A2(_06634_),
    .A1(net6027));
 sg13g2_a22oi_1 _16279_ (.Y(_06639_),
    .B1(_06637_),
    .B2(net5862),
    .A2(_06635_),
    .A1(net6099));
 sg13g2_a21oi_1 _16280_ (.A1(_06638_),
    .A2(_06639_),
    .Y(_06640_),
    .B1(net5834));
 sg13g2_nor3_2 _16281_ (.A(net6116),
    .B(_06633_),
    .C(_06640_),
    .Y(_06641_));
 sg13g2_o21ai_1 _16282_ (.B1(_06641_),
    .Y(_06642_),
    .A1(_06617_),
    .A2(_06626_));
 sg13g2_mux4_1 _16283_ (.S0(net6201),
    .A0(\top1.memory1.mem2[80][1] ),
    .A1(\top1.memory1.mem2[81][1] ),
    .A2(\top1.memory1.mem2[82][1] ),
    .A3(\top1.memory1.mem2[83][1] ),
    .S1(net6137),
    .X(_06643_));
 sg13g2_nor2_1 _16284_ (.A(\top1.memory1.mem2[85][1] ),
    .B(net5974),
    .Y(_06644_));
 sg13g2_nor2_1 _16285_ (.A(\top1.memory1.mem2[84][1] ),
    .B(net6040),
    .Y(_06645_));
 sg13g2_nor2_1 _16286_ (.A(\top1.memory1.mem2[87][1] ),
    .B(net5933),
    .Y(_06646_));
 sg13g2_o21ai_1 _16287_ (.B1(net6021),
    .Y(_06647_),
    .A1(\top1.memory1.mem2[86][1] ),
    .A2(net5895));
 sg13g2_nor4_1 _16288_ (.A(_06644_),
    .B(_06645_),
    .C(_06646_),
    .D(_06647_),
    .Y(_06648_));
 sg13g2_mux4_1 _16289_ (.S0(net6202),
    .A0(\top1.memory1.mem2[92][1] ),
    .A1(\top1.memory1.mem2[93][1] ),
    .A2(\top1.memory1.mem2[94][1] ),
    .A3(\top1.memory1.mem2[95][1] ),
    .S1(net6137),
    .X(_06649_));
 sg13g2_nand2_1 _16290_ (.Y(_06650_),
    .A(net5852),
    .B(_06649_));
 sg13g2_mux4_1 _16291_ (.S0(net6201),
    .A0(\top1.memory1.mem2[88][1] ),
    .A1(\top1.memory1.mem2[89][1] ),
    .A2(\top1.memory1.mem2[90][1] ),
    .A3(\top1.memory1.mem2[91][1] ),
    .S1(net6137),
    .X(_06651_));
 sg13g2_a22oi_1 _16292_ (.Y(_06652_),
    .B1(_06651_),
    .B2(net6083),
    .A2(_06643_),
    .A1(net5874));
 sg13g2_nand2_1 _16293_ (.Y(_06653_),
    .A(_06650_),
    .B(_06652_));
 sg13g2_o21ai_1 _16294_ (.B1(_05516_),
    .Y(_06654_),
    .A1(_06648_),
    .A2(_06653_));
 sg13g2_mux4_1 _16295_ (.S0(net6197),
    .A0(\top1.memory1.mem2[76][1] ),
    .A1(\top1.memory1.mem2[77][1] ),
    .A2(\top1.memory1.mem2[78][1] ),
    .A3(\top1.memory1.mem2[79][1] ),
    .S1(net6133),
    .X(_06655_));
 sg13g2_nor3_1 _16296_ (.A(net6200),
    .B(net6136),
    .C(\top1.memory1.mem2[68][1] ),
    .Y(_06656_));
 sg13g2_a21oi_1 _16297_ (.A1(_03901_),
    .A2(net5903),
    .Y(_06657_),
    .B1(net6011));
 sg13g2_a221oi_1 _16298_ (.B2(_03902_),
    .C1(_06656_),
    .B1(net5944),
    .A1(_03900_),
    .Y(_06658_),
    .A2(net5983));
 sg13g2_mux4_1 _16299_ (.S0(net6197),
    .A0(\top1.memory1.mem2[64][1] ),
    .A1(\top1.memory1.mem2[65][1] ),
    .A2(\top1.memory1.mem2[66][1] ),
    .A3(\top1.memory1.mem2[67][1] ),
    .S1(net6133),
    .X(_06659_));
 sg13g2_mux4_1 _16300_ (.S0(net6200),
    .A0(\top1.memory1.mem2[72][1] ),
    .A1(\top1.memory1.mem2[73][1] ),
    .A2(\top1.memory1.mem2[74][1] ),
    .A3(\top1.memory1.mem2[75][1] ),
    .S1(net6136),
    .X(_06660_));
 sg13g2_a22oi_1 _16301_ (.Y(_06661_),
    .B1(_06659_),
    .B2(net5873),
    .A2(_06655_),
    .A1(net5850));
 sg13g2_a22oi_1 _16302_ (.Y(_06662_),
    .B1(_06660_),
    .B2(net6086),
    .A2(_06658_),
    .A1(_06657_));
 sg13g2_a21o_2 _16303_ (.A2(_06662_),
    .A1(_06661_),
    .B1(_03977_),
    .X(_06663_));
 sg13g2_mux4_1 _16304_ (.S0(net6246),
    .A0(\top1.memory1.mem2[112][1] ),
    .A1(\top1.memory1.mem2[113][1] ),
    .A2(\top1.memory1.mem2[114][1] ),
    .A3(\top1.memory1.mem2[115][1] ),
    .S1(net6181),
    .X(_06664_));
 sg13g2_mux4_1 _16305_ (.S0(net6237),
    .A0(\top1.memory1.mem2[116][1] ),
    .A1(\top1.memory1.mem2[117][1] ),
    .A2(\top1.memory1.mem2[118][1] ),
    .A3(\top1.memory1.mem2[119][1] ),
    .S1(net6172),
    .X(_06665_));
 sg13g2_a22oi_1 _16306_ (.Y(_06666_),
    .B1(_06665_),
    .B2(net6030),
    .A2(_06664_),
    .A1(net5884));
 sg13g2_mux4_1 _16307_ (.S0(net6237),
    .A0(\top1.memory1.mem2[124][1] ),
    .A1(\top1.memory1.mem2[125][1] ),
    .A2(\top1.memory1.mem2[126][1] ),
    .A3(\top1.memory1.mem2[127][1] ),
    .S1(net6172),
    .X(_06667_));
 sg13g2_mux4_1 _16308_ (.S0(net6240),
    .A0(\top1.memory1.mem2[120][1] ),
    .A1(\top1.memory1.mem2[121][1] ),
    .A2(\top1.memory1.mem2[122][1] ),
    .A3(\top1.memory1.mem2[123][1] ),
    .S1(net6175),
    .X(_06668_));
 sg13g2_a22oi_1 _16309_ (.Y(_06669_),
    .B1(_06668_),
    .B2(net6094),
    .A2(_06667_),
    .A1(net5859));
 sg13g2_a21oi_2 _16310_ (.B1(net5838),
    .Y(_06670_),
    .A2(_06669_),
    .A1(_06666_));
 sg13g2_mux4_1 _16311_ (.S0(net6238),
    .A0(\top1.memory1.mem2[104][1] ),
    .A1(\top1.memory1.mem2[105][1] ),
    .A2(\top1.memory1.mem2[106][1] ),
    .A3(\top1.memory1.mem2[107][1] ),
    .S1(net6173),
    .X(_06671_));
 sg13g2_a22oi_1 _16312_ (.Y(_06672_),
    .B1(net5926),
    .B2(\top1.memory1.mem2[102][1] ),
    .A2(net6070),
    .A1(\top1.memory1.mem2[100][1] ));
 sg13g2_a22oi_1 _16313_ (.Y(_06673_),
    .B1(net5966),
    .B2(\top1.memory1.mem2[103][1] ),
    .A2(net6006),
    .A1(\top1.memory1.mem2[101][1] ));
 sg13g2_a21oi_1 _16314_ (.A1(_06672_),
    .A2(_06673_),
    .Y(_06674_),
    .B1(net6014));
 sg13g2_mux4_1 _16315_ (.S0(net6236),
    .A0(\top1.memory1.mem2[108][1] ),
    .A1(\top1.memory1.mem2[109][1] ),
    .A2(\top1.memory1.mem2[110][1] ),
    .A3(\top1.memory1.mem2[111][1] ),
    .S1(net6171),
    .X(_06675_));
 sg13g2_mux4_1 _16316_ (.S0(net6227),
    .A0(\top1.memory1.mem2[96][1] ),
    .A1(\top1.memory1.mem2[97][1] ),
    .A2(\top1.memory1.mem2[98][1] ),
    .A3(\top1.memory1.mem2[99][1] ),
    .S1(net6162),
    .X(_06676_));
 sg13g2_nand2_1 _16317_ (.Y(_06677_),
    .A(net5880),
    .B(_06676_));
 sg13g2_a22oi_1 _16318_ (.Y(_06678_),
    .B1(_06675_),
    .B2(net5859),
    .A2(_06671_),
    .A1(net6093));
 sg13g2_nand2_1 _16319_ (.Y(_06679_),
    .A(_06677_),
    .B(_06678_));
 sg13g2_o21ai_1 _16320_ (.B1(_05443_),
    .Y(_06680_),
    .A1(_06674_),
    .A2(_06679_));
 sg13g2_nor2_2 _16321_ (.A(_03830_),
    .B(_06670_),
    .Y(_06681_));
 sg13g2_nand4_1 _16322_ (.B(_06663_),
    .C(_06680_),
    .A(_06654_),
    .Y(_06682_),
    .D(_06681_));
 sg13g2_a21oi_1 _16323_ (.A1(_06642_),
    .A2(_06682_),
    .Y(_06683_),
    .B1(net6111));
 sg13g2_a22oi_1 _16324_ (.Y(_06684_),
    .B1(net5913),
    .B2(\top1.memory1.mem2[154][1] ),
    .A2(net6059),
    .A1(\top1.memory1.mem2[152][1] ));
 sg13g2_a22oi_1 _16325_ (.Y(_06685_),
    .B1(net5953),
    .B2(\top1.memory1.mem2[155][1] ),
    .A2(net5997),
    .A1(\top1.memory1.mem2[153][1] ));
 sg13g2_a21oi_2 _16326_ (.B1(net6078),
    .Y(_06686_),
    .A2(_06685_),
    .A1(_06684_));
 sg13g2_nor2_1 _16327_ (.A(\top1.memory1.mem2[149][1] ),
    .B(net5975),
    .Y(_06687_));
 sg13g2_nor2_1 _16328_ (.A(\top1.memory1.mem2[151][1] ),
    .B(net5935),
    .Y(_06688_));
 sg13g2_nor2_1 _16329_ (.A(\top1.memory1.mem2[150][1] ),
    .B(net5896),
    .Y(_06689_));
 sg13g2_o21ai_1 _16330_ (.B1(net6020),
    .Y(_06690_),
    .A1(\top1.memory1.mem2[148][1] ),
    .A2(net6041));
 sg13g2_nor4_1 _16331_ (.A(_06687_),
    .B(_06688_),
    .C(_06689_),
    .D(_06690_),
    .Y(_06691_));
 sg13g2_a22oi_1 _16332_ (.Y(_06692_),
    .B1(net5948),
    .B2(\top1.memory1.mem2[159][1] ),
    .A2(net5989),
    .A1(\top1.memory1.mem2[157][1] ));
 sg13g2_a22oi_1 _16333_ (.Y(_06693_),
    .B1(net5908),
    .B2(\top1.memory1.mem2[158][1] ),
    .A2(net6053),
    .A1(\top1.memory1.mem2[156][1] ));
 sg13g2_nand2_1 _16334_ (.Y(_06694_),
    .A(_06692_),
    .B(_06693_));
 sg13g2_a22oi_1 _16335_ (.Y(_06695_),
    .B1(net5948),
    .B2(\top1.memory1.mem2[147][1] ),
    .A2(net6053),
    .A1(\top1.memory1.mem2[144][1] ));
 sg13g2_a22oi_1 _16336_ (.Y(_06696_),
    .B1(net5908),
    .B2(\top1.memory1.mem2[146][1] ),
    .A2(net5989),
    .A1(\top1.memory1.mem2[145][1] ));
 sg13g2_a21oi_1 _16337_ (.A1(_06695_),
    .A2(_06696_),
    .Y(_06697_),
    .B1(net5868));
 sg13g2_a21oi_1 _16338_ (.A1(net5851),
    .A2(_06694_),
    .Y(_06698_),
    .B1(net6105));
 sg13g2_nor3_1 _16339_ (.A(_06686_),
    .B(_06691_),
    .C(_06697_),
    .Y(_06699_));
 sg13g2_a22oi_1 _16340_ (.Y(_06700_),
    .B1(net5905),
    .B2(\top1.memory1.mem2[142][1] ),
    .A2(net5986),
    .A1(\top1.memory1.mem2[141][1] ));
 sg13g2_a22oi_1 _16341_ (.Y(_06701_),
    .B1(net5946),
    .B2(\top1.memory1.mem2[143][1] ),
    .A2(net6050),
    .A1(\top1.memory1.mem2[140][1] ));
 sg13g2_a21oi_1 _16342_ (.A1(_06700_),
    .A2(_06701_),
    .Y(_06702_),
    .B1(net5842));
 sg13g2_a22oi_1 _16343_ (.Y(_06703_),
    .B1(net5906),
    .B2(\top1.memory1.mem2[138][1] ),
    .A2(net5948),
    .A1(\top1.memory1.mem2[139][1] ));
 sg13g2_a22oi_1 _16344_ (.Y(_06704_),
    .B1(net5987),
    .B2(\top1.memory1.mem2[137][1] ),
    .A2(net6051),
    .A1(\top1.memory1.mem2[136][1] ));
 sg13g2_nand2_1 _16345_ (.Y(_06705_),
    .A(_06703_),
    .B(_06704_));
 sg13g2_a22oi_1 _16346_ (.Y(_06706_),
    .B1(net5905),
    .B2(\top1.memory1.mem2[130][1] ),
    .A2(net6050),
    .A1(\top1.memory1.mem2[128][1] ));
 sg13g2_a22oi_1 _16347_ (.Y(_06707_),
    .B1(net5946),
    .B2(\top1.memory1.mem2[131][1] ),
    .A2(net5986),
    .A1(\top1.memory1.mem2[129][1] ));
 sg13g2_a21oi_1 _16348_ (.A1(_06706_),
    .A2(_06707_),
    .Y(_06708_),
    .B1(net5867));
 sg13g2_nor2_1 _16349_ (.A(\top1.memory1.mem2[134][1] ),
    .B(net5891),
    .Y(_06709_));
 sg13g2_nor2_1 _16350_ (.A(\top1.memory1.mem2[132][1] ),
    .B(net6038),
    .Y(_06710_));
 sg13g2_nor2_1 _16351_ (.A(\top1.memory1.mem2[135][1] ),
    .B(net5931),
    .Y(_06711_));
 sg13g2_o21ai_1 _16352_ (.B1(net6019),
    .Y(_06712_),
    .A1(\top1.memory1.mem2[133][1] ),
    .A2(net5972));
 sg13g2_nor4_1 _16353_ (.A(_06709_),
    .B(_06710_),
    .C(_06711_),
    .D(_06712_),
    .Y(_06713_));
 sg13g2_a21oi_1 _16354_ (.A1(net6085),
    .A2(_06705_),
    .Y(_06714_),
    .B1(net6122));
 sg13g2_nor3_2 _16355_ (.A(_06702_),
    .B(_06708_),
    .C(_06713_),
    .Y(_06715_));
 sg13g2_a221oi_1 _16356_ (.B2(_06715_),
    .C1(net6119),
    .B1(_06714_),
    .A1(_06698_),
    .Y(_06716_),
    .A2(_06699_));
 sg13g2_a22oi_1 _16357_ (.Y(_06717_),
    .B1(net5927),
    .B2(\top1.memory1.mem2[190][1] ),
    .A2(net5967),
    .A1(\top1.memory1.mem2[191][1] ));
 sg13g2_a22oi_1 _16358_ (.Y(_06718_),
    .B1(net6007),
    .B2(\top1.memory1.mem2[189][1] ),
    .A2(net6071),
    .A1(\top1.memory1.mem2[188][1] ));
 sg13g2_a21oi_1 _16359_ (.A1(_06717_),
    .A2(_06718_),
    .Y(_06719_),
    .B1(net5848));
 sg13g2_a22oi_1 _16360_ (.Y(_06720_),
    .B1(net5923),
    .B2(\top1.memory1.mem2[186][1] ),
    .A2(net5963),
    .A1(\top1.memory1.mem2[187][1] ));
 sg13g2_a22oi_1 _16361_ (.Y(_06721_),
    .B1(net6004),
    .B2(\top1.memory1.mem2[185][1] ),
    .A2(net6066),
    .A1(\top1.memory1.mem2[184][1] ));
 sg13g2_a21oi_1 _16362_ (.A1(_06720_),
    .A2(_06721_),
    .Y(_06722_),
    .B1(net6080));
 sg13g2_a22oi_1 _16363_ (.Y(_06723_),
    .B1(net5927),
    .B2(\top1.memory1.mem2[182][1] ),
    .A2(net5967),
    .A1(\top1.memory1.mem2[183][1] ));
 sg13g2_a22oi_1 _16364_ (.Y(_06724_),
    .B1(net6005),
    .B2(\top1.memory1.mem2[181][1] ),
    .A2(net6067),
    .A1(\top1.memory1.mem2[180][1] ));
 sg13g2_a21oi_2 _16365_ (.B1(net6014),
    .Y(_06725_),
    .A2(_06724_),
    .A1(_06723_));
 sg13g2_a22oi_1 _16366_ (.Y(_06726_),
    .B1(net5927),
    .B2(\top1.memory1.mem2[178][1] ),
    .A2(net5967),
    .A1(\top1.memory1.mem2[179][1] ));
 sg13g2_a22oi_1 _16367_ (.Y(_06727_),
    .B1(net6007),
    .B2(\top1.memory1.mem2[177][1] ),
    .A2(net6071),
    .A1(\top1.memory1.mem2[176][1] ));
 sg13g2_a21oi_1 _16368_ (.A1(_06726_),
    .A2(_06727_),
    .Y(_06728_),
    .B1(net5871));
 sg13g2_nor4_2 _16369_ (.A(_06719_),
    .B(_06722_),
    .C(_06725_),
    .Y(_06729_),
    .D(_06728_));
 sg13g2_nor2_2 _16370_ (.A(net5837),
    .B(_06729_),
    .Y(_06730_));
 sg13g2_a22oi_1 _16371_ (.Y(_06731_),
    .B1(net5920),
    .B2(\top1.memory1.mem2[162][1] ),
    .A2(net5958),
    .A1(\top1.memory1.mem2[163][1] ));
 sg13g2_a22oi_1 _16372_ (.Y(_06732_),
    .B1(net5998),
    .B2(\top1.memory1.mem2[161][1] ),
    .A2(net6057),
    .A1(\top1.memory1.mem2[160][1] ));
 sg13g2_a21oi_1 _16373_ (.A1(_06731_),
    .A2(_06732_),
    .Y(_06733_),
    .B1(net5870));
 sg13g2_a22oi_1 _16374_ (.Y(_06734_),
    .B1(net5918),
    .B2(\top1.memory1.mem2[170][1] ),
    .A2(net5958),
    .A1(\top1.memory1.mem2[171][1] ));
 sg13g2_a22oi_1 _16375_ (.Y(_06735_),
    .B1(net5999),
    .B2(\top1.memory1.mem2[169][1] ),
    .A2(net6063),
    .A1(\top1.memory1.mem2[168][1] ));
 sg13g2_a21oi_1 _16376_ (.A1(_06734_),
    .A2(_06735_),
    .Y(_06736_),
    .B1(net6081));
 sg13g2_a22oi_1 _16377_ (.Y(_06737_),
    .B1(net5918),
    .B2(\top1.memory1.mem2[174][1] ),
    .A2(net5958),
    .A1(\top1.memory1.mem2[175][1] ));
 sg13g2_a22oi_1 _16378_ (.Y(_06738_),
    .B1(net5999),
    .B2(\top1.memory1.mem2[173][1] ),
    .A2(net6063),
    .A1(\top1.memory1.mem2[172][1] ));
 sg13g2_a21oi_2 _16379_ (.B1(net5847),
    .Y(_06739_),
    .A2(_06738_),
    .A1(_06737_));
 sg13g2_a22oi_1 _16380_ (.Y(_06740_),
    .B1(net5922),
    .B2(\top1.memory1.mem2[166][1] ),
    .A2(net5962),
    .A1(\top1.memory1.mem2[167][1] ));
 sg13g2_a22oi_1 _16381_ (.Y(_06741_),
    .B1(net6003),
    .B2(\top1.memory1.mem2[165][1] ),
    .A2(net6065),
    .A1(\top1.memory1.mem2[164][1] ));
 sg13g2_a21oi_2 _16382_ (.B1(net6012),
    .Y(_06742_),
    .A2(_06741_),
    .A1(_06740_));
 sg13g2_nor4_2 _16383_ (.A(_06733_),
    .B(_06736_),
    .C(_06739_),
    .Y(_06743_),
    .D(_06742_));
 sg13g2_o21ai_1 _16384_ (.B1(_05514_),
    .Y(_06744_),
    .A1(net5836),
    .A2(_06743_));
 sg13g2_nor3_1 _16385_ (.A(_06716_),
    .B(_06730_),
    .C(_06744_),
    .Y(_06745_));
 sg13g2_nor2_1 _16386_ (.A(\top1.memory1.mem2[193][1] ),
    .B(net5978),
    .Y(_06746_));
 sg13g2_nor2_1 _16387_ (.A(\top1.memory1.mem2[195][1] ),
    .B(net5939),
    .Y(_06747_));
 sg13g2_nor2_1 _16388_ (.A(\top1.memory1.mem2[192][1] ),
    .B(net6041),
    .Y(_06748_));
 sg13g2_nor3_1 _16389_ (.A(net6129),
    .B(_06747_),
    .C(_06748_),
    .Y(_06749_));
 sg13g2_o21ai_1 _16390_ (.B1(_06749_),
    .Y(_06750_),
    .A1(\top1.memory1.mem2[194][1] ),
    .A2(net5898));
 sg13g2_nor2_1 _16391_ (.A(\top1.memory1.mem2[199][1] ),
    .B(net5939),
    .Y(_06751_));
 sg13g2_nor2_1 _16392_ (.A(\top1.memory1.mem2[198][1] ),
    .B(net5898),
    .Y(_06752_));
 sg13g2_nor2_1 _16393_ (.A(\top1.memory1.mem2[196][1] ),
    .B(net6044),
    .Y(_06753_));
 sg13g2_o21ai_1 _16394_ (.B1(net6131),
    .Y(_06754_),
    .A1(\top1.memory1.mem2[197][1] ),
    .A2(net5978));
 sg13g2_nor4_1 _16395_ (.A(_06751_),
    .B(_06752_),
    .C(_06753_),
    .D(_06754_),
    .Y(_06755_));
 sg13g2_o21ai_1 _16396_ (.B1(_03978_),
    .Y(_06756_),
    .A1(_06746_),
    .A2(_06750_));
 sg13g2_o21ai_1 _16397_ (.B1(net6109),
    .Y(_06757_),
    .A1(_06755_),
    .A2(_06756_));
 sg13g2_or3_1 _16398_ (.A(_06683_),
    .B(_06745_),
    .C(_06757_),
    .X(_06758_));
 sg13g2_a22oi_1 _16399_ (.Y(_06759_),
    .B1(net5960),
    .B2(_03888_),
    .A2(net6001),
    .A1(_03886_));
 sg13g2_a221oi_1 _16400_ (.B2(_03887_),
    .C1(net6012),
    .B1(net5918),
    .A1(_03885_),
    .Y(_06760_),
    .A2(net6063));
 sg13g2_mux4_1 _16401_ (.S0(net6214),
    .A0(\top1.memory1.mem1[8][1] ),
    .A1(\top1.memory1.mem1[9][1] ),
    .A2(\top1.memory1.mem1[10][1] ),
    .A3(\top1.memory1.mem1[11][1] ),
    .S1(net6149),
    .X(_06761_));
 sg13g2_mux4_1 _16402_ (.S0(net6211),
    .A0(\top1.memory1.mem1[0][1] ),
    .A1(\top1.memory1.mem1[1][1] ),
    .A2(\top1.memory1.mem1[2][1] ),
    .A3(\top1.memory1.mem1[3][1] ),
    .S1(net6146),
    .X(_06762_));
 sg13g2_and2_1 _16403_ (.A(net5878),
    .B(_06762_),
    .X(_06763_));
 sg13g2_mux4_1 _16404_ (.S0(net6214),
    .A0(\top1.memory1.mem1[12][1] ),
    .A1(\top1.memory1.mem1[13][1] ),
    .A2(\top1.memory1.mem1[14][1] ),
    .A3(\top1.memory1.mem1[15][1] ),
    .S1(net6149),
    .X(_06764_));
 sg13g2_a21oi_1 _16405_ (.A1(net6090),
    .A2(_06761_),
    .Y(_06765_),
    .B1(net6124));
 sg13g2_a221oi_1 _16406_ (.B2(net5853),
    .C1(_06763_),
    .B1(_06764_),
    .A1(_06759_),
    .Y(_06766_),
    .A2(_06760_));
 sg13g2_mux4_1 _16407_ (.S0(net6229),
    .A0(\top1.memory1.mem1[16][1] ),
    .A1(\top1.memory1.mem1[17][1] ),
    .A2(\top1.memory1.mem1[18][1] ),
    .A3(\top1.memory1.mem1[19][1] ),
    .S1(net6164),
    .X(_06767_));
 sg13g2_mux4_1 _16408_ (.S0(net6232),
    .A0(\top1.memory1.mem1[24][1] ),
    .A1(\top1.memory1.mem1[25][1] ),
    .A2(\top1.memory1.mem1[26][1] ),
    .A3(\top1.memory1.mem1[27][1] ),
    .S1(net6167),
    .X(_06768_));
 sg13g2_a22oi_1 _16409_ (.Y(_06769_),
    .B1(net5960),
    .B2(_03892_),
    .A2(net6069),
    .A1(_03889_));
 sg13g2_a221oi_1 _16410_ (.B2(_03891_),
    .C1(net6012),
    .B1(net5920),
    .A1(_03890_),
    .Y(_06770_),
    .A2(net6000));
 sg13g2_mux4_1 _16411_ (.S0(net6222),
    .A0(\top1.memory1.mem1[28][1] ),
    .A1(\top1.memory1.mem1[29][1] ),
    .A2(\top1.memory1.mem1[30][1] ),
    .A3(\top1.memory1.mem1[31][1] ),
    .S1(net6157),
    .X(_06771_));
 sg13g2_a22oi_1 _16412_ (.Y(_06772_),
    .B1(_06768_),
    .B2(net6091),
    .A2(_06767_),
    .A1(net5882));
 sg13g2_a221oi_1 _16413_ (.B2(net5856),
    .C1(net6106),
    .B1(_06771_),
    .A1(_06769_),
    .Y(_06773_),
    .A2(_06770_));
 sg13g2_a221oi_1 _16414_ (.B2(_06773_),
    .C1(net6118),
    .B1(_06772_),
    .A1(_06765_),
    .Y(_06774_),
    .A2(_06766_));
 sg13g2_mux4_1 _16415_ (.S0(net6247),
    .A0(\top1.memory1.mem1[60][1] ),
    .A1(\top1.memory1.mem1[61][1] ),
    .A2(\top1.memory1.mem1[62][1] ),
    .A3(\top1.memory1.mem1[63][1] ),
    .S1(net6182),
    .X(_06775_));
 sg13g2_mux4_1 _16416_ (.S0(net6254),
    .A0(\top1.memory1.mem1[48][1] ),
    .A1(\top1.memory1.mem1[49][1] ),
    .A2(\top1.memory1.mem1[50][1] ),
    .A3(\top1.memory1.mem1[51][1] ),
    .S1(net6189),
    .X(_06776_));
 sg13g2_mux4_1 _16417_ (.S0(net6246),
    .A0(\top1.memory1.mem1[52][1] ),
    .A1(\top1.memory1.mem1[53][1] ),
    .A2(\top1.memory1.mem1[54][1] ),
    .A3(\top1.memory1.mem1[55][1] ),
    .S1(net6181),
    .X(_06777_));
 sg13g2_mux4_1 _16418_ (.S0(net6254),
    .A0(\top1.memory1.mem1[56][1] ),
    .A1(\top1.memory1.mem1[57][1] ),
    .A2(\top1.memory1.mem1[58][1] ),
    .A3(\top1.memory1.mem1[59][1] ),
    .S1(net6189),
    .X(_06778_));
 sg13g2_a22oi_1 _16419_ (.Y(_06779_),
    .B1(_06777_),
    .B2(net6032),
    .A2(_06775_),
    .A1(net5861));
 sg13g2_a22oi_1 _16420_ (.Y(_06780_),
    .B1(_06778_),
    .B2(net6097),
    .A2(_06776_),
    .A1(net5886));
 sg13g2_a21oi_1 _16421_ (.A1(_06779_),
    .A2(_06780_),
    .Y(_06781_),
    .B1(net5840));
 sg13g2_mux4_1 _16422_ (.S0(net6254),
    .A0(\top1.memory1.mem1[44][1] ),
    .A1(\top1.memory1.mem1[45][1] ),
    .A2(\top1.memory1.mem1[46][1] ),
    .A3(\top1.memory1.mem1[47][1] ),
    .S1(net6189),
    .X(_06782_));
 sg13g2_mux4_1 _16423_ (.S0(net6258),
    .A0(\top1.memory1.mem1[36][1] ),
    .A1(\top1.memory1.mem1[37][1] ),
    .A2(\top1.memory1.mem1[38][1] ),
    .A3(\top1.memory1.mem1[39][1] ),
    .S1(net6193),
    .X(_06783_));
 sg13g2_mux4_1 _16424_ (.S0(net6256),
    .A0(\top1.memory1.mem1[40][1] ),
    .A1(\top1.memory1.mem1[41][1] ),
    .A2(\top1.memory1.mem1[42][1] ),
    .A3(\top1.memory1.mem1[43][1] ),
    .S1(net6191),
    .X(_06784_));
 sg13g2_mux4_1 _16425_ (.S0(net6257),
    .A0(\top1.memory1.mem1[32][1] ),
    .A1(\top1.memory1.mem1[33][1] ),
    .A2(\top1.memory1.mem1[34][1] ),
    .A3(\top1.memory1.mem1[35][1] ),
    .S1(net6192),
    .X(_06785_));
 sg13g2_a22oi_1 _16426_ (.Y(_06786_),
    .B1(_06784_),
    .B2(net6097),
    .A2(_06782_),
    .A1(net5864));
 sg13g2_a22oi_1 _16427_ (.Y(_06787_),
    .B1(_06785_),
    .B2(net5886),
    .A2(_06783_),
    .A1(net6033));
 sg13g2_a21oi_1 _16428_ (.A1(_06786_),
    .A2(_06787_),
    .Y(_06788_),
    .B1(net5835));
 sg13g2_o21ai_1 _16429_ (.B1(net6021),
    .Y(_06789_),
    .A1(\top1.memory1.mem1[85][1] ),
    .A2(net5973));
 sg13g2_nor2_1 _16430_ (.A(\top1.memory1.mem1[86][1] ),
    .B(net5894),
    .Y(_06790_));
 sg13g2_nor2_1 _16431_ (.A(\top1.memory1.mem1[87][1] ),
    .B(net5937),
    .Y(_06791_));
 sg13g2_nor2_1 _16432_ (.A(\top1.memory1.mem1[84][1] ),
    .B(net6039),
    .Y(_06792_));
 sg13g2_or4_1 _16433_ (.A(_06789_),
    .B(_06790_),
    .C(_06791_),
    .D(_06792_),
    .X(_06793_));
 sg13g2_a22oi_1 _16434_ (.Y(_06794_),
    .B1(net5911),
    .B2(\top1.memory1.mem1[82][1] ),
    .A2(net5951),
    .A1(\top1.memory1.mem1[83][1] ));
 sg13g2_a22oi_1 _16435_ (.Y(_06795_),
    .B1(net5993),
    .B2(\top1.memory1.mem1[81][1] ),
    .A2(net6056),
    .A1(\top1.memory1.mem1[80][1] ));
 sg13g2_a21o_1 _16436_ (.A2(_06795_),
    .A1(_06794_),
    .B1(net5869),
    .X(_06796_));
 sg13g2_mux4_1 _16437_ (.S0(net6209),
    .A0(\top1.memory1.mem1[92][1] ),
    .A1(\top1.memory1.mem1[93][1] ),
    .A2(\top1.memory1.mem1[94][1] ),
    .A3(\top1.memory1.mem1[95][1] ),
    .S1(net6144),
    .X(_06797_));
 sg13g2_mux4_1 _16438_ (.S0(net6209),
    .A0(\top1.memory1.mem1[88][1] ),
    .A1(\top1.memory1.mem1[89][1] ),
    .A2(\top1.memory1.mem1[90][1] ),
    .A3(\top1.memory1.mem1[91][1] ),
    .S1(net6144),
    .X(_06798_));
 sg13g2_mux4_1 _16439_ (.S0(net6233),
    .A0(\top1.memory1.mem1[96][1] ),
    .A1(\top1.memory1.mem1[97][1] ),
    .A2(\top1.memory1.mem1[98][1] ),
    .A3(\top1.memory1.mem1[99][1] ),
    .S1(net6168),
    .X(_06799_));
 sg13g2_mux4_1 _16440_ (.S0(net6239),
    .A0(\top1.memory1.mem1[108][1] ),
    .A1(\top1.memory1.mem1[109][1] ),
    .A2(\top1.memory1.mem1[110][1] ),
    .A3(\top1.memory1.mem1[111][1] ),
    .S1(net6174),
    .X(_06800_));
 sg13g2_mux4_1 _16441_ (.S0(net6249),
    .A0(\top1.memory1.mem1[104][1] ),
    .A1(\top1.memory1.mem1[105][1] ),
    .A2(\top1.memory1.mem1[106][1] ),
    .A3(\top1.memory1.mem1[107][1] ),
    .S1(net6184),
    .X(_06801_));
 sg13g2_mux4_1 _16442_ (.S0(net6239),
    .A0(\top1.memory1.mem1[100][1] ),
    .A1(\top1.memory1.mem1[101][1] ),
    .A2(\top1.memory1.mem1[102][1] ),
    .A3(\top1.memory1.mem1[103][1] ),
    .S1(net6174),
    .X(_06802_));
 sg13g2_a22oi_1 _16443_ (.Y(_06803_),
    .B1(_06801_),
    .B2(net6099),
    .A2(_06799_),
    .A1(net5888));
 sg13g2_a22oi_1 _16444_ (.Y(_06804_),
    .B1(_06802_),
    .B2(net6031),
    .A2(_06800_),
    .A1(net5860));
 sg13g2_a21oi_1 _16445_ (.A1(_06803_),
    .A2(_06804_),
    .Y(_06805_),
    .B1(net5832));
 sg13g2_mux4_1 _16446_ (.S0(net6243),
    .A0(\top1.memory1.mem1[116][1] ),
    .A1(\top1.memory1.mem1[117][1] ),
    .A2(\top1.memory1.mem1[118][1] ),
    .A3(\top1.memory1.mem1[119][1] ),
    .S1(net6178),
    .X(_06806_));
 sg13g2_mux4_1 _16447_ (.S0(net6241),
    .A0(\top1.memory1.mem1[124][1] ),
    .A1(\top1.memory1.mem1[125][1] ),
    .A2(\top1.memory1.mem1[126][1] ),
    .A3(\top1.memory1.mem1[127][1] ),
    .S1(net6176),
    .X(_06807_));
 sg13g2_mux4_1 _16448_ (.S0(net6243),
    .A0(\top1.memory1.mem1[112][1] ),
    .A1(\top1.memory1.mem1[113][1] ),
    .A2(\top1.memory1.mem1[114][1] ),
    .A3(\top1.memory1.mem1[115][1] ),
    .S1(net6178),
    .X(_06808_));
 sg13g2_mux4_1 _16449_ (.S0(net6241),
    .A0(\top1.memory1.mem1[120][1] ),
    .A1(\top1.memory1.mem1[121][1] ),
    .A2(\top1.memory1.mem1[122][1] ),
    .A3(\top1.memory1.mem1[123][1] ),
    .S1(net6176),
    .X(_06809_));
 sg13g2_a22oi_1 _16450_ (.Y(_06810_),
    .B1(_06808_),
    .B2(net5884),
    .A2(_06806_),
    .A1(net6030));
 sg13g2_a22oi_1 _16451_ (.Y(_06811_),
    .B1(_06809_),
    .B2(net6094),
    .A2(_06807_),
    .A1(net5861));
 sg13g2_a21oi_2 _16452_ (.B1(net5838),
    .Y(_06812_),
    .A2(_06811_),
    .A1(_06810_));
 sg13g2_mux4_1 _16453_ (.S0(net6198),
    .A0(\top1.memory1.mem1[64][1] ),
    .A1(\top1.memory1.mem1[65][1] ),
    .A2(\top1.memory1.mem1[66][1] ),
    .A3(\top1.memory1.mem1[67][1] ),
    .S1(net6134),
    .X(_06813_));
 sg13g2_mux4_1 _16454_ (.S0(net6199),
    .A0(\top1.memory1.mem1[76][1] ),
    .A1(\top1.memory1.mem1[77][1] ),
    .A2(\top1.memory1.mem1[78][1] ),
    .A3(\top1.memory1.mem1[79][1] ),
    .S1(net6135),
    .X(_06814_));
 sg13g2_a22oi_1 _16455_ (.Y(_06815_),
    .B1(net5984),
    .B2(_03894_),
    .A2(net6049),
    .A1(_03893_));
 sg13g2_a221oi_1 _16456_ (.B2(_03895_),
    .C1(net6011),
    .B1(net5904),
    .A1(_03896_),
    .Y(_06816_),
    .A2(net5945));
 sg13g2_mux4_1 _16457_ (.S0(net6199),
    .A0(\top1.memory1.mem1[72][1] ),
    .A1(\top1.memory1.mem1[73][1] ),
    .A2(\top1.memory1.mem1[74][1] ),
    .A3(\top1.memory1.mem1[75][1] ),
    .S1(net6135),
    .X(_06817_));
 sg13g2_or2_2 _16458_ (.X(_06818_),
    .B(_06788_),
    .A(_06781_));
 sg13g2_o21ai_1 _16459_ (.B1(net6102),
    .Y(_06819_),
    .A1(_06774_),
    .A2(_06818_));
 sg13g2_or2_2 _16460_ (.X(_06820_),
    .B(_06812_),
    .A(_06805_));
 sg13g2_a221oi_1 _16461_ (.B2(net6087),
    .C1(net6104),
    .B1(_06798_),
    .A1(net5853),
    .Y(_06821_),
    .A2(_06797_));
 sg13g2_nand3_1 _16462_ (.B(_06796_),
    .C(_06821_),
    .A(_06793_),
    .Y(_06822_));
 sg13g2_a22oi_1 _16463_ (.Y(_06823_),
    .B1(_06817_),
    .B2(net6083),
    .A2(_06814_),
    .A1(net5850));
 sg13g2_a221oi_1 _16464_ (.B2(_06816_),
    .C1(net6121),
    .B1(_06815_),
    .A1(net5873),
    .Y(_06824_),
    .A2(_06813_));
 sg13g2_a21oi_2 _16465_ (.B1(_05479_),
    .Y(_06825_),
    .A2(_06824_),
    .A1(_06823_));
 sg13g2_a221oi_1 _16466_ (.B2(_06825_),
    .C1(net6111),
    .B1(_06822_),
    .A1(net6113),
    .Y(_06826_),
    .A2(_06820_));
 sg13g2_nor2_1 _16467_ (.A(\top1.memory1.mem1[133][1] ),
    .B(net5976),
    .Y(_06827_));
 sg13g2_nor2_1 _16468_ (.A(\top1.memory1.mem1[135][1] ),
    .B(net5930),
    .Y(_06828_));
 sg13g2_nor2_1 _16469_ (.A(\top1.memory1.mem1[132][1] ),
    .B(net6042),
    .Y(_06829_));
 sg13g2_o21ai_1 _16470_ (.B1(net6019),
    .Y(_06830_),
    .A1(\top1.memory1.mem1[134][1] ),
    .A2(net5891));
 sg13g2_nor4_2 _16471_ (.A(_06827_),
    .B(_06828_),
    .C(_06829_),
    .Y(_06831_),
    .D(_06830_));
 sg13g2_mux4_1 _16472_ (.S0(net6203),
    .A0(\top1.memory1.mem1[140][1] ),
    .A1(\top1.memory1.mem1[141][1] ),
    .A2(\top1.memory1.mem1[142][1] ),
    .A3(\top1.memory1.mem1[143][1] ),
    .S1(net6139),
    .X(_06832_));
 sg13g2_a22oi_1 _16473_ (.Y(_06833_),
    .B1(net5902),
    .B2(\top1.memory1.mem1[130][1] ),
    .A2(net6047),
    .A1(\top1.memory1.mem1[128][1] ));
 sg13g2_a22oi_1 _16474_ (.Y(_06834_),
    .B1(net5943),
    .B2(\top1.memory1.mem1[131][1] ),
    .A2(net5982),
    .A1(\top1.memory1.mem1[129][1] ));
 sg13g2_a21oi_1 _16475_ (.A1(_06833_),
    .A2(_06834_),
    .Y(_06835_),
    .B1(net5867));
 sg13g2_a22oi_1 _16476_ (.Y(_06836_),
    .B1(net5907),
    .B2(\top1.memory1.mem1[138][1] ),
    .A2(net5947),
    .A1(\top1.memory1.mem1[139][1] ));
 sg13g2_a22oi_1 _16477_ (.Y(_06837_),
    .B1(net5988),
    .B2(\top1.memory1.mem1[137][1] ),
    .A2(net6052),
    .A1(\top1.memory1.mem1[136][1] ));
 sg13g2_a21oi_1 _16478_ (.A1(_06836_),
    .A2(_06837_),
    .Y(_06838_),
    .B1(net6076));
 sg13g2_a21o_1 _16479_ (.A2(_06832_),
    .A1(net5851),
    .B1(net6122),
    .X(_06839_));
 sg13g2_nor4_2 _16480_ (.A(_06831_),
    .B(_06835_),
    .C(_06838_),
    .Y(_06840_),
    .D(_06839_));
 sg13g2_a22oi_1 _16481_ (.Y(_06841_),
    .B1(net5909),
    .B2(\top1.memory1.mem1[158][1] ),
    .A2(net5948),
    .A1(\top1.memory1.mem1[159][1] ));
 sg13g2_a22oi_1 _16482_ (.Y(_06842_),
    .B1(net5990),
    .B2(\top1.memory1.mem1[157][1] ),
    .A2(net6054),
    .A1(\top1.memory1.mem1[156][1] ));
 sg13g2_a21oi_2 _16483_ (.B1(net5842),
    .Y(_06843_),
    .A2(_06842_),
    .A1(_06841_));
 sg13g2_mux4_1 _16484_ (.S0(net6205),
    .A0(\top1.memory1.mem1[144][1] ),
    .A1(\top1.memory1.mem1[145][1] ),
    .A2(\top1.memory1.mem1[146][1] ),
    .A3(\top1.memory1.mem1[147][1] ),
    .S1(net6141),
    .X(_06844_));
 sg13g2_a22oi_1 _16485_ (.Y(_06845_),
    .B1(net5908),
    .B2(\top1.memory1.mem1[154][1] ),
    .A2(net6053),
    .A1(\top1.memory1.mem1[152][1] ));
 sg13g2_a22oi_1 _16486_ (.Y(_06846_),
    .B1(net5949),
    .B2(\top1.memory1.mem1[155][1] ),
    .A2(net5989),
    .A1(\top1.memory1.mem1[153][1] ));
 sg13g2_a21oi_1 _16487_ (.A1(_06845_),
    .A2(_06846_),
    .Y(_06847_),
    .B1(net6076));
 sg13g2_nor2_1 _16488_ (.A(\top1.memory1.mem1[148][1] ),
    .B(net6037),
    .Y(_06848_));
 sg13g2_nor2_1 _16489_ (.A(\top1.memory1.mem1[150][1] ),
    .B(net5890),
    .Y(_06849_));
 sg13g2_nor2_1 _16490_ (.A(\top1.memory1.mem1[149][1] ),
    .B(net5971),
    .Y(_06850_));
 sg13g2_o21ai_1 _16491_ (.B1(net6020),
    .Y(_06851_),
    .A1(\top1.memory1.mem1[151][1] ),
    .A2(net5934));
 sg13g2_nor4_2 _16492_ (.A(_06848_),
    .B(_06849_),
    .C(_06850_),
    .Y(_06852_),
    .D(_06851_));
 sg13g2_a21o_1 _16493_ (.A2(_06844_),
    .A1(net5875),
    .B1(net6105),
    .X(_06853_));
 sg13g2_nor4_1 _16494_ (.A(_06843_),
    .B(_06847_),
    .C(_06852_),
    .D(_06853_),
    .Y(_06854_));
 sg13g2_or3_2 _16495_ (.A(net6119),
    .B(_06840_),
    .C(_06854_),
    .X(_06855_));
 sg13g2_mux4_1 _16496_ (.S0(net6220),
    .A0(\top1.memory1.mem1[168][1] ),
    .A1(\top1.memory1.mem1[169][1] ),
    .A2(\top1.memory1.mem1[170][1] ),
    .A3(\top1.memory1.mem1[171][1] ),
    .S1(net6155),
    .X(_06856_));
 sg13g2_mux4_1 _16497_ (.S0(net6221),
    .A0(\top1.memory1.mem1[164][1] ),
    .A1(\top1.memory1.mem1[165][1] ),
    .A2(\top1.memory1.mem1[166][1] ),
    .A3(\top1.memory1.mem1[167][1] ),
    .S1(net6156),
    .X(_06857_));
 sg13g2_mux4_1 _16498_ (.S0(net6212),
    .A0(\top1.memory1.mem1[160][1] ),
    .A1(\top1.memory1.mem1[161][1] ),
    .A2(\top1.memory1.mem1[162][1] ),
    .A3(\top1.memory1.mem1[163][1] ),
    .S1(net6147),
    .X(_06858_));
 sg13g2_mux4_1 _16499_ (.S0(net6220),
    .A0(\top1.memory1.mem1[172][1] ),
    .A1(\top1.memory1.mem1[173][1] ),
    .A2(\top1.memory1.mem1[174][1] ),
    .A3(\top1.memory1.mem1[175][1] ),
    .S1(net6155),
    .X(_06859_));
 sg13g2_a22oi_1 _16500_ (.Y(_06860_),
    .B1(_06858_),
    .B2(net5881),
    .A2(_06856_),
    .A1(net6089));
 sg13g2_a22oi_1 _16501_ (.Y(_06861_),
    .B1(_06859_),
    .B2(net5856),
    .A2(_06857_),
    .A1(net6026));
 sg13g2_a21oi_2 _16502_ (.B1(net5836),
    .Y(_06862_),
    .A2(_06861_),
    .A1(_06860_));
 sg13g2_mux4_1 _16503_ (.S0(net6224),
    .A0(\top1.memory1.mem1[180][1] ),
    .A1(\top1.memory1.mem1[181][1] ),
    .A2(\top1.memory1.mem1[182][1] ),
    .A3(\top1.memory1.mem1[183][1] ),
    .S1(net6159),
    .X(_06863_));
 sg13g2_mux4_1 _16504_ (.S0(net6221),
    .A0(\top1.memory1.mem1[184][1] ),
    .A1(\top1.memory1.mem1[185][1] ),
    .A2(\top1.memory1.mem1[186][1] ),
    .A3(\top1.memory1.mem1[187][1] ),
    .S1(net6156),
    .X(_06864_));
 sg13g2_mux4_1 _16505_ (.S0(net6225),
    .A0(\top1.memory1.mem1[188][1] ),
    .A1(\top1.memory1.mem1[189][1] ),
    .A2(\top1.memory1.mem1[190][1] ),
    .A3(\top1.memory1.mem1[191][1] ),
    .S1(net6160),
    .X(_06865_));
 sg13g2_mux4_1 _16506_ (.S0(net6225),
    .A0(\top1.memory1.mem1[176][1] ),
    .A1(\top1.memory1.mem1[177][1] ),
    .A2(\top1.memory1.mem1[178][1] ),
    .A3(\top1.memory1.mem1[179][1] ),
    .S1(net6160),
    .X(_06866_));
 sg13g2_a22oi_1 _16507_ (.Y(_06867_),
    .B1(_06865_),
    .B2(net5857),
    .A2(_06863_),
    .A1(net6025));
 sg13g2_a22oi_1 _16508_ (.Y(_06868_),
    .B1(_06866_),
    .B2(net5881),
    .A2(_06864_),
    .A1(net6090));
 sg13g2_a21oi_2 _16509_ (.B1(net5837),
    .Y(_06869_),
    .A2(_06868_),
    .A1(_06867_));
 sg13g2_nor3_2 _16510_ (.A(net5831),
    .B(_06862_),
    .C(_06869_),
    .Y(_06870_));
 sg13g2_nor2_1 _16511_ (.A(\top1.memory1.mem1[193][1] ),
    .B(net5977),
    .Y(_06871_));
 sg13g2_or3_1 _16512_ (.A(net6210),
    .B(net6145),
    .C(\top1.memory1.mem1[192][1] ),
    .X(_06872_));
 sg13g2_o21ai_1 _16513_ (.B1(_06872_),
    .Y(_06873_),
    .A1(\top1.memory1.mem1[194][1] ),
    .A2(net5897));
 sg13g2_nor2_1 _16514_ (.A(\top1.memory1.mem1[195][1] ),
    .B(net5937),
    .Y(_06874_));
 sg13g2_nor4_1 _16515_ (.A(net6131),
    .B(_06871_),
    .C(_06873_),
    .D(_06874_),
    .Y(_06875_));
 sg13g2_o21ai_1 _16516_ (.B1(net6130),
    .Y(_06876_),
    .A1(\top1.memory1.mem1[198][1] ),
    .A2(net5894));
 sg13g2_nor2_1 _16517_ (.A(\top1.memory1.mem1[197][1] ),
    .B(net5973),
    .Y(_06877_));
 sg13g2_nor2_1 _16518_ (.A(\top1.memory1.mem1[196][1] ),
    .B(net6039),
    .Y(_06878_));
 sg13g2_nor2_1 _16519_ (.A(\top1.memory1.mem1[199][1] ),
    .B(net5937),
    .Y(_06879_));
 sg13g2_nor4_1 _16520_ (.A(_06876_),
    .B(_06877_),
    .C(_06878_),
    .D(_06879_),
    .Y(_06880_));
 sg13g2_nor3_1 _16521_ (.A(_03979_),
    .B(_06875_),
    .C(_06880_),
    .Y(_06881_));
 sg13g2_or2_1 _16522_ (.X(_06882_),
    .B(_06881_),
    .A(net6108));
 sg13g2_a221oi_1 _16523_ (.B2(_06870_),
    .C1(_06882_),
    .B1(_06855_),
    .A1(_06819_),
    .Y(_06883_),
    .A2(_06826_));
 sg13g2_nor2_1 _16524_ (.A(net6101),
    .B(_06883_),
    .Y(_06884_));
 sg13g2_a22oi_1 _16525_ (.Y(_01055_),
    .B1(_06758_),
    .B2(_06884_),
    .A2(_03852_),
    .A1(net6101));
 sg13g2_a22oi_1 _16526_ (.Y(_06885_),
    .B1(net5911),
    .B2(_03911_),
    .A2(net6056),
    .A1(_03909_));
 sg13g2_a221oi_1 _16527_ (.B2(_03912_),
    .C1(net6077),
    .B1(net5951),
    .A1(_03910_),
    .Y(_06886_),
    .A2(net5992));
 sg13g2_mux4_1 _16528_ (.S0(net6209),
    .A0(\top1.memory1.mem1[84][2] ),
    .A1(\top1.memory1.mem1[85][2] ),
    .A2(\top1.memory1.mem1[86][2] ),
    .A3(\top1.memory1.mem1[87][2] ),
    .S1(net6144),
    .X(_06887_));
 sg13g2_mux4_1 _16529_ (.S0(net6209),
    .A0(\top1.memory1.mem1[92][2] ),
    .A1(\top1.memory1.mem1[93][2] ),
    .A2(\top1.memory1.mem1[94][2] ),
    .A3(\top1.memory1.mem1[95][2] ),
    .S1(net6144),
    .X(_06888_));
 sg13g2_mux4_1 _16530_ (.S0(net6209),
    .A0(\top1.memory1.mem1[80][2] ),
    .A1(\top1.memory1.mem1[81][2] ),
    .A2(\top1.memory1.mem1[82][2] ),
    .A3(\top1.memory1.mem1[83][2] ),
    .S1(net6144),
    .X(_06889_));
 sg13g2_and2_1 _16531_ (.A(net5877),
    .B(_06889_),
    .X(_06890_));
 sg13g2_a21oi_1 _16532_ (.A1(net5853),
    .A2(_06888_),
    .Y(_06891_),
    .B1(net6104));
 sg13g2_a221oi_1 _16533_ (.B2(net6021),
    .C1(_06890_),
    .B1(_06887_),
    .A1(_06885_),
    .Y(_06892_),
    .A2(_06886_));
 sg13g2_mux4_1 _16534_ (.S0(net6199),
    .A0(\top1.memory1.mem1[68][2] ),
    .A1(\top1.memory1.mem1[69][2] ),
    .A2(\top1.memory1.mem1[70][2] ),
    .A3(\top1.memory1.mem1[71][2] ),
    .S1(net6135),
    .X(_06893_));
 sg13g2_a21o_1 _16535_ (.A2(_06893_),
    .A1(net6018),
    .B1(net6121),
    .X(_06894_));
 sg13g2_a22oi_1 _16536_ (.Y(_06895_),
    .B1(net5942),
    .B2(\top1.memory1.mem1[67][2] ),
    .A2(net6046),
    .A1(\top1.memory1.mem1[64][2] ));
 sg13g2_a22oi_1 _16537_ (.Y(_06896_),
    .B1(net5901),
    .B2(\top1.memory1.mem1[66][2] ),
    .A2(net5981),
    .A1(\top1.memory1.mem1[65][2] ));
 sg13g2_a21oi_1 _16538_ (.A1(_06895_),
    .A2(_06896_),
    .Y(_06897_),
    .B1(net5868));
 sg13g2_o21ai_1 _16539_ (.B1(net6083),
    .Y(_06898_),
    .A1(\top1.memory1.mem1[72][2] ),
    .A2(net6036));
 sg13g2_nor2_1 _16540_ (.A(\top1.memory1.mem1[73][2] ),
    .B(net5970),
    .Y(_06899_));
 sg13g2_nor2_1 _16541_ (.A(\top1.memory1.mem1[74][2] ),
    .B(net5890),
    .Y(_06900_));
 sg13g2_nor2_1 _16542_ (.A(\top1.memory1.mem1[75][2] ),
    .B(net5932),
    .Y(_06901_));
 sg13g2_nor4_1 _16543_ (.A(_06898_),
    .B(_06899_),
    .C(_06900_),
    .D(_06901_),
    .Y(_06902_));
 sg13g2_a22oi_1 _16544_ (.Y(_06903_),
    .B1(net5901),
    .B2(\top1.memory1.mem1[78][2] ),
    .A2(net6046),
    .A1(\top1.memory1.mem1[76][2] ));
 sg13g2_a22oi_1 _16545_ (.Y(_06904_),
    .B1(net5942),
    .B2(\top1.memory1.mem1[79][2] ),
    .A2(net5981),
    .A1(\top1.memory1.mem1[77][2] ));
 sg13g2_a21oi_1 _16546_ (.A1(_06903_),
    .A2(_06904_),
    .Y(_06905_),
    .B1(net5844));
 sg13g2_or4_2 _16547_ (.A(_06894_),
    .B(_06897_),
    .C(_06902_),
    .D(_06905_),
    .X(_06906_));
 sg13g2_mux4_1 _16548_ (.S0(net6243),
    .A0(\top1.memory1.mem1[116][2] ),
    .A1(\top1.memory1.mem1[117][2] ),
    .A2(\top1.memory1.mem1[118][2] ),
    .A3(\top1.memory1.mem1[119][2] ),
    .S1(net6178),
    .X(_06907_));
 sg13g2_mux4_1 _16549_ (.S0(net6241),
    .A0(\top1.memory1.mem1[120][2] ),
    .A1(\top1.memory1.mem1[121][2] ),
    .A2(\top1.memory1.mem1[122][2] ),
    .A3(\top1.memory1.mem1[123][2] ),
    .S1(net6176),
    .X(_06908_));
 sg13g2_a22oi_1 _16550_ (.Y(_06909_),
    .B1(_06908_),
    .B2(net6094),
    .A2(_06907_),
    .A1(net6030));
 sg13g2_mux4_1 _16551_ (.S0(net6245),
    .A0(\top1.memory1.mem1[124][2] ),
    .A1(\top1.memory1.mem1[125][2] ),
    .A2(\top1.memory1.mem1[126][2] ),
    .A3(\top1.memory1.mem1[127][2] ),
    .S1(net6180),
    .X(_06910_));
 sg13g2_mux4_1 _16552_ (.S0(net6245),
    .A0(\top1.memory1.mem1[112][2] ),
    .A1(\top1.memory1.mem1[113][2] ),
    .A2(\top1.memory1.mem1[114][2] ),
    .A3(\top1.memory1.mem1[115][2] ),
    .S1(net6180),
    .X(_06911_));
 sg13g2_a22oi_1 _16553_ (.Y(_06912_),
    .B1(_06911_),
    .B2(net5884),
    .A2(_06910_),
    .A1(net5861));
 sg13g2_a21oi_2 _16554_ (.B1(net5838),
    .Y(_06913_),
    .A2(_06912_),
    .A1(_06909_));
 sg13g2_mux4_1 _16555_ (.S0(net6249),
    .A0(\top1.memory1.mem1[104][2] ),
    .A1(\top1.memory1.mem1[105][2] ),
    .A2(\top1.memory1.mem1[106][2] ),
    .A3(\top1.memory1.mem1[107][2] ),
    .S1(net6184),
    .X(_06914_));
 sg13g2_mux4_1 _16556_ (.S0(net6225),
    .A0(\top1.memory1.mem1[100][2] ),
    .A1(\top1.memory1.mem1[101][2] ),
    .A2(\top1.memory1.mem1[102][2] ),
    .A3(\top1.memory1.mem1[103][2] ),
    .S1(net6160),
    .X(_06915_));
 sg13g2_mux4_1 _16557_ (.S0(net6239),
    .A0(\top1.memory1.mem1[108][2] ),
    .A1(\top1.memory1.mem1[109][2] ),
    .A2(\top1.memory1.mem1[110][2] ),
    .A3(\top1.memory1.mem1[111][2] ),
    .S1(net6174),
    .X(_06916_));
 sg13g2_mux4_1 _16558_ (.S0(net6226),
    .A0(\top1.memory1.mem1[96][2] ),
    .A1(\top1.memory1.mem1[97][2] ),
    .A2(\top1.memory1.mem1[98][2] ),
    .A3(\top1.memory1.mem1[99][2] ),
    .S1(net6161),
    .X(_06917_));
 sg13g2_a22oi_1 _16559_ (.Y(_06918_),
    .B1(_06916_),
    .B2(net5860),
    .A2(_06914_),
    .A1(net6093));
 sg13g2_a22oi_1 _16560_ (.Y(_06919_),
    .B1(_06917_),
    .B2(net5880),
    .A2(_06915_),
    .A1(net6029));
 sg13g2_a21oi_1 _16561_ (.A1(_06918_),
    .A2(_06919_),
    .Y(_06920_),
    .B1(net5832));
 sg13g2_mux4_1 _16562_ (.S0(net6231),
    .A0(\top1.memory1.mem1[16][2] ),
    .A1(\top1.memory1.mem1[17][2] ),
    .A2(\top1.memory1.mem1[18][2] ),
    .A3(\top1.memory1.mem1[19][2] ),
    .S1(net6166),
    .X(_06921_));
 sg13g2_a22oi_1 _16563_ (.Y(_06922_),
    .B1(net6005),
    .B2(_03906_),
    .A2(net6067),
    .A1(_03905_));
 sg13g2_a221oi_1 _16564_ (.B2(_03907_),
    .C1(net6081),
    .B1(net5924),
    .A1(_03908_),
    .Y(_06923_),
    .A2(net5964));
 sg13g2_a22oi_1 _16565_ (.Y(_06924_),
    .B1(_06922_),
    .B2(_06923_),
    .A2(_06921_),
    .A1(net5882));
 sg13g2_mux4_1 _16566_ (.S0(net6222),
    .A0(\top1.memory1.mem1[20][2] ),
    .A1(\top1.memory1.mem1[21][2] ),
    .A2(\top1.memory1.mem1[22][2] ),
    .A3(\top1.memory1.mem1[23][2] ),
    .S1(net6157),
    .X(_06925_));
 sg13g2_mux4_1 _16567_ (.S0(net6222),
    .A0(\top1.memory1.mem1[28][2] ),
    .A1(\top1.memory1.mem1[29][2] ),
    .A2(\top1.memory1.mem1[30][2] ),
    .A3(\top1.memory1.mem1[31][2] ),
    .S1(net6157),
    .X(_06926_));
 sg13g2_a22oi_1 _16568_ (.Y(_06927_),
    .B1(_06926_),
    .B2(net5856),
    .A2(_06925_),
    .A1(net6026));
 sg13g2_a21oi_1 _16569_ (.A1(_06924_),
    .A2(_06927_),
    .Y(_06928_),
    .B1(_05517_));
 sg13g2_mux4_1 _16570_ (.S0(net6258),
    .A0(\top1.memory1.mem1[32][2] ),
    .A1(\top1.memory1.mem1[33][2] ),
    .A2(\top1.memory1.mem1[34][2] ),
    .A3(\top1.memory1.mem1[35][2] ),
    .S1(net6193),
    .X(_06929_));
 sg13g2_mux4_1 _16571_ (.S0(net6257),
    .A0(\top1.memory1.mem1[40][2] ),
    .A1(\top1.memory1.mem1[41][2] ),
    .A2(\top1.memory1.mem1[42][2] ),
    .A3(\top1.memory1.mem1[43][2] ),
    .S1(net6192),
    .X(_06930_));
 sg13g2_a22oi_1 _16572_ (.Y(_06931_),
    .B1(_06930_),
    .B2(net6097),
    .A2(_06929_),
    .A1(net5887));
 sg13g2_mux4_1 _16573_ (.S0(net6259),
    .A0(\top1.memory1.mem1[36][2] ),
    .A1(\top1.memory1.mem1[37][2] ),
    .A2(\top1.memory1.mem1[38][2] ),
    .A3(\top1.memory1.mem1[39][2] ),
    .S1(net6194),
    .X(_06932_));
 sg13g2_mux4_1 _16574_ (.S0(net6256),
    .A0(\top1.memory1.mem1[44][2] ),
    .A1(\top1.memory1.mem1[45][2] ),
    .A2(\top1.memory1.mem1[46][2] ),
    .A3(\top1.memory1.mem1[47][2] ),
    .S1(net6191),
    .X(_06933_));
 sg13g2_a22oi_1 _16575_ (.Y(_06934_),
    .B1(_06933_),
    .B2(net5864),
    .A2(_06932_),
    .A1(net6033));
 sg13g2_a21oi_2 _16576_ (.B1(net5835),
    .Y(_06935_),
    .A2(_06934_),
    .A1(_06931_));
 sg13g2_mux4_1 _16577_ (.S0(net6211),
    .A0(\top1.memory1.mem1[0][2] ),
    .A1(\top1.memory1.mem1[1][2] ),
    .A2(\top1.memory1.mem1[2][2] ),
    .A3(\top1.memory1.mem1[3][2] ),
    .S1(net6146),
    .X(_06936_));
 sg13g2_nand2_1 _16578_ (.Y(_06937_),
    .A(net6211),
    .B(\top1.memory1.mem1[11][2] ));
 sg13g2_nand2b_1 _16579_ (.Y(_06938_),
    .B(\top1.memory1.mem1[10][2] ),
    .A_N(net6211));
 sg13g2_nand3_1 _16580_ (.B(_06937_),
    .C(_06938_),
    .A(net6146),
    .Y(_06939_));
 sg13g2_a221oi_1 _16581_ (.B2(_03904_),
    .C1(net6077),
    .B1(net5992),
    .A1(_03903_),
    .Y(_06940_),
    .A2(net6057));
 sg13g2_a22oi_1 _16582_ (.Y(_06941_),
    .B1(_06939_),
    .B2(_06940_),
    .A2(_06936_),
    .A1(net5877));
 sg13g2_mux4_1 _16583_ (.S0(net6213),
    .A0(\top1.memory1.mem1[12][2] ),
    .A1(\top1.memory1.mem1[13][2] ),
    .A2(\top1.memory1.mem1[14][2] ),
    .A3(\top1.memory1.mem1[15][2] ),
    .S1(net6146),
    .X(_06942_));
 sg13g2_mux4_1 _16584_ (.S0(net6214),
    .A0(\top1.memory1.mem1[4][2] ),
    .A1(\top1.memory1.mem1[5][2] ),
    .A2(\top1.memory1.mem1[6][2] ),
    .A3(\top1.memory1.mem1[7][2] ),
    .S1(net6149),
    .X(_06943_));
 sg13g2_a22oi_1 _16585_ (.Y(_06944_),
    .B1(_06943_),
    .B2(net6021),
    .A2(_06942_),
    .A1(net5853));
 sg13g2_a21oi_2 _16586_ (.B1(_03977_),
    .Y(_06945_),
    .A2(_06944_),
    .A1(_06941_));
 sg13g2_mux4_1 _16587_ (.S0(net6245),
    .A0(\top1.memory1.mem1[60][2] ),
    .A1(\top1.memory1.mem1[61][2] ),
    .A2(\top1.memory1.mem1[62][2] ),
    .A3(\top1.memory1.mem1[63][2] ),
    .S1(net6180),
    .X(_06946_));
 sg13g2_a22oi_1 _16588_ (.Y(_06947_),
    .B1(net5929),
    .B2(\top1.memory1.mem1[58][2] ),
    .A2(net5969),
    .A1(\top1.memory1.mem1[59][2] ));
 sg13g2_a22oi_1 _16589_ (.Y(_06948_),
    .B1(net6008),
    .B2(\top1.memory1.mem1[57][2] ),
    .A2(net6072),
    .A1(\top1.memory1.mem1[56][2] ));
 sg13g2_a21o_1 _16590_ (.A2(_06948_),
    .A1(_06947_),
    .B1(net6082),
    .X(_06949_));
 sg13g2_mux4_1 _16591_ (.S0(net6246),
    .A0(\top1.memory1.mem1[52][2] ),
    .A1(\top1.memory1.mem1[53][2] ),
    .A2(\top1.memory1.mem1[54][2] ),
    .A3(\top1.memory1.mem1[55][2] ),
    .S1(net6181),
    .X(_06950_));
 sg13g2_mux4_1 _16592_ (.S0(net6255),
    .A0(\top1.memory1.mem1[48][2] ),
    .A1(\top1.memory1.mem1[49][2] ),
    .A2(\top1.memory1.mem1[50][2] ),
    .A3(\top1.memory1.mem1[51][2] ),
    .S1(net6190),
    .X(_06951_));
 sg13g2_and2_1 _16593_ (.A(net5886),
    .B(_06951_),
    .X(_06952_));
 sg13g2_a221oi_1 _16594_ (.B2(net6033),
    .C1(_06952_),
    .B1(_06950_),
    .A1(net5864),
    .Y(_06953_),
    .A2(_06946_));
 sg13g2_a21oi_2 _16595_ (.B1(net5840),
    .Y(_06954_),
    .A2(_06953_),
    .A1(_06949_));
 sg13g2_nor4_2 _16596_ (.A(_06928_),
    .B(_06935_),
    .C(_06945_),
    .Y(_06955_),
    .D(_06954_));
 sg13g2_or2_2 _16597_ (.X(_06956_),
    .B(_06920_),
    .A(_06913_));
 sg13g2_a21oi_2 _16598_ (.B1(_05479_),
    .Y(_06957_),
    .A2(_06892_),
    .A1(_06891_));
 sg13g2_a221oi_1 _16599_ (.B2(_06906_),
    .C1(net6111),
    .B1(_06957_),
    .A1(net6113),
    .Y(_06958_),
    .A2(_06956_));
 sg13g2_o21ai_1 _16600_ (.B1(_06958_),
    .Y(_06959_),
    .A1(net6113),
    .A2(_06955_));
 sg13g2_o21ai_1 _16601_ (.B1(net6130),
    .Y(_06960_),
    .A1(\top1.memory1.mem1[196][2] ),
    .A2(net6039));
 sg13g2_nor2_1 _16602_ (.A(\top1.memory1.mem1[198][2] ),
    .B(net5894),
    .Y(_06961_));
 sg13g2_nor2_1 _16603_ (.A(\top1.memory1.mem1[197][2] ),
    .B(net5973),
    .Y(_06962_));
 sg13g2_nor2_1 _16604_ (.A(\top1.memory1.mem1[199][2] ),
    .B(net5933),
    .Y(_06963_));
 sg13g2_nor4_2 _16605_ (.A(_06960_),
    .B(_06961_),
    .C(_06962_),
    .Y(_06964_),
    .D(_06963_));
 sg13g2_nor2_1 _16606_ (.A(\top1.memory1.mem1[192][2] ),
    .B(net6043),
    .Y(_06965_));
 sg13g2_nor2_1 _16607_ (.A(\top1.memory1.mem1[194][2] ),
    .B(net5897),
    .Y(_06966_));
 sg13g2_nor2_1 _16608_ (.A(\top1.memory1.mem1[193][2] ),
    .B(net5977),
    .Y(_06967_));
 sg13g2_nor4_1 _16609_ (.A(net6131),
    .B(_06965_),
    .C(_06966_),
    .D(_06967_),
    .Y(_06968_));
 sg13g2_o21ai_1 _16610_ (.B1(_06968_),
    .Y(_06969_),
    .A1(\top1.memory1.mem1[195][2] ),
    .A2(net5938));
 sg13g2_nor2_1 _16611_ (.A(_03979_),
    .B(_06964_),
    .Y(_06970_));
 sg13g2_a21oi_1 _16612_ (.A1(_06969_),
    .A2(_06970_),
    .Y(_06971_),
    .B1(net6108));
 sg13g2_nor2_1 _16613_ (.A(\top1.memory1.mem1[154][2] ),
    .B(net5892),
    .Y(_06972_));
 sg13g2_nor2_1 _16614_ (.A(\top1.memory1.mem1[153][2] ),
    .B(net5972),
    .Y(_06973_));
 sg13g2_nor2_1 _16615_ (.A(\top1.memory1.mem1[155][2] ),
    .B(net5935),
    .Y(_06974_));
 sg13g2_o21ai_1 _16616_ (.B1(net6085),
    .Y(_06975_),
    .A1(\top1.memory1.mem1[152][2] ),
    .A2(net6038));
 sg13g2_nor4_1 _16617_ (.A(_06972_),
    .B(_06973_),
    .C(_06974_),
    .D(_06975_),
    .Y(_06976_));
 sg13g2_a22oi_1 _16618_ (.Y(_06977_),
    .B1(net5904),
    .B2(\top1.memory1.mem1[150][2] ),
    .A2(net5945),
    .A1(\top1.memory1.mem1[151][2] ));
 sg13g2_a22oi_1 _16619_ (.Y(_06978_),
    .B1(net5984),
    .B2(\top1.memory1.mem1[149][2] ),
    .A2(net6049),
    .A1(\top1.memory1.mem1[148][2] ));
 sg13g2_a21oi_1 _16620_ (.A1(_06977_),
    .A2(_06978_),
    .Y(_06979_),
    .B1(net6011));
 sg13g2_a22oi_1 _16621_ (.Y(_06980_),
    .B1(net5908),
    .B2(\top1.memory1.mem1[146][2] ),
    .A2(net5949),
    .A1(\top1.memory1.mem1[147][2] ));
 sg13g2_a22oi_1 _16622_ (.Y(_06981_),
    .B1(net5989),
    .B2(\top1.memory1.mem1[145][2] ),
    .A2(net6053),
    .A1(\top1.memory1.mem1[144][2] ));
 sg13g2_a21oi_1 _16623_ (.A1(_06980_),
    .A2(_06981_),
    .Y(_06982_),
    .B1(net5867));
 sg13g2_a22oi_1 _16624_ (.Y(_06983_),
    .B1(net5909),
    .B2(\top1.memory1.mem1[158][2] ),
    .A2(net6054),
    .A1(\top1.memory1.mem1[156][2] ));
 sg13g2_a22oi_1 _16625_ (.Y(_06984_),
    .B1(net5949),
    .B2(\top1.memory1.mem1[159][2] ),
    .A2(net5990),
    .A1(\top1.memory1.mem1[157][2] ));
 sg13g2_a21oi_2 _16626_ (.B1(net5842),
    .Y(_06985_),
    .A2(_06984_),
    .A1(_06983_));
 sg13g2_nor4_2 _16627_ (.A(_06976_),
    .B(_06979_),
    .C(_06982_),
    .Y(_06986_),
    .D(_06985_));
 sg13g2_nand2b_2 _16628_ (.Y(_06987_),
    .B(_05516_),
    .A_N(_06986_));
 sg13g2_a22oi_1 _16629_ (.Y(_06988_),
    .B1(net5907),
    .B2(\top1.memory1.mem1[134][2] ),
    .A2(net5947),
    .A1(\top1.memory1.mem1[135][2] ));
 sg13g2_a22oi_1 _16630_ (.Y(_06989_),
    .B1(net5982),
    .B2(\top1.memory1.mem1[133][2] ),
    .A2(net6047),
    .A1(\top1.memory1.mem1[132][2] ));
 sg13g2_a21oi_1 _16631_ (.A1(_06988_),
    .A2(_06989_),
    .Y(_06990_),
    .B1(net6015));
 sg13g2_a22oi_1 _16632_ (.Y(_06991_),
    .B1(net5982),
    .B2(\top1.memory1.mem1[129][2] ),
    .A2(net6047),
    .A1(\top1.memory1.mem1[128][2] ));
 sg13g2_a22oi_1 _16633_ (.Y(_06992_),
    .B1(net5902),
    .B2(\top1.memory1.mem1[130][2] ),
    .A2(net5943),
    .A1(\top1.memory1.mem1[131][2] ));
 sg13g2_a21oi_1 _16634_ (.A1(_06991_),
    .A2(_06992_),
    .Y(_06993_),
    .B1(net5868));
 sg13g2_a22oi_1 _16635_ (.Y(_06994_),
    .B1(net5907),
    .B2(\top1.memory1.mem1[142][2] ),
    .A2(net5947),
    .A1(\top1.memory1.mem1[143][2] ));
 sg13g2_a22oi_1 _16636_ (.Y(_06995_),
    .B1(net5988),
    .B2(\top1.memory1.mem1[141][2] ),
    .A2(net6052),
    .A1(\top1.memory1.mem1[140][2] ));
 sg13g2_a21oi_1 _16637_ (.A1(_06994_),
    .A2(_06995_),
    .Y(_06996_),
    .B1(net5842));
 sg13g2_nor2_1 _16638_ (.A(\top1.memory1.mem1[136][2] ),
    .B(net6036),
    .Y(_06997_));
 sg13g2_nor2_1 _16639_ (.A(\top1.memory1.mem1[139][2] ),
    .B(net5931),
    .Y(_06998_));
 sg13g2_nor2_1 _16640_ (.A(\top1.memory1.mem1[138][2] ),
    .B(net5891),
    .Y(_06999_));
 sg13g2_o21ai_1 _16641_ (.B1(net6084),
    .Y(_07000_),
    .A1(\top1.memory1.mem1[137][2] ),
    .A2(net5970));
 sg13g2_nor4_1 _16642_ (.A(_06997_),
    .B(_06998_),
    .C(_06999_),
    .D(_07000_),
    .Y(_07001_));
 sg13g2_or4_2 _16643_ (.A(_06990_),
    .B(_06993_),
    .C(_06996_),
    .D(_07001_),
    .X(_07002_));
 sg13g2_a22oi_1 _16644_ (.Y(_07003_),
    .B1(net5926),
    .B2(\top1.memory1.mem1[178][2] ),
    .A2(net5966),
    .A1(\top1.memory1.mem1[179][2] ));
 sg13g2_a22oi_1 _16645_ (.Y(_07004_),
    .B1(net6006),
    .B2(\top1.memory1.mem1[177][2] ),
    .A2(net6070),
    .A1(\top1.memory1.mem1[176][2] ));
 sg13g2_a21oi_1 _16646_ (.A1(_07003_),
    .A2(_07004_),
    .Y(_07005_),
    .B1(net5871));
 sg13g2_a22oi_1 _16647_ (.Y(_07006_),
    .B1(net5926),
    .B2(\top1.memory1.mem1[182][2] ),
    .A2(net5966),
    .A1(\top1.memory1.mem1[183][2] ));
 sg13g2_a22oi_1 _16648_ (.Y(_07007_),
    .B1(net6006),
    .B2(\top1.memory1.mem1[181][2] ),
    .A2(net6070),
    .A1(\top1.memory1.mem1[180][2] ));
 sg13g2_a21oi_2 _16649_ (.B1(net6014),
    .Y(_07008_),
    .A2(_07007_),
    .A1(_07006_));
 sg13g2_a22oi_1 _16650_ (.Y(_07009_),
    .B1(net5926),
    .B2(\top1.memory1.mem1[190][2] ),
    .A2(net5966),
    .A1(\top1.memory1.mem1[191][2] ));
 sg13g2_a22oi_1 _16651_ (.Y(_07010_),
    .B1(net6006),
    .B2(\top1.memory1.mem1[189][2] ),
    .A2(net6070),
    .A1(\top1.memory1.mem1[188][2] ));
 sg13g2_a21oi_1 _16652_ (.A1(_07009_),
    .A2(_07010_),
    .Y(_07011_),
    .B1(net5848));
 sg13g2_nor2_1 _16653_ (.A(\top1.memory1.mem1[186][2] ),
    .B(net5899),
    .Y(_07012_));
 sg13g2_nor2_1 _16654_ (.A(\top1.memory1.mem1[187][2] ),
    .B(net5940),
    .Y(_07013_));
 sg13g2_nor2_1 _16655_ (.A(\top1.memory1.mem1[184][2] ),
    .B(net6045),
    .Y(_07014_));
 sg13g2_o21ai_1 _16656_ (.B1(net6089),
    .Y(_07015_),
    .A1(\top1.memory1.mem1[185][2] ),
    .A2(net5979));
 sg13g2_nor4_2 _16657_ (.A(_07012_),
    .B(_07013_),
    .C(_07014_),
    .Y(_07016_),
    .D(_07015_));
 sg13g2_nor4_2 _16658_ (.A(_07005_),
    .B(_07008_),
    .C(_07011_),
    .Y(_07017_),
    .D(_07016_));
 sg13g2_nand2b_1 _16659_ (.Y(_07018_),
    .B(_05452_),
    .A_N(_07017_));
 sg13g2_nor2_1 _16660_ (.A(\top1.memory1.mem1[170][2] ),
    .B(net5900),
    .Y(_07019_));
 sg13g2_nor2_1 _16661_ (.A(\top1.memory1.mem1[169][2] ),
    .B(net5980),
    .Y(_07020_));
 sg13g2_nor2_1 _16662_ (.A(\top1.memory1.mem1[168][2] ),
    .B(net6045),
    .Y(_07021_));
 sg13g2_o21ai_1 _16663_ (.B1(net6089),
    .Y(_07022_),
    .A1(\top1.memory1.mem1[171][2] ),
    .A2(net5941));
 sg13g2_nor4_1 _16664_ (.A(_07019_),
    .B(_07020_),
    .C(_07021_),
    .D(_07022_),
    .Y(_07023_));
 sg13g2_a22oi_1 _16665_ (.Y(_07024_),
    .B1(net5919),
    .B2(\top1.memory1.mem1[166][2] ),
    .A2(net6064),
    .A1(\top1.memory1.mem1[164][2] ));
 sg13g2_a22oi_1 _16666_ (.Y(_07025_),
    .B1(net5959),
    .B2(\top1.memory1.mem1[167][2] ),
    .A2(net6000),
    .A1(\top1.memory1.mem1[165][2] ));
 sg13g2_a21oi_1 _16667_ (.A1(_07024_),
    .A2(_07025_),
    .Y(_07026_),
    .B1(net6012));
 sg13g2_a22oi_1 _16668_ (.Y(_07027_),
    .B1(net5918),
    .B2(\top1.memory1.mem1[174][2] ),
    .A2(net6063),
    .A1(\top1.memory1.mem1[172][2] ));
 sg13g2_a22oi_1 _16669_ (.Y(_07028_),
    .B1(net5958),
    .B2(\top1.memory1.mem1[175][2] ),
    .A2(net5999),
    .A1(\top1.memory1.mem1[173][2] ));
 sg13g2_a21oi_1 _16670_ (.A1(_07027_),
    .A2(_07028_),
    .Y(_07029_),
    .B1(net5847));
 sg13g2_a22oi_1 _16671_ (.Y(_07030_),
    .B1(net5918),
    .B2(\top1.memory1.mem1[162][2] ),
    .A2(net5958),
    .A1(\top1.memory1.mem1[163][2] ));
 sg13g2_a22oi_1 _16672_ (.Y(_07031_),
    .B1(net5999),
    .B2(\top1.memory1.mem1[161][2] ),
    .A2(net6063),
    .A1(\top1.memory1.mem1[160][2] ));
 sg13g2_a21oi_1 _16673_ (.A1(_07030_),
    .A2(_07031_),
    .Y(_07032_),
    .B1(net5870));
 sg13g2_or4_2 _16674_ (.A(_07023_),
    .B(_07026_),
    .C(_07029_),
    .D(_07032_),
    .X(_07033_));
 sg13g2_a22oi_1 _16675_ (.Y(_07034_),
    .B1(_07033_),
    .B2(_05443_),
    .A2(_07002_),
    .A1(_03976_));
 sg13g2_nand4_1 _16676_ (.B(_06987_),
    .C(_07018_),
    .A(_05514_),
    .Y(_07035_),
    .D(_07034_));
 sg13g2_nand3_1 _16677_ (.B(_06971_),
    .C(_07035_),
    .A(_06959_),
    .Y(_07036_));
 sg13g2_mux4_1 _16678_ (.S0(net6237),
    .A0(\top1.memory1.mem2[124][2] ),
    .A1(\top1.memory1.mem2[125][2] ),
    .A2(\top1.memory1.mem2[126][2] ),
    .A3(\top1.memory1.mem2[127][2] ),
    .S1(net6172),
    .X(_07037_));
 sg13g2_mux4_1 _16679_ (.S0(net6240),
    .A0(\top1.memory1.mem2[112][2] ),
    .A1(\top1.memory1.mem2[113][2] ),
    .A2(\top1.memory1.mem2[114][2] ),
    .A3(\top1.memory1.mem2[115][2] ),
    .S1(net6175),
    .X(_07038_));
 sg13g2_mux4_1 _16680_ (.S0(net6237),
    .A0(\top1.memory1.mem2[116][2] ),
    .A1(\top1.memory1.mem2[117][2] ),
    .A2(\top1.memory1.mem2[118][2] ),
    .A3(\top1.memory1.mem2[119][2] ),
    .S1(net6172),
    .X(_07039_));
 sg13g2_mux4_1 _16681_ (.S0(net6240),
    .A0(\top1.memory1.mem2[120][2] ),
    .A1(\top1.memory1.mem2[121][2] ),
    .A2(\top1.memory1.mem2[122][2] ),
    .A3(\top1.memory1.mem2[123][2] ),
    .S1(net6175),
    .X(_07040_));
 sg13g2_a22oi_1 _16682_ (.Y(_07041_),
    .B1(_07039_),
    .B2(net6031),
    .A2(_07037_),
    .A1(net5859));
 sg13g2_a22oi_1 _16683_ (.Y(_07042_),
    .B1(_07040_),
    .B2(net6095),
    .A2(_07038_),
    .A1(net5885));
 sg13g2_a21oi_2 _16684_ (.B1(net5838),
    .Y(_07043_),
    .A2(_07042_),
    .A1(_07041_));
 sg13g2_mux4_1 _16685_ (.S0(net6223),
    .A0(\top1.memory1.mem2[100][2] ),
    .A1(\top1.memory1.mem2[101][2] ),
    .A2(\top1.memory1.mem2[102][2] ),
    .A3(\top1.memory1.mem2[103][2] ),
    .S1(net6158),
    .X(_07044_));
 sg13g2_mux4_1 _16686_ (.S0(net6227),
    .A0(\top1.memory1.mem2[96][2] ),
    .A1(\top1.memory1.mem2[97][2] ),
    .A2(\top1.memory1.mem2[98][2] ),
    .A3(\top1.memory1.mem2[99][2] ),
    .S1(net6162),
    .X(_07045_));
 sg13g2_a22oi_1 _16687_ (.Y(_07046_),
    .B1(_07045_),
    .B2(net5880),
    .A2(_07044_),
    .A1(net6025));
 sg13g2_mux4_1 _16688_ (.S0(net6236),
    .A0(\top1.memory1.mem2[104][2] ),
    .A1(\top1.memory1.mem2[105][2] ),
    .A2(\top1.memory1.mem2[106][2] ),
    .A3(\top1.memory1.mem2[107][2] ),
    .S1(net6171),
    .X(_07047_));
 sg13g2_mux4_1 _16689_ (.S0(net6236),
    .A0(\top1.memory1.mem2[108][2] ),
    .A1(\top1.memory1.mem2[109][2] ),
    .A2(\top1.memory1.mem2[110][2] ),
    .A3(\top1.memory1.mem2[111][2] ),
    .S1(net6171),
    .X(_07048_));
 sg13g2_a22oi_1 _16690_ (.Y(_07049_),
    .B1(_07048_),
    .B2(net5859),
    .A2(_07047_),
    .A1(net6093));
 sg13g2_a21oi_1 _16691_ (.A1(_07046_),
    .A2(_07049_),
    .Y(_07050_),
    .B1(net5832));
 sg13g2_mux4_1 _16692_ (.S0(net6198),
    .A0(\top1.memory1.mem2[64][2] ),
    .A1(\top1.memory1.mem2[65][2] ),
    .A2(\top1.memory1.mem2[66][2] ),
    .A3(\top1.memory1.mem2[67][2] ),
    .S1(net6134),
    .X(_07051_));
 sg13g2_mux4_1 _16693_ (.S0(net6197),
    .A0(\top1.memory1.mem2[76][2] ),
    .A1(\top1.memory1.mem2[77][2] ),
    .A2(\top1.memory1.mem2[78][2] ),
    .A3(\top1.memory1.mem2[79][2] ),
    .S1(net6133),
    .X(_07052_));
 sg13g2_a22oi_1 _16694_ (.Y(_07053_),
    .B1(net5903),
    .B2(_03921_),
    .A2(net6048),
    .A1(_03919_));
 sg13g2_a221oi_1 _16695_ (.B2(_03922_),
    .C1(net6075),
    .B1(net5944),
    .A1(_03920_),
    .Y(_07054_),
    .A2(net5983));
 sg13g2_mux4_1 _16696_ (.S0(net6200),
    .A0(\top1.memory1.mem2[68][2] ),
    .A1(\top1.memory1.mem2[69][2] ),
    .A2(\top1.memory1.mem2[70][2] ),
    .A3(\top1.memory1.mem2[71][2] ),
    .S1(net6136),
    .X(_07055_));
 sg13g2_mux4_1 _16697_ (.S0(net6201),
    .A0(\top1.memory1.mem2[80][2] ),
    .A1(\top1.memory1.mem2[81][2] ),
    .A2(\top1.memory1.mem2[82][2] ),
    .A3(\top1.memory1.mem2[83][2] ),
    .S1(net6137),
    .X(_07056_));
 sg13g2_a22oi_1 _16698_ (.Y(_07057_),
    .B1(net5911),
    .B2(\top1.memory1.mem2[94][2] ),
    .A2(net5951),
    .A1(\top1.memory1.mem2[95][2] ));
 sg13g2_a22oi_1 _16699_ (.Y(_07058_),
    .B1(net5993),
    .B2(\top1.memory1.mem2[93][2] ),
    .A2(net6056),
    .A1(\top1.memory1.mem2[92][2] ));
 sg13g2_a21o_1 _16700_ (.A2(_07058_),
    .A1(_07057_),
    .B1(net5845),
    .X(_07059_));
 sg13g2_mux4_1 _16701_ (.S0(net6202),
    .A0(\top1.memory1.mem2[84][2] ),
    .A1(\top1.memory1.mem2[85][2] ),
    .A2(\top1.memory1.mem2[86][2] ),
    .A3(\top1.memory1.mem2[87][2] ),
    .S1(net6138),
    .X(_07060_));
 sg13g2_nor2_1 _16702_ (.A(\top1.memory1.mem2[91][2] ),
    .B(net5933),
    .Y(_07061_));
 sg13g2_nor2_1 _16703_ (.A(\top1.memory1.mem2[90][2] ),
    .B(net5895),
    .Y(_07062_));
 sg13g2_nor2_1 _16704_ (.A(\top1.memory1.mem2[89][2] ),
    .B(net5974),
    .Y(_07063_));
 sg13g2_o21ai_1 _16705_ (.B1(net6083),
    .Y(_07064_),
    .A1(\top1.memory1.mem2[88][2] ),
    .A2(net6040));
 sg13g2_or4_1 _16706_ (.A(_07061_),
    .B(_07062_),
    .C(_07063_),
    .D(_07064_),
    .X(_07065_));
 sg13g2_a21oi_1 _16707_ (.A1(_03914_),
    .A2(net5915),
    .Y(_07066_),
    .B1(net6077));
 sg13g2_nor3_1 _16708_ (.A(net6216),
    .B(net6151),
    .C(\top1.memory1.mem2[8][2] ),
    .Y(_07067_));
 sg13g2_a221oi_1 _16709_ (.B2(_03915_),
    .C1(_07067_),
    .B1(net5955),
    .A1(_03913_),
    .Y(_07068_),
    .A2(net5996));
 sg13g2_mux4_1 _16710_ (.S0(net6216),
    .A0(\top1.memory1.mem2[4][2] ),
    .A1(\top1.memory1.mem2[5][2] ),
    .A2(\top1.memory1.mem2[6][2] ),
    .A3(\top1.memory1.mem2[7][2] ),
    .S1(net6151),
    .X(_07069_));
 sg13g2_mux4_1 _16711_ (.S0(net6215),
    .A0(\top1.memory1.mem2[12][2] ),
    .A1(\top1.memory1.mem2[13][2] ),
    .A2(\top1.memory1.mem2[14][2] ),
    .A3(\top1.memory1.mem2[15][2] ),
    .S1(net6150),
    .X(_07070_));
 sg13g2_a22oi_1 _16712_ (.Y(_07071_),
    .B1(net5921),
    .B2(\top1.memory1.mem2[2][2] ),
    .A2(net6065),
    .A1(\top1.memory1.mem2[0][2] ));
 sg13g2_a22oi_1 _16713_ (.Y(_07072_),
    .B1(net5961),
    .B2(\top1.memory1.mem2[3][2] ),
    .A2(net6002),
    .A1(\top1.memory1.mem2[1][2] ));
 sg13g2_a21o_1 _16714_ (.A2(_07072_),
    .A1(_07071_),
    .B1(net5871),
    .X(_07073_));
 sg13g2_a21o_1 _16715_ (.A2(_07070_),
    .A1(net5854),
    .B1(net6125),
    .X(_07074_));
 sg13g2_a221oi_1 _16716_ (.B2(net6023),
    .C1(_07074_),
    .B1(_07069_),
    .A1(_07066_),
    .Y(_07075_),
    .A2(_07068_));
 sg13g2_a21oi_1 _16717_ (.A1(_03918_),
    .A2(net5963),
    .Y(_07076_),
    .B1(net6080));
 sg13g2_nor3_1 _16718_ (.A(net6230),
    .B(net6165),
    .C(\top1.memory1.mem2[24][2] ),
    .Y(_07077_));
 sg13g2_a221oi_1 _16719_ (.B2(_03917_),
    .C1(_07077_),
    .B1(net5923),
    .A1(_03916_),
    .Y(_07078_),
    .A2(net6004));
 sg13g2_mux4_1 _16720_ (.S0(net6230),
    .A0(\top1.memory1.mem2[20][2] ),
    .A1(\top1.memory1.mem2[21][2] ),
    .A2(\top1.memory1.mem2[22][2] ),
    .A3(\top1.memory1.mem2[23][2] ),
    .S1(net6165),
    .X(_07079_));
 sg13g2_mux4_1 _16721_ (.S0(net6216),
    .A0(\top1.memory1.mem2[28][2] ),
    .A1(\top1.memory1.mem2[29][2] ),
    .A2(\top1.memory1.mem2[30][2] ),
    .A3(\top1.memory1.mem2[31][2] ),
    .S1(net6151),
    .X(_07080_));
 sg13g2_mux4_1 _16722_ (.S0(net6231),
    .A0(\top1.memory1.mem2[16][2] ),
    .A1(\top1.memory1.mem2[17][2] ),
    .A2(\top1.memory1.mem2[18][2] ),
    .A3(\top1.memory1.mem2[19][2] ),
    .S1(net6166),
    .X(_07081_));
 sg13g2_and2_1 _16723_ (.A(net5882),
    .B(_07081_),
    .X(_07082_));
 sg13g2_a21oi_1 _16724_ (.A1(net5854),
    .A2(_07080_),
    .Y(_07083_),
    .B1(net6106));
 sg13g2_a221oi_1 _16725_ (.B2(net6027),
    .C1(_07082_),
    .B1(_07079_),
    .A1(_07076_),
    .Y(_07084_),
    .A2(_07078_));
 sg13g2_a221oi_1 _16726_ (.B2(_07084_),
    .C1(net6119),
    .B1(_07083_),
    .A1(_07073_),
    .Y(_07085_),
    .A2(_07075_));
 sg13g2_mux4_1 _16727_ (.S0(net6252),
    .A0(\top1.memory1.mem2[60][2] ),
    .A1(\top1.memory1.mem2[61][2] ),
    .A2(\top1.memory1.mem2[62][2] ),
    .A3(\top1.memory1.mem2[63][2] ),
    .S1(net6187),
    .X(_07086_));
 sg13g2_mux4_1 _16728_ (.S0(net6253),
    .A0(\top1.memory1.mem2[48][2] ),
    .A1(\top1.memory1.mem2[49][2] ),
    .A2(\top1.memory1.mem2[50][2] ),
    .A3(\top1.memory1.mem2[51][2] ),
    .S1(net6188),
    .X(_07087_));
 sg13g2_mux4_1 _16729_ (.S0(net6250),
    .A0(\top1.memory1.mem2[56][2] ),
    .A1(\top1.memory1.mem2[57][2] ),
    .A2(\top1.memory1.mem2[58][2] ),
    .A3(\top1.memory1.mem2[59][2] ),
    .S1(net6185),
    .X(_07088_));
 sg13g2_mux4_1 _16730_ (.S0(net6251),
    .A0(\top1.memory1.mem2[52][2] ),
    .A1(\top1.memory1.mem2[53][2] ),
    .A2(\top1.memory1.mem2[54][2] ),
    .A3(\top1.memory1.mem2[55][2] ),
    .S1(net6186),
    .X(_07089_));
 sg13g2_a22oi_1 _16731_ (.Y(_07090_),
    .B1(_07088_),
    .B2(net6097),
    .A2(_07086_),
    .A1(net5862));
 sg13g2_a22oi_1 _16732_ (.Y(_07091_),
    .B1(_07089_),
    .B2(net6034),
    .A2(_07087_),
    .A1(net5888));
 sg13g2_a21oi_1 _16733_ (.A1(_07090_),
    .A2(_07091_),
    .Y(_07092_),
    .B1(net5840));
 sg13g2_mux4_1 _16734_ (.S0(net6249),
    .A0(\top1.memory1.mem2[40][2] ),
    .A1(\top1.memory1.mem2[41][2] ),
    .A2(\top1.memory1.mem2[42][2] ),
    .A3(\top1.memory1.mem2[43][2] ),
    .S1(net6184),
    .X(_07093_));
 sg13g2_mux4_1 _16735_ (.S0(net6234),
    .A0(\top1.memory1.mem2[44][2] ),
    .A1(\top1.memory1.mem2[45][2] ),
    .A2(\top1.memory1.mem2[46][2] ),
    .A3(\top1.memory1.mem2[47][2] ),
    .S1(net6169),
    .X(_07094_));
 sg13g2_mux4_1 _16736_ (.S0(net6232),
    .A0(\top1.memory1.mem2[32][2] ),
    .A1(\top1.memory1.mem2[33][2] ),
    .A2(\top1.memory1.mem2[34][2] ),
    .A3(\top1.memory1.mem2[35][2] ),
    .S1(net6167),
    .X(_07095_));
 sg13g2_mux4_1 _16737_ (.S0(net6234),
    .A0(\top1.memory1.mem2[36][2] ),
    .A1(\top1.memory1.mem2[37][2] ),
    .A2(\top1.memory1.mem2[38][2] ),
    .A3(\top1.memory1.mem2[39][2] ),
    .S1(net6169),
    .X(_07096_));
 sg13g2_a22oi_1 _16738_ (.Y(_07097_),
    .B1(_07095_),
    .B2(net5883),
    .A2(_07093_),
    .A1(net6099));
 sg13g2_a22oi_1 _16739_ (.Y(_07098_),
    .B1(_07096_),
    .B2(net6027),
    .A2(_07094_),
    .A1(net5858));
 sg13g2_a21oi_1 _16740_ (.A1(_07097_),
    .A2(_07098_),
    .Y(_07099_),
    .B1(net5834));
 sg13g2_or2_2 _16741_ (.X(_07100_),
    .B(_07099_),
    .A(_07092_));
 sg13g2_o21ai_1 _16742_ (.B1(net6102),
    .Y(_07101_),
    .A1(_07085_),
    .A2(_07100_));
 sg13g2_a221oi_1 _16743_ (.B2(net6017),
    .C1(net6104),
    .B1(_07060_),
    .A1(net5874),
    .Y(_07102_),
    .A2(_07056_));
 sg13g2_nand3_1 _16744_ (.B(_07065_),
    .C(_07102_),
    .A(_07059_),
    .Y(_07103_));
 sg13g2_a22oi_1 _16745_ (.Y(_07104_),
    .B1(_07053_),
    .B2(_07054_),
    .A2(_07051_),
    .A1(net5873));
 sg13g2_a221oi_1 _16746_ (.B2(net6017),
    .C1(net6120),
    .B1(_07055_),
    .A1(net5850),
    .Y(_07105_),
    .A2(_07052_));
 sg13g2_a21oi_2 _16747_ (.B1(_05479_),
    .Y(_07106_),
    .A2(_07105_),
    .A1(_07104_));
 sg13g2_or2_2 _16748_ (.X(_07107_),
    .B(_07050_),
    .A(_07043_));
 sg13g2_a221oi_1 _16749_ (.B2(net6113),
    .C1(net6111),
    .B1(_07107_),
    .A1(_07103_),
    .Y(_07108_),
    .A2(_07106_));
 sg13g2_mux4_1 _16750_ (.S0(net6232),
    .A0(\top1.memory1.mem2[180][2] ),
    .A1(\top1.memory1.mem2[181][2] ),
    .A2(\top1.memory1.mem2[182][2] ),
    .A3(\top1.memory1.mem2[183][2] ),
    .S1(net6167),
    .X(_07109_));
 sg13g2_mux4_1 _16751_ (.S0(net6234),
    .A0(\top1.memory1.mem2[176][2] ),
    .A1(\top1.memory1.mem2[177][2] ),
    .A2(\top1.memory1.mem2[178][2] ),
    .A3(\top1.memory1.mem2[179][2] ),
    .S1(net6169),
    .X(_07110_));
 sg13g2_mux4_1 _16752_ (.S0(net6232),
    .A0(\top1.memory1.mem2[188][2] ),
    .A1(\top1.memory1.mem2[189][2] ),
    .A2(\top1.memory1.mem2[190][2] ),
    .A3(\top1.memory1.mem2[191][2] ),
    .S1(net6167),
    .X(_07111_));
 sg13g2_mux4_1 _16753_ (.S0(net6230),
    .A0(\top1.memory1.mem2[184][2] ),
    .A1(\top1.memory1.mem2[185][2] ),
    .A2(\top1.memory1.mem2[186][2] ),
    .A3(\top1.memory1.mem2[187][2] ),
    .S1(net6165),
    .X(_07112_));
 sg13g2_a22oi_1 _16754_ (.Y(_07113_),
    .B1(_07111_),
    .B2(net5858),
    .A2(_07109_),
    .A1(net6027));
 sg13g2_a22oi_1 _16755_ (.Y(_07114_),
    .B1(_07112_),
    .B2(net6091),
    .A2(_07110_),
    .A1(net5882));
 sg13g2_a21oi_2 _16756_ (.B1(net5837),
    .Y(_07115_),
    .A2(_07114_),
    .A1(_07113_));
 sg13g2_nor2_1 _16757_ (.A(net5831),
    .B(_07115_),
    .Y(_07116_));
 sg13g2_mux4_1 _16758_ (.S0(net6217),
    .A0(\top1.memory1.mem2[164][2] ),
    .A1(\top1.memory1.mem2[165][2] ),
    .A2(\top1.memory1.mem2[166][2] ),
    .A3(\top1.memory1.mem2[167][2] ),
    .S1(net6152),
    .X(_07117_));
 sg13g2_mux4_1 _16759_ (.S0(net6229),
    .A0(\top1.memory1.mem2[168][2] ),
    .A1(\top1.memory1.mem2[169][2] ),
    .A2(\top1.memory1.mem2[170][2] ),
    .A3(\top1.memory1.mem2[171][2] ),
    .S1(net6164),
    .X(_07118_));
 sg13g2_a22oi_1 _16760_ (.Y(_07119_),
    .B1(net5915),
    .B2(\top1.memory1.mem2[162][2] ),
    .A2(net5955),
    .A1(\top1.memory1.mem2[163][2] ));
 sg13g2_a22oi_1 _16761_ (.Y(_07120_),
    .B1(net5995),
    .B2(\top1.memory1.mem2[161][2] ),
    .A2(net6060),
    .A1(\top1.memory1.mem2[160][2] ));
 sg13g2_a21o_1 _16762_ (.A2(_07120_),
    .A1(_07119_),
    .B1(net5869),
    .X(_07121_));
 sg13g2_mux4_1 _16763_ (.S0(net6214),
    .A0(\top1.memory1.mem2[172][2] ),
    .A1(\top1.memory1.mem2[173][2] ),
    .A2(\top1.memory1.mem2[174][2] ),
    .A3(\top1.memory1.mem2[175][2] ),
    .S1(net6149),
    .X(_07122_));
 sg13g2_and2_1 _16764_ (.A(net5853),
    .B(_07122_),
    .X(_07123_));
 sg13g2_a221oi_1 _16765_ (.B2(net6091),
    .C1(_07123_),
    .B1(_07118_),
    .A1(net6023),
    .Y(_07124_),
    .A2(_07117_));
 sg13g2_a21oi_2 _16766_ (.B1(net5836),
    .Y(_07125_),
    .A2(_07124_),
    .A1(_07121_));
 sg13g2_a22oi_1 _16767_ (.Y(_07126_),
    .B1(net5905),
    .B2(\top1.memory1.mem2[130][2] ),
    .A2(net6050),
    .A1(\top1.memory1.mem2[128][2] ));
 sg13g2_a22oi_1 _16768_ (.Y(_07127_),
    .B1(net5946),
    .B2(\top1.memory1.mem2[131][2] ),
    .A2(net5986),
    .A1(\top1.memory1.mem2[129][2] ));
 sg13g2_a21oi_1 _16769_ (.A1(_07126_),
    .A2(_07127_),
    .Y(_07128_),
    .B1(net5867));
 sg13g2_nor2_1 _16770_ (.A(\top1.memory1.mem2[137][2] ),
    .B(net5972),
    .Y(_07129_));
 sg13g2_nor2_1 _16771_ (.A(\top1.memory1.mem2[138][2] ),
    .B(net5891),
    .Y(_07130_));
 sg13g2_nor2_1 _16772_ (.A(\top1.memory1.mem2[136][2] ),
    .B(net6038),
    .Y(_07131_));
 sg13g2_o21ai_1 _16773_ (.B1(net6084),
    .Y(_07132_),
    .A1(\top1.memory1.mem2[139][2] ),
    .A2(net5930));
 sg13g2_nor4_1 _16774_ (.A(_07129_),
    .B(_07130_),
    .C(_07131_),
    .D(_07132_),
    .Y(_07133_));
 sg13g2_a22oi_1 _16775_ (.Y(_07134_),
    .B1(net5905),
    .B2(\top1.memory1.mem2[142][2] ),
    .A2(net5946),
    .A1(\top1.memory1.mem2[143][2] ));
 sg13g2_a22oi_1 _16776_ (.Y(_07135_),
    .B1(net5986),
    .B2(\top1.memory1.mem2[141][2] ),
    .A2(net6050),
    .A1(\top1.memory1.mem2[140][2] ));
 sg13g2_a21oi_1 _16777_ (.A1(_07134_),
    .A2(_07135_),
    .Y(_07136_),
    .B1(net5842));
 sg13g2_a22oi_1 _16778_ (.Y(_07137_),
    .B1(net5950),
    .B2(\top1.memory1.mem2[135][2] ),
    .A2(net5987),
    .A1(\top1.memory1.mem2[133][2] ));
 sg13g2_a22oi_1 _16779_ (.Y(_07138_),
    .B1(net5906),
    .B2(\top1.memory1.mem2[134][2] ),
    .A2(net6051),
    .A1(\top1.memory1.mem2[132][2] ));
 sg13g2_a21oi_1 _16780_ (.A1(_07137_),
    .A2(_07138_),
    .Y(_07139_),
    .B1(net6011));
 sg13g2_or4_2 _16781_ (.A(_07128_),
    .B(_07133_),
    .C(_07136_),
    .D(_07139_),
    .X(_07140_));
 sg13g2_a22oi_1 _16782_ (.Y(_07141_),
    .B1(net5914),
    .B2(\top1.memory1.mem2[150][2] ),
    .A2(net5954),
    .A1(\top1.memory1.mem2[151][2] ));
 sg13g2_a22oi_1 _16783_ (.Y(_07142_),
    .B1(net5994),
    .B2(\top1.memory1.mem2[149][2] ),
    .A2(net6058),
    .A1(\top1.memory1.mem2[148][2] ));
 sg13g2_a21oi_1 _16784_ (.A1(_07141_),
    .A2(_07142_),
    .Y(_07143_),
    .B1(net6015));
 sg13g2_nor2_1 _16785_ (.A(\top1.memory1.mem2[154][2] ),
    .B(net5896),
    .Y(_07144_));
 sg13g2_nor2_1 _16786_ (.A(\top1.memory1.mem2[153][2] ),
    .B(net5975),
    .Y(_07145_));
 sg13g2_nor2_1 _16787_ (.A(\top1.memory1.mem2[155][2] ),
    .B(net5939),
    .Y(_07146_));
 sg13g2_o21ai_1 _16788_ (.B1(net6088),
    .Y(_07147_),
    .A1(\top1.memory1.mem2[152][2] ),
    .A2(net6042));
 sg13g2_nor4_1 _16789_ (.A(_07144_),
    .B(_07145_),
    .C(_07146_),
    .D(_07147_),
    .Y(_07148_));
 sg13g2_a22oi_1 _16790_ (.Y(_07149_),
    .B1(net5913),
    .B2(\top1.memory1.mem2[158][2] ),
    .A2(net6058),
    .A1(\top1.memory1.mem2[156][2] ));
 sg13g2_a22oi_1 _16791_ (.Y(_07150_),
    .B1(net5953),
    .B2(\top1.memory1.mem2[159][2] ),
    .A2(net5994),
    .A1(\top1.memory1.mem2[157][2] ));
 sg13g2_a21oi_1 _16792_ (.A1(_07149_),
    .A2(_07150_),
    .Y(_07151_),
    .B1(net5845));
 sg13g2_a22oi_1 _16793_ (.Y(_07152_),
    .B1(net5953),
    .B2(\top1.memory1.mem2[147][2] ),
    .A2(net5994),
    .A1(\top1.memory1.mem2[145][2] ));
 sg13g2_a22oi_1 _16794_ (.Y(_07153_),
    .B1(net5913),
    .B2(\top1.memory1.mem2[146][2] ),
    .A2(net6058),
    .A1(\top1.memory1.mem2[144][2] ));
 sg13g2_a21oi_1 _16795_ (.A1(_07152_),
    .A2(_07153_),
    .Y(_07154_),
    .B1(net5869));
 sg13g2_or4_1 _16796_ (.A(_07143_),
    .B(_07148_),
    .C(_07151_),
    .D(_07154_),
    .X(_07155_));
 sg13g2_a221oi_1 _16797_ (.B2(_05516_),
    .C1(_07125_),
    .B1(_07155_),
    .A1(_03976_),
    .Y(_07156_),
    .A2(_07140_));
 sg13g2_o21ai_1 _16798_ (.B1(net6132),
    .Y(_07157_),
    .A1(\top1.memory1.mem2[199][2] ),
    .A2(net5939));
 sg13g2_nor2_1 _16799_ (.A(\top1.memory1.mem2[198][2] ),
    .B(net5898),
    .Y(_07158_));
 sg13g2_nor2_1 _16800_ (.A(\top1.memory1.mem2[197][2] ),
    .B(net5978),
    .Y(_07159_));
 sg13g2_nor2_1 _16801_ (.A(\top1.memory1.mem2[196][2] ),
    .B(net6044),
    .Y(_07160_));
 sg13g2_nor4_1 _16802_ (.A(_07157_),
    .B(_07158_),
    .C(_07159_),
    .D(_07160_),
    .Y(_07161_));
 sg13g2_a21oi_1 _16803_ (.A1(_03923_),
    .A2(net5915),
    .Y(_07162_),
    .B1(net6131));
 sg13g2_nand2b_1 _16804_ (.Y(_07163_),
    .B(net5954),
    .A_N(\top1.memory1.mem2[195][2] ));
 sg13g2_o21ai_1 _16805_ (.B1(_07163_),
    .Y(_07164_),
    .A1(\top1.memory1.mem2[192][2] ),
    .A2(net6041));
 sg13g2_o21ai_1 _16806_ (.B1(_07162_),
    .Y(_07165_),
    .A1(\top1.memory1.mem2[193][2] ),
    .A2(net5979));
 sg13g2_o21ai_1 _16807_ (.B1(_03978_),
    .Y(_07166_),
    .A1(_07164_),
    .A2(_07165_));
 sg13g2_o21ai_1 _16808_ (.B1(net6108),
    .Y(_07167_),
    .A1(_07161_),
    .A2(_07166_));
 sg13g2_a221oi_1 _16809_ (.B2(_07156_),
    .C1(_07167_),
    .B1(_07116_),
    .A1(_07101_),
    .Y(_07168_),
    .A2(_07108_));
 sg13g2_nor2_1 _16810_ (.A(_03832_),
    .B(_07168_),
    .Y(_07169_));
 sg13g2_a22oi_1 _16811_ (.Y(_01056_),
    .B1(_07036_),
    .B2(_07169_),
    .A2(_03853_),
    .A1(net6101));
 sg13g2_nand3_1 _16812_ (.B(net7075),
    .C(net7223),
    .A(net7286),
    .Y(_07170_));
 sg13g2_nand2_1 _16813_ (.Y(_07171_),
    .A(net2648),
    .B(net6350));
 sg13g2_o21ai_1 _16814_ (.B1(_07171_),
    .Y(_01057_),
    .A1(net7357),
    .A2(net6350));
 sg13g2_nand2_1 _16815_ (.Y(_07172_),
    .A(net3141),
    .B(net6351));
 sg13g2_o21ai_1 _16816_ (.B1(_07172_),
    .Y(_01058_),
    .A1(net7554),
    .A2(net6351));
 sg13g2_nand2_1 _16817_ (.Y(_07173_),
    .A(net3360),
    .B(net6350));
 sg13g2_o21ai_1 _16818_ (.B1(_07173_),
    .Y(_01059_),
    .A1(net7714),
    .A2(net6350));
 sg13g2_nand3_1 _16819_ (.B(net7100),
    .C(net7216),
    .A(net7282),
    .Y(_07174_));
 sg13g2_nand2_1 _16820_ (.Y(_07175_),
    .A(net4046),
    .B(net6349));
 sg13g2_o21ai_1 _16821_ (.B1(_07175_),
    .Y(_01060_),
    .A1(net7343),
    .A2(net6349));
 sg13g2_nand2_1 _16822_ (.Y(_07176_),
    .A(net3834),
    .B(net6349));
 sg13g2_o21ai_1 _16823_ (.B1(_07176_),
    .Y(_01061_),
    .A1(net7541),
    .A2(net6348));
 sg13g2_nand2_1 _16824_ (.Y(_07177_),
    .A(net4267),
    .B(net6348));
 sg13g2_o21ai_1 _16825_ (.B1(_07177_),
    .Y(_01062_),
    .A1(net7686),
    .A2(net6348));
 sg13g2_nand3_1 _16826_ (.B(net7100),
    .C(net7216),
    .A(net7362),
    .Y(_07178_));
 sg13g2_nand2_1 _16827_ (.Y(_07179_),
    .A(net3114),
    .B(net6347));
 sg13g2_o21ai_1 _16828_ (.B1(_07179_),
    .Y(_01063_),
    .A1(net7343),
    .A2(net6347));
 sg13g2_nand2_1 _16829_ (.Y(_07180_),
    .A(net3170),
    .B(net6347));
 sg13g2_o21ai_1 _16830_ (.B1(_07180_),
    .Y(_01064_),
    .A1(net7541),
    .A2(net6346));
 sg13g2_nand2_1 _16831_ (.Y(_07181_),
    .A(net2881),
    .B(net6346));
 sg13g2_o21ai_1 _16832_ (.B1(_07181_),
    .Y(_01065_),
    .A1(net7686),
    .A2(net6346));
 sg13g2_nor3_2 _16833_ (.A(net7107),
    .B(net7097),
    .C(net7202),
    .Y(_07182_));
 sg13g2_nor2_1 _16834_ (.A(net4201),
    .B(net6345),
    .Y(_07183_));
 sg13g2_a21oi_1 _16835_ (.A1(net7343),
    .A2(net6345),
    .Y(_01066_),
    .B1(_07183_));
 sg13g2_nor2_1 _16836_ (.A(net3921),
    .B(net6345),
    .Y(_07184_));
 sg13g2_a21oi_1 _16837_ (.A1(net7541),
    .A2(net6345),
    .Y(_01067_),
    .B1(_07184_));
 sg13g2_nor2_1 _16838_ (.A(net4627),
    .B(net6344),
    .Y(_07185_));
 sg13g2_a21oi_1 _16839_ (.A1(net7686),
    .A2(net6344),
    .Y(_01068_),
    .B1(_07185_));
 sg13g2_nor3_2 _16840_ (.A(net7267),
    .B(net7246),
    .C(net7200),
    .Y(_07186_));
 sg13g2_nor2_1 _16841_ (.A(net4175),
    .B(net6818),
    .Y(_07187_));
 sg13g2_a21oi_1 _16842_ (.A1(net7311),
    .A2(net6818),
    .Y(_01069_),
    .B1(_07187_));
 sg13g2_nor2_1 _16843_ (.A(net4237),
    .B(net6818),
    .Y(_07188_));
 sg13g2_a21oi_1 _16844_ (.A1(net7509),
    .A2(net6818),
    .Y(_01070_),
    .B1(_07188_));
 sg13g2_nor2_1 _16845_ (.A(net4834),
    .B(net6817),
    .Y(_07189_));
 sg13g2_a21oi_1 _16846_ (.A1(net7666),
    .A2(net6817),
    .Y(_01071_),
    .B1(_07189_));
 sg13g2_nand3_1 _16847_ (.B(net7240),
    .C(net7213),
    .A(net7066),
    .Y(_07190_));
 sg13g2_nand2_1 _16848_ (.Y(_07191_),
    .A(net3073),
    .B(net6342));
 sg13g2_o21ai_1 _16849_ (.B1(_07191_),
    .Y(_01072_),
    .A1(net7337),
    .A2(net6342));
 sg13g2_nand2_1 _16850_ (.Y(_07192_),
    .A(net3102),
    .B(net6343));
 sg13g2_o21ai_1 _16851_ (.B1(_07192_),
    .Y(_01073_),
    .A1(net7534),
    .A2(net6342));
 sg13g2_nand2_1 _16852_ (.Y(_07193_),
    .A(net4271),
    .B(net6342));
 sg13g2_o21ai_1 _16853_ (.B1(_07193_),
    .Y(_01074_),
    .A1(net7690),
    .A2(net6342));
 sg13g2_nand3_1 _16854_ (.B(net7240),
    .C(net7213),
    .A(net7102),
    .Y(_07194_));
 sg13g2_nand2_1 _16855_ (.Y(_07195_),
    .A(net3745),
    .B(net6340));
 sg13g2_o21ai_1 _16856_ (.B1(_07195_),
    .Y(_01075_),
    .A1(net7336),
    .A2(net6340));
 sg13g2_nand2_1 _16857_ (.Y(_07196_),
    .A(net2690),
    .B(net6341));
 sg13g2_o21ai_1 _16858_ (.B1(_07196_),
    .Y(_01076_),
    .A1(net7534),
    .A2(net6340));
 sg13g2_nand2_1 _16859_ (.Y(_07197_),
    .A(net4221),
    .B(net6340));
 sg13g2_o21ai_1 _16860_ (.B1(_07197_),
    .Y(_01077_),
    .A1(net7690),
    .A2(net6340));
 sg13g2_nand3_1 _16861_ (.B(net7240),
    .C(net7227),
    .A(net7083),
    .Y(_07198_));
 sg13g2_nand2_1 _16862_ (.Y(_07199_),
    .A(net2995),
    .B(net6338));
 sg13g2_o21ai_1 _16863_ (.B1(_07199_),
    .Y(_01078_),
    .A1(net7336),
    .A2(net6338));
 sg13g2_nand2_1 _16864_ (.Y(_07200_),
    .A(net3837),
    .B(net6339));
 sg13g2_o21ai_1 _16865_ (.B1(_07200_),
    .Y(_01079_),
    .A1(net7534),
    .A2(net6338));
 sg13g2_nand2_1 _16866_ (.Y(_07201_),
    .A(net3329),
    .B(net6338));
 sg13g2_o21ai_1 _16867_ (.B1(_07201_),
    .Y(_01080_),
    .A1(net7690),
    .A2(net6338));
 sg13g2_nor2_1 _16868_ (.A(net7559),
    .B(_03995_),
    .Y(_01081_));
 sg13g2_o21ai_1 _16869_ (.B1(net4625),
    .Y(_07202_),
    .A1(\top1.mem_ctl.state_reg[1] ),
    .A2(_03991_));
 sg13g2_inv_1 _16870_ (.Y(_01082_),
    .A(net4626));
 sg13g2_nand3_1 _16871_ (.B(net7083),
    .C(net7226),
    .A(net7101),
    .Y(_07203_));
 sg13g2_nand2_1 _16872_ (.Y(_07204_),
    .A(net3300),
    .B(net6336));
 sg13g2_o21ai_1 _16873_ (.B1(_07204_),
    .Y(_01083_),
    .A1(net7354),
    .A2(net6336));
 sg13g2_nand2_1 _16874_ (.Y(_07205_),
    .A(net2645),
    .B(net6336));
 sg13g2_o21ai_1 _16875_ (.B1(_07205_),
    .Y(_01084_),
    .A1(net7551),
    .A2(net6336));
 sg13g2_nand2_1 _16876_ (.Y(_07206_),
    .A(net2947),
    .B(net6337));
 sg13g2_o21ai_1 _16877_ (.B1(_07206_),
    .Y(_01085_),
    .A1(net7709),
    .A2(net6337));
 sg13g2_nand3_1 _16878_ (.B(net7101),
    .C(net7226),
    .A(net7102),
    .Y(_07207_));
 sg13g2_nand2_1 _16879_ (.Y(_07208_),
    .A(net3392),
    .B(net6334));
 sg13g2_o21ai_1 _16880_ (.B1(_07208_),
    .Y(_01086_),
    .A1(net7354),
    .A2(net6334));
 sg13g2_nand2_1 _16881_ (.Y(_07209_),
    .A(net3304),
    .B(net6334));
 sg13g2_o21ai_1 _16882_ (.B1(_07209_),
    .Y(_01087_),
    .A1(net7551),
    .A2(net6334));
 sg13g2_nand2_1 _16883_ (.Y(_07210_),
    .A(net3653),
    .B(net6335));
 sg13g2_o21ai_1 _16884_ (.B1(_07210_),
    .Y(_01088_),
    .A1(net7709),
    .A2(net6335));
 sg13g2_nand3_1 _16885_ (.B(net7100),
    .C(net7220),
    .A(net7405),
    .Y(_07211_));
 sg13g2_nand2_1 _16886_ (.Y(_07212_),
    .A(net2737),
    .B(net6332));
 sg13g2_o21ai_1 _16887_ (.B1(_07212_),
    .Y(_01089_),
    .A1(net7343),
    .A2(net6332));
 sg13g2_nand2_1 _16888_ (.Y(_07213_),
    .A(net3607),
    .B(net6332));
 sg13g2_o21ai_1 _16889_ (.B1(_07213_),
    .Y(_01090_),
    .A1(net7542),
    .A2(net6332));
 sg13g2_nand2_1 _16890_ (.Y(_07214_),
    .A(net2684),
    .B(net6332));
 sg13g2_o21ai_1 _16891_ (.B1(_07214_),
    .Y(_01091_),
    .A1(net7702),
    .A2(net6332));
 sg13g2_nand3_1 _16892_ (.B(net7238),
    .C(net7220),
    .A(net7100),
    .Y(_07215_));
 sg13g2_nand2_1 _16893_ (.Y(_07216_),
    .A(net3620),
    .B(net6330));
 sg13g2_o21ai_1 _16894_ (.B1(_07216_),
    .Y(_01092_),
    .A1(net7343),
    .A2(net6330));
 sg13g2_nand2_1 _16895_ (.Y(_07217_),
    .A(net3672),
    .B(net6330));
 sg13g2_o21ai_1 _16896_ (.B1(_07217_),
    .Y(_01093_),
    .A1(net7541),
    .A2(net6330));
 sg13g2_nand2_1 _16897_ (.Y(_07218_),
    .A(net3161),
    .B(net6330));
 sg13g2_o21ai_1 _16898_ (.B1(_07218_),
    .Y(_01094_),
    .A1(net7702),
    .A2(net6330));
 sg13g2_nor3_1 _16899_ (.A(_04101_),
    .B(net7267),
    .C(net7199),
    .Y(_07219_));
 sg13g2_nor2_1 _16900_ (.A(net4699),
    .B(net6816),
    .Y(_07220_));
 sg13g2_a21oi_1 _16901_ (.A1(net7309),
    .A2(net6816),
    .Y(_01095_),
    .B1(_07220_));
 sg13g2_nor2_1 _16902_ (.A(net4592),
    .B(net6815),
    .Y(_07221_));
 sg13g2_a21oi_1 _16903_ (.A1(net7511),
    .A2(net6815),
    .Y(_01096_),
    .B1(_07221_));
 sg13g2_nor2_1 _16904_ (.A(net3828),
    .B(net6815),
    .Y(_07222_));
 sg13g2_a21oi_1 _16905_ (.A1(net7666),
    .A2(net6815),
    .Y(_01097_),
    .B1(_07222_));
 sg13g2_nand3_1 _16906_ (.B(net7235),
    .C(net7220),
    .A(net7100),
    .Y(_07223_));
 sg13g2_nand2_1 _16907_ (.Y(_07224_),
    .A(net3316),
    .B(net6328));
 sg13g2_o21ai_1 _16908_ (.B1(_07224_),
    .Y(_01098_),
    .A1(net7343),
    .A2(net6328));
 sg13g2_nand2_1 _16909_ (.Y(_07225_),
    .A(net3124),
    .B(net6328));
 sg13g2_o21ai_1 _16910_ (.B1(_07225_),
    .Y(_01099_),
    .A1(net7541),
    .A2(net6328));
 sg13g2_nand2_1 _16911_ (.Y(_07226_),
    .A(net2844),
    .B(net6328));
 sg13g2_o21ai_1 _16912_ (.B1(_07226_),
    .Y(_01100_),
    .A1(net7702),
    .A2(net6328));
 sg13g2_nand3_1 _16913_ (.B(net7066),
    .C(net7226),
    .A(net7100),
    .Y(_07227_));
 sg13g2_nand2_1 _16914_ (.Y(_07228_),
    .A(net3695),
    .B(net6326));
 sg13g2_o21ai_1 _16915_ (.B1(_07228_),
    .Y(_01101_),
    .A1(net7354),
    .A2(net6326));
 sg13g2_nand2_1 _16916_ (.Y(_07229_),
    .A(net3704),
    .B(net6326));
 sg13g2_o21ai_1 _16917_ (.B1(_07229_),
    .Y(_01102_),
    .A1(net7551),
    .A2(net6326));
 sg13g2_nand2_1 _16918_ (.Y(_07230_),
    .A(net3874),
    .B(net6327));
 sg13g2_o21ai_1 _16919_ (.B1(_07230_),
    .Y(_01103_),
    .A1(net7709),
    .A2(net6327));
 sg13g2_nand3_1 _16920_ (.B(net7247),
    .C(net7218),
    .A(net7117),
    .Y(_07231_));
 sg13g2_nand2_1 _16921_ (.Y(_07232_),
    .A(net3639),
    .B(net6325));
 sg13g2_o21ai_1 _16922_ (.B1(_07232_),
    .Y(_01104_),
    .A1(net7348),
    .A2(net6325));
 sg13g2_nand2_1 _16923_ (.Y(_07233_),
    .A(net2592),
    .B(net6324));
 sg13g2_o21ai_1 _16924_ (.B1(_07233_),
    .Y(_01105_),
    .A1(net7545),
    .A2(net6324));
 sg13g2_nand2_1 _16925_ (.Y(_07234_),
    .A(net4306),
    .B(net6325));
 sg13g2_o21ai_1 _16926_ (.B1(_07234_),
    .Y(_01106_),
    .A1(net7705),
    .A2(net6325));
 sg13g2_nand3_1 _16927_ (.B(net7277),
    .C(net7218),
    .A(net7117),
    .Y(_07235_));
 sg13g2_nand2_1 _16928_ (.Y(_07236_),
    .A(net3042),
    .B(net6323));
 sg13g2_o21ai_1 _16929_ (.B1(_07236_),
    .Y(_01107_),
    .A1(net7348),
    .A2(net6323));
 sg13g2_nand2_1 _16930_ (.Y(_07237_),
    .A(net3409),
    .B(net6322));
 sg13g2_o21ai_1 _16931_ (.B1(_07237_),
    .Y(_01108_),
    .A1(net7545),
    .A2(net6322));
 sg13g2_nand2_1 _16932_ (.Y(_07238_),
    .A(net2771),
    .B(net6323));
 sg13g2_o21ai_1 _16933_ (.B1(_07238_),
    .Y(_01109_),
    .A1(net7705),
    .A2(net6323));
 sg13g2_nor3_2 _16934_ (.A(net7098),
    .B(_04291_),
    .C(net7202),
    .Y(_07239_));
 sg13g2_nor2_1 _16935_ (.A(net4641),
    .B(net6320),
    .Y(_07240_));
 sg13g2_a21oi_1 _16936_ (.A1(net7354),
    .A2(net6320),
    .Y(_01110_),
    .B1(_07240_));
 sg13g2_nor2_1 _16937_ (.A(net4674),
    .B(net6320),
    .Y(_07241_));
 sg13g2_a21oi_1 _16938_ (.A1(net7551),
    .A2(net6320),
    .Y(_01111_),
    .B1(_07241_));
 sg13g2_nor2_1 _16939_ (.A(net4574),
    .B(net6321),
    .Y(_07242_));
 sg13g2_a21oi_1 _16940_ (.A1(net7709),
    .A2(net6321),
    .Y(_01112_),
    .B1(_07242_));
 sg13g2_nand3_1 _16941_ (.B(net7100),
    .C(net7216),
    .A(net7408),
    .Y(_07243_));
 sg13g2_nand2_1 _16942_ (.Y(_07244_),
    .A(net2625),
    .B(net6319));
 sg13g2_o21ai_1 _16943_ (.B1(_07244_),
    .Y(_01113_),
    .A1(net7343),
    .A2(net6319));
 sg13g2_nand2_1 _16944_ (.Y(_07245_),
    .A(net3699),
    .B(net6319));
 sg13g2_o21ai_1 _16945_ (.B1(_07245_),
    .Y(_01114_),
    .A1(net7541),
    .A2(net6318));
 sg13g2_nand2_1 _16946_ (.Y(_07246_),
    .A(net3117),
    .B(net6318));
 sg13g2_o21ai_1 _16947_ (.B1(_07246_),
    .Y(_01115_),
    .A1(net7686),
    .A2(net6318));
 sg13g2_nand3_1 _16948_ (.B(net7102),
    .C(net7217),
    .A(net7116),
    .Y(_07247_));
 sg13g2_nand2_1 _16949_ (.Y(_07248_),
    .A(net2957),
    .B(net6317));
 sg13g2_o21ai_1 _16950_ (.B1(_07248_),
    .Y(_01116_),
    .A1(net7347),
    .A2(net6317));
 sg13g2_nand2_1 _16951_ (.Y(_07249_),
    .A(net3923),
    .B(net6316));
 sg13g2_o21ai_1 _16952_ (.B1(_07249_),
    .Y(_01117_),
    .A1(net7544),
    .A2(net6316));
 sg13g2_nand2_1 _16953_ (.Y(_07250_),
    .A(net3550),
    .B(net6316));
 sg13g2_o21ai_1 _16954_ (.B1(_07250_),
    .Y(_01118_),
    .A1(net7703),
    .A2(net6316));
 sg13g2_nand3_1 _16955_ (.B(net7083),
    .C(net7217),
    .A(net7116),
    .Y(_07251_));
 sg13g2_nand2_1 _16956_ (.Y(_07252_),
    .A(net3136),
    .B(net6315));
 sg13g2_o21ai_1 _16957_ (.B1(_07252_),
    .Y(_01119_),
    .A1(net7347),
    .A2(net6315));
 sg13g2_nand2_1 _16958_ (.Y(_07253_),
    .A(net2785),
    .B(net6314));
 sg13g2_o21ai_1 _16959_ (.B1(_07253_),
    .Y(_01120_),
    .A1(net7544),
    .A2(net6314));
 sg13g2_nand2_1 _16960_ (.Y(_07254_),
    .A(net3065),
    .B(net6314));
 sg13g2_o21ai_1 _16961_ (.B1(_07254_),
    .Y(_01121_),
    .A1(net7703),
    .A2(net6314));
 sg13g2_nand3_1 _16962_ (.B(net7042),
    .C(net7217),
    .A(net7116),
    .Y(_07255_));
 sg13g2_nand2_1 _16963_ (.Y(_07256_),
    .A(net2582),
    .B(net6313));
 sg13g2_o21ai_1 _16964_ (.B1(_07256_),
    .Y(_01122_),
    .A1(net7347),
    .A2(net6313));
 sg13g2_nand2_1 _16965_ (.Y(_07257_),
    .A(net3019),
    .B(net6312));
 sg13g2_o21ai_1 _16966_ (.B1(_07257_),
    .Y(_01123_),
    .A1(net7544),
    .A2(net6312));
 sg13g2_nand2_1 _16967_ (.Y(_07258_),
    .A(net2789),
    .B(net6312));
 sg13g2_o21ai_1 _16968_ (.B1(_07258_),
    .Y(_01124_),
    .A1(net7703),
    .A2(net6312));
 sg13g2_nand3_1 _16969_ (.B(net7065),
    .C(net7211),
    .A(_04129_),
    .Y(_07259_));
 sg13g2_nand2_1 _16970_ (.Y(_07260_),
    .A(net3450),
    .B(net6311));
 sg13g2_o21ai_1 _16971_ (.B1(_07260_),
    .Y(_01125_),
    .A1(net7309),
    .A2(net6311));
 sg13g2_nand2_1 _16972_ (.Y(_07261_),
    .A(net3361),
    .B(net6311));
 sg13g2_o21ai_1 _16973_ (.B1(_07261_),
    .Y(_01126_),
    .A1(net7511),
    .A2(net6310));
 sg13g2_nand2_1 _16974_ (.Y(_07262_),
    .A(net2669),
    .B(net6310));
 sg13g2_o21ai_1 _16975_ (.B1(_07262_),
    .Y(_01127_),
    .A1(net7666),
    .A2(net6310));
 sg13g2_nand3_1 _16976_ (.B(net7273),
    .C(net7218),
    .A(net7117),
    .Y(_07263_));
 sg13g2_nand2_1 _16977_ (.Y(_07264_),
    .A(net3011),
    .B(net6309));
 sg13g2_o21ai_1 _16978_ (.B1(_07264_),
    .Y(_01128_),
    .A1(net7348),
    .A2(net6309));
 sg13g2_nand2_1 _16979_ (.Y(_07265_),
    .A(net3384),
    .B(net6308));
 sg13g2_o21ai_1 _16980_ (.B1(_07265_),
    .Y(_01129_),
    .A1(net7545),
    .A2(net6308));
 sg13g2_nand2_1 _16981_ (.Y(_07266_),
    .A(net3742),
    .B(net6309));
 sg13g2_o21ai_1 _16982_ (.B1(_07266_),
    .Y(_01130_),
    .A1(net7705),
    .A2(net6309));
 sg13g2_nand3_1 _16983_ (.B(net7081),
    .C(net7209),
    .A(net7361),
    .Y(_07267_));
 sg13g2_nand2_1 _16984_ (.Y(_07268_),
    .A(net2677),
    .B(net6306));
 sg13g2_o21ai_1 _16985_ (.B1(_07268_),
    .Y(_01131_),
    .A1(net7325),
    .A2(net6306));
 sg13g2_nand2_1 _16986_ (.Y(_07269_),
    .A(net2519),
    .B(net6306));
 sg13g2_o21ai_1 _16987_ (.B1(_07269_),
    .Y(_01132_),
    .A1(net7524),
    .A2(net6306));
 sg13g2_nand2_1 _16988_ (.Y(_07270_),
    .A(net2492),
    .B(net6306));
 sg13g2_o21ai_1 _16989_ (.B1(_07270_),
    .Y(_01133_),
    .A1(net7681),
    .A2(net6306));
 sg13g2_nor3_1 _16990_ (.A(net7272),
    .B(_04154_),
    .C(net7201),
    .Y(_07271_));
 sg13g2_nor2_1 _16991_ (.A(net4293),
    .B(net6814),
    .Y(_07272_));
 sg13g2_a21oi_1 _16992_ (.A1(net7310),
    .A2(net6814),
    .Y(_01134_),
    .B1(_07272_));
 sg13g2_nor2_1 _16993_ (.A(net4821),
    .B(net6813),
    .Y(_07273_));
 sg13g2_a21oi_1 _16994_ (.A1(net7509),
    .A2(net6813),
    .Y(_01135_),
    .B1(_07273_));
 sg13g2_nor2_1 _16995_ (.A(net4531),
    .B(net6814),
    .Y(_07274_));
 sg13g2_a21oi_1 _16996_ (.A1(net7668),
    .A2(net6814),
    .Y(_01136_),
    .B1(_07274_));
 sg13g2_nor3_1 _16997_ (.A(net7276),
    .B(_04154_),
    .C(net7200),
    .Y(_07275_));
 sg13g2_nor2_1 _16998_ (.A(net4382),
    .B(net6812),
    .Y(_07276_));
 sg13g2_a21oi_1 _16999_ (.A1(net7310),
    .A2(net6812),
    .Y(_01137_),
    .B1(_07276_));
 sg13g2_nor2_1 _17000_ (.A(net4193),
    .B(net6811),
    .Y(_07277_));
 sg13g2_a21oi_1 _17001_ (.A1(net7509),
    .A2(net6811),
    .Y(_01138_),
    .B1(_07277_));
 sg13g2_nor2_1 _17002_ (.A(net4546),
    .B(net6812),
    .Y(_07278_));
 sg13g2_a21oi_1 _17003_ (.A1(net7668),
    .A2(net6812),
    .Y(_01139_),
    .B1(_07278_));
 sg13g2_nor2_2 _17004_ (.A(_03962_),
    .B(_03971_),
    .Y(_07279_));
 sg13g2_a21oi_1 _17005_ (.A1(net6110),
    .A2(_00063_),
    .Y(_07280_),
    .B1(_03971_));
 sg13g2_o21ai_1 _17006_ (.B1(_03966_),
    .Y(_07281_),
    .A1(\top1.fsm.state_reg[2] ),
    .A2(_03967_));
 sg13g2_o21ai_1 _17007_ (.B1(\top1.fsm.sending_data ),
    .Y(_07282_),
    .A1(_03949_),
    .A2(_07281_));
 sg13g2_o21ai_1 _17008_ (.B1(_07282_),
    .Y(_01140_),
    .A1(_03949_),
    .A2(_07280_));
 sg13g2_nor2_1 _17009_ (.A(\top1.fsm.sending_pending ),
    .B(_03987_),
    .Y(_07283_));
 sg13g2_nor2_1 _17010_ (.A(_03972_),
    .B(_07283_),
    .Y(_07284_));
 sg13g2_nor2_1 _17011_ (.A(\top1.fsm.state_reg[2] ),
    .B(_00063_),
    .Y(_07285_));
 sg13g2_a21o_1 _17012_ (.A2(_07285_),
    .A1(_03958_),
    .B1(_03953_),
    .X(_07286_));
 sg13g2_a21oi_1 _17013_ (.A1(_03955_),
    .A2(_07286_),
    .Y(_07287_),
    .B1(_07284_));
 sg13g2_o21ai_1 _17014_ (.B1(_07287_),
    .Y(_07288_),
    .A1(\top1.fsm.sending_pending ),
    .A2(net7560));
 sg13g2_inv_1 _17015_ (.Y(_01141_),
    .A(_07288_));
 sg13g2_nor3_1 _17016_ (.A(_04154_),
    .B(net7246),
    .C(net7200),
    .Y(_07289_));
 sg13g2_nor2_1 _17017_ (.A(net4215),
    .B(net6809),
    .Y(_07290_));
 sg13g2_a21oi_1 _17018_ (.A1(net7310),
    .A2(net6809),
    .Y(_01142_),
    .B1(_07290_));
 sg13g2_nor2_1 _17019_ (.A(net4064),
    .B(net6809),
    .Y(_07291_));
 sg13g2_a21oi_1 _17020_ (.A1(net7509),
    .A2(net6809),
    .Y(_01143_),
    .B1(_07291_));
 sg13g2_nor2_1 _17021_ (.A(net4226),
    .B(net6810),
    .Y(_07292_));
 sg13g2_a21oi_1 _17022_ (.A1(net7668),
    .A2(net6809),
    .Y(_01144_),
    .B1(_07292_));
 sg13g2_nand2b_1 _17023_ (.Y(_07293_),
    .B(_07287_),
    .A_N(_03960_));
 sg13g2_a22oi_1 _17024_ (.Y(_01145_),
    .B1(_07293_),
    .B2(_03833_),
    .A2(_07287_),
    .A1(net7560));
 sg13g2_nand3b_1 _17025_ (.B(_03972_),
    .C(_03952_),
    .Y(_07294_),
    .A_N(_04017_));
 sg13g2_nand4_1 _17026_ (.B(\top1.fsm.cpt[2] ),
    .C(\top1.fsm.cpt[3] ),
    .A(\top1.fsm.cpt[4] ),
    .Y(_07295_),
    .D(_03943_));
 sg13g2_a21oi_1 _17027_ (.A1(_03953_),
    .A2(_07295_),
    .Y(_07296_),
    .B1(_03946_));
 sg13g2_o21ai_1 _17028_ (.B1(_07296_),
    .Y(_07297_),
    .A1(_03962_),
    .A2(_07294_));
 sg13g2_nor3_1 _17029_ (.A(_03942_),
    .B(_03947_),
    .C(net5931),
    .Y(_07298_));
 sg13g2_nand4_1 _17030_ (.B(_03980_),
    .C(net6019),
    .A(\top1.fsm.state_reg[0] ),
    .Y(_07299_),
    .D(_07298_));
 sg13g2_nand3_1 _17031_ (.B(_03941_),
    .C(_04025_),
    .A(\top1.fsm.sending_pending ),
    .Y(_07300_));
 sg13g2_nor2_1 _17032_ (.A(\top1.fsm.cpt[4] ),
    .B(_07300_),
    .Y(_07301_));
 sg13g2_nor2_1 _17033_ (.A(_00065_),
    .B(_07301_),
    .Y(_07302_));
 sg13g2_or2_1 _17034_ (.X(_07303_),
    .B(_07302_),
    .A(_03985_));
 sg13g2_a22oi_1 _17035_ (.Y(_07304_),
    .B1(_07303_),
    .B2(_03968_),
    .A2(_07299_),
    .A1(_03951_));
 sg13g2_a21oi_1 _17036_ (.A1(_03992_),
    .A2(_07304_),
    .Y(_07305_),
    .B1(_07297_));
 sg13g2_a21o_1 _17037_ (.A2(_07297_),
    .A1(\top1.fsm.re ),
    .B1(_07305_),
    .X(_01146_));
 sg13g2_nand3_1 _17038_ (.B(net7074),
    .C(net7222),
    .A(net7362),
    .Y(_07306_));
 sg13g2_nand2_1 _17039_ (.Y(_07307_),
    .A(net3111),
    .B(net6304));
 sg13g2_o21ai_1 _17040_ (.B1(_07307_),
    .Y(_01147_),
    .A1(net7358),
    .A2(net6304));
 sg13g2_nand2_1 _17041_ (.Y(_07308_),
    .A(net3997),
    .B(net6304));
 sg13g2_o21ai_1 _17042_ (.B1(_07308_),
    .Y(_01148_),
    .A1(net7555),
    .A2(net6304));
 sg13g2_nand2_1 _17043_ (.Y(_07309_),
    .A(net3931),
    .B(net6305));
 sg13g2_o21ai_1 _17044_ (.B1(_07309_),
    .Y(_01149_),
    .A1(net7715),
    .A2(net6304));
 sg13g2_nand3_1 _17045_ (.B(net7081),
    .C(net7209),
    .A(net7280),
    .Y(_07310_));
 sg13g2_nand2_1 _17046_ (.Y(_07311_),
    .A(net2612),
    .B(net6302));
 sg13g2_o21ai_1 _17047_ (.B1(_07311_),
    .Y(_01150_),
    .A1(net7325),
    .A2(net6302));
 sg13g2_nand2_1 _17048_ (.Y(_07312_),
    .A(net2954),
    .B(net6302));
 sg13g2_o21ai_1 _17049_ (.B1(_07312_),
    .Y(_01151_),
    .A1(net7524),
    .A2(net6302));
 sg13g2_nand2_1 _17050_ (.Y(_07313_),
    .A(net3168),
    .B(net6302));
 sg13g2_o21ai_1 _17051_ (.B1(_07313_),
    .Y(_01152_),
    .A1(net7681),
    .A2(net6302));
 sg13g2_nor3_1 _17052_ (.A(net7107),
    .B(net7250),
    .C(net7197),
    .Y(_07314_));
 sg13g2_nor2_1 _17053_ (.A(net4394),
    .B(net6301),
    .Y(_07315_));
 sg13g2_a21oi_1 _17054_ (.A1(net7301),
    .A2(net6301),
    .Y(_01153_),
    .B1(_07315_));
 sg13g2_nor2_1 _17055_ (.A(net4169),
    .B(net6300),
    .Y(_07316_));
 sg13g2_a21oi_1 _17056_ (.A1(net7496),
    .A2(net6300),
    .Y(_01154_),
    .B1(_07316_));
 sg13g2_nor2_1 _17057_ (.A(net4542),
    .B(net6301),
    .Y(_07317_));
 sg13g2_a21oi_1 _17058_ (.A1(net7656),
    .A2(net6300),
    .Y(_01155_),
    .B1(_07317_));
 sg13g2_o21ai_1 _17059_ (.B1(_03968_),
    .Y(_07318_),
    .A1(_03944_),
    .A2(_03985_));
 sg13g2_a221oi_1 _17060_ (.B2(\top1.fsm.state_reg[1] ),
    .C1(_03962_),
    .B1(_03965_),
    .A1(net6110),
    .Y(_07319_),
    .A2(_00067_));
 sg13g2_nand4_1 _17061_ (.B(_03952_),
    .C(_03969_),
    .A(_03945_),
    .Y(_07320_),
    .D(_07319_));
 sg13g2_nand3b_1 _17062_ (.B(_07318_),
    .C(_07320_),
    .Y(_07321_),
    .A_N(_03949_));
 sg13g2_or2_2 _17063_ (.X(_07322_),
    .B(net5824),
    .A(_07279_));
 sg13g2_nand2_1 _17064_ (.Y(_07323_),
    .A(net6215),
    .B(net5824));
 sg13g2_o21ai_1 _17065_ (.B1(_07323_),
    .Y(_01156_),
    .A1(net6215),
    .A2(_07322_));
 sg13g2_nor3_1 _17066_ (.A(net6059),
    .B(net5954),
    .C(_07322_),
    .Y(_07324_));
 sg13g2_a21o_1 _17067_ (.A2(net5824),
    .A1(net6150),
    .B1(_07324_),
    .X(_01157_));
 sg13g2_nand2_1 _17068_ (.Y(_07325_),
    .A(net6128),
    .B(net5824));
 sg13g2_nor2_1 _17069_ (.A(_00073_),
    .B(net5935),
    .Y(_07326_));
 sg13g2_xnor2_1 _17070_ (.Y(_07327_),
    .A(_00073_),
    .B(net5935));
 sg13g2_o21ai_1 _17071_ (.B1(_07325_),
    .Y(_01158_),
    .A1(_07322_),
    .A2(_07327_));
 sg13g2_nand2_1 _17072_ (.Y(_07328_),
    .A(\top1.addr_out[3] ),
    .B(net5824));
 sg13g2_xor2_1 _17073_ (.B(_07326_),
    .A(_00072_),
    .X(_07329_));
 sg13g2_o21ai_1 _17074_ (.B1(_07328_),
    .Y(_01159_),
    .A1(_07322_),
    .A2(_07329_));
 sg13g2_nand2_1 _17075_ (.Y(_07330_),
    .A(net6123),
    .B(_07321_));
 sg13g2_nor3_1 _17076_ (.A(_00071_),
    .B(net5935),
    .C(net5843),
    .Y(_07331_));
 sg13g2_o21ai_1 _17077_ (.B1(_00071_),
    .Y(_07332_),
    .A1(net5935),
    .A2(net5843));
 sg13g2_nand2b_1 _17078_ (.Y(_07333_),
    .B(_07332_),
    .A_N(_07331_));
 sg13g2_o21ai_1 _17079_ (.B1(_07330_),
    .Y(_01160_),
    .A1(_07322_),
    .A2(_07333_));
 sg13g2_nand2_1 _17080_ (.Y(_07334_),
    .A(net6117),
    .B(net5824));
 sg13g2_xor2_1 _17081_ (.B(_07331_),
    .A(_00070_),
    .X(_07335_));
 sg13g2_o21ai_1 _17082_ (.B1(_07334_),
    .Y(_01161_),
    .A1(_07322_),
    .A2(_07335_));
 sg13g2_nand2_1 _17083_ (.Y(_07336_),
    .A(net6113),
    .B(net5824));
 sg13g2_nand3_1 _17084_ (.B(net5854),
    .C(_05452_),
    .A(net5955),
    .Y(_07337_));
 sg13g2_nor2_1 _17085_ (.A(_00069_),
    .B(_07337_),
    .Y(_07338_));
 sg13g2_xnor2_1 _17086_ (.Y(_07339_),
    .A(_00069_),
    .B(_07337_));
 sg13g2_o21ai_1 _17087_ (.B1(_07336_),
    .Y(_01162_),
    .A1(_07322_),
    .A2(_07339_));
 sg13g2_nand2_1 _17088_ (.Y(_07340_),
    .A(net6112),
    .B(net5824));
 sg13g2_xor2_1 _17089_ (.B(_07338_),
    .A(_00068_),
    .X(_07341_));
 sg13g2_o21ai_1 _17090_ (.B1(_07340_),
    .Y(_01163_),
    .A1(_07322_),
    .A2(_07341_));
 sg13g2_nand3_1 _17091_ (.B(net7079),
    .C(net7208),
    .A(net7285),
    .Y(_07342_));
 sg13g2_nand2_1 _17092_ (.Y(_07343_),
    .A(net3072),
    .B(net6299));
 sg13g2_o21ai_1 _17093_ (.B1(_07343_),
    .Y(_01164_),
    .A1(net7309),
    .A2(net6299));
 sg13g2_nand2_1 _17094_ (.Y(_07344_),
    .A(net4211),
    .B(net6298));
 sg13g2_o21ai_1 _17095_ (.B1(_07344_),
    .Y(_01165_),
    .A1(net7509),
    .A2(net6298));
 sg13g2_nand2_1 _17096_ (.Y(_07345_),
    .A(net3051),
    .B(net6299));
 sg13g2_o21ai_1 _17097_ (.B1(_07345_),
    .Y(_01166_),
    .A1(net7668),
    .A2(net6299));
 sg13g2_nand3_1 _17098_ (.B(net7235),
    .C(net7218),
    .A(net7117),
    .Y(_07346_));
 sg13g2_nand2_1 _17099_ (.Y(_07347_),
    .A(net2657),
    .B(net6296));
 sg13g2_o21ai_1 _17100_ (.B1(_07347_),
    .Y(_01167_),
    .A1(net7348),
    .A2(net6296));
 sg13g2_nand2_1 _17101_ (.Y(_07348_),
    .A(net3177),
    .B(net6296));
 sg13g2_o21ai_1 _17102_ (.B1(_07348_),
    .Y(_01168_),
    .A1(net7547),
    .A2(net6296));
 sg13g2_nand2_1 _17103_ (.Y(_07349_),
    .A(net3338),
    .B(net6297));
 sg13g2_o21ai_1 _17104_ (.B1(_07349_),
    .Y(_01169_),
    .A1(net7705),
    .A2(net6297));
 sg13g2_nand3_1 _17105_ (.B(net7247),
    .C(net7222),
    .A(net7075),
    .Y(_07350_));
 sg13g2_nand2_1 _17106_ (.Y(_07351_),
    .A(net2784),
    .B(net6295));
 sg13g2_o21ai_1 _17107_ (.B1(_07351_),
    .Y(_01170_),
    .A1(net7357),
    .A2(net6294));
 sg13g2_nand2_1 _17108_ (.Y(_07352_),
    .A(net2730),
    .B(net6295));
 sg13g2_o21ai_1 _17109_ (.B1(_07352_),
    .Y(_01171_),
    .A1(net7554),
    .A2(net6295));
 sg13g2_nand2_1 _17110_ (.Y(_07353_),
    .A(net2738),
    .B(net6294));
 sg13g2_o21ai_1 _17111_ (.B1(_07353_),
    .Y(_01172_),
    .A1(net7714),
    .A2(net6294));
 sg13g2_nand3_1 _17112_ (.B(net7066),
    .C(net7217),
    .A(net7116),
    .Y(_07354_));
 sg13g2_nand2_1 _17113_ (.Y(_07355_),
    .A(net3807),
    .B(net6293));
 sg13g2_o21ai_1 _17114_ (.B1(_07355_),
    .Y(_01173_),
    .A1(net7347),
    .A2(net6293));
 sg13g2_nand2_1 _17115_ (.Y(_07356_),
    .A(net3567),
    .B(net6292));
 sg13g2_o21ai_1 _17116_ (.B1(_07356_),
    .Y(_01174_),
    .A1(net7544),
    .A2(net6292));
 sg13g2_nand2_1 _17117_ (.Y(_07357_),
    .A(net4297),
    .B(net6292));
 sg13g2_o21ai_1 _17118_ (.B1(_07357_),
    .Y(_01175_),
    .A1(net7703),
    .A2(net6292));
 sg13g2_nor3_1 _17119_ (.A(net7402),
    .B(net7267),
    .C(net7198),
    .Y(_07358_));
 sg13g2_nor2_1 _17120_ (.A(net4374),
    .B(net6808),
    .Y(_07359_));
 sg13g2_a21oi_1 _17121_ (.A1(net7310),
    .A2(net6808),
    .Y(_01176_),
    .B1(_07359_));
 sg13g2_nor2_1 _17122_ (.A(net4207),
    .B(net6807),
    .Y(_07360_));
 sg13g2_a21oi_1 _17123_ (.A1(net7510),
    .A2(net6807),
    .Y(_01177_),
    .B1(_07360_));
 sg13g2_nor2_1 _17124_ (.A(net4847),
    .B(net6807),
    .Y(_07361_));
 sg13g2_a21oi_1 _17125_ (.A1(net7667),
    .A2(net6807),
    .Y(_01178_),
    .B1(_07361_));
 sg13g2_nand3_1 _17126_ (.B(net7237),
    .C(net7207),
    .A(net7254),
    .Y(_07362_));
 sg13g2_nand2_1 _17127_ (.Y(_07363_),
    .A(net2485),
    .B(net6805));
 sg13g2_o21ai_1 _17128_ (.B1(_07363_),
    .Y(_01179_),
    .A1(net7304),
    .A2(net6805));
 sg13g2_nand2_1 _17129_ (.Y(_07364_),
    .A(net3076),
    .B(net6805));
 sg13g2_o21ai_1 _17130_ (.B1(_07364_),
    .Y(_01180_),
    .A1(net7502),
    .A2(net6805));
 sg13g2_nand2_1 _17131_ (.Y(_07365_),
    .A(net3748),
    .B(net6806));
 sg13g2_o21ai_1 _17132_ (.B1(_07365_),
    .Y(_01181_),
    .A1(net7661),
    .A2(net6806));
 sg13g2_nand3_1 _17133_ (.B(net7282),
    .C(net7217),
    .A(net7116),
    .Y(_07366_));
 sg13g2_nand2_1 _17134_ (.Y(_07367_),
    .A(net3626),
    .B(net6290));
 sg13g2_o21ai_1 _17135_ (.B1(_07367_),
    .Y(_01182_),
    .A1(net7347),
    .A2(net6290));
 sg13g2_nand2_1 _17136_ (.Y(_07368_),
    .A(net4292),
    .B(net6291));
 sg13g2_o21ai_1 _17137_ (.B1(_07368_),
    .Y(_01183_),
    .A1(net7545),
    .A2(net6291));
 sg13g2_nand2_1 _17138_ (.Y(_07369_),
    .A(net3862),
    .B(net6290));
 sg13g2_o21ai_1 _17139_ (.B1(_07369_),
    .Y(_01184_),
    .A1(net7704),
    .A2(net6290));
 sg13g2_nand3_1 _17140_ (.B(net7362),
    .C(net7217),
    .A(net7116),
    .Y(_07370_));
 sg13g2_nand2_1 _17141_ (.Y(_07371_),
    .A(net3298),
    .B(net6288));
 sg13g2_o21ai_1 _17142_ (.B1(_07371_),
    .Y(_01185_),
    .A1(net7347),
    .A2(net6288));
 sg13g2_nand2_1 _17143_ (.Y(_07372_),
    .A(net3498),
    .B(net6289));
 sg13g2_o21ai_1 _17144_ (.B1(_07372_),
    .Y(_01186_),
    .A1(net7545),
    .A2(net6289));
 sg13g2_nand2_1 _17145_ (.Y(_07373_),
    .A(net3404),
    .B(net6288));
 sg13g2_o21ai_1 _17146_ (.B1(_07373_),
    .Y(_01187_),
    .A1(net7704),
    .A2(net6288));
 sg13g2_nand3_1 _17147_ (.B(net7279),
    .C(net7219),
    .A(net7116),
    .Y(_07374_));
 sg13g2_nand2_1 _17148_ (.Y(_07375_),
    .A(net3293),
    .B(net6286));
 sg13g2_o21ai_1 _17149_ (.B1(_07375_),
    .Y(_01188_),
    .A1(net7347),
    .A2(net6286));
 sg13g2_nand2_1 _17150_ (.Y(_07376_),
    .A(net3851),
    .B(net6287));
 sg13g2_o21ai_1 _17151_ (.B1(_07376_),
    .Y(_01189_),
    .A1(net7545),
    .A2(net6287));
 sg13g2_nand2_1 _17152_ (.Y(_07377_),
    .A(net2867),
    .B(net6286));
 sg13g2_o21ai_1 _17153_ (.B1(_07377_),
    .Y(_01190_),
    .A1(net7704),
    .A2(net6286));
 sg13g2_nand3_1 _17154_ (.B(net7254),
    .C(net7206),
    .A(net7264),
    .Y(_07378_));
 sg13g2_nand2_1 _17155_ (.Y(_07379_),
    .A(net2911),
    .B(net6803));
 sg13g2_o21ai_1 _17156_ (.B1(_07379_),
    .Y(_01191_),
    .A1(net7304),
    .A2(net6803));
 sg13g2_nand2_1 _17157_ (.Y(_07380_),
    .A(net2536),
    .B(net6803));
 sg13g2_o21ai_1 _17158_ (.B1(_07380_),
    .Y(_01192_),
    .A1(net7502),
    .A2(net6803));
 sg13g2_nand2_1 _17159_ (.Y(_07381_),
    .A(net3354),
    .B(net6804));
 sg13g2_o21ai_1 _17160_ (.B1(_07381_),
    .Y(_01193_),
    .A1(net7661),
    .A2(net6804));
 sg13g2_nand3_1 _17161_ (.B(net7286),
    .C(net7217),
    .A(net7116),
    .Y(_07382_));
 sg13g2_nand2_1 _17162_ (.Y(_07383_),
    .A(net3407),
    .B(net6285));
 sg13g2_o21ai_1 _17163_ (.B1(_07383_),
    .Y(_01194_),
    .A1(net7348),
    .A2(net6285));
 sg13g2_nand2_1 _17164_ (.Y(_07384_),
    .A(net3366),
    .B(net6284));
 sg13g2_o21ai_1 _17165_ (.B1(_07384_),
    .Y(_01195_),
    .A1(net7545),
    .A2(net6284));
 sg13g2_nand2_1 _17166_ (.Y(_07385_),
    .A(net3940),
    .B(net6285));
 sg13g2_o21ai_1 _17167_ (.B1(_07385_),
    .Y(_01196_),
    .A1(net7705),
    .A2(net6285));
 sg13g2_nand3_1 _17168_ (.B(net7236),
    .C(net7206),
    .A(net7254),
    .Y(_07386_));
 sg13g2_nand2_1 _17169_ (.Y(_07387_),
    .A(net4354),
    .B(net6801));
 sg13g2_o21ai_1 _17170_ (.B1(_07387_),
    .Y(_01197_),
    .A1(net7304),
    .A2(net6801));
 sg13g2_nand2_1 _17171_ (.Y(_07388_),
    .A(net3716),
    .B(net6801));
 sg13g2_o21ai_1 _17172_ (.B1(_07388_),
    .Y(_01198_),
    .A1(net7502),
    .A2(net6801));
 sg13g2_nand2_1 _17173_ (.Y(_07389_),
    .A(net3553),
    .B(net6802));
 sg13g2_o21ai_1 _17174_ (.B1(_07389_),
    .Y(_01199_),
    .A1(net7661),
    .A2(net6802));
 sg13g2_nand3_1 _17175_ (.B(net7065),
    .C(net7206),
    .A(net7257),
    .Y(_07390_));
 sg13g2_nand2_1 _17176_ (.Y(_07391_),
    .A(net2585),
    .B(net6282));
 sg13g2_o21ai_1 _17177_ (.B1(_07391_),
    .Y(_01200_),
    .A1(net7301),
    .A2(net6282));
 sg13g2_nand2_1 _17178_ (.Y(_07392_),
    .A(net2573),
    .B(net6282));
 sg13g2_o21ai_1 _17179_ (.B1(_07392_),
    .Y(_01201_),
    .A1(net7500),
    .A2(net6282));
 sg13g2_nand2_1 _17180_ (.Y(_07393_),
    .A(net2921),
    .B(net6283));
 sg13g2_o21ai_1 _17181_ (.B1(_07393_),
    .Y(_01202_),
    .A1(net7660),
    .A2(net6283));
 sg13g2_nand3_1 _17182_ (.B(net7257),
    .C(net7206),
    .A(net7104),
    .Y(_07394_));
 sg13g2_nand2_1 _17183_ (.Y(_07395_),
    .A(net3444),
    .B(net6280));
 sg13g2_o21ai_1 _17184_ (.B1(_07395_),
    .Y(_01203_),
    .A1(net7301),
    .A2(net6280));
 sg13g2_nand2_1 _17185_ (.Y(_07396_),
    .A(net3090),
    .B(net6280));
 sg13g2_o21ai_1 _17186_ (.B1(_07396_),
    .Y(_01204_),
    .A1(net7500),
    .A2(net6280));
 sg13g2_nand2_1 _17187_ (.Y(_07397_),
    .A(net4396),
    .B(net6281));
 sg13g2_o21ai_1 _17188_ (.B1(_07397_),
    .Y(_01205_),
    .A1(net7660),
    .A2(net6281));
 sg13g2_nand3_1 _17189_ (.B(net7257),
    .C(net7206),
    .A(net7085),
    .Y(_07398_));
 sg13g2_nand2_1 _17190_ (.Y(_07399_),
    .A(net3311),
    .B(net6278));
 sg13g2_o21ai_1 _17191_ (.B1(_07399_),
    .Y(_01206_),
    .A1(net7301),
    .A2(net6278));
 sg13g2_nand2_1 _17192_ (.Y(_07400_),
    .A(net2528),
    .B(net6278));
 sg13g2_o21ai_1 _17193_ (.B1(_07400_),
    .Y(_01207_),
    .A1(net7500),
    .A2(net6278));
 sg13g2_nand2_1 _17194_ (.Y(_07401_),
    .A(net4043),
    .B(net6279));
 sg13g2_o21ai_1 _17195_ (.B1(_07401_),
    .Y(_01208_),
    .A1(net7660),
    .A2(net6279));
 sg13g2_nand3_1 _17196_ (.B(net7043),
    .C(net7206),
    .A(net7257),
    .Y(_07402_));
 sg13g2_nand2_1 _17197_ (.Y(_07403_),
    .A(net2696),
    .B(net6276));
 sg13g2_o21ai_1 _17198_ (.B1(_07403_),
    .Y(_01209_),
    .A1(net7301),
    .A2(net6276));
 sg13g2_nand2_1 _17199_ (.Y(_07404_),
    .A(net2508),
    .B(net6276));
 sg13g2_o21ai_1 _17200_ (.B1(_07404_),
    .Y(_01210_),
    .A1(net7500),
    .A2(net6276));
 sg13g2_nand2_1 _17201_ (.Y(_07405_),
    .A(net3288),
    .B(net6277));
 sg13g2_o21ai_1 _17202_ (.B1(_07405_),
    .Y(_01211_),
    .A1(net7660),
    .A2(net6277));
 sg13g2_nand3_1 _17203_ (.B(net7257),
    .C(net7206),
    .A(net7406),
    .Y(_07406_));
 sg13g2_nand2_1 _17204_ (.Y(_07407_),
    .A(net3766),
    .B(net6799));
 sg13g2_o21ai_1 _17205_ (.B1(_07407_),
    .Y(_01212_),
    .A1(net7295),
    .A2(net6799));
 sg13g2_nand2_1 _17206_ (.Y(_07408_),
    .A(net3044),
    .B(net6799));
 sg13g2_o21ai_1 _17207_ (.B1(_07408_),
    .Y(_01213_),
    .A1(net7493),
    .A2(net6799));
 sg13g2_nand2_1 _17208_ (.Y(_07409_),
    .A(net3237),
    .B(net6800));
 sg13g2_o21ai_1 _17209_ (.B1(_07409_),
    .Y(_01214_),
    .A1(net7652),
    .A2(net6800));
 sg13g2_nand3_1 _17210_ (.B(net7257),
    .C(net7205),
    .A(net7281),
    .Y(_07410_));
 sg13g2_nand2_1 _17211_ (.Y(_07411_),
    .A(net3209),
    .B(net6797));
 sg13g2_o21ai_1 _17212_ (.B1(_07411_),
    .Y(_01215_),
    .A1(net7295),
    .A2(net6797));
 sg13g2_nand2_1 _17213_ (.Y(_07412_),
    .A(net2621),
    .B(net6797));
 sg13g2_o21ai_1 _17214_ (.B1(_07412_),
    .Y(_01216_),
    .A1(net7500),
    .A2(net6797));
 sg13g2_nand2_1 _17215_ (.Y(_07413_),
    .A(net3902),
    .B(net6798));
 sg13g2_o21ai_1 _17216_ (.B1(_07413_),
    .Y(_01217_),
    .A1(net7652),
    .A2(net6797));
 sg13g2_nand3_1 _17217_ (.B(net7239),
    .C(net7210),
    .A(net7242),
    .Y(_07414_));
 sg13g2_nand2_1 _17218_ (.Y(_07415_),
    .A(net3614),
    .B(net6795));
 sg13g2_o21ai_1 _17219_ (.B1(_07415_),
    .Y(_01218_),
    .A1(net7326),
    .A2(net6795));
 sg13g2_nand2_1 _17220_ (.Y(_07416_),
    .A(net3182),
    .B(net6795));
 sg13g2_o21ai_1 _17221_ (.B1(_07416_),
    .Y(_01219_),
    .A1(net7525),
    .A2(net6795));
 sg13g2_nand2_1 _17222_ (.Y(_07417_),
    .A(net3757),
    .B(net6795));
 sg13g2_o21ai_1 _17223_ (.B1(_07417_),
    .Y(_01220_),
    .A1(net7682),
    .A2(net6795));
 sg13g2_nand3_1 _17224_ (.B(net7237),
    .C(net7211),
    .A(_04129_),
    .Y(_07418_));
 sg13g2_nand2_1 _17225_ (.Y(_07419_),
    .A(net2460),
    .B(net6794));
 sg13g2_o21ai_1 _17226_ (.B1(_07419_),
    .Y(_01221_),
    .A1(net7309),
    .A2(net6794));
 sg13g2_nand2_1 _17227_ (.Y(_07420_),
    .A(net3606),
    .B(net6793));
 sg13g2_o21ai_1 _17228_ (.B1(_07420_),
    .Y(_01222_),
    .A1(net7510),
    .A2(net6793));
 sg13g2_nand2_1 _17229_ (.Y(_07421_),
    .A(net2987),
    .B(net6793));
 sg13g2_o21ai_1 _17230_ (.B1(_07421_),
    .Y(_01223_),
    .A1(net7667),
    .A2(net6793));
 sg13g2_nand3_1 _17231_ (.B(net7257),
    .C(net7205),
    .A(net7280),
    .Y(_07422_));
 sg13g2_nand2_1 _17232_ (.Y(_07423_),
    .A(net3516),
    .B(net6791));
 sg13g2_o21ai_1 _17233_ (.B1(_07423_),
    .Y(_01224_),
    .A1(net7295),
    .A2(net6791));
 sg13g2_nand2_1 _17234_ (.Y(_07424_),
    .A(net2773),
    .B(net6791));
 sg13g2_o21ai_1 _17235_ (.B1(_07424_),
    .Y(_01225_),
    .A1(net7493),
    .A2(net6791));
 sg13g2_nand2_1 _17236_ (.Y(_07425_),
    .A(net3558),
    .B(net6792));
 sg13g2_o21ai_1 _17237_ (.B1(_07425_),
    .Y(_01226_),
    .A1(net7652),
    .A2(net6792));
 sg13g2_nand3_1 _17238_ (.B(net7255),
    .C(net7206),
    .A(net7285),
    .Y(_07426_));
 sg13g2_nand2_1 _17239_ (.Y(_07427_),
    .A(net2767),
    .B(net6789));
 sg13g2_o21ai_1 _17240_ (.B1(_07427_),
    .Y(_01227_),
    .A1(net7301),
    .A2(net6789));
 sg13g2_nand2_1 _17241_ (.Y(_07428_),
    .A(net2576),
    .B(net6789));
 sg13g2_o21ai_1 _17242_ (.B1(_07428_),
    .Y(_01228_),
    .A1(net7502),
    .A2(net6789));
 sg13g2_nand2_1 _17243_ (.Y(_07429_),
    .A(net2647),
    .B(net6790));
 sg13g2_o21ai_1 _17244_ (.B1(_07429_),
    .Y(_01229_),
    .A1(net7660),
    .A2(net6790));
 sg13g2_nor3_1 _17245_ (.A(net7271),
    .B(_04165_),
    .C(net7197),
    .Y(_07430_));
 sg13g2_nor2_1 _17246_ (.A(net4749),
    .B(net6787),
    .Y(_07431_));
 sg13g2_a21oi_1 _17247_ (.A1(net7301),
    .A2(net6787),
    .Y(_01230_),
    .B1(_07431_));
 sg13g2_nor2_1 _17248_ (.A(net4536),
    .B(net6787),
    .Y(_07432_));
 sg13g2_a21oi_1 _17249_ (.A1(net7500),
    .A2(net6787),
    .Y(_01231_),
    .B1(_07432_));
 sg13g2_nor2_1 _17250_ (.A(net4427),
    .B(net6788),
    .Y(_07433_));
 sg13g2_a21oi_1 _17251_ (.A1(net7660),
    .A2(net6788),
    .Y(_01232_),
    .B1(_07433_));
 sg13g2_nor3_1 _17252_ (.A(net7275),
    .B(_04165_),
    .C(net7197),
    .Y(_07434_));
 sg13g2_nor2_1 _17253_ (.A(net4414),
    .B(net6785),
    .Y(_07435_));
 sg13g2_a21oi_1 _17254_ (.A1(net7302),
    .A2(net6785),
    .Y(_01233_),
    .B1(_07435_));
 sg13g2_nor2_1 _17255_ (.A(net4823),
    .B(net6785),
    .Y(_07436_));
 sg13g2_a21oi_1 _17256_ (.A1(net7500),
    .A2(net6785),
    .Y(_01234_),
    .B1(_07436_));
 sg13g2_nor2_1 _17257_ (.A(net4609),
    .B(net6786),
    .Y(_07437_));
 sg13g2_a21oi_1 _17258_ (.A1(net7660),
    .A2(net6786),
    .Y(_01235_),
    .B1(_07437_));
 sg13g2_nor3_1 _17259_ (.A(_04165_),
    .B(net7245),
    .C(net7197),
    .Y(_07438_));
 sg13g2_nor2_1 _17260_ (.A(net4391),
    .B(net6783),
    .Y(_07439_));
 sg13g2_a21oi_1 _17261_ (.A1(net7302),
    .A2(net6783),
    .Y(_01236_),
    .B1(_07439_));
 sg13g2_nor2_1 _17262_ (.A(net4771),
    .B(net6783),
    .Y(_07440_));
 sg13g2_a21oi_1 _17263_ (.A1(net7500),
    .A2(net6783),
    .Y(_01237_),
    .B1(_07440_));
 sg13g2_nor2_1 _17264_ (.A(net3885),
    .B(net6784),
    .Y(_07441_));
 sg13g2_a21oi_1 _17265_ (.A1(net7660),
    .A2(net6784),
    .Y(_01238_),
    .B1(_07441_));
 sg13g2_nor3_1 _17266_ (.A(net7402),
    .B(net7249),
    .C(net7194),
    .Y(_07442_));
 sg13g2_nor2_1 _17267_ (.A(net4504),
    .B(net6781),
    .Y(_07443_));
 sg13g2_a21oi_1 _17268_ (.A1(net7297),
    .A2(net6782),
    .Y(_01239_),
    .B1(_07443_));
 sg13g2_nor2_1 _17269_ (.A(net4080),
    .B(net6782),
    .Y(_07444_));
 sg13g2_a21oi_1 _17270_ (.A1(net7495),
    .A2(net6781),
    .Y(_01240_),
    .B1(_07444_));
 sg13g2_nor2_1 _17271_ (.A(net4085),
    .B(net6781),
    .Y(_07445_));
 sg13g2_a21oi_1 _17272_ (.A1(net7655),
    .A2(net6781),
    .Y(_01241_),
    .B1(_07445_));
 sg13g2_nor3_1 _17273_ (.A(net7249),
    .B(_04217_),
    .C(net7194),
    .Y(_07446_));
 sg13g2_nor2_1 _17274_ (.A(net3772),
    .B(net6779),
    .Y(_07447_));
 sg13g2_a21oi_1 _17275_ (.A1(net7297),
    .A2(net6779),
    .Y(_01242_),
    .B1(_07447_));
 sg13g2_nor2_1 _17276_ (.A(net4632),
    .B(net6779),
    .Y(_07448_));
 sg13g2_a21oi_1 _17277_ (.A1(net7495),
    .A2(net6779),
    .Y(_01243_),
    .B1(_07448_));
 sg13g2_nor2_1 _17278_ (.A(net4747),
    .B(net6780),
    .Y(_07449_));
 sg13g2_a21oi_1 _17279_ (.A1(net7655),
    .A2(net6780),
    .Y(_01244_),
    .B1(_07449_));
 sg13g2_nand3_1 _17280_ (.B(net7042),
    .C(net7213),
    .A(net7240),
    .Y(_07450_));
 sg13g2_nand2_1 _17281_ (.Y(_07451_),
    .A(net3104),
    .B(net6274));
 sg13g2_o21ai_1 _17282_ (.B1(_07451_),
    .Y(_01245_),
    .A1(net7336),
    .A2(net6274));
 sg13g2_nand2_1 _17283_ (.Y(_07452_),
    .A(net4136),
    .B(net6275));
 sg13g2_o21ai_1 _17284_ (.B1(_07452_),
    .Y(_01246_),
    .A1(net7534),
    .A2(net6275));
 sg13g2_nand2_1 _17285_ (.Y(_07453_),
    .A(net2618),
    .B(net6274));
 sg13g2_o21ai_1 _17286_ (.B1(_07453_),
    .Y(_01247_),
    .A1(net7690),
    .A2(net6274));
 sg13g2_nand3_1 _17287_ (.B(net7074),
    .C(net7223),
    .A(net7279),
    .Y(_07454_));
 sg13g2_nand2_1 _17288_ (.Y(_07455_),
    .A(net2491),
    .B(net6273));
 sg13g2_o21ai_1 _17289_ (.B1(_07455_),
    .Y(_01248_),
    .A1(net7358),
    .A2(net6272));
 sg13g2_nand2_1 _17290_ (.Y(_07456_),
    .A(net4496),
    .B(net6272));
 sg13g2_o21ai_1 _17291_ (.B1(_07456_),
    .Y(_01249_),
    .A1(net7555),
    .A2(net6272));
 sg13g2_nand2_1 _17292_ (.Y(_07457_),
    .A(net3481),
    .B(net6273));
 sg13g2_o21ai_1 _17293_ (.B1(_07457_),
    .Y(_01250_),
    .A1(net7715),
    .A2(net6272));
 sg13g2_nor3_1 _17294_ (.A(_04141_),
    .B(net7249),
    .C(net7194),
    .Y(_07458_));
 sg13g2_nor2_1 _17295_ (.A(net4272),
    .B(net6777),
    .Y(_07459_));
 sg13g2_a21oi_1 _17296_ (.A1(net7297),
    .A2(net6777),
    .Y(_01251_),
    .B1(_07459_));
 sg13g2_nor2_1 _17297_ (.A(net4829),
    .B(net6777),
    .Y(_07460_));
 sg13g2_a21oi_1 _17298_ (.A1(net7495),
    .A2(net6777),
    .Y(_01252_),
    .B1(_07460_));
 sg13g2_nor2_1 _17299_ (.A(net4507),
    .B(net6778),
    .Y(_07461_));
 sg13g2_a21oi_1 _17300_ (.A1(net7655),
    .A2(net6778),
    .Y(_01253_),
    .B1(_07461_));
 sg13g2_nor3_1 _17301_ (.A(net7249),
    .B(_04235_),
    .C(net7194),
    .Y(_02528_));
 sg13g2_nor2_1 _17302_ (.A(net3988),
    .B(net6775),
    .Y(_02529_));
 sg13g2_a21oi_1 _17303_ (.A1(net7297),
    .A2(net6775),
    .Y(_01254_),
    .B1(_02529_));
 sg13g2_nor2_1 _17304_ (.A(net4367),
    .B(net6775),
    .Y(_02530_));
 sg13g2_a21oi_1 _17305_ (.A1(net7495),
    .A2(net6775),
    .Y(_01255_),
    .B1(_02530_));
 sg13g2_nor2_1 _17306_ (.A(net4122),
    .B(net6776),
    .Y(_02531_));
 sg13g2_a21oi_1 _17307_ (.A1(net7655),
    .A2(net6776),
    .Y(_01256_),
    .B1(_02531_));
 sg13g2_nand3_1 _17308_ (.B(net7264),
    .C(net7211),
    .A(_04129_),
    .Y(_02532_));
 sg13g2_nand2_1 _17309_ (.Y(_02533_),
    .A(net2533),
    .B(net6774));
 sg13g2_o21ai_1 _17310_ (.B1(_02533_),
    .Y(_01257_),
    .A1(net7309),
    .A2(net6774));
 sg13g2_nand2_1 _17311_ (.Y(_02534_),
    .A(net3798),
    .B(net6773));
 sg13g2_o21ai_1 _17312_ (.B1(_02534_),
    .Y(_01258_),
    .A1(net7510),
    .A2(net6773));
 sg13g2_nand2_1 _17313_ (.Y(_02535_),
    .A(net3919),
    .B(net6773));
 sg13g2_o21ai_1 _17314_ (.B1(_02535_),
    .Y(_01259_),
    .A1(net7667),
    .A2(net6773));
 sg13g2_nand3_1 _17315_ (.B(net7240),
    .C(net7213),
    .A(net7408),
    .Y(_02536_));
 sg13g2_nand2_1 _17316_ (.Y(_02537_),
    .A(net2661),
    .B(net6771));
 sg13g2_o21ai_1 _17317_ (.B1(_02537_),
    .Y(_01260_),
    .A1(net7326),
    .A2(net6771));
 sg13g2_nand2_1 _17318_ (.Y(_02538_),
    .A(net2910),
    .B(net6771));
 sg13g2_o21ai_1 _17319_ (.B1(_02538_),
    .Y(_01261_),
    .A1(net7525),
    .A2(net6771));
 sg13g2_nand2_1 _17320_ (.Y(_02539_),
    .A(net3660),
    .B(net6772));
 sg13g2_o21ai_1 _17321_ (.B1(_02539_),
    .Y(_01262_),
    .A1(net7683),
    .A2(net6772));
 sg13g2_nor3_1 _17322_ (.A(_04101_),
    .B(net7250),
    .C(net7195),
    .Y(_02540_));
 sg13g2_nor2_1 _17323_ (.A(net4537),
    .B(net6770),
    .Y(_02541_));
 sg13g2_a21oi_1 _17324_ (.A1(net7297),
    .A2(net6770),
    .Y(_01263_),
    .B1(_02541_));
 sg13g2_nor2_1 _17325_ (.A(net3916),
    .B(net6770),
    .Y(_02542_));
 sg13g2_a21oi_1 _17326_ (.A1(net7496),
    .A2(net6770),
    .Y(_01264_),
    .B1(_02542_));
 sg13g2_nor2_1 _17327_ (.A(net4663),
    .B(net6769),
    .Y(_02543_));
 sg13g2_a21oi_1 _17328_ (.A1(net7655),
    .A2(net6769),
    .Y(_01265_),
    .B1(_02543_));
 sg13g2_nand3_1 _17329_ (.B(net7240),
    .C(net7210),
    .A(net7281),
    .Y(_02544_));
 sg13g2_nand2_1 _17330_ (.Y(_02545_),
    .A(net4186),
    .B(net6767));
 sg13g2_o21ai_1 _17331_ (.B1(_02545_),
    .Y(_01266_),
    .A1(net7326),
    .A2(net6767));
 sg13g2_nand2_1 _17332_ (.Y(_02546_),
    .A(net2933),
    .B(net6767));
 sg13g2_o21ai_1 _17333_ (.B1(_02546_),
    .Y(_01267_),
    .A1(net7525),
    .A2(net6767));
 sg13g2_nand2_1 _17334_ (.Y(_02547_),
    .A(net2668),
    .B(net6767));
 sg13g2_o21ai_1 _17335_ (.B1(_02547_),
    .Y(_01268_),
    .A1(net7682),
    .A2(net6767));
 sg13g2_nor3_1 _17336_ (.A(_04152_),
    .B(net7250),
    .C(net7195),
    .Y(_02548_));
 sg13g2_nor2_1 _17337_ (.A(net3928),
    .B(net6766),
    .Y(_02549_));
 sg13g2_a21oi_1 _17338_ (.A1(net7297),
    .A2(net6766),
    .Y(_01269_),
    .B1(_02549_));
 sg13g2_nor2_1 _17339_ (.A(net4685),
    .B(net6766),
    .Y(_02550_));
 sg13g2_a21oi_1 _17340_ (.A1(net7496),
    .A2(net6766),
    .Y(_01270_),
    .B1(_02550_));
 sg13g2_nor2_1 _17341_ (.A(net4358),
    .B(net6765),
    .Y(_02551_));
 sg13g2_a21oi_1 _17342_ (.A1(net7655),
    .A2(net6765),
    .Y(_01271_),
    .B1(_02551_));
 sg13g2_nor3_1 _17343_ (.A(net7250),
    .B(net7234),
    .C(net7195),
    .Y(_02552_));
 sg13g2_nor2_1 _17344_ (.A(net4853),
    .B(net6764),
    .Y(_02553_));
 sg13g2_a21oi_1 _17345_ (.A1(net7297),
    .A2(net6764),
    .Y(_01272_),
    .B1(_02553_));
 sg13g2_nor2_1 _17346_ (.A(net3655),
    .B(net6764),
    .Y(_02554_));
 sg13g2_a21oi_1 _17347_ (.A1(net7496),
    .A2(net6764),
    .Y(_01273_),
    .B1(_02554_));
 sg13g2_nor2_1 _17348_ (.A(net4526),
    .B(net6763),
    .Y(_02555_));
 sg13g2_a21oi_1 _17349_ (.A1(net7655),
    .A2(net6763),
    .Y(_01274_),
    .B1(_02555_));
 sg13g2_nor3_1 _17350_ (.A(_04040_),
    .B(net7250),
    .C(net7195),
    .Y(_02556_));
 sg13g2_nor2_1 _17351_ (.A(net4256),
    .B(net6271),
    .Y(_02557_));
 sg13g2_a21oi_1 _17352_ (.A1(net7300),
    .A2(net6271),
    .Y(_01275_),
    .B1(_02557_));
 sg13g2_nor2_1 _17353_ (.A(net4015),
    .B(net6270),
    .Y(_02558_));
 sg13g2_a21oi_1 _17354_ (.A1(net7496),
    .A2(net6270),
    .Y(_01276_),
    .B1(_02558_));
 sg13g2_nor2_1 _17355_ (.A(net4288),
    .B(net6271),
    .Y(_02559_));
 sg13g2_a21oi_1 _17356_ (.A1(net7656),
    .A2(net6270),
    .Y(_01277_),
    .B1(_02559_));
 sg13g2_nand3_1 _17357_ (.B(net7240),
    .C(net7213),
    .A(net7362),
    .Y(_02560_));
 sg13g2_nand2_1 _17358_ (.Y(_02561_),
    .A(net3303),
    .B(net6761));
 sg13g2_o21ai_1 _17359_ (.B1(_02561_),
    .Y(_01278_),
    .A1(net7332),
    .A2(net6761));
 sg13g2_nand2_1 _17360_ (.Y(_02562_),
    .A(net3265),
    .B(net6761));
 sg13g2_o21ai_1 _17361_ (.B1(_02562_),
    .Y(_01279_),
    .A1(net7525),
    .A2(net6761));
 sg13g2_nand2_1 _17362_ (.Y(_02563_),
    .A(net3123),
    .B(net6762));
 sg13g2_o21ai_1 _17363_ (.B1(_02563_),
    .Y(_01280_),
    .A1(net7682),
    .A2(net6762));
 sg13g2_nor3_1 _17364_ (.A(_04087_),
    .B(net7250),
    .C(net7195),
    .Y(_02564_));
 sg13g2_nor2_1 _17365_ (.A(net4320),
    .B(net6268),
    .Y(_02565_));
 sg13g2_a21oi_1 _17366_ (.A1(net7300),
    .A2(net6268),
    .Y(_01281_),
    .B1(_02565_));
 sg13g2_nor2_1 _17367_ (.A(net4811),
    .B(net6269),
    .Y(_02566_));
 sg13g2_a21oi_1 _17368_ (.A1(net7496),
    .A2(net6269),
    .Y(_01282_),
    .B1(_02566_));
 sg13g2_nor2_1 _17369_ (.A(net4732),
    .B(net6269),
    .Y(_02567_));
 sg13g2_a21oi_1 _17370_ (.A1(net7656),
    .A2(net6269),
    .Y(_01283_),
    .B1(_02567_));
 sg13g2_nor3_2 _17371_ (.A(net7369),
    .B(net7269),
    .C(_04152_),
    .Y(_02568_));
 sg13g2_a21oi_1 _17372_ (.A1(net9),
    .A2(_03924_),
    .Y(_02569_),
    .B1(net11));
 sg13g2_o21ai_1 _17373_ (.B1(_03925_),
    .Y(_02570_),
    .A1(net12),
    .A2(_02569_));
 sg13g2_a21oi_1 _17374_ (.A1(_03926_),
    .A2(_02570_),
    .Y(_02571_),
    .B1(net15));
 sg13g2_nor2_1 _17375_ (.A(net4388),
    .B(net6760),
    .Y(_02572_));
 sg13g2_a21oi_1 _17376_ (.A1(net6760),
    .A2(net7149),
    .Y(_01284_),
    .B1(_02572_));
 sg13g2_nor2_1 _17377_ (.A(net10),
    .B(net11),
    .Y(_02573_));
 sg13g2_nor3_1 _17378_ (.A(net12),
    .B(net13),
    .C(_02573_),
    .Y(_02574_));
 sg13g2_nor3_2 _17379_ (.A(net14),
    .B(net15),
    .C(_02574_),
    .Y(_02575_));
 sg13g2_nor2_1 _17380_ (.A(net4089),
    .B(net6760),
    .Y(_02576_));
 sg13g2_a21oi_1 _17381_ (.A1(net6759),
    .A2(net7445),
    .Y(_01285_),
    .B1(_02576_));
 sg13g2_nor4_2 _17382_ (.A(net12),
    .B(net13),
    .C(net14),
    .Y(_02577_),
    .D(net15));
 sg13g2_nor2_1 _17383_ (.A(net4164),
    .B(net6759),
    .Y(_02578_));
 sg13g2_a21oi_1 _17384_ (.A1(net6759),
    .A2(net7599),
    .Y(_01286_),
    .B1(_02578_));
 sg13g2_nor3_1 _17385_ (.A(_04065_),
    .B(net7250),
    .C(net7197),
    .Y(_02579_));
 sg13g2_nor2_1 _17386_ (.A(net4086),
    .B(net6267),
    .Y(_02580_));
 sg13g2_a21oi_1 _17387_ (.A1(net7301),
    .A2(net6267),
    .Y(_01287_),
    .B1(_02580_));
 sg13g2_nor2_1 _17388_ (.A(net4273),
    .B(net6266),
    .Y(_02581_));
 sg13g2_a21oi_1 _17389_ (.A1(net7496),
    .A2(net6266),
    .Y(_01288_),
    .B1(_02581_));
 sg13g2_nor2_1 _17390_ (.A(net3918),
    .B(net6267),
    .Y(_02582_));
 sg13g2_a21oi_1 _17391_ (.A1(net7656),
    .A2(net6266),
    .Y(_01289_),
    .B1(_02582_));
 sg13g2_nor3_1 _17392_ (.A(net7284),
    .B(net7249),
    .C(net7194),
    .Y(_02583_));
 sg13g2_nor2_1 _17393_ (.A(net4000),
    .B(net6757),
    .Y(_02584_));
 sg13g2_a21oi_1 _17394_ (.A1(net7289),
    .A2(net6757),
    .Y(_01290_),
    .B1(_02584_));
 sg13g2_nor2_1 _17395_ (.A(net4357),
    .B(net6758),
    .Y(_02585_));
 sg13g2_a21oi_1 _17396_ (.A1(net7495),
    .A2(net6758),
    .Y(_01291_),
    .B1(_02585_));
 sg13g2_nor2_1 _17397_ (.A(net3858),
    .B(net6758),
    .Y(_02586_));
 sg13g2_a21oi_1 _17398_ (.A1(net7647),
    .A2(net6758),
    .Y(_01292_),
    .B1(_02586_));
 sg13g2_nor3_1 _17399_ (.A(net7271),
    .B(net7249),
    .C(net7194),
    .Y(_02587_));
 sg13g2_nor2_1 _17400_ (.A(net4615),
    .B(net6755),
    .Y(_02588_));
 sg13g2_a21oi_1 _17401_ (.A1(net7289),
    .A2(net6755),
    .Y(_01293_),
    .B1(_02588_));
 sg13g2_nor2_1 _17402_ (.A(net4570),
    .B(net6756),
    .Y(_02589_));
 sg13g2_a21oi_1 _17403_ (.A1(net7495),
    .A2(net6756),
    .Y(_01294_),
    .B1(_02589_));
 sg13g2_nor2_1 _17404_ (.A(net4548),
    .B(net6756),
    .Y(_02590_));
 sg13g2_a21oi_1 _17405_ (.A1(net7647),
    .A2(net6756),
    .Y(_01295_),
    .B1(_02590_));
 sg13g2_nor3_1 _17406_ (.A(net7267),
    .B(_04235_),
    .C(net7198),
    .Y(_02591_));
 sg13g2_nor2_1 _17407_ (.A(net4671),
    .B(net6753),
    .Y(_02592_));
 sg13g2_a21oi_1 _17408_ (.A1(net7309),
    .A2(net6754),
    .Y(_01296_),
    .B1(_02592_));
 sg13g2_nor2_1 _17409_ (.A(net3816),
    .B(net6753),
    .Y(_02593_));
 sg13g2_a21oi_1 _17410_ (.A1(net7513),
    .A2(net6753),
    .Y(_01297_),
    .B1(_02593_));
 sg13g2_nor2_1 _17411_ (.A(net4721),
    .B(net6753),
    .Y(_02594_));
 sg13g2_a21oi_1 _17412_ (.A1(net7667),
    .A2(net6753),
    .Y(_01298_),
    .B1(_02594_));
 sg13g2_nand3_1 _17413_ (.B(net7240),
    .C(net7213),
    .A(net7279),
    .Y(_02595_));
 sg13g2_nand2_1 _17414_ (.Y(_02596_),
    .A(net2812),
    .B(net6751));
 sg13g2_o21ai_1 _17415_ (.B1(_02596_),
    .Y(_01299_),
    .A1(net7326),
    .A2(net6751));
 sg13g2_nand2_1 _17416_ (.Y(_02597_),
    .A(net2636),
    .B(net6751));
 sg13g2_o21ai_1 _17417_ (.B1(_02597_),
    .Y(_01300_),
    .A1(net7525),
    .A2(net6751));
 sg13g2_nand2_1 _17418_ (.Y(_02598_),
    .A(net4432),
    .B(net6752));
 sg13g2_o21ai_1 _17419_ (.B1(_02598_),
    .Y(_01301_),
    .A1(net7682),
    .A2(net6752));
 sg13g2_nor3_2 _17420_ (.A(net7276),
    .B(net7267),
    .C(net7200),
    .Y(_02599_));
 sg13g2_nor2_1 _17421_ (.A(net4690),
    .B(net6750),
    .Y(_02600_));
 sg13g2_a21oi_1 _17422_ (.A1(net7311),
    .A2(net6750),
    .Y(_01302_),
    .B1(_02600_));
 sg13g2_nor2_1 _17423_ (.A(net4549),
    .B(net6750),
    .Y(_02601_));
 sg13g2_a21oi_1 _17424_ (.A1(net7509),
    .A2(net6750),
    .Y(_01303_),
    .B1(_02601_));
 sg13g2_nor2_1 _17425_ (.A(net4298),
    .B(net6749),
    .Y(_02602_));
 sg13g2_a21oi_1 _17426_ (.A1(net7666),
    .A2(net6749),
    .Y(_01304_),
    .B1(_02602_));
 sg13g2_nor2_1 _17427_ (.A(_04041_),
    .B(net7198),
    .Y(_02603_));
 sg13g2_nor2_1 _17428_ (.A(net4693),
    .B(net6264),
    .Y(_02604_));
 sg13g2_a21oi_1 _17429_ (.A1(net7316),
    .A2(net6264),
    .Y(_01305_),
    .B1(_02604_));
 sg13g2_nor2_1 _17430_ (.A(net4275),
    .B(net6265),
    .Y(_02605_));
 sg13g2_a21oi_1 _17431_ (.A1(net7507),
    .A2(net6265),
    .Y(_01306_),
    .B1(_02605_));
 sg13g2_nor2_1 _17432_ (.A(net4633),
    .B(net6264),
    .Y(_02606_));
 sg13g2_a21oi_1 _17433_ (.A1(net7670),
    .A2(net6264),
    .Y(_01307_),
    .B1(_02606_));
 sg13g2_nand2b_1 _17434_ (.Y(_02607_),
    .B(_04135_),
    .A_N(net7559));
 sg13g2_mux2_1 _17435_ (.A0(\top1.addr_in[8] ),
    .A1(net4851),
    .S(_02607_),
    .X(_01308_));
 sg13g2_a21o_1 _17436_ (.A2(_03990_),
    .A1(_03975_),
    .B1(_03945_),
    .X(_02608_));
 sg13g2_nand3_1 _17437_ (.B(_07318_),
    .C(_02608_),
    .A(_04017_),
    .Y(_02609_));
 sg13g2_mux2_1 _17438_ (.A0(_00006_),
    .A1(\top1.addr_out[8] ),
    .S(_02609_),
    .X(_01309_));
 sg13g2_nor2_1 _17439_ (.A(net4858),
    .B(net4851),
    .Y(_02610_));
 sg13g2_nor2_1 _17440_ (.A(_04135_),
    .B(_02610_),
    .Y(_01310_));
 sg13g2_nor2_1 _17441_ (.A(\top1.mem_ctl.signal_detected ),
    .B(_04042_),
    .Y(_02611_));
 sg13g2_mux2_1 _17442_ (.A0(net4482),
    .A1(net7565),
    .S(net6263),
    .X(_01311_));
 sg13g2_mux2_1 _17443_ (.A0(net4585),
    .A1(net7564),
    .S(net6263),
    .X(_01312_));
 sg13g2_nor2_1 _17444_ (.A(net4675),
    .B(net6263),
    .Y(_02612_));
 sg13g2_a21oi_1 _17445_ (.A1(_03845_),
    .A2(net6262),
    .Y(_01313_),
    .B1(_02612_));
 sg13g2_mux2_1 _17446_ (.A0(net4589),
    .A1(\top1.addr_in[3] ),
    .S(net6263),
    .X(_01314_));
 sg13g2_nor2_1 _17447_ (.A(net4739),
    .B(net6262),
    .Y(_02613_));
 sg13g2_a21oi_1 _17448_ (.A1(_03846_),
    .A2(net6262),
    .Y(_01315_),
    .B1(_02613_));
 sg13g2_mux2_1 _17449_ (.A0(net4713),
    .A1(net7563),
    .S(net6262),
    .X(_01316_));
 sg13g2_nor2_1 _17450_ (.A(net4705),
    .B(net6262),
    .Y(_02614_));
 sg13g2_a21oi_1 _17451_ (.A1(_03847_),
    .A2(net6262),
    .Y(_01317_),
    .B1(_02614_));
 sg13g2_nor2_1 _17452_ (.A(net4303),
    .B(net6262),
    .Y(_02615_));
 sg13g2_a21oi_1 _17453_ (.A1(_03848_),
    .A2(net6262),
    .Y(_01318_),
    .B1(_02615_));
 sg13g2_nor2_1 _17454_ (.A(net4860),
    .B(\top1.addr_in[8] ),
    .Y(_02616_));
 sg13g2_nor2_1 _17455_ (.A(_04135_),
    .B(net4861),
    .Y(_01319_));
 sg13g2_nand2_1 _17456_ (.Y(_02617_),
    .A(\top1.event_time[22] ),
    .B(_05042_));
 sg13g2_xnor2_1 _17457_ (.Y(_01320_),
    .A(\top1.event_time[22] ),
    .B(net6897));
 sg13g2_xnor2_1 _17458_ (.Y(_01321_),
    .A(\top1.event_time[23] ),
    .B(_02617_));
 sg13g2_nand3_1 _17459_ (.B(\top1.event_time[22] ),
    .C(_05042_),
    .A(\top1.event_time[23] ),
    .Y(_02618_));
 sg13g2_xnor2_1 _17460_ (.Y(_01322_),
    .A(\top1.event_time[24] ),
    .B(_02618_));
 sg13g2_or3_1 _17461_ (.A(\top1.event_time[26] ),
    .B(_05035_),
    .C(net6897),
    .X(_02619_));
 sg13g2_nor3_1 _17462_ (.A(_03834_),
    .B(_05035_),
    .C(net6897),
    .Y(_02620_));
 sg13g2_a21oi_1 _17463_ (.A1(_03834_),
    .A2(_02619_),
    .Y(_01323_),
    .B1(_02620_));
 sg13g2_nor2_1 _17464_ (.A(\top1.event_time[26] ),
    .B(_02620_),
    .Y(_02621_));
 sg13g2_nor2_1 _17465_ (.A(_05044_),
    .B(_02621_),
    .Y(_01324_));
 sg13g2_nand3_1 _17466_ (.B(net7258),
    .C(net7214),
    .A(net7286),
    .Y(_02622_));
 sg13g2_nand2_1 _17467_ (.Y(_02623_),
    .A(net3262),
    .B(net6747));
 sg13g2_o21ai_1 _17468_ (.B1(_02623_),
    .Y(_01325_),
    .A1(net7329),
    .A2(net6747));
 sg13g2_nand2_1 _17469_ (.Y(_02624_),
    .A(net3488),
    .B(net6747));
 sg13g2_o21ai_1 _17470_ (.B1(_02624_),
    .Y(_01326_),
    .A1(net7528),
    .A2(net6747));
 sg13g2_nand2_1 _17471_ (.Y(_02625_),
    .A(net2597),
    .B(net6748));
 sg13g2_o21ai_1 _17472_ (.B1(_02625_),
    .Y(_01327_),
    .A1(net7686),
    .A2(net6748));
 sg13g2_nor2_1 _17473_ (.A(net4242),
    .B(net6759),
    .Y(_02626_));
 sg13g2_a21oi_1 _17474_ (.A1(net7319),
    .A2(net6759),
    .Y(_01328_),
    .B1(_02626_));
 sg13g2_nor2_1 _17475_ (.A(net4520),
    .B(net6759),
    .Y(_02627_));
 sg13g2_a21oi_1 _17476_ (.A1(net7514),
    .A2(net6759),
    .Y(_01329_),
    .B1(_02627_));
 sg13g2_nor2_1 _17477_ (.A(net4023),
    .B(net6759),
    .Y(_02628_));
 sg13g2_a21oi_1 _17478_ (.A1(net7675),
    .A2(net6760),
    .Y(_01330_),
    .B1(_02628_));
 sg13g2_nand2_1 _17479_ (.Y(_02629_),
    .A(net3254),
    .B(net6823));
 sg13g2_o21ai_1 _17480_ (.B1(_02629_),
    .Y(_01331_),
    .A1(net6823),
    .A2(net7165));
 sg13g2_nand2_1 _17481_ (.Y(_02630_),
    .A(net3402),
    .B(net6823));
 sg13g2_o21ai_1 _17482_ (.B1(_02630_),
    .Y(_01332_),
    .A1(net6823),
    .A2(net7461));
 sg13g2_nand2_1 _17483_ (.Y(_02631_),
    .A(net3593),
    .B(net6823));
 sg13g2_o21ai_1 _17484_ (.B1(_02631_),
    .Y(_01333_),
    .A1(net6823),
    .A2(net7616));
 sg13g2_nand2_1 _17485_ (.Y(_02632_),
    .A(net2927),
    .B(net6899));
 sg13g2_o21ai_1 _17486_ (.B1(_02632_),
    .Y(_01334_),
    .A1(net6899),
    .A2(net7156));
 sg13g2_nand2_1 _17487_ (.Y(_02633_),
    .A(net3281),
    .B(net6899));
 sg13g2_o21ai_1 _17488_ (.B1(_02633_),
    .Y(_01335_),
    .A1(net6899),
    .A2(net7451));
 sg13g2_nand2_1 _17489_ (.Y(_02634_),
    .A(net3823),
    .B(net6898));
 sg13g2_o21ai_1 _17490_ (.B1(_02634_),
    .Y(_01336_),
    .A1(net6898),
    .A2(net7610));
 sg13g2_nand2_1 _17491_ (.Y(_02635_),
    .A(net3171),
    .B(net6458));
 sg13g2_o21ai_1 _17492_ (.B1(_02635_),
    .Y(_01337_),
    .A1(net6458),
    .A2(net7187));
 sg13g2_nand2_1 _17493_ (.Y(_02636_),
    .A(net4299),
    .B(net6459));
 sg13g2_o21ai_1 _17494_ (.B1(_02636_),
    .Y(_01338_),
    .A1(net6458),
    .A2(net7484));
 sg13g2_nand2_1 _17495_ (.Y(_02637_),
    .A(net3832),
    .B(net6458));
 sg13g2_o21ai_1 _17496_ (.B1(_02637_),
    .Y(_01339_),
    .A1(net6459),
    .A2(net7642));
 sg13g2_nand2_1 _17497_ (.Y(_02638_),
    .A(net3729),
    .B(net6873));
 sg13g2_o21ai_1 _17498_ (.B1(_02638_),
    .Y(_01340_),
    .A1(net6873),
    .A2(net7188));
 sg13g2_nand2_1 _17499_ (.Y(_02639_),
    .A(net3121),
    .B(net6874));
 sg13g2_o21ai_1 _17500_ (.B1(_02639_),
    .Y(_01341_),
    .A1(net6874),
    .A2(net7485));
 sg13g2_nand2_1 _17501_ (.Y(_02640_),
    .A(net3477),
    .B(net6874));
 sg13g2_o21ai_1 _17502_ (.B1(_02640_),
    .Y(_01342_),
    .A1(net6874),
    .A2(net7641));
 sg13g2_nand2_1 _17503_ (.Y(_02641_),
    .A(net4489),
    .B(net6424));
 sg13g2_o21ai_1 _17504_ (.B1(_02641_),
    .Y(_01343_),
    .A1(net6424),
    .A2(net7181));
 sg13g2_nand2_1 _17505_ (.Y(_02642_),
    .A(net2660),
    .B(net6424));
 sg13g2_o21ai_1 _17506_ (.B1(_02642_),
    .Y(_01344_),
    .A1(net6424),
    .A2(net7478));
 sg13g2_nand2_1 _17507_ (.Y(_02643_),
    .A(net3482),
    .B(net6424));
 sg13g2_o21ai_1 _17508_ (.B1(_02643_),
    .Y(_01345_),
    .A1(net6424),
    .A2(net7639));
 sg13g2_nor2_1 _17509_ (.A(net4392),
    .B(net6416),
    .Y(_02644_));
 sg13g2_a21oi_1 _17510_ (.A1(net6416),
    .A2(net7122),
    .Y(_01346_),
    .B1(_02644_));
 sg13g2_nor2_1 _17511_ (.A(net4540),
    .B(net6417),
    .Y(_02645_));
 sg13g2_a21oi_1 _17512_ (.A1(net6416),
    .A2(net7420),
    .Y(_01347_),
    .B1(_02645_));
 sg13g2_nor2_1 _17513_ (.A(net4407),
    .B(net6416),
    .Y(_02646_));
 sg13g2_a21oi_1 _17514_ (.A1(net6416),
    .A2(net7575),
    .Y(_01348_),
    .B1(_02646_));
 sg13g2_nor2_1 _17515_ (.A(net4731),
    .B(net6406),
    .Y(_02647_));
 sg13g2_a21oi_1 _17516_ (.A1(net6407),
    .A2(net7120),
    .Y(_01349_),
    .B1(_02647_));
 sg13g2_nor2_1 _17517_ (.A(net4635),
    .B(net6406),
    .Y(_02648_));
 sg13g2_a21oi_1 _17518_ (.A1(net6406),
    .A2(net7415),
    .Y(_01350_),
    .B1(_02648_));
 sg13g2_nor2_1 _17519_ (.A(net4527),
    .B(net6406),
    .Y(_02649_));
 sg13g2_a21oi_1 _17520_ (.A1(net6407),
    .A2(net7575),
    .Y(_01351_),
    .B1(_02649_));
 sg13g2_nand2_1 _17521_ (.Y(_02650_),
    .A(net2489),
    .B(net6405));
 sg13g2_o21ai_1 _17522_ (.B1(_02650_),
    .Y(_01352_),
    .A1(net6405),
    .A2(net7137));
 sg13g2_nand2_1 _17523_ (.Y(_02651_),
    .A(net2605),
    .B(net6404));
 sg13g2_o21ai_1 _17524_ (.B1(_02651_),
    .Y(_01353_),
    .A1(net6404),
    .A2(net7431));
 sg13g2_nand2_1 _17525_ (.Y(_02652_),
    .A(net2616),
    .B(net6404));
 sg13g2_o21ai_1 _17526_ (.B1(_02652_),
    .Y(_01354_),
    .A1(net6404),
    .A2(net7591));
 sg13g2_nor2_1 _17527_ (.A(net4815),
    .B(net6388),
    .Y(_02653_));
 sg13g2_a21oi_1 _17528_ (.A1(net6389),
    .A2(net7160),
    .Y(_01355_),
    .B1(_02653_));
 sg13g2_nor2_1 _17529_ (.A(net4668),
    .B(net6388),
    .Y(_02654_));
 sg13g2_a21oi_1 _17530_ (.A1(net6388),
    .A2(net7457),
    .Y(_01356_),
    .B1(_02654_));
 sg13g2_nor2_1 _17531_ (.A(net4359),
    .B(net6389),
    .Y(_02655_));
 sg13g2_a21oi_1 _17532_ (.A1(net6389),
    .A2(net7620),
    .Y(_01357_),
    .B1(_02655_));
 sg13g2_nand2_1 _17533_ (.Y(_02656_),
    .A(net2946),
    .B(net6387));
 sg13g2_o21ai_1 _17534_ (.B1(_02656_),
    .Y(_01358_),
    .A1(net6387),
    .A2(net7173));
 sg13g2_nand2_1 _17535_ (.Y(_02657_),
    .A(net3749),
    .B(net6387));
 sg13g2_o21ai_1 _17536_ (.B1(_02657_),
    .Y(_01359_),
    .A1(net6386),
    .A2(net7469));
 sg13g2_nand2_1 _17537_ (.Y(_02658_),
    .A(net4153),
    .B(net6387));
 sg13g2_o21ai_1 _17538_ (.B1(_02658_),
    .Y(_01360_),
    .A1(net6386),
    .A2(net7628));
 sg13g2_nand2_1 _17539_ (.Y(_02659_),
    .A(net3125),
    .B(net6470));
 sg13g2_o21ai_1 _17540_ (.B1(_02659_),
    .Y(_01361_),
    .A1(net6470),
    .A2(net7176));
 sg13g2_nand2_1 _17541_ (.Y(_02660_),
    .A(net2751),
    .B(net6470));
 sg13g2_o21ai_1 _17542_ (.B1(_02660_),
    .Y(_01362_),
    .A1(net6471),
    .A2(net7472));
 sg13g2_nand2_1 _17543_ (.Y(_02661_),
    .A(net2975),
    .B(net6470));
 sg13g2_o21ai_1 _17544_ (.B1(_02661_),
    .Y(_01363_),
    .A1(net6471),
    .A2(net7632));
 sg13g2_nor2_1 _17545_ (.A(net4429),
    .B(net6904),
    .Y(_02662_));
 sg13g2_a21oi_1 _17546_ (.A1(net6904),
    .A2(net7121),
    .Y(_01364_),
    .B1(_02662_));
 sg13g2_nor2_1 _17547_ (.A(net4765),
    .B(net6904),
    .Y(_02663_));
 sg13g2_a21oi_1 _17548_ (.A1(net6904),
    .A2(net7416),
    .Y(_01365_),
    .B1(_02663_));
 sg13g2_nor2_1 _17549_ (.A(net4541),
    .B(net6904),
    .Y(_02664_));
 sg13g2_a21oi_1 _17550_ (.A1(net6904),
    .A2(net7581),
    .Y(_01366_),
    .B1(_02664_));
 sg13g2_nor2_1 _17551_ (.A(net4722),
    .B(net6902),
    .Y(_02665_));
 sg13g2_a21oi_1 _17552_ (.A1(net6902),
    .A2(net7127),
    .Y(_01367_),
    .B1(_02665_));
 sg13g2_nor2_1 _17553_ (.A(net4301),
    .B(net6902),
    .Y(_02666_));
 sg13g2_a21oi_1 _17554_ (.A1(net6902),
    .A2(net7423),
    .Y(_01368_),
    .B1(_02666_));
 sg13g2_nor2_1 _17555_ (.A(net4445),
    .B(net6902),
    .Y(_02667_));
 sg13g2_a21oi_1 _17556_ (.A1(net6902),
    .A2(net7582),
    .Y(_01369_),
    .B1(_02667_));
 sg13g2_nand2_1 _17557_ (.Y(_02668_),
    .A(net3286),
    .B(net6911));
 sg13g2_o21ai_1 _17558_ (.B1(_02668_),
    .Y(_01370_),
    .A1(net6911),
    .A2(net7126));
 sg13g2_nand2_1 _17559_ (.Y(_02669_),
    .A(net3356),
    .B(net6910));
 sg13g2_o21ai_1 _17560_ (.B1(_02669_),
    .Y(_01371_),
    .A1(net6910),
    .A2(net7420));
 sg13g2_nand2_1 _17561_ (.Y(_02670_),
    .A(net3307),
    .B(net6910));
 sg13g2_o21ai_1 _17562_ (.B1(_02670_),
    .Y(_01372_),
    .A1(net6910),
    .A2(net7578));
 sg13g2_nand2_1 _17563_ (.Y(_02671_),
    .A(net2472),
    .B(net6909));
 sg13g2_o21ai_1 _17564_ (.B1(_02671_),
    .Y(_01373_),
    .A1(net6909),
    .A2(net7133));
 sg13g2_nand2_1 _17565_ (.Y(_02672_),
    .A(net3230),
    .B(net6908));
 sg13g2_o21ai_1 _17566_ (.B1(_02672_),
    .Y(_01374_),
    .A1(net6908),
    .A2(net7428));
 sg13g2_nand2_1 _17567_ (.Y(_02673_),
    .A(net3595),
    .B(net6908));
 sg13g2_o21ai_1 _17568_ (.B1(_02673_),
    .Y(_01375_),
    .A1(net6908),
    .A2(net7588));
 sg13g2_nand2_1 _17569_ (.Y(_02674_),
    .A(net2892),
    .B(net6491));
 sg13g2_o21ai_1 _17570_ (.B1(_02674_),
    .Y(_01376_),
    .A1(net6490),
    .A2(net7153));
 sg13g2_nand2_1 _17571_ (.Y(_02675_),
    .A(net2961),
    .B(net6491));
 sg13g2_o21ai_1 _17572_ (.B1(_02675_),
    .Y(_01377_),
    .A1(net6491),
    .A2(net7449));
 sg13g2_nand2_1 _17573_ (.Y(_02676_),
    .A(net2588),
    .B(net6491));
 sg13g2_o21ai_1 _17574_ (.B1(_02676_),
    .Y(_01378_),
    .A1(net6490),
    .A2(net7608));
 sg13g2_nand2_1 _17575_ (.Y(_02677_),
    .A(net3373),
    .B(net6748));
 sg13g2_o21ai_1 _17576_ (.B1(_02677_),
    .Y(_01379_),
    .A1(net7159),
    .A2(net6748));
 sg13g2_nand2_1 _17577_ (.Y(_02678_),
    .A(net4258),
    .B(net6747));
 sg13g2_o21ai_1 _17578_ (.B1(_02678_),
    .Y(_01380_),
    .A1(net7453),
    .A2(net6747));
 sg13g2_nand2_1 _17579_ (.Y(_02679_),
    .A(net2574),
    .B(net6747));
 sg13g2_o21ai_1 _17580_ (.B1(_02679_),
    .Y(_01381_),
    .A1(net7614),
    .A2(net6747));
 sg13g2_nand2_1 _17581_ (.Y(_02680_),
    .A(net3995),
    .B(net6825));
 sg13g2_o21ai_1 _17582_ (.B1(_02680_),
    .Y(_01382_),
    .A1(net6825),
    .A2(net7155));
 sg13g2_nand2_1 _17583_ (.Y(_02681_),
    .A(net3835),
    .B(net6825));
 sg13g2_o21ai_1 _17584_ (.B1(_02681_),
    .Y(_01383_),
    .A1(net6825),
    .A2(net7451));
 sg13g2_nand2_1 _17585_ (.Y(_02682_),
    .A(net3964),
    .B(net6826));
 sg13g2_o21ai_1 _17586_ (.B1(_02682_),
    .Y(_01384_),
    .A1(net6826),
    .A2(net7614));
 sg13g2_nor2_1 _17587_ (.A(net4657),
    .B(net6264),
    .Y(_02683_));
 sg13g2_a21oi_1 _17588_ (.A1(net7145),
    .A2(net6264),
    .Y(_01385_),
    .B1(_02683_));
 sg13g2_nor2_1 _17589_ (.A(net4694),
    .B(net6264),
    .Y(_02684_));
 sg13g2_a21oi_1 _17590_ (.A1(net7438),
    .A2(net6264),
    .Y(_01386_),
    .B1(_02684_));
 sg13g2_nor2_1 _17591_ (.A(net4282),
    .B(net6265),
    .Y(_02685_));
 sg13g2_a21oi_1 _17592_ (.A1(net7592),
    .A2(net6265),
    .Y(_01387_),
    .B1(_02685_));
 sg13g2_nor2_1 _17593_ (.A(net4679),
    .B(net6749),
    .Y(_02686_));
 sg13g2_a21oi_1 _17594_ (.A1(net7140),
    .A2(net6749),
    .Y(_01388_),
    .B1(_02686_));
 sg13g2_nor2_1 _17595_ (.A(net4623),
    .B(net6749),
    .Y(_02687_));
 sg13g2_a21oi_1 _17596_ (.A1(net7434),
    .A2(net6749),
    .Y(_01389_),
    .B1(_02687_));
 sg13g2_nor2_1 _17597_ (.A(net4457),
    .B(net6749),
    .Y(_02688_));
 sg13g2_a21oi_1 _17598_ (.A1(net7596),
    .A2(net6749),
    .Y(_01390_),
    .B1(_02688_));
 sg13g2_nand2_1 _17599_ (.Y(_02689_),
    .A(net2566),
    .B(net6752));
 sg13g2_o21ai_1 _17600_ (.B1(_02689_),
    .Y(_01391_),
    .A1(net7156),
    .A2(net6752));
 sg13g2_nand2_1 _17601_ (.Y(_02690_),
    .A(net3116),
    .B(net6751));
 sg13g2_o21ai_1 _17602_ (.B1(_02690_),
    .Y(_01392_),
    .A1(net7451),
    .A2(net6751));
 sg13g2_nand2_1 _17603_ (.Y(_02691_),
    .A(net3103),
    .B(net6751));
 sg13g2_o21ai_1 _17604_ (.B1(_02691_),
    .Y(_01393_),
    .A1(net7611),
    .A2(net6751));
 sg13g2_nand2_1 _17605_ (.Y(_02692_),
    .A(net3973),
    .B(net6762));
 sg13g2_o21ai_1 _17606_ (.B1(_02692_),
    .Y(_01394_),
    .A1(net6762),
    .A2(net7156));
 sg13g2_nand2_1 _17607_ (.Y(_02693_),
    .A(net2899),
    .B(net6761));
 sg13g2_o21ai_1 _17608_ (.B1(_02693_),
    .Y(_01395_),
    .A1(net6761),
    .A2(net7452));
 sg13g2_nand2_1 _17609_ (.Y(_02694_),
    .A(net2542),
    .B(net6761));
 sg13g2_o21ai_1 _17610_ (.B1(_02694_),
    .Y(_01396_),
    .A1(net6761),
    .A2(net7610));
 sg13g2_nand2_1 _17611_ (.Y(_02695_),
    .A(net2556),
    .B(net6768));
 sg13g2_o21ai_1 _17612_ (.B1(_02695_),
    .Y(_01397_),
    .A1(net6768),
    .A2(net7155));
 sg13g2_nand2_1 _17613_ (.Y(_02696_),
    .A(net3762),
    .B(net6768));
 sg13g2_o21ai_1 _17614_ (.B1(_02696_),
    .Y(_01398_),
    .A1(net6767),
    .A2(net7452));
 sg13g2_nand2_1 _17615_ (.Y(_02697_),
    .A(net2879),
    .B(net6767));
 sg13g2_o21ai_1 _17616_ (.B1(_02697_),
    .Y(_01399_),
    .A1(net6768),
    .A2(net7611));
 sg13g2_nand2_1 _17617_ (.Y(_02698_),
    .A(net3670),
    .B(net6772));
 sg13g2_o21ai_1 _17618_ (.B1(_02698_),
    .Y(_01400_),
    .A1(net6772),
    .A2(net7155));
 sg13g2_nand2_1 _17619_ (.Y(_02699_),
    .A(net3622),
    .B(net6771));
 sg13g2_o21ai_1 _17620_ (.B1(_02699_),
    .Y(_01401_),
    .A1(net6771),
    .A2(net7451));
 sg13g2_nand2_1 _17621_ (.Y(_02700_),
    .A(net4018),
    .B(net6771));
 sg13g2_o21ai_1 _17622_ (.B1(_02700_),
    .Y(_01402_),
    .A1(net6771),
    .A2(net7610));
 sg13g2_nand2_1 _17623_ (.Y(_02701_),
    .A(net2575),
    .B(net6274));
 sg13g2_o21ai_1 _17624_ (.B1(_02701_),
    .Y(_01403_),
    .A1(net6274),
    .A2(net7155));
 sg13g2_nand2_1 _17625_ (.Y(_02702_),
    .A(net4083),
    .B(net6275));
 sg13g2_o21ai_1 _17626_ (.B1(_02702_),
    .Y(_01404_),
    .A1(net6275),
    .A2(net7462));
 sg13g2_nand2_1 _17627_ (.Y(_02703_),
    .A(net3492),
    .B(net6274));
 sg13g2_o21ai_1 _17628_ (.B1(_02703_),
    .Y(_01405_),
    .A1(net6274),
    .A2(net7610));
 sg13g2_nand2_1 _17629_ (.Y(_02704_),
    .A(net3418),
    .B(net6338));
 sg13g2_o21ai_1 _17630_ (.B1(_02704_),
    .Y(_01406_),
    .A1(net6338),
    .A2(net7155));
 sg13g2_nand2_1 _17631_ (.Y(_02705_),
    .A(net3511),
    .B(net6339));
 sg13g2_o21ai_1 _17632_ (.B1(_02705_),
    .Y(_01407_),
    .A1(net6339),
    .A2(net7462));
 sg13g2_nand2_1 _17633_ (.Y(_02706_),
    .A(net4323),
    .B(net6338));
 sg13g2_o21ai_1 _17634_ (.B1(_02706_),
    .Y(_01408_),
    .A1(net6339),
    .A2(net7610));
 sg13g2_nand2_1 _17635_ (.Y(_02707_),
    .A(net3018),
    .B(net6340));
 sg13g2_o21ai_1 _17636_ (.B1(_02707_),
    .Y(_01409_),
    .A1(net6340),
    .A2(net7155));
 sg13g2_nand2_1 _17637_ (.Y(_02708_),
    .A(net3333),
    .B(net6341));
 sg13g2_o21ai_1 _17638_ (.B1(_02708_),
    .Y(_01410_),
    .A1(net6340),
    .A2(net7462));
 sg13g2_nand2_1 _17639_ (.Y(_02709_),
    .A(net3438),
    .B(net6341));
 sg13g2_o21ai_1 _17640_ (.B1(_02709_),
    .Y(_01411_),
    .A1(net6341),
    .A2(net7615));
 sg13g2_nand2_1 _17641_ (.Y(_02710_),
    .A(net2763),
    .B(net6342));
 sg13g2_o21ai_1 _17642_ (.B1(_02710_),
    .Y(_01412_),
    .A1(net6342),
    .A2(net7155));
 sg13g2_nand2_1 _17643_ (.Y(_02711_),
    .A(net3093),
    .B(net6343));
 sg13g2_o21ai_1 _17644_ (.B1(_02711_),
    .Y(_01413_),
    .A1(net6342),
    .A2(net7462));
 sg13g2_nand2_1 _17645_ (.Y(_02712_),
    .A(net3448),
    .B(net6343));
 sg13g2_o21ai_1 _17646_ (.B1(_02712_),
    .Y(_01414_),
    .A1(net6343),
    .A2(net7615));
 sg13g2_nand2_1 _17647_ (.Y(_02713_),
    .A(net2759),
    .B(net6820));
 sg13g2_o21ai_1 _17648_ (.B1(_02713_),
    .Y(_01415_),
    .A1(net6820),
    .A2(net7156));
 sg13g2_nand2_1 _17649_ (.Y(_02714_),
    .A(net3364),
    .B(net6820));
 sg13g2_o21ai_1 _17650_ (.B1(_02714_),
    .Y(_01416_),
    .A1(net6820),
    .A2(net7451));
 sg13g2_nand2_1 _17651_ (.Y(_02715_),
    .A(net3551),
    .B(net6819));
 sg13g2_o21ai_1 _17652_ (.B1(_02715_),
    .Y(_01417_),
    .A1(net6819),
    .A2(net7610));
 sg13g2_nor2_1 _17653_ (.A(net4110),
    .B(net6821),
    .Y(_02716_));
 sg13g2_a21oi_1 _17654_ (.A1(net6821),
    .A2(net7140),
    .Y(_01418_),
    .B1(_02716_));
 sg13g2_nor2_1 _17655_ (.A(net4691),
    .B(net6821),
    .Y(_02717_));
 sg13g2_a21oi_1 _17656_ (.A1(net6821),
    .A2(net7434),
    .Y(_01419_),
    .B1(_02717_));
 sg13g2_nor2_1 _17657_ (.A(net4576),
    .B(net6821),
    .Y(_02718_));
 sg13g2_a21oi_1 _17658_ (.A1(net6821),
    .A2(net7596),
    .Y(_01420_),
    .B1(_02718_));
 sg13g2_nand2_1 _17659_ (.Y(_02719_),
    .A(net3193),
    .B(net6796));
 sg13g2_o21ai_1 _17660_ (.B1(_02719_),
    .Y(_01421_),
    .A1(net6796),
    .A2(net7156));
 sg13g2_nand2_1 _17661_ (.Y(_02720_),
    .A(net3947),
    .B(net6796));
 sg13g2_o21ai_1 _17662_ (.B1(_02720_),
    .Y(_01422_),
    .A1(net6796),
    .A2(net7451));
 sg13g2_nand2_1 _17663_ (.Y(_02721_),
    .A(net3680),
    .B(net6795));
 sg13g2_o21ai_1 _17664_ (.B1(_02721_),
    .Y(_01423_),
    .A1(net6795),
    .A2(net7610));
 sg13g2_nand2_1 _17665_ (.Y(_02722_),
    .A(net3777),
    .B(net6828));
 sg13g2_o21ai_1 _17666_ (.B1(_02722_),
    .Y(_01424_),
    .A1(net6828),
    .A2(net7156));
 sg13g2_nand2_1 _17667_ (.Y(_02723_),
    .A(net2826),
    .B(net6828));
 sg13g2_o21ai_1 _17668_ (.B1(_02723_),
    .Y(_01425_),
    .A1(net6828),
    .A2(net7451));
 sg13g2_nand2_1 _17669_ (.Y(_02724_),
    .A(net3860),
    .B(net6827));
 sg13g2_o21ai_1 _17670_ (.B1(_02724_),
    .Y(_01426_),
    .A1(net6827),
    .A2(net7610));
 sg13g2_nand2_1 _17671_ (.Y(_02725_),
    .A(net3332),
    .B(net6294));
 sg13g2_o21ai_1 _17672_ (.B1(_02725_),
    .Y(_01427_),
    .A1(net6294),
    .A2(net7186));
 sg13g2_nand2_1 _17673_ (.Y(_02726_),
    .A(net2615),
    .B(net6294));
 sg13g2_o21ai_1 _17674_ (.B1(_02726_),
    .Y(_01428_),
    .A1(net6294),
    .A2(net7483));
 sg13g2_nand2_1 _17675_ (.Y(_02727_),
    .A(net2522),
    .B(net6294));
 sg13g2_o21ai_1 _17676_ (.B1(_02727_),
    .Y(_01429_),
    .A1(net6295),
    .A2(net7641));
 sg13g2_nand2_1 _17677_ (.Y(_02728_),
    .A(net3467),
    .B(net6360));
 sg13g2_o21ai_1 _17678_ (.B1(_02728_),
    .Y(_01430_),
    .A1(net6361),
    .A2(net7186));
 sg13g2_nand2_1 _17679_ (.Y(_02729_),
    .A(net3933),
    .B(net6360));
 sg13g2_o21ai_1 _17680_ (.B1(_02729_),
    .Y(_01431_),
    .A1(net6360),
    .A2(net7483));
 sg13g2_nand2_1 _17681_ (.Y(_02730_),
    .A(net2827),
    .B(net6360));
 sg13g2_o21ai_1 _17682_ (.B1(_02730_),
    .Y(_01432_),
    .A1(net6361),
    .A2(net7641));
 sg13g2_nand2_1 _17683_ (.Y(_02731_),
    .A(net2823),
    .B(net6358));
 sg13g2_o21ai_1 _17684_ (.B1(_02731_),
    .Y(_01433_),
    .A1(net6359),
    .A2(net7186));
 sg13g2_nand2_1 _17685_ (.Y(_02732_),
    .A(net2937),
    .B(net6358));
 sg13g2_o21ai_1 _17686_ (.B1(_02732_),
    .Y(_01434_),
    .A1(net6358),
    .A2(net7483));
 sg13g2_nand2_1 _17687_ (.Y(_02733_),
    .A(net3068),
    .B(net6358));
 sg13g2_o21ai_1 _17688_ (.B1(_02733_),
    .Y(_01435_),
    .A1(net6359),
    .A2(net7642));
 sg13g2_nand2_1 _17689_ (.Y(_02734_),
    .A(net3532),
    .B(net6350));
 sg13g2_o21ai_1 _17690_ (.B1(_02734_),
    .Y(_01436_),
    .A1(net6351),
    .A2(net7186));
 sg13g2_nand2_1 _17691_ (.Y(_02735_),
    .A(net2929),
    .B(net6350));
 sg13g2_o21ai_1 _17692_ (.B1(_02735_),
    .Y(_01437_),
    .A1(net6350),
    .A2(net7483));
 sg13g2_nand2_1 _17693_ (.Y(_02736_),
    .A(net2503),
    .B(net6350));
 sg13g2_o21ai_1 _17694_ (.B1(_02736_),
    .Y(_01438_),
    .A1(net6351),
    .A2(net7642));
 sg13g2_nand2_1 _17695_ (.Y(_02737_),
    .A(net3153),
    .B(net6272));
 sg13g2_o21ai_1 _17696_ (.B1(_02737_),
    .Y(_01439_),
    .A1(net6272),
    .A2(net7187));
 sg13g2_nand2_1 _17697_ (.Y(_02738_),
    .A(net3503),
    .B(net6273));
 sg13g2_o21ai_1 _17698_ (.B1(_02738_),
    .Y(_01440_),
    .A1(net6272),
    .A2(net7484));
 sg13g2_nand2_1 _17699_ (.Y(_02739_),
    .A(net3681),
    .B(net6272));
 sg13g2_o21ai_1 _17700_ (.B1(_02739_),
    .Y(_01441_),
    .A1(net6273),
    .A2(net7642));
 sg13g2_nand2_1 _17701_ (.Y(_02740_),
    .A(net3664),
    .B(net6304));
 sg13g2_o21ai_1 _17702_ (.B1(_02740_),
    .Y(_01442_),
    .A1(net6304),
    .A2(net7187));
 sg13g2_nand2_1 _17703_ (.Y(_02741_),
    .A(net3225),
    .B(net6305));
 sg13g2_o21ai_1 _17704_ (.B1(_02741_),
    .Y(_01443_),
    .A1(net6305),
    .A2(net7484));
 sg13g2_nand2_1 _17705_ (.Y(_02742_),
    .A(net3836),
    .B(net6304));
 sg13g2_o21ai_1 _17706_ (.B1(_02742_),
    .Y(_01444_),
    .A1(net6305),
    .A2(net7641));
 sg13g2_nand2_1 _17707_ (.Y(_02743_),
    .A(net3610),
    .B(net6456));
 sg13g2_o21ai_1 _17708_ (.B1(_02743_),
    .Y(_01445_),
    .A1(net6456),
    .A2(net7187));
 sg13g2_nand2_1 _17709_ (.Y(_02744_),
    .A(net3708),
    .B(net6457));
 sg13g2_o21ai_1 _17710_ (.B1(_02744_),
    .Y(_01446_),
    .A1(net6456),
    .A2(net7484));
 sg13g2_nand2_1 _17711_ (.Y(_02745_),
    .A(net3719),
    .B(net6456));
 sg13g2_o21ai_1 _17712_ (.B1(_02745_),
    .Y(_01447_),
    .A1(net6457),
    .A2(net7641));
 sg13g2_nor2_1 _17713_ (.A(net3971),
    .B(net6895),
    .Y(_02746_));
 sg13g2_a21oi_1 _17714_ (.A1(net6895),
    .A2(net7140),
    .Y(_01448_),
    .B1(_02746_));
 sg13g2_nor2_1 _17715_ (.A(net4754),
    .B(net6895),
    .Y(_02747_));
 sg13g2_a21oi_1 _17716_ (.A1(net6895),
    .A2(net7434),
    .Y(_01449_),
    .B1(_02747_));
 sg13g2_nor2_1 _17717_ (.A(net4839),
    .B(net6895),
    .Y(_02748_));
 sg13g2_a21oi_1 _17718_ (.A1(net6895),
    .A2(net7596),
    .Y(_01450_),
    .B1(_02748_));
 sg13g2_nand2_1 _17719_ (.Y(_02749_),
    .A(net3868),
    .B(net6454));
 sg13g2_o21ai_1 _17720_ (.B1(_02749_),
    .Y(_01451_),
    .A1(net6454),
    .A2(net7186));
 sg13g2_nand2_1 _17721_ (.Y(_02750_),
    .A(net3229),
    .B(net6455));
 sg13g2_o21ai_1 _17722_ (.B1(_02750_),
    .Y(_01452_),
    .A1(net6455),
    .A2(net7483));
 sg13g2_nand2_1 _17723_ (.Y(_02751_),
    .A(net3207),
    .B(net6454));
 sg13g2_o21ai_1 _17724_ (.B1(_02751_),
    .Y(_01453_),
    .A1(net6454),
    .A2(net7640));
 sg13g2_nand2_1 _17725_ (.Y(_02752_),
    .A(net3202),
    .B(net6452));
 sg13g2_o21ai_1 _17726_ (.B1(_02752_),
    .Y(_01454_),
    .A1(net6452),
    .A2(net7186));
 sg13g2_nand2_1 _17727_ (.Y(_02753_),
    .A(net3308),
    .B(net6453));
 sg13g2_o21ai_1 _17728_ (.B1(_02753_),
    .Y(_01455_),
    .A1(net6453),
    .A2(net7483));
 sg13g2_nand2_1 _17729_ (.Y(_02754_),
    .A(net3347),
    .B(net6452));
 sg13g2_o21ai_1 _17730_ (.B1(_02754_),
    .Y(_01456_),
    .A1(net6452),
    .A2(net7640));
 sg13g2_nand2_1 _17731_ (.Y(_02755_),
    .A(net3335),
    .B(net6450));
 sg13g2_o21ai_1 _17732_ (.B1(_02755_),
    .Y(_01457_),
    .A1(net6450),
    .A2(net7186));
 sg13g2_nand2_1 _17733_ (.Y(_02756_),
    .A(net3217),
    .B(net6451));
 sg13g2_o21ai_1 _17734_ (.B1(_02756_),
    .Y(_01458_),
    .A1(net6451),
    .A2(net7483));
 sg13g2_nand2_1 _17735_ (.Y(_02757_),
    .A(net3747),
    .B(net6450));
 sg13g2_o21ai_1 _17736_ (.B1(_02757_),
    .Y(_01459_),
    .A1(net6450),
    .A2(net7639));
 sg13g2_nand2_1 _17737_ (.Y(_02758_),
    .A(net4239),
    .B(net6448));
 sg13g2_o21ai_1 _17738_ (.B1(_02758_),
    .Y(_01460_),
    .A1(net6448),
    .A2(net7186));
 sg13g2_nand2_1 _17739_ (.Y(_02759_),
    .A(net3629),
    .B(net6449));
 sg13g2_o21ai_1 _17740_ (.B1(_02759_),
    .Y(_01461_),
    .A1(net6449),
    .A2(net7483));
 sg13g2_nand2_1 _17741_ (.Y(_02760_),
    .A(net4368),
    .B(net6448));
 sg13g2_o21ai_1 _17742_ (.B1(_02760_),
    .Y(_01462_),
    .A1(net6448),
    .A2(net7639));
 sg13g2_nand2_1 _17743_ (.Y(_02761_),
    .A(net3081),
    .B(net6446));
 sg13g2_o21ai_1 _17744_ (.B1(_02761_),
    .Y(_01463_),
    .A1(net6446),
    .A2(net7188));
 sg13g2_nand2_1 _17745_ (.Y(_02762_),
    .A(net3559),
    .B(net6446));
 sg13g2_o21ai_1 _17746_ (.B1(_02762_),
    .Y(_01464_),
    .A1(net6447),
    .A2(net7485));
 sg13g2_nand2_1 _17747_ (.Y(_02763_),
    .A(net2463),
    .B(net6447));
 sg13g2_o21ai_1 _17748_ (.B1(_02763_),
    .Y(_01465_),
    .A1(net6446),
    .A2(net7640));
 sg13g2_nand2_1 _17749_ (.Y(_02764_),
    .A(net3127),
    .B(net6444));
 sg13g2_o21ai_1 _17750_ (.B1(_02764_),
    .Y(_01466_),
    .A1(net6444),
    .A2(net7188));
 sg13g2_nand2_1 _17751_ (.Y(_02765_),
    .A(net2965),
    .B(net6445));
 sg13g2_o21ai_1 _17752_ (.B1(_02765_),
    .Y(_01467_),
    .A1(net6444),
    .A2(net7485));
 sg13g2_nand2_1 _17753_ (.Y(_02766_),
    .A(net3535),
    .B(net6445));
 sg13g2_o21ai_1 _17754_ (.B1(_02766_),
    .Y(_01468_),
    .A1(net6444),
    .A2(net7640));
 sg13g2_nand2_1 _17755_ (.Y(_02767_),
    .A(net3715),
    .B(net6442));
 sg13g2_o21ai_1 _17756_ (.B1(_02767_),
    .Y(_01469_),
    .A1(net6442),
    .A2(net7188));
 sg13g2_nand2_1 _17757_ (.Y(_02768_),
    .A(net2935),
    .B(net6443));
 sg13g2_o21ai_1 _17758_ (.B1(_02768_),
    .Y(_01470_),
    .A1(net6442),
    .A2(net7485));
 sg13g2_nand2_1 _17759_ (.Y(_02769_),
    .A(net2863),
    .B(net6443));
 sg13g2_o21ai_1 _17760_ (.B1(_02769_),
    .Y(_01471_),
    .A1(net6442),
    .A2(net7640));
 sg13g2_nand2_1 _17761_ (.Y(_02770_),
    .A(net2732),
    .B(net6440));
 sg13g2_o21ai_1 _17762_ (.B1(_02770_),
    .Y(_01472_),
    .A1(net6440),
    .A2(net7188));
 sg13g2_nand2_1 _17763_ (.Y(_02771_),
    .A(net2529),
    .B(net6440));
 sg13g2_o21ai_1 _17764_ (.B1(_02771_),
    .Y(_01473_),
    .A1(net6440),
    .A2(net7485));
 sg13g2_nand2_1 _17765_ (.Y(_02772_),
    .A(net2904),
    .B(net6441));
 sg13g2_o21ai_1 _17766_ (.B1(_02772_),
    .Y(_01474_),
    .A1(net6441),
    .A2(net7640));
 sg13g2_nand2_1 _17767_ (.Y(_02773_),
    .A(net2772),
    .B(net6894));
 sg13g2_o21ai_1 _17768_ (.B1(_02773_),
    .Y(_01475_),
    .A1(net6893),
    .A2(net7188));
 sg13g2_nand2_1 _17769_ (.Y(_02774_),
    .A(net3415),
    .B(net6894));
 sg13g2_o21ai_1 _17770_ (.B1(_02774_),
    .Y(_01476_),
    .A1(net6893),
    .A2(net7485));
 sg13g2_nand2_1 _17771_ (.Y(_02775_),
    .A(net3256),
    .B(net6894));
 sg13g2_o21ai_1 _17772_ (.B1(_02775_),
    .Y(_01477_),
    .A1(net6894),
    .A2(net7641));
 sg13g2_nor2_1 _17773_ (.A(net4692),
    .B(net6439),
    .Y(_02776_));
 sg13g2_a21oi_1 _17774_ (.A1(net6438),
    .A2(net7142),
    .Y(_01478_),
    .B1(_02776_));
 sg13g2_nor2_1 _17775_ (.A(net4339),
    .B(net6438),
    .Y(_02777_));
 sg13g2_a21oi_1 _17776_ (.A1(net6438),
    .A2(net7436),
    .Y(_01479_),
    .B1(_02777_));
 sg13g2_nor2_1 _17777_ (.A(net4602),
    .B(net6438),
    .Y(_02778_));
 sg13g2_a21oi_1 _17778_ (.A1(net6438),
    .A2(net7598),
    .Y(_01480_),
    .B1(_02778_));
 sg13g2_nand2_1 _17779_ (.Y(_02779_),
    .A(net3924),
    .B(net6891));
 sg13g2_o21ai_1 _17780_ (.B1(_02779_),
    .Y(_01481_),
    .A1(net6891),
    .A2(net7188));
 sg13g2_nand2_1 _17781_ (.Y(_02780_),
    .A(net3913),
    .B(net6892));
 sg13g2_o21ai_1 _17782_ (.B1(_02780_),
    .Y(_01482_),
    .A1(net6892),
    .A2(net7485));
 sg13g2_nand2_1 _17783_ (.Y(_02781_),
    .A(net3322),
    .B(net6892));
 sg13g2_o21ai_1 _17784_ (.B1(_02781_),
    .Y(_01483_),
    .A1(net6892),
    .A2(net7641));
 sg13g2_nand2_1 _17785_ (.Y(_02782_),
    .A(net3842),
    .B(net6889));
 sg13g2_o21ai_1 _17786_ (.B1(_02782_),
    .Y(_01484_),
    .A1(net6889),
    .A2(net7188));
 sg13g2_nand2_1 _17787_ (.Y(_02783_),
    .A(net4003),
    .B(net6890));
 sg13g2_o21ai_1 _17788_ (.B1(_02783_),
    .Y(_01485_),
    .A1(net6890),
    .A2(net7485));
 sg13g2_nand2_1 _17789_ (.Y(_02784_),
    .A(net4508),
    .B(net6890));
 sg13g2_o21ai_1 _17790_ (.B1(_02784_),
    .Y(_01486_),
    .A1(net6890),
    .A2(net7640));
 sg13g2_nand2_1 _17791_ (.Y(_02785_),
    .A(net2516),
    .B(net6887));
 sg13g2_o21ai_1 _17792_ (.B1(_02785_),
    .Y(_01487_),
    .A1(net6887),
    .A2(net7173));
 sg13g2_nand2_1 _17793_ (.Y(_02786_),
    .A(net3750),
    .B(net6887));
 sg13g2_o21ai_1 _17794_ (.B1(_02786_),
    .Y(_01488_),
    .A1(net6887),
    .A2(net7469));
 sg13g2_nand2_1 _17795_ (.Y(_02787_),
    .A(net3061),
    .B(net6887));
 sg13g2_o21ai_1 _17796_ (.B1(_02787_),
    .Y(_01489_),
    .A1(net6888),
    .A2(net7634));
 sg13g2_nand2_1 _17797_ (.Y(_02788_),
    .A(net2722),
    .B(net6885));
 sg13g2_o21ai_1 _17798_ (.B1(_02788_),
    .Y(_01490_),
    .A1(net6885),
    .A2(net7179));
 sg13g2_nand2_1 _17799_ (.Y(_02789_),
    .A(net3091),
    .B(net6885));
 sg13g2_o21ai_1 _17800_ (.B1(_02789_),
    .Y(_01491_),
    .A1(net6885),
    .A2(net7474));
 sg13g2_nand2_1 _17801_ (.Y(_02790_),
    .A(net3387),
    .B(net6885));
 sg13g2_o21ai_1 _17802_ (.B1(_02790_),
    .Y(_01492_),
    .A1(net6885),
    .A2(net7639));
 sg13g2_nand2_1 _17803_ (.Y(_02791_),
    .A(net3543),
    .B(net6883));
 sg13g2_o21ai_1 _17804_ (.B1(_02791_),
    .Y(_01493_),
    .A1(net6883),
    .A2(net7179));
 sg13g2_nand2_1 _17805_ (.Y(_02792_),
    .A(net3954),
    .B(net6883));
 sg13g2_o21ai_1 _17806_ (.B1(_02792_),
    .Y(_01494_),
    .A1(net6883),
    .A2(net7474));
 sg13g2_nand2_1 _17807_ (.Y(_02793_),
    .A(net3723),
    .B(net6883));
 sg13g2_o21ai_1 _17808_ (.B1(_02793_),
    .Y(_01495_),
    .A1(net6883),
    .A2(net7639));
 sg13g2_nand2_1 _17809_ (.Y(_02794_),
    .A(net2988),
    .B(net6881));
 sg13g2_o21ai_1 _17810_ (.B1(_02794_),
    .Y(_01496_),
    .A1(net6881),
    .A2(net7179));
 sg13g2_nand2_1 _17811_ (.Y(_02795_),
    .A(net2734),
    .B(net6881));
 sg13g2_o21ai_1 _17812_ (.B1(_02795_),
    .Y(_01497_),
    .A1(net6881),
    .A2(net7474));
 sg13g2_nand2_1 _17813_ (.Y(_02796_),
    .A(net4360),
    .B(net6881));
 sg13g2_o21ai_1 _17814_ (.B1(_02796_),
    .Y(_01498_),
    .A1(net6881),
    .A2(net7639));
 sg13g2_nand2_1 _17815_ (.Y(_02797_),
    .A(net2861),
    .B(net6436));
 sg13g2_o21ai_1 _17816_ (.B1(_02797_),
    .Y(_01499_),
    .A1(net6436),
    .A2(net7181));
 sg13g2_nand2_1 _17817_ (.Y(_02798_),
    .A(net2906),
    .B(net6436));
 sg13g2_o21ai_1 _17818_ (.B1(_02798_),
    .Y(_01500_),
    .A1(net6436),
    .A2(net7478));
 sg13g2_nand2_1 _17819_ (.Y(_02799_),
    .A(net2514),
    .B(net6436));
 sg13g2_o21ai_1 _17820_ (.B1(_02799_),
    .Y(_01501_),
    .A1(net6436),
    .A2(net7636));
 sg13g2_nand2_1 _17821_ (.Y(_02800_),
    .A(net3154),
    .B(net6434));
 sg13g2_o21ai_1 _17822_ (.B1(_02800_),
    .Y(_01502_),
    .A1(net6434),
    .A2(net7181));
 sg13g2_nand2_1 _17823_ (.Y(_02801_),
    .A(net2982),
    .B(net6434));
 sg13g2_o21ai_1 _17824_ (.B1(_02801_),
    .Y(_01503_),
    .A1(net6434),
    .A2(net7478));
 sg13g2_nand2_1 _17825_ (.Y(_02802_),
    .A(net2909),
    .B(net6434));
 sg13g2_o21ai_1 _17826_ (.B1(_02802_),
    .Y(_01504_),
    .A1(net6434),
    .A2(net7639));
 sg13g2_nand2_1 _17827_ (.Y(_02803_),
    .A(net3496),
    .B(net6432));
 sg13g2_o21ai_1 _17828_ (.B1(_02803_),
    .Y(_01505_),
    .A1(net6432),
    .A2(net7181));
 sg13g2_nand2_1 _17829_ (.Y(_02804_),
    .A(net3711),
    .B(net6432));
 sg13g2_o21ai_1 _17830_ (.B1(_02804_),
    .Y(_01506_),
    .A1(net6432),
    .A2(net7478));
 sg13g2_nand2_1 _17831_ (.Y(_02805_),
    .A(net3082),
    .B(net6432));
 sg13g2_o21ai_1 _17832_ (.B1(_02805_),
    .Y(_01507_),
    .A1(net6432),
    .A2(net7639));
 sg13g2_nor2_1 _17833_ (.A(net4002),
    .B(net6431),
    .Y(_02806_));
 sg13g2_a21oi_1 _17834_ (.A1(net6430),
    .A2(net7142),
    .Y(_01508_),
    .B1(_02806_));
 sg13g2_nor2_1 _17835_ (.A(net4223),
    .B(net6430),
    .Y(_02807_));
 sg13g2_a21oi_1 _17836_ (.A1(net6430),
    .A2(net7436),
    .Y(_01509_),
    .B1(_02807_));
 sg13g2_nor2_1 _17837_ (.A(net4599),
    .B(net6430),
    .Y(_02808_));
 sg13g2_a21oi_1 _17838_ (.A1(net6430),
    .A2(net7598),
    .Y(_01510_),
    .B1(_02808_));
 sg13g2_nand2_1 _17839_ (.Y(_02809_),
    .A(net2629),
    .B(net6880));
 sg13g2_o21ai_1 _17840_ (.B1(_02809_),
    .Y(_01511_),
    .A1(net6879),
    .A2(net7180));
 sg13g2_nand2_1 _17841_ (.Y(_02810_),
    .A(net3900),
    .B(net6880));
 sg13g2_o21ai_1 _17842_ (.B1(_02810_),
    .Y(_01512_),
    .A1(net6880),
    .A2(net7474));
 sg13g2_nand2_1 _17843_ (.Y(_02811_),
    .A(net2512),
    .B(net6879));
 sg13g2_o21ai_1 _17844_ (.B1(_02811_),
    .Y(_01513_),
    .A1(net6879),
    .A2(net7634));
 sg13g2_nand2_1 _17845_ (.Y(_02812_),
    .A(net3630),
    .B(net6878));
 sg13g2_o21ai_1 _17846_ (.B1(_02812_),
    .Y(_01514_),
    .A1(net6877),
    .A2(net7179));
 sg13g2_nand2_1 _17847_ (.Y(_02813_),
    .A(net2458),
    .B(net6878));
 sg13g2_o21ai_1 _17848_ (.B1(_02813_),
    .Y(_01515_),
    .A1(net6878),
    .A2(net7474));
 sg13g2_nand2_1 _17849_ (.Y(_02814_),
    .A(net2956),
    .B(net6878));
 sg13g2_o21ai_1 _17850_ (.B1(_02814_),
    .Y(_01516_),
    .A1(net6877),
    .A2(net7634));
 sg13g2_nand2_1 _17851_ (.Y(_02815_),
    .A(net4096),
    .B(net6876));
 sg13g2_o21ai_1 _17852_ (.B1(_02815_),
    .Y(_01517_),
    .A1(net6875),
    .A2(net7179));
 sg13g2_nand2_1 _17853_ (.Y(_02816_),
    .A(net2513),
    .B(net6876));
 sg13g2_o21ai_1 _17854_ (.B1(_02816_),
    .Y(_01518_),
    .A1(net6876),
    .A2(net7474));
 sg13g2_nand2_1 _17855_ (.Y(_02817_),
    .A(net3350),
    .B(net6876));
 sg13g2_o21ai_1 _17856_ (.B1(_02817_),
    .Y(_01519_),
    .A1(net6875),
    .A2(net7634));
 sg13g2_nand2_1 _17857_ (.Y(_02818_),
    .A(net4161),
    .B(net6868));
 sg13g2_o21ai_1 _17858_ (.B1(_02818_),
    .Y(_01520_),
    .A1(net6867),
    .A2(net7179));
 sg13g2_nand2_1 _17859_ (.Y(_02819_),
    .A(net3352),
    .B(net6868));
 sg13g2_o21ai_1 _17860_ (.B1(_02819_),
    .Y(_01521_),
    .A1(net6868),
    .A2(net7474));
 sg13g2_nand2_1 _17861_ (.Y(_02820_),
    .A(net3677),
    .B(net6868));
 sg13g2_o21ai_1 _17862_ (.B1(_02820_),
    .Y(_01522_),
    .A1(net6867),
    .A2(net7634));
 sg13g2_nor2_1 _17863_ (.A(net4219),
    .B(net6428),
    .Y(_02821_));
 sg13g2_a21oi_1 _17864_ (.A1(net6428),
    .A2(net7119),
    .Y(_01523_),
    .B1(_02821_));
 sg13g2_nor2_1 _17865_ (.A(net4819),
    .B(net6428),
    .Y(_02822_));
 sg13g2_a21oi_1 _17866_ (.A1(net6428),
    .A2(net7413),
    .Y(_01524_),
    .B1(_02822_));
 sg13g2_nor2_1 _17867_ (.A(net3853),
    .B(net6428),
    .Y(_02823_));
 sg13g2_a21oi_1 _17868_ (.A1(net6428),
    .A2(net7574),
    .Y(_01525_),
    .B1(_02823_));
 sg13g2_nor2_1 _17869_ (.A(net4605),
    .B(net6426),
    .Y(_02824_));
 sg13g2_a21oi_1 _17870_ (.A1(net6426),
    .A2(net7119),
    .Y(_01526_),
    .B1(_02824_));
 sg13g2_nor2_1 _17871_ (.A(net4503),
    .B(net6426),
    .Y(_02825_));
 sg13g2_a21oi_1 _17872_ (.A1(net6426),
    .A2(net7413),
    .Y(_01527_),
    .B1(_02825_));
 sg13g2_nor2_1 _17873_ (.A(net4369),
    .B(net6426),
    .Y(_02826_));
 sg13g2_a21oi_1 _17874_ (.A1(net6426),
    .A2(net7574),
    .Y(_01528_),
    .B1(_02826_));
 sg13g2_nor2_1 _17875_ (.A(net3712),
    .B(net6422),
    .Y(_02827_));
 sg13g2_a21oi_1 _17876_ (.A1(net6422),
    .A2(net7119),
    .Y(_01529_),
    .B1(_02827_));
 sg13g2_nor2_1 _17877_ (.A(net4774),
    .B(net6422),
    .Y(_02828_));
 sg13g2_a21oi_1 _17878_ (.A1(net6422),
    .A2(net7413),
    .Y(_01530_),
    .B1(_02828_));
 sg13g2_nor2_1 _17879_ (.A(net4335),
    .B(net6422),
    .Y(_02829_));
 sg13g2_a21oi_1 _17880_ (.A1(net6422),
    .A2(net7574),
    .Y(_01531_),
    .B1(_02829_));
 sg13g2_nor2_1 _17881_ (.A(net4416),
    .B(net6420),
    .Y(_02830_));
 sg13g2_a21oi_1 _17882_ (.A1(net6420),
    .A2(net7119),
    .Y(_01532_),
    .B1(_02830_));
 sg13g2_nor2_1 _17883_ (.A(net4516),
    .B(net6420),
    .Y(_02831_));
 sg13g2_a21oi_1 _17884_ (.A1(net6420),
    .A2(net7414),
    .Y(_01533_),
    .B1(_02831_));
 sg13g2_nor2_1 _17885_ (.A(net4174),
    .B(net6420),
    .Y(_02832_));
 sg13g2_a21oi_1 _17886_ (.A1(net6420),
    .A2(net7574),
    .Y(_01534_),
    .B1(_02832_));
 sg13g2_nor2_1 _17887_ (.A(net4557),
    .B(net6418),
    .Y(_02833_));
 sg13g2_a21oi_1 _17888_ (.A1(net6418),
    .A2(net7122),
    .Y(_01535_),
    .B1(_02833_));
 sg13g2_nor2_1 _17889_ (.A(net4053),
    .B(net6419),
    .Y(_02834_));
 sg13g2_a21oi_1 _17890_ (.A1(net6419),
    .A2(net7419),
    .Y(_01536_),
    .B1(_02834_));
 sg13g2_nor2_1 _17891_ (.A(net4408),
    .B(net6418),
    .Y(_02835_));
 sg13g2_a21oi_1 _17892_ (.A1(net6418),
    .A2(net7575),
    .Y(_01537_),
    .B1(_02835_));
 sg13g2_nor2_1 _17893_ (.A(net4718),
    .B(net6415),
    .Y(_02836_));
 sg13g2_a21oi_1 _17894_ (.A1(net6414),
    .A2(net7142),
    .Y(_01538_),
    .B1(_02836_));
 sg13g2_nor2_1 _17895_ (.A(net4439),
    .B(net6414),
    .Y(_02837_));
 sg13g2_a21oi_1 _17896_ (.A1(net6414),
    .A2(net7436),
    .Y(_01539_),
    .B1(_02837_));
 sg13g2_nor2_1 _17897_ (.A(net4748),
    .B(net6414),
    .Y(_02838_));
 sg13g2_a21oi_1 _17898_ (.A1(net6414),
    .A2(net7597),
    .Y(_01540_),
    .B1(_02838_));
 sg13g2_nor2_1 _17899_ (.A(net4670),
    .B(net6412),
    .Y(_02839_));
 sg13g2_a21oi_1 _17900_ (.A1(net6412),
    .A2(net7122),
    .Y(_01541_),
    .B1(_02839_));
 sg13g2_nor2_1 _17901_ (.A(net4543),
    .B(net6413),
    .Y(_02840_));
 sg13g2_a21oi_1 _17902_ (.A1(net6413),
    .A2(net7419),
    .Y(_01542_),
    .B1(_02840_));
 sg13g2_nor2_1 _17903_ (.A(net4509),
    .B(net6412),
    .Y(_02841_));
 sg13g2_a21oi_1 _17904_ (.A1(net6412),
    .A2(net7575),
    .Y(_01543_),
    .B1(_02841_));
 sg13g2_nand2_1 _17905_ (.Y(_02842_),
    .A(net3812),
    .B(net6410));
 sg13g2_o21ai_1 _17906_ (.B1(_02842_),
    .Y(_01544_),
    .A1(net6410),
    .A2(net7122));
 sg13g2_nand2_1 _17907_ (.Y(_02843_),
    .A(net2569),
    .B(net6411));
 sg13g2_o21ai_1 _17908_ (.B1(_02843_),
    .Y(_01545_),
    .A1(net6411),
    .A2(net7419));
 sg13g2_nand2_1 _17909_ (.Y(_02844_),
    .A(net2678),
    .B(net6410));
 sg13g2_o21ai_1 _17910_ (.B1(_02844_),
    .Y(_01546_),
    .A1(net6410),
    .A2(net7576));
 sg13g2_nor2_1 _17911_ (.A(net3882),
    .B(net6408),
    .Y(_02845_));
 sg13g2_a21oi_1 _17912_ (.A1(net6408),
    .A2(net7120),
    .Y(_01547_),
    .B1(_02845_));
 sg13g2_nor2_1 _17913_ (.A(net4535),
    .B(net6408),
    .Y(_02846_));
 sg13g2_a21oi_1 _17914_ (.A1(net6408),
    .A2(net7415),
    .Y(_01548_),
    .B1(_02846_));
 sg13g2_nor2_1 _17915_ (.A(net3696),
    .B(net6408),
    .Y(_02847_));
 sg13g2_a21oi_1 _17916_ (.A1(net6408),
    .A2(net7575),
    .Y(_01549_),
    .B1(_02847_));
 sg13g2_nor2_1 _17917_ (.A(net4716),
    .B(net6398),
    .Y(_02848_));
 sg13g2_a21oi_1 _17918_ (.A1(net6398),
    .A2(net7120),
    .Y(_01550_),
    .B1(_02848_));
 sg13g2_nor2_1 _17919_ (.A(net4547),
    .B(net6398),
    .Y(_02849_));
 sg13g2_a21oi_1 _17920_ (.A1(net6398),
    .A2(net7415),
    .Y(_01551_),
    .B1(_02849_));
 sg13g2_nor2_1 _17921_ (.A(net4493),
    .B(net6398),
    .Y(_02850_));
 sg13g2_a21oi_1 _17922_ (.A1(net6398),
    .A2(net7576),
    .Y(_01552_),
    .B1(_02850_));
 sg13g2_nor2_1 _17923_ (.A(net4415),
    .B(net6394),
    .Y(_02851_));
 sg13g2_a21oi_1 _17924_ (.A1(net6394),
    .A2(net7121),
    .Y(_01553_),
    .B1(_02851_));
 sg13g2_nor2_1 _17925_ (.A(net4650),
    .B(net6394),
    .Y(_02852_));
 sg13g2_a21oi_1 _17926_ (.A1(net6394),
    .A2(net7415),
    .Y(_01554_),
    .B1(_02852_));
 sg13g2_nor2_1 _17927_ (.A(net4571),
    .B(net6394),
    .Y(_02853_));
 sg13g2_a21oi_1 _17928_ (.A1(net6394),
    .A2(net7575),
    .Y(_01555_),
    .B1(_02853_));
 sg13g2_nor2_1 _17929_ (.A(net3449),
    .B(net6392),
    .Y(_02854_));
 sg13g2_a21oi_1 _17930_ (.A1(net6392),
    .A2(net7121),
    .Y(_01556_),
    .B1(_02854_));
 sg13g2_nor2_1 _17931_ (.A(net3817),
    .B(net6392),
    .Y(_02855_));
 sg13g2_a21oi_1 _17932_ (.A1(net6392),
    .A2(net7415),
    .Y(_01557_),
    .B1(_02855_));
 sg13g2_nor2_1 _17933_ (.A(net4387),
    .B(net6392),
    .Y(_02856_));
 sg13g2_a21oi_1 _17934_ (.A1(net6392),
    .A2(net7576),
    .Y(_01558_),
    .B1(_02856_));
 sg13g2_nor2_1 _17935_ (.A(net3612),
    .B(net6469),
    .Y(_02857_));
 sg13g2_a21oi_1 _17936_ (.A1(net6469),
    .A2(net7120),
    .Y(_01559_),
    .B1(_02857_));
 sg13g2_nor2_1 _17937_ (.A(net4785),
    .B(net6468),
    .Y(_02858_));
 sg13g2_a21oi_1 _17938_ (.A1(net6468),
    .A2(net7415),
    .Y(_01560_),
    .B1(_02858_));
 sg13g2_nor2_1 _17939_ (.A(net4444),
    .B(net6468),
    .Y(_02859_));
 sg13g2_a21oi_1 _17940_ (.A1(net6468),
    .A2(net7574),
    .Y(_01561_),
    .B1(_02859_));
 sg13g2_nor2_1 _17941_ (.A(net4584),
    .B(net6467),
    .Y(_02860_));
 sg13g2_a21oi_1 _17942_ (.A1(net6467),
    .A2(net7120),
    .Y(_01562_),
    .B1(_02860_));
 sg13g2_nor2_1 _17943_ (.A(net4655),
    .B(net6466),
    .Y(_02861_));
 sg13g2_a21oi_1 _17944_ (.A1(net6466),
    .A2(net7415),
    .Y(_01563_),
    .B1(_02861_));
 sg13g2_nor2_1 _17945_ (.A(net4420),
    .B(net6466),
    .Y(_02862_));
 sg13g2_a21oi_1 _17946_ (.A1(net6466),
    .A2(net7575),
    .Y(_01564_),
    .B1(_02862_));
 sg13g2_nor2_1 _17947_ (.A(net4701),
    .B(net6465),
    .Y(_02863_));
 sg13g2_a21oi_1 _17948_ (.A1(net6465),
    .A2(net7120),
    .Y(_01565_),
    .B1(_02863_));
 sg13g2_nor2_1 _17949_ (.A(net4450),
    .B(net6464),
    .Y(_02864_));
 sg13g2_a21oi_1 _17950_ (.A1(net6464),
    .A2(net7415),
    .Y(_01566_),
    .B1(_02864_));
 sg13g2_nor2_1 _17951_ (.A(net4331),
    .B(net6464),
    .Y(_02865_));
 sg13g2_a21oi_1 _17952_ (.A1(net6464),
    .A2(net7575),
    .Y(_01567_),
    .B1(_02865_));
 sg13g2_nand2_1 _17953_ (.Y(_02866_),
    .A(net3510),
    .B(net6901));
 sg13g2_o21ai_1 _17954_ (.B1(_02866_),
    .Y(_01568_),
    .A1(net6900),
    .A2(net7142));
 sg13g2_nand2_1 _17955_ (.Y(_02867_),
    .A(net2952),
    .B(net6900));
 sg13g2_o21ai_1 _17956_ (.B1(_02867_),
    .Y(_01569_),
    .A1(net6900),
    .A2(net7436));
 sg13g2_nand2_1 _17957_ (.Y(_02868_),
    .A(net3569),
    .B(net6900));
 sg13g2_o21ai_1 _17958_ (.B1(_02868_),
    .Y(_01570_),
    .A1(net6900),
    .A2(net7597));
 sg13g2_nor2_1 _17959_ (.A(net4715),
    .B(net6463),
    .Y(_02869_));
 sg13g2_a21oi_1 _17960_ (.A1(net6463),
    .A2(net7136),
    .Y(_01571_),
    .B1(_02869_));
 sg13g2_nor2_1 _17961_ (.A(net4733),
    .B(net6462),
    .Y(_02870_));
 sg13g2_a21oi_1 _17962_ (.A1(net6462),
    .A2(net7430),
    .Y(_01572_),
    .B1(_02870_));
 sg13g2_nor2_1 _17963_ (.A(net4060),
    .B(net6462),
    .Y(_02871_));
 sg13g2_a21oi_1 _17964_ (.A1(net6462),
    .A2(net7590),
    .Y(_01573_),
    .B1(_02871_));
 sg13g2_nor2_1 _17965_ (.A(net4343),
    .B(net6461),
    .Y(_02872_));
 sg13g2_a21oi_1 _17966_ (.A1(net6461),
    .A2(net7136),
    .Y(_01574_),
    .B1(_02872_));
 sg13g2_nor2_1 _17967_ (.A(net4381),
    .B(net6460),
    .Y(_02873_));
 sg13g2_a21oi_1 _17968_ (.A1(net6460),
    .A2(net7430),
    .Y(_01575_),
    .B1(_02873_));
 sg13g2_nor2_1 _17969_ (.A(net4471),
    .B(net6460),
    .Y(_02874_));
 sg13g2_a21oi_1 _17970_ (.A1(net6460),
    .A2(net7590),
    .Y(_01576_),
    .B1(_02874_));
 sg13g2_nor2_1 _17971_ (.A(net4544),
    .B(net6485),
    .Y(_02875_));
 sg13g2_a21oi_1 _17972_ (.A1(net6485),
    .A2(net7136),
    .Y(_01577_),
    .B1(_02875_));
 sg13g2_nor2_1 _17973_ (.A(net4375),
    .B(net6484),
    .Y(_02876_));
 sg13g2_a21oi_1 _17974_ (.A1(net6484),
    .A2(net7430),
    .Y(_01578_),
    .B1(_02876_));
 sg13g2_nor2_1 _17975_ (.A(net4337),
    .B(net6484),
    .Y(_02877_));
 sg13g2_a21oi_1 _17976_ (.A1(net6484),
    .A2(net7590),
    .Y(_01579_),
    .B1(_02877_));
 sg13g2_nor2_1 _17977_ (.A(net4553),
    .B(net6483),
    .Y(_02878_));
 sg13g2_a21oi_1 _17978_ (.A1(net6483),
    .A2(net7136),
    .Y(_01580_),
    .B1(_02878_));
 sg13g2_nor2_1 _17979_ (.A(net4130),
    .B(net6482),
    .Y(_02879_));
 sg13g2_a21oi_1 _17980_ (.A1(net6482),
    .A2(net7430),
    .Y(_01581_),
    .B1(_02879_));
 sg13g2_nor2_1 _17981_ (.A(net4475),
    .B(net6482),
    .Y(_02880_));
 sg13g2_a21oi_1 _17982_ (.A1(net6482),
    .A2(net7590),
    .Y(_01582_),
    .B1(_02880_));
 sg13g2_nor2_1 _17983_ (.A(net4624),
    .B(net6481),
    .Y(_02881_));
 sg13g2_a21oi_1 _17984_ (.A1(net6481),
    .A2(net7138),
    .Y(_01583_),
    .B1(_02881_));
 sg13g2_nor2_1 _17985_ (.A(net4313),
    .B(net6480),
    .Y(_02882_));
 sg13g2_a21oi_1 _17986_ (.A1(net6480),
    .A2(net7432),
    .Y(_01584_),
    .B1(_02882_));
 sg13g2_nor2_1 _17987_ (.A(net4734),
    .B(net6480),
    .Y(_02883_));
 sg13g2_a21oi_1 _17988_ (.A1(net6480),
    .A2(net7592),
    .Y(_01585_),
    .B1(_02883_));
 sg13g2_nand2_1 _17989_ (.Y(_02884_),
    .A(net2641),
    .B(net6479));
 sg13g2_o21ai_1 _17990_ (.B1(_02884_),
    .Y(_01586_),
    .A1(net6479),
    .A2(net7138));
 sg13g2_nand2_1 _17991_ (.Y(_02885_),
    .A(net3799),
    .B(net6478));
 sg13g2_o21ai_1 _17992_ (.B1(_02885_),
    .Y(_01587_),
    .A1(net6478),
    .A2(net7432));
 sg13g2_nand2_1 _17993_ (.Y(_02886_),
    .A(net4227),
    .B(net6478));
 sg13g2_o21ai_1 _17994_ (.B1(_02886_),
    .Y(_01588_),
    .A1(net6478),
    .A2(net7592));
 sg13g2_nand2_1 _17995_ (.Y(_02887_),
    .A(net3214),
    .B(net6477));
 sg13g2_o21ai_1 _17996_ (.B1(_02887_),
    .Y(_01589_),
    .A1(net6477),
    .A2(net7138));
 sg13g2_nand2_1 _17997_ (.Y(_02888_),
    .A(net2838),
    .B(net6477));
 sg13g2_o21ai_1 _17998_ (.B1(_02888_),
    .Y(_01590_),
    .A1(net6477),
    .A2(net7432));
 sg13g2_nand2_1 _17999_ (.Y(_02889_),
    .A(net2640),
    .B(net6476));
 sg13g2_o21ai_1 _18000_ (.B1(_02889_),
    .Y(_01591_),
    .A1(net6476),
    .A2(net7592));
 sg13g2_nand2_1 _18001_ (.Y(_02890_),
    .A(net3021),
    .B(net6475));
 sg13g2_o21ai_1 _18002_ (.B1(_02890_),
    .Y(_01592_),
    .A1(net6475),
    .A2(net7138));
 sg13g2_nand2_1 _18003_ (.Y(_02891_),
    .A(net3992),
    .B(net6474));
 sg13g2_o21ai_1 _18004_ (.B1(_02891_),
    .Y(_01593_),
    .A1(net6474),
    .A2(net7432));
 sg13g2_nand2_1 _18005_ (.Y(_02892_),
    .A(net2831),
    .B(net6474));
 sg13g2_o21ai_1 _18006_ (.B1(_02892_),
    .Y(_01594_),
    .A1(net6474),
    .A2(net7592));
 sg13g2_nor2_1 _18007_ (.A(net4636),
    .B(net6473),
    .Y(_02893_));
 sg13g2_a21oi_1 _18008_ (.A1(net6473),
    .A2(net7137),
    .Y(_01595_),
    .B1(_02893_));
 sg13g2_nor2_1 _18009_ (.A(net4566),
    .B(net6472),
    .Y(_02894_));
 sg13g2_a21oi_1 _18010_ (.A1(net6472),
    .A2(net7431),
    .Y(_01596_),
    .B1(_02894_));
 sg13g2_nor2_1 _18011_ (.A(net3977),
    .B(net6472),
    .Y(_02895_));
 sg13g2_a21oi_1 _18012_ (.A1(net6472),
    .A2(net7591),
    .Y(_01597_),
    .B1(_02895_));
 sg13g2_nor2_1 _18013_ (.A(net4517),
    .B(net6906),
    .Y(_02896_));
 sg13g2_a21oi_1 _18014_ (.A1(net6906),
    .A2(net7142),
    .Y(_01598_),
    .B1(_02896_));
 sg13g2_nor2_1 _18015_ (.A(net4684),
    .B(net6906),
    .Y(_02897_));
 sg13g2_a21oi_1 _18016_ (.A1(net6906),
    .A2(net7436),
    .Y(_01599_),
    .B1(_02897_));
 sg13g2_nor2_1 _18017_ (.A(net4254),
    .B(net6907),
    .Y(_02898_));
 sg13g2_a21oi_1 _18018_ (.A1(net6907),
    .A2(net7595),
    .Y(_01600_),
    .B1(_02898_));
 sg13g2_nand2_1 _18019_ (.Y(_02899_),
    .A(net2604),
    .B(net6487));
 sg13g2_o21ai_1 _18020_ (.B1(_02899_),
    .Y(_01601_),
    .A1(net6486),
    .A2(net7137));
 sg13g2_nand2_1 _18021_ (.Y(_02900_),
    .A(net2655),
    .B(net6486));
 sg13g2_o21ai_1 _18022_ (.B1(_02900_),
    .Y(_01602_),
    .A1(net6486),
    .A2(net7431));
 sg13g2_nand2_1 _18023_ (.Y(_02901_),
    .A(net2836),
    .B(net6486));
 sg13g2_o21ai_1 _18024_ (.B1(_02901_),
    .Y(_01603_),
    .A1(net6486),
    .A2(net7591));
 sg13g2_nand2_1 _18025_ (.Y(_02902_),
    .A(net2705),
    .B(net6489));
 sg13g2_o21ai_1 _18026_ (.B1(_02902_),
    .Y(_01604_),
    .A1(net6489),
    .A2(net7136));
 sg13g2_nand2_1 _18027_ (.Y(_02903_),
    .A(net3309),
    .B(net6488));
 sg13g2_o21ai_1 _18028_ (.B1(_02903_),
    .Y(_01605_),
    .A1(net6488),
    .A2(net7431));
 sg13g2_nand2_1 _18029_ (.Y(_02904_),
    .A(net2662),
    .B(net6488));
 sg13g2_o21ai_1 _18030_ (.B1(_02904_),
    .Y(_01606_),
    .A1(net6488),
    .A2(net7590));
 sg13g2_nand2_1 _18031_ (.Y(_02905_),
    .A(net2567),
    .B(net6499));
 sg13g2_o21ai_1 _18032_ (.B1(_02905_),
    .Y(_01607_),
    .A1(net6499),
    .A2(net7137));
 sg13g2_nand2_1 _18033_ (.Y(_02906_),
    .A(net2760),
    .B(net6498));
 sg13g2_o21ai_1 _18034_ (.B1(_02906_),
    .Y(_01608_),
    .A1(net6498),
    .A2(net7430));
 sg13g2_nand2_1 _18035_ (.Y(_02907_),
    .A(net2925),
    .B(net6498));
 sg13g2_o21ai_1 _18036_ (.B1(_02907_),
    .Y(_01609_),
    .A1(net6498),
    .A2(net7591));
 sg13g2_nand2_1 _18037_ (.Y(_02908_),
    .A(net3972),
    .B(net6497));
 sg13g2_o21ai_1 _18038_ (.B1(_02908_),
    .Y(_01610_),
    .A1(net6497),
    .A2(net7136));
 sg13g2_nand2_1 _18039_ (.Y(_02909_),
    .A(net2973),
    .B(net6496));
 sg13g2_o21ai_1 _18040_ (.B1(_02909_),
    .Y(_01611_),
    .A1(net6496),
    .A2(net7430));
 sg13g2_nand2_1 _18041_ (.Y(_02910_),
    .A(net3442),
    .B(net6496));
 sg13g2_o21ai_1 _18042_ (.B1(_02910_),
    .Y(_01612_),
    .A1(net6496),
    .A2(net7590));
 sg13g2_nand2_1 _18043_ (.Y(_02911_),
    .A(net3079),
    .B(net6495));
 sg13g2_o21ai_1 _18044_ (.B1(_02911_),
    .Y(_01613_),
    .A1(net6495),
    .A2(net7136));
 sg13g2_nand2_1 _18045_ (.Y(_02912_),
    .A(net3585),
    .B(net6494));
 sg13g2_o21ai_1 _18046_ (.B1(_02912_),
    .Y(_01614_),
    .A1(net6494),
    .A2(net7430));
 sg13g2_nand2_1 _18047_ (.Y(_02913_),
    .A(net3126),
    .B(net6494));
 sg13g2_o21ai_1 _18048_ (.B1(_02913_),
    .Y(_01615_),
    .A1(net6494),
    .A2(net7590));
 sg13g2_nand2_1 _18049_ (.Y(_02914_),
    .A(net3578),
    .B(net6493));
 sg13g2_o21ai_1 _18050_ (.B1(_02914_),
    .Y(_01616_),
    .A1(net6493),
    .A2(net7136));
 sg13g2_nand2_1 _18051_ (.Y(_02915_),
    .A(net2854),
    .B(net6492));
 sg13g2_o21ai_1 _18052_ (.B1(_02915_),
    .Y(_01617_),
    .A1(net6492),
    .A2(net7430));
 sg13g2_nand2_1 _18053_ (.Y(_02916_),
    .A(net2473),
    .B(net6492));
 sg13g2_o21ai_1 _18054_ (.B1(_02916_),
    .Y(_01618_),
    .A1(net6492),
    .A2(net7590));
 sg13g2_nor2_1 _18055_ (.A(net4405),
    .B(net6352),
    .Y(_02917_));
 sg13g2_a21oi_1 _18056_ (.A1(net6353),
    .A2(net7160),
    .Y(_01619_),
    .B1(_02917_));
 sg13g2_nor2_1 _18057_ (.A(net3840),
    .B(net6352),
    .Y(_02918_));
 sg13g2_a21oi_1 _18058_ (.A1(net6352),
    .A2(net7457),
    .Y(_01620_),
    .B1(_02918_));
 sg13g2_nor2_1 _18059_ (.A(net4216),
    .B(net6353),
    .Y(_02919_));
 sg13g2_a21oi_1 _18060_ (.A1(net6353),
    .A2(net7620),
    .Y(_01621_),
    .B1(_02919_));
 sg13g2_nor2_1 _18061_ (.A(net4449),
    .B(net6354),
    .Y(_02920_));
 sg13g2_a21oi_1 _18062_ (.A1(net6355),
    .A2(net7160),
    .Y(_01622_),
    .B1(_02920_));
 sg13g2_nor2_1 _18063_ (.A(net4490),
    .B(net6354),
    .Y(_02921_));
 sg13g2_a21oi_1 _18064_ (.A1(net6354),
    .A2(net7457),
    .Y(_01623_),
    .B1(_02921_));
 sg13g2_nor2_1 _18065_ (.A(net4072),
    .B(net6355),
    .Y(_02922_));
 sg13g2_a21oi_1 _18066_ (.A1(net6355),
    .A2(net7620),
    .Y(_01624_),
    .B1(_02922_));
 sg13g2_nor2_1 _18067_ (.A(net4773),
    .B(net6356),
    .Y(_02923_));
 sg13g2_a21oi_1 _18068_ (.A1(net6357),
    .A2(net7160),
    .Y(_01625_),
    .B1(_02923_));
 sg13g2_nor2_1 _18069_ (.A(net4485),
    .B(net6356),
    .Y(_02924_));
 sg13g2_a21oi_1 _18070_ (.A1(net6356),
    .A2(net7456),
    .Y(_01626_),
    .B1(_02924_));
 sg13g2_nor2_1 _18071_ (.A(net4154),
    .B(net6357),
    .Y(_02925_));
 sg13g2_a21oi_1 _18072_ (.A1(net6357),
    .A2(net7620),
    .Y(_01627_),
    .B1(_02925_));
 sg13g2_nor2_1 _18073_ (.A(net4443),
    .B(net6817),
    .Y(_02926_));
 sg13g2_a21oi_1 _18074_ (.A1(net6817),
    .A2(net7140),
    .Y(_01628_),
    .B1(_02926_));
 sg13g2_nor2_1 _18075_ (.A(net4746),
    .B(net6817),
    .Y(_02927_));
 sg13g2_a21oi_1 _18076_ (.A1(net6817),
    .A2(net7434),
    .Y(_01629_),
    .B1(_02927_));
 sg13g2_nor2_1 _18077_ (.A(net4506),
    .B(net6817),
    .Y(_02928_));
 sg13g2_a21oi_1 _18078_ (.A1(net6817),
    .A2(net7596),
    .Y(_01630_),
    .B1(_02928_));
 sg13g2_nor2_1 _18079_ (.A(net4158),
    .B(net6344),
    .Y(_02929_));
 sg13g2_a21oi_1 _18080_ (.A1(net6344),
    .A2(net7160),
    .Y(_01631_),
    .B1(_02929_));
 sg13g2_nor2_1 _18081_ (.A(net4312),
    .B(net6344),
    .Y(_02930_));
 sg13g2_a21oi_1 _18082_ (.A1(net6344),
    .A2(net7456),
    .Y(_01632_),
    .B1(_02930_));
 sg13g2_nor2_1 _18083_ (.A(net4233),
    .B(net6344),
    .Y(_02931_));
 sg13g2_a21oi_1 _18084_ (.A1(net6344),
    .A2(net7628),
    .Y(_01633_),
    .B1(_02931_));
 sg13g2_nand2_1 _18085_ (.Y(_02932_),
    .A(net2811),
    .B(net6346));
 sg13g2_o21ai_1 _18086_ (.B1(_02932_),
    .Y(_01634_),
    .A1(net6346),
    .A2(net7160));
 sg13g2_nand2_1 _18087_ (.Y(_02933_),
    .A(net4399),
    .B(net6346));
 sg13g2_o21ai_1 _18088_ (.B1(_02933_),
    .Y(_01635_),
    .A1(net6346),
    .A2(net7456));
 sg13g2_nand2_1 _18089_ (.Y(_02934_),
    .A(net3617),
    .B(net6346));
 sg13g2_o21ai_1 _18090_ (.B1(_02934_),
    .Y(_01636_),
    .A1(net6347),
    .A2(net7628));
 sg13g2_nand2_1 _18091_ (.Y(_02935_),
    .A(net2731),
    .B(net6348));
 sg13g2_o21ai_1 _18092_ (.B1(_02935_),
    .Y(_01637_),
    .A1(net6348),
    .A2(net7159));
 sg13g2_nand2_1 _18093_ (.Y(_02936_),
    .A(net2701),
    .B(net6348));
 sg13g2_o21ai_1 _18094_ (.B1(_02936_),
    .Y(_01638_),
    .A1(net6348),
    .A2(net7456));
 sg13g2_nand2_1 _18095_ (.Y(_02937_),
    .A(net4129),
    .B(net6348));
 sg13g2_o21ai_1 _18096_ (.B1(_02937_),
    .Y(_01639_),
    .A1(net6349),
    .A2(net7628));
 sg13g2_nand2_1 _18097_ (.Y(_02938_),
    .A(net2596),
    .B(net6318));
 sg13g2_o21ai_1 _18098_ (.B1(_02938_),
    .Y(_01640_),
    .A1(net6318),
    .A2(net7159));
 sg13g2_nand2_1 _18099_ (.Y(_02939_),
    .A(net4351),
    .B(net6318));
 sg13g2_o21ai_1 _18100_ (.B1(_02939_),
    .Y(_01641_),
    .A1(net6318),
    .A2(net7456));
 sg13g2_nand2_1 _18101_ (.Y(_02940_),
    .A(net2845),
    .B(net6318));
 sg13g2_o21ai_1 _18102_ (.B1(_02940_),
    .Y(_01642_),
    .A1(net6319),
    .A2(net7628));
 sg13g2_nor2_1 _18103_ (.A(net3915),
    .B(net6321),
    .Y(_02941_));
 sg13g2_a21oi_1 _18104_ (.A1(net6321),
    .A2(net7181),
    .Y(_01643_),
    .B1(_02941_));
 sg13g2_nor2_1 _18105_ (.A(net4782),
    .B(net6320),
    .Y(_02942_));
 sg13g2_a21oi_1 _18106_ (.A1(net6320),
    .A2(net7477),
    .Y(_01644_),
    .B1(_02942_));
 sg13g2_nor2_1 _18107_ (.A(net4678),
    .B(net6320),
    .Y(_02943_));
 sg13g2_a21oi_1 _18108_ (.A1(net6320),
    .A2(net7636),
    .Y(_01645_),
    .B1(_02943_));
 sg13g2_nand2_1 _18109_ (.Y(_02944_),
    .A(net3876),
    .B(net6337));
 sg13g2_o21ai_1 _18110_ (.B1(_02944_),
    .Y(_01646_),
    .A1(net6337),
    .A2(net7181));
 sg13g2_nand2_1 _18111_ (.Y(_02945_),
    .A(net2887),
    .B(net6336));
 sg13g2_o21ai_1 _18112_ (.B1(_02945_),
    .Y(_01647_),
    .A1(net6336),
    .A2(net7477));
 sg13g2_nand2_1 _18113_ (.Y(_02946_),
    .A(net4016),
    .B(net6336));
 sg13g2_o21ai_1 _18114_ (.B1(_02946_),
    .Y(_01648_),
    .A1(net6336),
    .A2(net7636));
 sg13g2_nand2_1 _18115_ (.Y(_02947_),
    .A(net3688),
    .B(net6335));
 sg13g2_o21ai_1 _18116_ (.B1(_02947_),
    .Y(_01649_),
    .A1(net6335),
    .A2(net7181));
 sg13g2_nand2_1 _18117_ (.Y(_02948_),
    .A(net3529),
    .B(net6334));
 sg13g2_o21ai_1 _18118_ (.B1(_02948_),
    .Y(_01650_),
    .A1(net6334),
    .A2(net7477));
 sg13g2_nand2_1 _18119_ (.Y(_02949_),
    .A(net3724),
    .B(net6334));
 sg13g2_o21ai_1 _18120_ (.B1(_02949_),
    .Y(_01651_),
    .A1(net6334),
    .A2(net7636));
 sg13g2_nand2_1 _18121_ (.Y(_02950_),
    .A(net3608),
    .B(net6327));
 sg13g2_o21ai_1 _18122_ (.B1(_02950_),
    .Y(_01652_),
    .A1(net6327),
    .A2(net7181));
 sg13g2_nand2_1 _18123_ (.Y(_02951_),
    .A(net3943),
    .B(net6326));
 sg13g2_o21ai_1 _18124_ (.B1(_02951_),
    .Y(_01653_),
    .A1(net6326),
    .A2(net7477));
 sg13g2_nand2_1 _18125_ (.Y(_02952_),
    .A(net3261),
    .B(net6326));
 sg13g2_o21ai_1 _18126_ (.B1(_02952_),
    .Y(_01654_),
    .A1(net6326),
    .A2(net7636));
 sg13g2_nand2_1 _18127_ (.Y(_02953_),
    .A(net3164),
    .B(net6329));
 sg13g2_o21ai_1 _18128_ (.B1(_02953_),
    .Y(_01655_),
    .A1(net6329),
    .A2(net7174));
 sg13g2_nand2_1 _18129_ (.Y(_02954_),
    .A(net3736),
    .B(net6329));
 sg13g2_o21ai_1 _18130_ (.B1(_02954_),
    .Y(_01656_),
    .A1(net6328),
    .A2(net7469));
 sg13g2_nand2_1 _18131_ (.Y(_02955_),
    .A(net3095),
    .B(net6329));
 sg13g2_o21ai_1 _18132_ (.B1(_02955_),
    .Y(_01657_),
    .A1(net6328),
    .A2(net7628));
 sg13g2_nor2_1 _18133_ (.A(net4855),
    .B(net6815),
    .Y(_02956_));
 sg13g2_a21oi_1 _18134_ (.A1(net6815),
    .A2(net7142),
    .Y(_01658_),
    .B1(_02956_));
 sg13g2_nor2_1 _18135_ (.A(net4736),
    .B(net6815),
    .Y(_02957_));
 sg13g2_a21oi_1 _18136_ (.A1(net6815),
    .A2(net7436),
    .Y(_01659_),
    .B1(_02957_));
 sg13g2_nor2_1 _18137_ (.A(net4662),
    .B(net6816),
    .Y(_02958_));
 sg13g2_a21oi_1 _18138_ (.A1(net6816),
    .A2(net7595),
    .Y(_01660_),
    .B1(_02958_));
 sg13g2_nand2_1 _18139_ (.Y(_02959_),
    .A(net3271),
    .B(net6331));
 sg13g2_o21ai_1 _18140_ (.B1(_02959_),
    .Y(_01661_),
    .A1(net6331),
    .A2(net7173));
 sg13g2_nand2_1 _18141_ (.Y(_02960_),
    .A(net3174),
    .B(net6331));
 sg13g2_o21ai_1 _18142_ (.B1(_02960_),
    .Y(_01662_),
    .A1(net6330),
    .A2(net7469));
 sg13g2_nand2_1 _18143_ (.Y(_02961_),
    .A(net4430),
    .B(net6331));
 sg13g2_o21ai_1 _18144_ (.B1(_02961_),
    .Y(_01663_),
    .A1(net6330),
    .A2(net7628));
 sg13g2_nand2_1 _18145_ (.Y(_02962_),
    .A(net3534),
    .B(net6333));
 sg13g2_o21ai_1 _18146_ (.B1(_02962_),
    .Y(_01664_),
    .A1(net6333),
    .A2(net7173));
 sg13g2_nand2_1 _18147_ (.Y(_02963_),
    .A(net2859),
    .B(net6332));
 sg13g2_o21ai_1 _18148_ (.B1(_02963_),
    .Y(_01665_),
    .A1(net6332),
    .A2(net7469));
 sg13g2_nand2_1 _18149_ (.Y(_02964_),
    .A(net3233),
    .B(net6333));
 sg13g2_o21ai_1 _18150_ (.B1(_02964_),
    .Y(_01666_),
    .A1(net6333),
    .A2(net7628));
 sg13g2_nand2_1 _18151_ (.Y(_02965_),
    .A(net3385),
    .B(net6324));
 sg13g2_o21ai_1 _18152_ (.B1(_02965_),
    .Y(_01667_),
    .A1(net6324),
    .A2(net7177));
 sg13g2_nand2_1 _18153_ (.Y(_02966_),
    .A(net2808),
    .B(net6324));
 sg13g2_o21ai_1 _18154_ (.B1(_02966_),
    .Y(_01668_),
    .A1(net6324),
    .A2(net7475));
 sg13g2_nand2_1 _18155_ (.Y(_02967_),
    .A(net3218),
    .B(net6324));
 sg13g2_o21ai_1 _18156_ (.B1(_02967_),
    .Y(_01669_),
    .A1(net6324),
    .A2(net7631));
 sg13g2_nand2_1 _18157_ (.Y(_02968_),
    .A(net3536),
    .B(net6322));
 sg13g2_o21ai_1 _18158_ (.B1(_02968_),
    .Y(_01670_),
    .A1(net6322),
    .A2(net7177));
 sg13g2_nand2_1 _18159_ (.Y(_02969_),
    .A(net3976),
    .B(net6322));
 sg13g2_o21ai_1 _18160_ (.B1(_02969_),
    .Y(_01671_),
    .A1(net6322),
    .A2(net7475));
 sg13g2_nand2_1 _18161_ (.Y(_02970_),
    .A(net3289),
    .B(net6322));
 sg13g2_o21ai_1 _18162_ (.B1(_02970_),
    .Y(_01672_),
    .A1(net6322),
    .A2(net7631));
 sg13g2_nand2_1 _18163_ (.Y(_02971_),
    .A(net3395),
    .B(net6308));
 sg13g2_o21ai_1 _18164_ (.B1(_02971_),
    .Y(_01673_),
    .A1(net6308),
    .A2(net7177));
 sg13g2_nand2_1 _18165_ (.Y(_02972_),
    .A(net4326),
    .B(net6308));
 sg13g2_o21ai_1 _18166_ (.B1(_02972_),
    .Y(_01674_),
    .A1(net6308),
    .A2(net7475));
 sg13g2_nand2_1 _18167_ (.Y(_02973_),
    .A(net2499),
    .B(net6308));
 sg13g2_o21ai_1 _18168_ (.B1(_02973_),
    .Y(_01675_),
    .A1(net6308),
    .A2(net7631));
 sg13g2_nand2_1 _18169_ (.Y(_02974_),
    .A(net3016),
    .B(net6284));
 sg13g2_o21ai_1 _18170_ (.B1(_02974_),
    .Y(_01676_),
    .A1(net6284),
    .A2(net7177));
 sg13g2_nand2_1 _18171_ (.Y(_02975_),
    .A(net2865),
    .B(net6284));
 sg13g2_o21ai_1 _18172_ (.B1(_02975_),
    .Y(_01677_),
    .A1(net6284),
    .A2(net7475));
 sg13g2_nand2_1 _18173_ (.Y(_02976_),
    .A(net2866),
    .B(net6284));
 sg13g2_o21ai_1 _18174_ (.B1(_02976_),
    .Y(_01678_),
    .A1(net6284),
    .A2(net7631));
 sg13g2_nand2_1 _18175_ (.Y(_02977_),
    .A(net3826),
    .B(net6286));
 sg13g2_o21ai_1 _18176_ (.B1(_02977_),
    .Y(_01679_),
    .A1(net6286),
    .A2(net7176));
 sg13g2_nand2_1 _18177_ (.Y(_02978_),
    .A(net3521),
    .B(net6286));
 sg13g2_o21ai_1 _18178_ (.B1(_02978_),
    .Y(_01680_),
    .A1(net6287),
    .A2(net7472));
 sg13g2_nand2_1 _18179_ (.Y(_02979_),
    .A(net3421),
    .B(net6286));
 sg13g2_o21ai_1 _18180_ (.B1(_02979_),
    .Y(_01681_),
    .A1(net6287),
    .A2(net7632));
 sg13g2_nand2_1 _18181_ (.Y(_02980_),
    .A(net3881),
    .B(net6288));
 sg13g2_o21ai_1 _18182_ (.B1(_02980_),
    .Y(_01682_),
    .A1(net6288),
    .A2(net7176));
 sg13g2_nand2_1 _18183_ (.Y(_02981_),
    .A(net2623),
    .B(net6288));
 sg13g2_o21ai_1 _18184_ (.B1(_02981_),
    .Y(_01683_),
    .A1(net6289),
    .A2(net7472));
 sg13g2_nand2_1 _18185_ (.Y(_02982_),
    .A(net3967),
    .B(net6288));
 sg13g2_o21ai_1 _18186_ (.B1(_02982_),
    .Y(_01684_),
    .A1(net6289),
    .A2(net7632));
 sg13g2_nand2_1 _18187_ (.Y(_02983_),
    .A(net3804),
    .B(net6290));
 sg13g2_o21ai_1 _18188_ (.B1(_02983_),
    .Y(_01685_),
    .A1(net6290),
    .A2(net7176));
 sg13g2_nand2_1 _18189_ (.Y(_02984_),
    .A(net3250),
    .B(net6290));
 sg13g2_o21ai_1 _18190_ (.B1(_02984_),
    .Y(_01686_),
    .A1(net6291),
    .A2(net7472));
 sg13g2_nand2_1 _18191_ (.Y(_02985_),
    .A(net3394),
    .B(net6290));
 sg13g2_o21ai_1 _18192_ (.B1(_02985_),
    .Y(_01687_),
    .A1(net6291),
    .A2(net7632));
 sg13g2_nand2_1 _18193_ (.Y(_02986_),
    .A(net2743),
    .B(net6310));
 sg13g2_o21ai_1 _18194_ (.B1(_02986_),
    .Y(_01688_),
    .A1(net6310),
    .A2(net7142));
 sg13g2_nand2_1 _18195_ (.Y(_02987_),
    .A(net2884),
    .B(net6310));
 sg13g2_o21ai_1 _18196_ (.B1(_02987_),
    .Y(_01689_),
    .A1(net6310),
    .A2(net7436));
 sg13g2_nand2_1 _18197_ (.Y(_02988_),
    .A(net3143),
    .B(net6310));
 sg13g2_o21ai_1 _18198_ (.B1(_02988_),
    .Y(_01690_),
    .A1(net6311),
    .A2(net7595));
 sg13g2_nand2_1 _18199_ (.Y(_02989_),
    .A(net2970),
    .B(net6312));
 sg13g2_o21ai_1 _18200_ (.B1(_02989_),
    .Y(_01691_),
    .A1(net6312),
    .A2(net7175));
 sg13g2_nand2_1 _18201_ (.Y(_02990_),
    .A(net3453),
    .B(net6313));
 sg13g2_o21ai_1 _18202_ (.B1(_02990_),
    .Y(_01692_),
    .A1(net6313),
    .A2(net7471));
 sg13g2_nand2_1 _18203_ (.Y(_02991_),
    .A(net2985),
    .B(net6312));
 sg13g2_o21ai_1 _18204_ (.B1(_02991_),
    .Y(_01693_),
    .A1(net6312),
    .A2(net7631));
 sg13g2_nand2_1 _18205_ (.Y(_02992_),
    .A(net4014),
    .B(net6314));
 sg13g2_o21ai_1 _18206_ (.B1(_02992_),
    .Y(_01694_),
    .A1(net6314),
    .A2(net7175));
 sg13g2_nand2_1 _18207_ (.Y(_02993_),
    .A(net2791),
    .B(net6315));
 sg13g2_o21ai_1 _18208_ (.B1(_02993_),
    .Y(_01695_),
    .A1(net6315),
    .A2(net7471));
 sg13g2_nand2_1 _18209_ (.Y(_02994_),
    .A(net3818),
    .B(net6314));
 sg13g2_o21ai_1 _18210_ (.B1(_02994_),
    .Y(_01696_),
    .A1(net6314),
    .A2(net7631));
 sg13g2_nand2_1 _18211_ (.Y(_02995_),
    .A(net2450),
    .B(net6316));
 sg13g2_o21ai_1 _18212_ (.B1(_02995_),
    .Y(_01697_),
    .A1(net6316),
    .A2(net7175));
 sg13g2_nand2_1 _18213_ (.Y(_02996_),
    .A(net4580),
    .B(net6317));
 sg13g2_o21ai_1 _18214_ (.B1(_02996_),
    .Y(_01698_),
    .A1(net6317),
    .A2(net7471));
 sg13g2_nand2_1 _18215_ (.Y(_02997_),
    .A(net3938),
    .B(net6316));
 sg13g2_o21ai_1 _18216_ (.B1(_02997_),
    .Y(_01699_),
    .A1(net6316),
    .A2(net7631));
 sg13g2_nand2_1 _18217_ (.Y(_02998_),
    .A(net3993),
    .B(net6292));
 sg13g2_o21ai_1 _18218_ (.B1(_02998_),
    .Y(_01700_),
    .A1(net6292),
    .A2(net7175));
 sg13g2_nand2_1 _18219_ (.Y(_02999_),
    .A(net2834),
    .B(net6293));
 sg13g2_o21ai_1 _18220_ (.B1(_02999_),
    .Y(_01701_),
    .A1(net6293),
    .A2(net7471));
 sg13g2_nand2_1 _18221_ (.Y(_03000_),
    .A(net3867),
    .B(net6292));
 sg13g2_o21ai_1 _18222_ (.B1(_03000_),
    .Y(_01702_),
    .A1(net6292),
    .A2(net7631));
 sg13g2_nand2_1 _18223_ (.Y(_03001_),
    .A(net3635),
    .B(net6296));
 sg13g2_o21ai_1 _18224_ (.B1(_03001_),
    .Y(_01703_),
    .A1(net6296),
    .A2(net7176));
 sg13g2_nand2_1 _18225_ (.Y(_03002_),
    .A(net3945),
    .B(net6296));
 sg13g2_o21ai_1 _18226_ (.B1(_03002_),
    .Y(_01704_),
    .A1(net6296),
    .A2(net7473));
 sg13g2_nand2_1 _18227_ (.Y(_03003_),
    .A(net3149),
    .B(net6297));
 sg13g2_o21ai_1 _18228_ (.B1(_03003_),
    .Y(_01705_),
    .A1(net6297),
    .A2(net7633));
 sg13g2_nand2_1 _18229_ (.Y(_03004_),
    .A(net3960),
    .B(net6362));
 sg13g2_o21ai_1 _18230_ (.B1(_03004_),
    .Y(_01706_),
    .A1(net6362),
    .A2(net7176));
 sg13g2_nand2_1 _18231_ (.Y(_03005_),
    .A(net2938),
    .B(net6362));
 sg13g2_o21ai_1 _18232_ (.B1(_03005_),
    .Y(_01707_),
    .A1(net6362),
    .A2(net7473));
 sg13g2_nand2_1 _18233_ (.Y(_03006_),
    .A(net3064),
    .B(net6363));
 sg13g2_o21ai_1 _18234_ (.B1(_03006_),
    .Y(_01708_),
    .A1(net6363),
    .A2(net7633));
 sg13g2_nand2_1 _18235_ (.Y(_03007_),
    .A(net2720),
    .B(net6364));
 sg13g2_o21ai_1 _18236_ (.B1(_03007_),
    .Y(_01709_),
    .A1(net6364),
    .A2(net7176));
 sg13g2_nand2_1 _18237_ (.Y(_03008_),
    .A(net3275),
    .B(net6364));
 sg13g2_o21ai_1 _18238_ (.B1(_03008_),
    .Y(_01710_),
    .A1(net6364),
    .A2(net7473));
 sg13g2_nand2_1 _18239_ (.Y(_03009_),
    .A(net3996),
    .B(net6365));
 sg13g2_o21ai_1 _18240_ (.B1(_03009_),
    .Y(_01711_),
    .A1(net6365),
    .A2(net7633));
 sg13g2_nor2_1 _18241_ (.A(net4426),
    .B(net6366),
    .Y(_03010_));
 sg13g2_a21oi_1 _18242_ (.A1(net6367),
    .A2(net7176),
    .Y(_01712_),
    .B1(_03010_));
 sg13g2_nor2_1 _18243_ (.A(net3897),
    .B(net6366),
    .Y(_03011_));
 sg13g2_a21oi_1 _18244_ (.A1(net6366),
    .A2(net7473),
    .Y(_01713_),
    .B1(_03011_));
 sg13g2_nor2_1 _18245_ (.A(net4180),
    .B(net6366),
    .Y(_03012_));
 sg13g2_a21oi_1 _18246_ (.A1(net6366),
    .A2(net7633),
    .Y(_01714_),
    .B1(_03012_));
 sg13g2_nor2_1 _18247_ (.A(net3441),
    .B(net6829),
    .Y(_03013_));
 sg13g2_a21oi_1 _18248_ (.A1(net6829),
    .A2(net7121),
    .Y(_01715_),
    .B1(_03013_));
 sg13g2_nor2_1 _18249_ (.A(net4274),
    .B(net6829),
    .Y(_03014_));
 sg13g2_a21oi_1 _18250_ (.A1(net6829),
    .A2(net7416),
    .Y(_01716_),
    .B1(_03014_));
 sg13g2_nor2_1 _18251_ (.A(net4826),
    .B(net6829),
    .Y(_03015_));
 sg13g2_a21oi_1 _18252_ (.A1(net6829),
    .A2(net7581),
    .Y(_01717_),
    .B1(_03015_));
 sg13g2_nor2_1 _18253_ (.A(net4194),
    .B(net6753),
    .Y(_03016_));
 sg13g2_a21oi_1 _18254_ (.A1(net7141),
    .A2(net6753),
    .Y(_01718_),
    .B1(_03016_));
 sg13g2_nor2_1 _18255_ (.A(net4259),
    .B(net6754),
    .Y(_03017_));
 sg13g2_a21oi_1 _18256_ (.A1(net7435),
    .A2(net6754),
    .Y(_01719_),
    .B1(_03017_));
 sg13g2_nor2_1 _18257_ (.A(net4152),
    .B(net6754),
    .Y(_03018_));
 sg13g2_a21oi_1 _18258_ (.A1(net7596),
    .A2(net6753),
    .Y(_01720_),
    .B1(_03018_));
 sg13g2_nor2_1 _18259_ (.A(net4775),
    .B(net6755),
    .Y(_03019_));
 sg13g2_a21oi_1 _18260_ (.A1(net7120),
    .A2(net6755),
    .Y(_01721_),
    .B1(_03019_));
 sg13g2_nor2_1 _18261_ (.A(net4479),
    .B(net6755),
    .Y(_03020_));
 sg13g2_a21oi_1 _18262_ (.A1(net7416),
    .A2(net6755),
    .Y(_01722_),
    .B1(_03020_));
 sg13g2_nor2_1 _18263_ (.A(net4772),
    .B(net6755),
    .Y(_03021_));
 sg13g2_a21oi_1 _18264_ (.A1(net7581),
    .A2(net6755),
    .Y(_01723_),
    .B1(_03021_));
 sg13g2_nor2_1 _18265_ (.A(net4240),
    .B(net6757),
    .Y(_03022_));
 sg13g2_a21oi_1 _18266_ (.A1(net7120),
    .A2(net6757),
    .Y(_01724_),
    .B1(_03022_));
 sg13g2_nor2_1 _18267_ (.A(net4562),
    .B(net6757),
    .Y(_03023_));
 sg13g2_a21oi_1 _18268_ (.A1(net7416),
    .A2(net6757),
    .Y(_01725_),
    .B1(_03023_));
 sg13g2_nor2_1 _18269_ (.A(net3984),
    .B(net6757),
    .Y(_03024_));
 sg13g2_a21oi_1 _18270_ (.A1(net7581),
    .A2(net6757),
    .Y(_01726_),
    .B1(_03024_));
 sg13g2_nor2_1 _18271_ (.A(net4652),
    .B(net6300),
    .Y(_03025_));
 sg13g2_a21oi_1 _18272_ (.A1(net6300),
    .A2(net7128),
    .Y(_01727_),
    .B1(_03025_));
 sg13g2_nor2_1 _18273_ (.A(net4040),
    .B(net6300),
    .Y(_03026_));
 sg13g2_a21oi_1 _18274_ (.A1(net6300),
    .A2(net7422),
    .Y(_01728_),
    .B1(_03026_));
 sg13g2_nor2_1 _18275_ (.A(net4210),
    .B(net6301),
    .Y(_03027_));
 sg13g2_a21oi_1 _18276_ (.A1(net6300),
    .A2(net7582),
    .Y(_01729_),
    .B1(_03027_));
 sg13g2_nor2_1 _18277_ (.A(net4413),
    .B(net6266),
    .Y(_03028_));
 sg13g2_a21oi_1 _18278_ (.A1(net7128),
    .A2(net6266),
    .Y(_01730_),
    .B1(_03028_));
 sg13g2_nor2_1 _18279_ (.A(net3926),
    .B(net6267),
    .Y(_03029_));
 sg13g2_a21oi_1 _18280_ (.A1(net7422),
    .A2(net6266),
    .Y(_01731_),
    .B1(_03029_));
 sg13g2_nor2_1 _18281_ (.A(net4196),
    .B(net6266),
    .Y(_03030_));
 sg13g2_a21oi_1 _18282_ (.A1(net7582),
    .A2(net6266),
    .Y(_01732_),
    .B1(_03030_));
 sg13g2_nor2_1 _18283_ (.A(net4353),
    .B(net6268),
    .Y(_03031_));
 sg13g2_a21oi_1 _18284_ (.A1(net6268),
    .A2(net7128),
    .Y(_01733_),
    .B1(_03031_));
 sg13g2_nor2_1 _18285_ (.A(net4789),
    .B(net6268),
    .Y(_03032_));
 sg13g2_a21oi_1 _18286_ (.A1(net6268),
    .A2(net7422),
    .Y(_01734_),
    .B1(_03032_));
 sg13g2_nor2_1 _18287_ (.A(net4463),
    .B(net6268),
    .Y(_03033_));
 sg13g2_a21oi_1 _18288_ (.A1(net6268),
    .A2(net7582),
    .Y(_01735_),
    .B1(_03033_));
 sg13g2_nor2_1 _18289_ (.A(net4435),
    .B(net6270),
    .Y(_03034_));
 sg13g2_a21oi_1 _18290_ (.A1(net6270),
    .A2(net7128),
    .Y(_01736_),
    .B1(_03034_));
 sg13g2_nor2_1 _18291_ (.A(net4581),
    .B(net6271),
    .Y(_03035_));
 sg13g2_a21oi_1 _18292_ (.A1(net6270),
    .A2(net7422),
    .Y(_01737_),
    .B1(_03035_));
 sg13g2_nor2_1 _18293_ (.A(net4135),
    .B(net6270),
    .Y(_03036_));
 sg13g2_a21oi_1 _18294_ (.A1(net6270),
    .A2(net7582),
    .Y(_01738_),
    .B1(_03036_));
 sg13g2_nor2_1 _18295_ (.A(net3714),
    .B(net6763),
    .Y(_03037_));
 sg13g2_a21oi_1 _18296_ (.A1(net6763),
    .A2(net7127),
    .Y(_01739_),
    .B1(_03037_));
 sg13g2_nor2_1 _18297_ (.A(net4197),
    .B(net6763),
    .Y(_03038_));
 sg13g2_a21oi_1 _18298_ (.A1(net6763),
    .A2(net7423),
    .Y(_01740_),
    .B1(_03038_));
 sg13g2_nor2_1 _18299_ (.A(net3470),
    .B(net6763),
    .Y(_03039_));
 sg13g2_a21oi_1 _18300_ (.A1(net6763),
    .A2(net7582),
    .Y(_01741_),
    .B1(_03039_));
 sg13g2_nor2_1 _18301_ (.A(net4567),
    .B(net6765),
    .Y(_03040_));
 sg13g2_a21oi_1 _18302_ (.A1(net6765),
    .A2(net7127),
    .Y(_01742_),
    .B1(_03040_));
 sg13g2_nor2_1 _18303_ (.A(net4166),
    .B(net6765),
    .Y(_03041_));
 sg13g2_a21oi_1 _18304_ (.A1(net6765),
    .A2(net7423),
    .Y(_01743_),
    .B1(_03041_));
 sg13g2_nor2_1 _18305_ (.A(net4004),
    .B(net6765),
    .Y(_03042_));
 sg13g2_a21oi_1 _18306_ (.A1(net6765),
    .A2(net7582),
    .Y(_01744_),
    .B1(_03042_));
 sg13g2_nor2_1 _18307_ (.A(net3920),
    .B(net6769),
    .Y(_03043_));
 sg13g2_a21oi_1 _18308_ (.A1(net6769),
    .A2(net7127),
    .Y(_01745_),
    .B1(_03043_));
 sg13g2_nor2_1 _18309_ (.A(net4478),
    .B(net6769),
    .Y(_03044_));
 sg13g2_a21oi_1 _18310_ (.A1(net6769),
    .A2(net7423),
    .Y(_01746_),
    .B1(_03044_));
 sg13g2_nor2_1 _18311_ (.A(net4411),
    .B(net6769),
    .Y(_03045_));
 sg13g2_a21oi_1 _18312_ (.A1(net6769),
    .A2(net7582),
    .Y(_01747_),
    .B1(_03045_));
 sg13g2_nand2_1 _18313_ (.Y(_03046_),
    .A(net2817),
    .B(net6773));
 sg13g2_o21ai_1 _18314_ (.B1(_03046_),
    .Y(_01748_),
    .A1(net6773),
    .A2(net7140));
 sg13g2_nand2_1 _18315_ (.Y(_03047_),
    .A(net4232),
    .B(net6773));
 sg13g2_o21ai_1 _18316_ (.B1(_03047_),
    .Y(_01749_),
    .A1(net6773),
    .A2(net7434));
 sg13g2_nand2_1 _18317_ (.Y(_03048_),
    .A(net3633),
    .B(net6774));
 sg13g2_o21ai_1 _18318_ (.B1(_03048_),
    .Y(_01750_),
    .A1(net6774),
    .A2(net7596));
 sg13g2_nor2_1 _18319_ (.A(net3327),
    .B(net6776),
    .Y(_03049_));
 sg13g2_a21oi_1 _18320_ (.A1(net6776),
    .A2(net7127),
    .Y(_01751_),
    .B1(_03049_));
 sg13g2_nor2_1 _18321_ (.A(net4397),
    .B(net6775),
    .Y(_03050_));
 sg13g2_a21oi_1 _18322_ (.A1(net6775),
    .A2(net7422),
    .Y(_01752_),
    .B1(_03050_));
 sg13g2_nor2_1 _18323_ (.A(net4145),
    .B(net6775),
    .Y(_03051_));
 sg13g2_a21oi_1 _18324_ (.A1(net6775),
    .A2(net7581),
    .Y(_01753_),
    .B1(_03051_));
 sg13g2_nor2_1 _18325_ (.A(net4112),
    .B(net6778),
    .Y(_03052_));
 sg13g2_a21oi_1 _18326_ (.A1(net6778),
    .A2(net7127),
    .Y(_01754_),
    .B1(_03052_));
 sg13g2_nor2_1 _18327_ (.A(net3755),
    .B(net6777),
    .Y(_03053_));
 sg13g2_a21oi_1 _18328_ (.A1(net6777),
    .A2(net7422),
    .Y(_01755_),
    .B1(_03053_));
 sg13g2_nor2_1 _18329_ (.A(net4131),
    .B(net6777),
    .Y(_03054_));
 sg13g2_a21oi_1 _18330_ (.A1(net6777),
    .A2(net7581),
    .Y(_01756_),
    .B1(_03054_));
 sg13g2_nor2_1 _18331_ (.A(net4564),
    .B(net6780),
    .Y(_03055_));
 sg13g2_a21oi_1 _18332_ (.A1(net6780),
    .A2(net7127),
    .Y(_01757_),
    .B1(_03055_));
 sg13g2_nor2_1 _18333_ (.A(net4181),
    .B(net6779),
    .Y(_03056_));
 sg13g2_a21oi_1 _18334_ (.A1(net6779),
    .A2(net7422),
    .Y(_01758_),
    .B1(_03056_));
 sg13g2_nor2_1 _18335_ (.A(net4620),
    .B(net6779),
    .Y(_03057_));
 sg13g2_a21oi_1 _18336_ (.A1(net6779),
    .A2(net7581),
    .Y(_01759_),
    .B1(_03057_));
 sg13g2_nor2_1 _18337_ (.A(net4472),
    .B(net6782),
    .Y(_03058_));
 sg13g2_a21oi_1 _18338_ (.A1(net6782),
    .A2(net7127),
    .Y(_01760_),
    .B1(_03058_));
 sg13g2_nor2_1 _18339_ (.A(net4505),
    .B(net6781),
    .Y(_03059_));
 sg13g2_a21oi_1 _18340_ (.A1(net6781),
    .A2(net7422),
    .Y(_01761_),
    .B1(_03059_));
 sg13g2_nor2_1 _18341_ (.A(net3570),
    .B(net6781),
    .Y(_03060_));
 sg13g2_a21oi_1 _18342_ (.A1(net6781),
    .A2(net7581),
    .Y(_01762_),
    .B1(_03060_));
 sg13g2_nor2_1 _18343_ (.A(net4781),
    .B(net6784),
    .Y(_03061_));
 sg13g2_a21oi_1 _18344_ (.A1(net6784),
    .A2(net7134),
    .Y(_01763_),
    .B1(_03061_));
 sg13g2_nor2_1 _18345_ (.A(net4827),
    .B(net6783),
    .Y(_03062_));
 sg13g2_a21oi_1 _18346_ (.A1(net6783),
    .A2(net7427),
    .Y(_01764_),
    .B1(_03062_));
 sg13g2_nor2_1 _18347_ (.A(net4098),
    .B(net6783),
    .Y(_03063_));
 sg13g2_a21oi_1 _18348_ (.A1(net6783),
    .A2(net7586),
    .Y(_01765_),
    .B1(_03063_));
 sg13g2_nor2_1 _18349_ (.A(net4474),
    .B(net6786),
    .Y(_03064_));
 sg13g2_a21oi_1 _18350_ (.A1(net6786),
    .A2(net7134),
    .Y(_01766_),
    .B1(_03064_));
 sg13g2_nor2_1 _18351_ (.A(net4841),
    .B(net6785),
    .Y(_03065_));
 sg13g2_a21oi_1 _18352_ (.A1(net6785),
    .A2(net7427),
    .Y(_01767_),
    .B1(_03065_));
 sg13g2_nor2_1 _18353_ (.A(net4491),
    .B(net6785),
    .Y(_03066_));
 sg13g2_a21oi_1 _18354_ (.A1(net6785),
    .A2(net7586),
    .Y(_01768_),
    .B1(_03066_));
 sg13g2_nor2_1 _18355_ (.A(net4575),
    .B(net6788),
    .Y(_03067_));
 sg13g2_a21oi_1 _18356_ (.A1(net6788),
    .A2(net7134),
    .Y(_01769_),
    .B1(_03067_));
 sg13g2_nor2_1 _18357_ (.A(net4647),
    .B(net6787),
    .Y(_03068_));
 sg13g2_a21oi_1 _18358_ (.A1(net6787),
    .A2(net7427),
    .Y(_01770_),
    .B1(_03068_));
 sg13g2_nor2_1 _18359_ (.A(net4597),
    .B(net6787),
    .Y(_03069_));
 sg13g2_a21oi_1 _18360_ (.A1(net6787),
    .A2(net7586),
    .Y(_01771_),
    .B1(_03069_));
 sg13g2_nand2_1 _18361_ (.Y(_03070_),
    .A(net2864),
    .B(net6790));
 sg13g2_o21ai_1 _18362_ (.B1(_03070_),
    .Y(_01772_),
    .A1(net6790),
    .A2(net7134));
 sg13g2_nand2_1 _18363_ (.Y(_03071_),
    .A(net2819),
    .B(net6789));
 sg13g2_o21ai_1 _18364_ (.B1(_03071_),
    .Y(_01773_),
    .A1(net6789),
    .A2(net7428));
 sg13g2_nand2_1 _18365_ (.Y(_03072_),
    .A(net2446),
    .B(net6789));
 sg13g2_o21ai_1 _18366_ (.B1(_03072_),
    .Y(_01774_),
    .A1(net6789),
    .A2(net7586));
 sg13g2_nand2_1 _18367_ (.Y(_03073_),
    .A(net2558),
    .B(net6792));
 sg13g2_o21ai_1 _18368_ (.B1(_03073_),
    .Y(_01775_),
    .A1(net6792),
    .A2(net7125));
 sg13g2_nand2_1 _18369_ (.Y(_03074_),
    .A(net3160),
    .B(net6791));
 sg13g2_o21ai_1 _18370_ (.B1(_03074_),
    .Y(_01776_),
    .A1(net6791),
    .A2(net7419));
 sg13g2_nand2_1 _18371_ (.Y(_03075_),
    .A(net3591),
    .B(net6791));
 sg13g2_o21ai_1 _18372_ (.B1(_03075_),
    .Y(_01777_),
    .A1(net6791),
    .A2(net7578));
 sg13g2_nand2_1 _18373_ (.Y(_03076_),
    .A(net2809),
    .B(net6793));
 sg13g2_o21ai_1 _18374_ (.B1(_03076_),
    .Y(_01778_),
    .A1(net6793),
    .A2(net7140));
 sg13g2_nand2_1 _18375_ (.Y(_03077_),
    .A(net3861),
    .B(net6793));
 sg13g2_o21ai_1 _18376_ (.B1(_03077_),
    .Y(_01779_),
    .A1(net6793),
    .A2(net7434));
 sg13g2_nand2_1 _18377_ (.Y(_03078_),
    .A(net2704),
    .B(net6794));
 sg13g2_o21ai_1 _18378_ (.B1(_03078_),
    .Y(_01780_),
    .A1(net6794),
    .A2(net7596));
 sg13g2_nand2_1 _18379_ (.Y(_03079_),
    .A(net2521),
    .B(net6797));
 sg13g2_o21ai_1 _18380_ (.B1(_03079_),
    .Y(_01781_),
    .A1(net6798),
    .A2(net7125));
 sg13g2_nand2_1 _18381_ (.Y(_03080_),
    .A(net3346),
    .B(net6798));
 sg13g2_o21ai_1 _18382_ (.B1(_03080_),
    .Y(_01782_),
    .A1(net6798),
    .A2(net7420));
 sg13g2_nand2_1 _18383_ (.Y(_03081_),
    .A(net3100),
    .B(net6797));
 sg13g2_o21ai_1 _18384_ (.B1(_03081_),
    .Y(_01783_),
    .A1(net6797),
    .A2(net7578));
 sg13g2_nand2_1 _18385_ (.Y(_03082_),
    .A(net3733),
    .B(net6800));
 sg13g2_o21ai_1 _18386_ (.B1(_03082_),
    .Y(_01784_),
    .A1(net6800),
    .A2(net7125));
 sg13g2_nand2_1 _18387_ (.Y(_03083_),
    .A(net3050),
    .B(net6799));
 sg13g2_o21ai_1 _18388_ (.B1(_03083_),
    .Y(_01785_),
    .A1(net6799),
    .A2(net7420));
 sg13g2_nand2_1 _18389_ (.Y(_03084_),
    .A(net3458),
    .B(net6799));
 sg13g2_o21ai_1 _18390_ (.B1(_03084_),
    .Y(_01786_),
    .A1(net6799),
    .A2(net7578));
 sg13g2_nand2_1 _18391_ (.Y(_03085_),
    .A(net3113),
    .B(net6277));
 sg13g2_o21ai_1 _18392_ (.B1(_03085_),
    .Y(_01787_),
    .A1(net6277),
    .A2(net7134));
 sg13g2_nand2_1 _18393_ (.Y(_03086_),
    .A(net3831),
    .B(net6276));
 sg13g2_o21ai_1 _18394_ (.B1(_03086_),
    .Y(_01788_),
    .A1(net6276),
    .A2(net7427));
 sg13g2_nand2_1 _18395_ (.Y(_03087_),
    .A(net3015),
    .B(net6276));
 sg13g2_o21ai_1 _18396_ (.B1(_03087_),
    .Y(_01789_),
    .A1(net6276),
    .A2(net7586));
 sg13g2_nand2_1 _18397_ (.Y(_03088_),
    .A(net3683),
    .B(net6279));
 sg13g2_o21ai_1 _18398_ (.B1(_03088_),
    .Y(_01790_),
    .A1(net6279),
    .A2(net7134));
 sg13g2_nand2_1 _18399_ (.Y(_03089_),
    .A(net3754),
    .B(net6278));
 sg13g2_o21ai_1 _18400_ (.B1(_03089_),
    .Y(_01791_),
    .A1(net6278),
    .A2(net7427));
 sg13g2_nand2_1 _18401_ (.Y(_03090_),
    .A(net3158),
    .B(net6278));
 sg13g2_o21ai_1 _18402_ (.B1(_03090_),
    .Y(_01792_),
    .A1(net6278),
    .A2(net7586));
 sg13g2_nand2_1 _18403_ (.Y(_03091_),
    .A(net3003),
    .B(net6281));
 sg13g2_o21ai_1 _18404_ (.B1(_03091_),
    .Y(_01793_),
    .A1(net6281),
    .A2(net7134));
 sg13g2_nand2_1 _18405_ (.Y(_03092_),
    .A(net3601),
    .B(net6280));
 sg13g2_o21ai_1 _18406_ (.B1(_03092_),
    .Y(_01794_),
    .A1(net6280),
    .A2(net7427));
 sg13g2_nand2_1 _18407_ (.Y(_03093_),
    .A(net4150),
    .B(net6280));
 sg13g2_o21ai_1 _18408_ (.B1(_03093_),
    .Y(_01795_),
    .A1(net6280),
    .A2(net7586));
 sg13g2_nand2_1 _18409_ (.Y(_03094_),
    .A(net2671),
    .B(net6283));
 sg13g2_o21ai_1 _18410_ (.B1(_03094_),
    .Y(_01796_),
    .A1(net6283),
    .A2(net7134));
 sg13g2_nand2_1 _18411_ (.Y(_03095_),
    .A(net3315),
    .B(net6282));
 sg13g2_o21ai_1 _18412_ (.B1(_03095_),
    .Y(_01797_),
    .A1(net6282),
    .A2(net7427));
 sg13g2_nand2_1 _18413_ (.Y(_03096_),
    .A(net2680),
    .B(net6282));
 sg13g2_o21ai_1 _18414_ (.B1(_03096_),
    .Y(_01798_),
    .A1(net6282),
    .A2(net7586));
 sg13g2_nand2_1 _18415_ (.Y(_03097_),
    .A(net2440),
    .B(net6802));
 sg13g2_o21ai_1 _18416_ (.B1(_03097_),
    .Y(_01799_),
    .A1(net6802),
    .A2(net7133));
 sg13g2_nand2_1 _18417_ (.Y(_03098_),
    .A(net4140),
    .B(net6801));
 sg13g2_o21ai_1 _18418_ (.B1(_03098_),
    .Y(_01800_),
    .A1(net6801),
    .A2(net7427));
 sg13g2_nand2_1 _18419_ (.Y(_03099_),
    .A(net3613),
    .B(net6801));
 sg13g2_o21ai_1 _18420_ (.B1(_03099_),
    .Y(_01801_),
    .A1(net6801),
    .A2(net7588));
 sg13g2_nand2_1 _18421_ (.Y(_03100_),
    .A(net3806),
    .B(net6804));
 sg13g2_o21ai_1 _18422_ (.B1(_03100_),
    .Y(_01802_),
    .A1(net6804),
    .A2(net7133));
 sg13g2_nand2_1 _18423_ (.Y(_03101_),
    .A(net4008),
    .B(net6803));
 sg13g2_o21ai_1 _18424_ (.B1(_03101_),
    .Y(_01803_),
    .A1(net6803),
    .A2(net7428));
 sg13g2_nand2_1 _18425_ (.Y(_03102_),
    .A(net3398),
    .B(net6803));
 sg13g2_o21ai_1 _18426_ (.B1(_03102_),
    .Y(_01804_),
    .A1(net6803),
    .A2(net7588));
 sg13g2_nand2_1 _18427_ (.Y(_03103_),
    .A(net3692),
    .B(net6806));
 sg13g2_o21ai_1 _18428_ (.B1(_03103_),
    .Y(_01805_),
    .A1(net6806),
    .A2(net7133));
 sg13g2_nand2_1 _18429_ (.Y(_03104_),
    .A(net3501),
    .B(net6805));
 sg13g2_o21ai_1 _18430_ (.B1(_03104_),
    .Y(_01806_),
    .A1(net6805),
    .A2(net7428));
 sg13g2_nand2_1 _18431_ (.Y(_03105_),
    .A(net3284),
    .B(net6805));
 sg13g2_o21ai_1 _18432_ (.B1(_03105_),
    .Y(_01807_),
    .A1(net6805),
    .A2(net7588));
 sg13g2_nor2_1 _18433_ (.A(net3785),
    .B(net6807),
    .Y(_03106_));
 sg13g2_a21oi_1 _18434_ (.A1(net6807),
    .A2(net7140),
    .Y(_01808_),
    .B1(_03106_));
 sg13g2_nor2_1 _18435_ (.A(net4824),
    .B(net6807),
    .Y(_03107_));
 sg13g2_a21oi_1 _18436_ (.A1(net6807),
    .A2(net7434),
    .Y(_01809_),
    .B1(_03107_));
 sg13g2_nor2_1 _18437_ (.A(net4212),
    .B(net6808),
    .Y(_03108_));
 sg13g2_a21oi_1 _18438_ (.A1(net6808),
    .A2(net7597),
    .Y(_01810_),
    .B1(_03108_));
 sg13g2_nor2_1 _18439_ (.A(net4783),
    .B(net6809),
    .Y(_03109_));
 sg13g2_a21oi_1 _18440_ (.A1(net6809),
    .A2(net7141),
    .Y(_01811_),
    .B1(_03109_));
 sg13g2_nor2_1 _18441_ (.A(net4039),
    .B(net6810),
    .Y(_03110_));
 sg13g2_a21oi_1 _18442_ (.A1(net6810),
    .A2(net7435),
    .Y(_01812_),
    .B1(_03110_));
 sg13g2_nor2_1 _18443_ (.A(net4191),
    .B(net6810),
    .Y(_03111_));
 sg13g2_a21oi_1 _18444_ (.A1(net6809),
    .A2(net7595),
    .Y(_01813_),
    .B1(_03111_));
 sg13g2_nor2_1 _18445_ (.A(net3673),
    .B(net6811),
    .Y(_03112_));
 sg13g2_a21oi_1 _18446_ (.A1(net6811),
    .A2(net7141),
    .Y(_01814_),
    .B1(_03112_));
 sg13g2_nor2_1 _18447_ (.A(net4502),
    .B(net6811),
    .Y(_03113_));
 sg13g2_a21oi_1 _18448_ (.A1(net6811),
    .A2(net7435),
    .Y(_01815_),
    .B1(_03113_));
 sg13g2_nor2_1 _18449_ (.A(net4498),
    .B(net6811),
    .Y(_03114_));
 sg13g2_a21oi_1 _18450_ (.A1(net6811),
    .A2(net7595),
    .Y(_01816_),
    .B1(_03114_));
 sg13g2_nor2_1 _18451_ (.A(net4452),
    .B(net6813),
    .Y(_03115_));
 sg13g2_a21oi_1 _18452_ (.A1(net6813),
    .A2(net7141),
    .Y(_01817_),
    .B1(_03115_));
 sg13g2_nor2_1 _18453_ (.A(net4448),
    .B(net6813),
    .Y(_03116_));
 sg13g2_a21oi_1 _18454_ (.A1(net6813),
    .A2(net7435),
    .Y(_01818_),
    .B1(_03116_));
 sg13g2_nor2_1 _18455_ (.A(net4767),
    .B(net6813),
    .Y(_03117_));
 sg13g2_a21oi_1 _18456_ (.A1(net6813),
    .A2(net7595),
    .Y(_01819_),
    .B1(_03117_));
 sg13g2_nand2_1 _18457_ (.Y(_03118_),
    .A(net2634),
    .B(net6298));
 sg13g2_o21ai_1 _18458_ (.B1(_03118_),
    .Y(_01820_),
    .A1(net6298),
    .A2(net7141));
 sg13g2_nand2_1 _18459_ (.Y(_03119_),
    .A(net2758),
    .B(net6298));
 sg13g2_o21ai_1 _18460_ (.B1(_03119_),
    .Y(_01821_),
    .A1(net6298),
    .A2(net7435));
 sg13g2_nand2_1 _18461_ (.Y(_03120_),
    .A(net3763),
    .B(net6298));
 sg13g2_o21ai_1 _18462_ (.B1(_03120_),
    .Y(_01822_),
    .A1(net6298),
    .A2(net7595));
 sg13g2_nand2_1 _18463_ (.Y(_03121_),
    .A(net3052),
    .B(net6303));
 sg13g2_o21ai_1 _18464_ (.B1(_03121_),
    .Y(_01823_),
    .A1(net6303),
    .A2(net7154));
 sg13g2_nand2_1 _18465_ (.Y(_03122_),
    .A(net4281),
    .B(net6303));
 sg13g2_o21ai_1 _18466_ (.B1(_03122_),
    .Y(_01824_),
    .A1(net6303),
    .A2(net7450));
 sg13g2_nand2_1 _18467_ (.Y(_03123_),
    .A(net3312),
    .B(net6302));
 sg13g2_o21ai_1 _18468_ (.B1(_03123_),
    .Y(_01825_),
    .A1(net6302),
    .A2(net7609));
 sg13g2_nand2_1 _18469_ (.Y(_03124_),
    .A(net2885),
    .B(net6307));
 sg13g2_o21ai_1 _18470_ (.B1(_03124_),
    .Y(_01826_),
    .A1(net6307),
    .A2(net7154));
 sg13g2_nand2_1 _18471_ (.Y(_03125_),
    .A(net3485),
    .B(net6307));
 sg13g2_o21ai_1 _18472_ (.B1(_03125_),
    .Y(_01827_),
    .A1(net6307),
    .A2(net7450));
 sg13g2_nand2_1 _18473_ (.Y(_03126_),
    .A(net3166),
    .B(net6306));
 sg13g2_o21ai_1 _18474_ (.B1(_03126_),
    .Y(_01828_),
    .A1(net6306),
    .A2(net7609));
 sg13g2_nand2_1 _18475_ (.Y(_03127_),
    .A(net4055),
    .B(net6369));
 sg13g2_o21ai_1 _18476_ (.B1(_03127_),
    .Y(_01829_),
    .A1(net6369),
    .A2(net7154));
 sg13g2_nand2_1 _18477_ (.Y(_03128_),
    .A(net3942),
    .B(net6369));
 sg13g2_o21ai_1 _18478_ (.B1(_03128_),
    .Y(_01830_),
    .A1(net6369),
    .A2(net7450));
 sg13g2_nand2_1 _18479_ (.Y(_03129_),
    .A(net4347),
    .B(net6368));
 sg13g2_o21ai_1 _18480_ (.B1(_03129_),
    .Y(_01831_),
    .A1(net6368),
    .A2(net7609));
 sg13g2_nand2_1 _18481_ (.Y(_03130_),
    .A(net4123),
    .B(net6371));
 sg13g2_o21ai_1 _18482_ (.B1(_03130_),
    .Y(_01832_),
    .A1(net6371),
    .A2(net7154));
 sg13g2_nand2_1 _18483_ (.Y(_03131_),
    .A(net4057),
    .B(net6370));
 sg13g2_o21ai_1 _18484_ (.B1(_03131_),
    .Y(_01833_),
    .A1(net6370),
    .A2(net7450));
 sg13g2_nand2_1 _18485_ (.Y(_03132_),
    .A(net2934),
    .B(net6370));
 sg13g2_o21ai_1 _18486_ (.B1(_03132_),
    .Y(_01834_),
    .A1(net6371),
    .A2(net7609));
 sg13g2_nand2_1 _18487_ (.Y(_03133_),
    .A(net3491),
    .B(net6372));
 sg13g2_o21ai_1 _18488_ (.B1(_03133_),
    .Y(_01835_),
    .A1(net6372),
    .A2(net7153));
 sg13g2_nand2_1 _18489_ (.Y(_03134_),
    .A(net3379),
    .B(net6373));
 sg13g2_o21ai_1 _18490_ (.B1(_03134_),
    .Y(_01836_),
    .A1(net6373),
    .A2(net7449));
 sg13g2_nand2_1 _18491_ (.Y(_03135_),
    .A(net3351),
    .B(net6373));
 sg13g2_o21ai_1 _18492_ (.B1(_03135_),
    .Y(_01837_),
    .A1(net6373),
    .A2(net7608));
 sg13g2_nand2_1 _18493_ (.Y(_03136_),
    .A(net3780),
    .B(net6831));
 sg13g2_o21ai_1 _18494_ (.B1(_03136_),
    .Y(_01838_),
    .A1(net6831),
    .A2(net7165));
 sg13g2_nand2_1 _18495_ (.Y(_03137_),
    .A(net2487),
    .B(net6832));
 sg13g2_o21ai_1 _18496_ (.B1(_03137_),
    .Y(_01839_),
    .A1(net6831),
    .A2(net7461));
 sg13g2_nand2_1 _18497_ (.Y(_03138_),
    .A(net3478),
    .B(net6831));
 sg13g2_o21ai_1 _18498_ (.B1(_03138_),
    .Y(_01840_),
    .A1(net6831),
    .A2(net7616));
 sg13g2_nand2_1 _18499_ (.Y(_03139_),
    .A(net3439),
    .B(net6375));
 sg13g2_o21ai_1 _18500_ (.B1(_03139_),
    .Y(_01841_),
    .A1(net6374),
    .A2(net7153));
 sg13g2_nand2_1 _18501_ (.Y(_03140_),
    .A(net2551),
    .B(net6374));
 sg13g2_o21ai_1 _18502_ (.B1(_03140_),
    .Y(_01842_),
    .A1(net6375),
    .A2(net7449));
 sg13g2_nand2_1 _18503_ (.Y(_03141_),
    .A(net2768),
    .B(net6375));
 sg13g2_o21ai_1 _18504_ (.B1(_03141_),
    .Y(_01843_),
    .A1(net6375),
    .A2(net7608));
 sg13g2_nand2_1 _18505_ (.Y(_03142_),
    .A(net2476),
    .B(net6376));
 sg13g2_o21ai_1 _18506_ (.B1(_03142_),
    .Y(_01844_),
    .A1(net6377),
    .A2(net7153));
 sg13g2_nand2_1 _18507_ (.Y(_03143_),
    .A(net3211),
    .B(net6377));
 sg13g2_o21ai_1 _18508_ (.B1(_03143_),
    .Y(_01845_),
    .A1(net6376),
    .A2(net7449));
 sg13g2_nand2_1 _18509_ (.Y(_03144_),
    .A(net2886),
    .B(net6377));
 sg13g2_o21ai_1 _18510_ (.B1(_03144_),
    .Y(_01846_),
    .A1(net6377),
    .A2(net7608));
 sg13g2_nand2_1 _18511_ (.Y(_03145_),
    .A(net3651),
    .B(net6378));
 sg13g2_o21ai_1 _18512_ (.B1(_03145_),
    .Y(_01847_),
    .A1(net6378),
    .A2(net7153));
 sg13g2_nand2_1 _18513_ (.Y(_03146_),
    .A(net3726),
    .B(net6379));
 sg13g2_o21ai_1 _18514_ (.B1(_03146_),
    .Y(_01848_),
    .A1(net6379),
    .A2(net7449));
 sg13g2_nand2_1 _18515_ (.Y(_03147_),
    .A(net3138),
    .B(net6378));
 sg13g2_o21ai_1 _18516_ (.B1(_03147_),
    .Y(_01849_),
    .A1(net6378),
    .A2(net7608));
 sg13g2_nand2_1 _18517_ (.Y(_03148_),
    .A(net4022),
    .B(net6380));
 sg13g2_o21ai_1 _18518_ (.B1(_03148_),
    .Y(_01850_),
    .A1(net6380),
    .A2(net7153));
 sg13g2_nand2_1 _18519_ (.Y(_03149_),
    .A(net3155),
    .B(net6381));
 sg13g2_o21ai_1 _18520_ (.B1(_03149_),
    .Y(_01851_),
    .A1(net6381),
    .A2(net7449));
 sg13g2_nand2_1 _18521_ (.Y(_03150_),
    .A(net3987),
    .B(net6380));
 sg13g2_o21ai_1 _18522_ (.B1(_03150_),
    .Y(_01852_),
    .A1(net6380),
    .A2(net7608));
 sg13g2_nand2_1 _18523_ (.Y(_03151_),
    .A(net3641),
    .B(net6382));
 sg13g2_o21ai_1 _18524_ (.B1(_03151_),
    .Y(_01853_),
    .A1(net6382),
    .A2(net7153));
 sg13g2_nand2_1 _18525_ (.Y(_03152_),
    .A(net4151),
    .B(net6383));
 sg13g2_o21ai_1 _18526_ (.B1(_03152_),
    .Y(_01854_),
    .A1(net6383),
    .A2(net7449));
 sg13g2_nand2_1 _18527_ (.Y(_03153_),
    .A(net3958),
    .B(net6382));
 sg13g2_o21ai_1 _18528_ (.B1(_03153_),
    .Y(_01855_),
    .A1(net6382),
    .A2(net7608));
 sg13g2_nand2_1 _18529_ (.Y(_03154_),
    .A(net3317),
    .B(net6384));
 sg13g2_o21ai_1 _18530_ (.B1(_03154_),
    .Y(_01856_),
    .A1(net6384),
    .A2(net7153));
 sg13g2_nand2_1 _18531_ (.Y(_03155_),
    .A(net2795),
    .B(net6385));
 sg13g2_o21ai_1 _18532_ (.B1(_03155_),
    .Y(_01857_),
    .A1(net6385),
    .A2(net7449));
 sg13g2_nand2_1 _18533_ (.Y(_03156_),
    .A(net2595),
    .B(net6384));
 sg13g2_o21ai_1 _18534_ (.B1(_03156_),
    .Y(_01858_),
    .A1(net6384),
    .A2(net7608));
 sg13g2_nand2_1 _18535_ (.Y(_03157_),
    .A(net2896),
    .B(net6834));
 sg13g2_o21ai_1 _18536_ (.B1(_03157_),
    .Y(_01859_),
    .A1(net6834),
    .A2(net7159));
 sg13g2_nand2_1 _18537_ (.Y(_03158_),
    .A(net3462),
    .B(net6833));
 sg13g2_o21ai_1 _18538_ (.B1(_03158_),
    .Y(_01860_),
    .A1(net6833),
    .A2(net7453));
 sg13g2_nand2_1 _18539_ (.Y(_03159_),
    .A(net2790),
    .B(net6833));
 sg13g2_o21ai_1 _18540_ (.B1(_03159_),
    .Y(_01861_),
    .A1(net6833),
    .A2(net7614));
 sg13g2_nand2_1 _18541_ (.Y(_03160_),
    .A(net3280),
    .B(net6836));
 sg13g2_o21ai_1 _18542_ (.B1(_03160_),
    .Y(_01862_),
    .A1(net6836),
    .A2(net7159));
 sg13g2_nand2_1 _18543_ (.Y(_03161_),
    .A(net3637),
    .B(net6835));
 sg13g2_o21ai_1 _18544_ (.B1(_03161_),
    .Y(_01863_),
    .A1(net6835),
    .A2(net7456));
 sg13g2_nand2_1 _18545_ (.Y(_03162_),
    .A(net2610),
    .B(net6835));
 sg13g2_o21ai_1 _18546_ (.B1(_03162_),
    .Y(_01864_),
    .A1(net6835),
    .A2(net7614));
 sg13g2_nand2_1 _18547_ (.Y(_03163_),
    .A(net3059),
    .B(net6838));
 sg13g2_o21ai_1 _18548_ (.B1(_03163_),
    .Y(_01865_),
    .A1(net6838),
    .A2(net7159));
 sg13g2_nand2_1 _18549_ (.Y(_03164_),
    .A(net4068),
    .B(net6837));
 sg13g2_o21ai_1 _18550_ (.B1(_03164_),
    .Y(_01866_),
    .A1(net6837),
    .A2(net7453));
 sg13g2_nand2_1 _18551_ (.Y(_03165_),
    .A(net3669),
    .B(net6837));
 sg13g2_o21ai_1 _18552_ (.B1(_03165_),
    .Y(_01867_),
    .A1(net6837),
    .A2(net7614));
 sg13g2_nand2_1 _18553_ (.Y(_03166_),
    .A(net2822),
    .B(net6839));
 sg13g2_o21ai_1 _18554_ (.B1(_03166_),
    .Y(_01868_),
    .A1(net6839),
    .A2(net7165));
 sg13g2_nand2_1 _18555_ (.Y(_03167_),
    .A(net2962),
    .B(net6840));
 sg13g2_o21ai_1 _18556_ (.B1(_03167_),
    .Y(_01869_),
    .A1(net6839),
    .A2(net7461));
 sg13g2_nand2_1 _18557_ (.Y(_03168_),
    .A(net4300),
    .B(net6839));
 sg13g2_o21ai_1 _18558_ (.B1(_03168_),
    .Y(_01870_),
    .A1(net6839),
    .A2(net7616));
 sg13g2_nand2_1 _18559_ (.Y(_03169_),
    .A(net2889),
    .B(net6842));
 sg13g2_o21ai_1 _18560_ (.B1(_03169_),
    .Y(_01871_),
    .A1(net6842),
    .A2(net7157));
 sg13g2_nand2_1 _18561_ (.Y(_03170_),
    .A(net2715),
    .B(net6842));
 sg13g2_o21ai_1 _18562_ (.B1(_03170_),
    .Y(_01872_),
    .A1(net6841),
    .A2(net7453));
 sg13g2_nand2_1 _18563_ (.Y(_03171_),
    .A(net2449),
    .B(net6841));
 sg13g2_o21ai_1 _18564_ (.B1(_03171_),
    .Y(_01873_),
    .A1(net6842),
    .A2(net7613));
 sg13g2_nand2_1 _18565_ (.Y(_03172_),
    .A(net2749),
    .B(net6844));
 sg13g2_o21ai_1 _18566_ (.B1(_03172_),
    .Y(_01874_),
    .A1(net6844),
    .A2(net7157));
 sg13g2_nand2_1 _18567_ (.Y(_03173_),
    .A(net2796),
    .B(net6844));
 sg13g2_o21ai_1 _18568_ (.B1(_03173_),
    .Y(_01875_),
    .A1(net6843),
    .A2(net7453));
 sg13g2_nand2_1 _18569_ (.Y(_03174_),
    .A(net3274),
    .B(net6843));
 sg13g2_o21ai_1 _18570_ (.B1(_03174_),
    .Y(_01876_),
    .A1(net6844),
    .A2(net7613));
 sg13g2_nand2_1 _18571_ (.Y(_03175_),
    .A(net2670),
    .B(net6846));
 sg13g2_o21ai_1 _18572_ (.B1(_03175_),
    .Y(_01877_),
    .A1(net6846),
    .A2(net7157));
 sg13g2_nand2_1 _18573_ (.Y(_03176_),
    .A(net3658),
    .B(net6845));
 sg13g2_o21ai_1 _18574_ (.B1(_03176_),
    .Y(_01878_),
    .A1(net6845),
    .A2(net7453));
 sg13g2_nand2_1 _18575_ (.Y(_03177_),
    .A(net3278),
    .B(net6845));
 sg13g2_o21ai_1 _18576_ (.B1(_03177_),
    .Y(_01879_),
    .A1(net6845),
    .A2(net7613));
 sg13g2_nand2_1 _18577_ (.Y(_03178_),
    .A(net2814),
    .B(net6848));
 sg13g2_o21ai_1 _18578_ (.B1(_03178_),
    .Y(_01880_),
    .A1(net6848),
    .A2(net7157));
 sg13g2_nand2_1 _18579_ (.Y(_03179_),
    .A(net4056),
    .B(net6847));
 sg13g2_o21ai_1 _18580_ (.B1(_03179_),
    .Y(_01881_),
    .A1(net6847),
    .A2(net7453));
 sg13g2_nand2_1 _18581_ (.Y(_03180_),
    .A(net4291),
    .B(net6847));
 sg13g2_o21ai_1 _18582_ (.B1(_03180_),
    .Y(_01882_),
    .A1(net6847),
    .A2(net7613));
 sg13g2_nand2_1 _18583_ (.Y(_03181_),
    .A(net4067),
    .B(net6390));
 sg13g2_o21ai_1 _18584_ (.B1(_03181_),
    .Y(_01883_),
    .A1(net6390),
    .A2(net7154));
 sg13g2_nand2_1 _18585_ (.Y(_03182_),
    .A(net3966),
    .B(net6391));
 sg13g2_o21ai_1 _18586_ (.B1(_03182_),
    .Y(_01884_),
    .A1(net6391),
    .A2(net7454));
 sg13g2_nand2_1 _18587_ (.Y(_03183_),
    .A(net4345),
    .B(net6391));
 sg13g2_o21ai_1 _18588_ (.B1(_03183_),
    .Y(_01885_),
    .A1(net6390),
    .A2(net7613));
 sg13g2_nand2_1 _18589_ (.Y(_03184_),
    .A(net3752),
    .B(net6396));
 sg13g2_o21ai_1 _18590_ (.B1(_03184_),
    .Y(_01886_),
    .A1(net6396),
    .A2(net7154));
 sg13g2_nand2_1 _18591_ (.Y(_03185_),
    .A(net3009),
    .B(net6397));
 sg13g2_o21ai_1 _18592_ (.B1(_03185_),
    .Y(_01887_),
    .A1(net6397),
    .A2(net7454));
 sg13g2_nand2_1 _18593_ (.Y(_03186_),
    .A(net2976),
    .B(net6396));
 sg13g2_o21ai_1 _18594_ (.B1(_03186_),
    .Y(_01888_),
    .A1(net6396),
    .A2(net7613));
 sg13g2_nand2_1 _18595_ (.Y(_03187_),
    .A(net3216),
    .B(net6400));
 sg13g2_o21ai_1 _18596_ (.B1(_03187_),
    .Y(_01889_),
    .A1(net6400),
    .A2(net7154));
 sg13g2_nand2_1 _18597_ (.Y(_03188_),
    .A(net4045),
    .B(net6401));
 sg13g2_o21ai_1 _18598_ (.B1(_03188_),
    .Y(_01890_),
    .A1(net6401),
    .A2(net7454));
 sg13g2_nand2_1 _18599_ (.Y(_03189_),
    .A(net4031),
    .B(net6401));
 sg13g2_o21ai_1 _18600_ (.B1(_03189_),
    .Y(_01891_),
    .A1(net6400),
    .A2(net7613));
 sg13g2_nand2_1 _18601_ (.Y(_03190_),
    .A(net2504),
    .B(net6402));
 sg13g2_o21ai_1 _18602_ (.B1(_03190_),
    .Y(_01892_),
    .A1(net6402),
    .A2(net7154));
 sg13g2_nand2_1 _18603_ (.Y(_03191_),
    .A(net3359),
    .B(net6403));
 sg13g2_o21ai_1 _18604_ (.B1(_03191_),
    .Y(_01893_),
    .A1(net6403),
    .A2(net7453));
 sg13g2_nand2_1 _18605_ (.Y(_03192_),
    .A(net2663),
    .B(net6402));
 sg13g2_o21ai_1 _18606_ (.B1(_03192_),
    .Y(_01894_),
    .A1(net6402),
    .A2(net7613));
 sg13g2_nand2_1 _18607_ (.Y(_03193_),
    .A(net3440),
    .B(net6849));
 sg13g2_o21ai_1 _18608_ (.B1(_03193_),
    .Y(_01895_),
    .A1(net6849),
    .A2(net7155));
 sg13g2_nand2_1 _18609_ (.Y(_03194_),
    .A(net3355),
    .B(net6849));
 sg13g2_o21ai_1 _18610_ (.B1(_03194_),
    .Y(_01896_),
    .A1(net6849),
    .A2(net7451));
 sg13g2_nand2_1 _18611_ (.Y(_03195_),
    .A(net3768),
    .B(net6850));
 sg13g2_o21ai_1 _18612_ (.B1(_03195_),
    .Y(_01897_),
    .A1(net6850),
    .A2(net7614));
 sg13g2_nand2_1 _18613_ (.Y(_03196_),
    .A(net3433),
    .B(net6851));
 sg13g2_o21ai_1 _18614_ (.B1(_03196_),
    .Y(_01898_),
    .A1(net6851),
    .A2(net7165));
 sg13g2_nand2_1 _18615_ (.Y(_03197_),
    .A(net3328),
    .B(net6851));
 sg13g2_o21ai_1 _18616_ (.B1(_03197_),
    .Y(_01899_),
    .A1(net6851),
    .A2(net7461));
 sg13g2_nand2_1 _18617_ (.Y(_03198_),
    .A(net3321),
    .B(net6851));
 sg13g2_o21ai_1 _18618_ (.B1(_03198_),
    .Y(_01900_),
    .A1(net6851),
    .A2(net7616));
 sg13g2_nand2_1 _18619_ (.Y(_03199_),
    .A(net3775),
    .B(net6854));
 sg13g2_o21ai_1 _18620_ (.B1(_03199_),
    .Y(_01901_),
    .A1(net6854),
    .A2(net7159));
 sg13g2_nand2_1 _18621_ (.Y(_03200_),
    .A(net2659),
    .B(net6853));
 sg13g2_o21ai_1 _18622_ (.B1(_03200_),
    .Y(_01902_),
    .A1(net6853),
    .A2(net7456));
 sg13g2_nand2_1 _18623_ (.Y(_03201_),
    .A(net4078),
    .B(net6853));
 sg13g2_o21ai_1 _18624_ (.B1(_03201_),
    .Y(_01903_),
    .A1(net6853),
    .A2(net7614));
 sg13g2_nand2_1 _18625_ (.Y(_03202_),
    .A(net2525),
    .B(net6856));
 sg13g2_o21ai_1 _18626_ (.B1(_03202_),
    .Y(_01904_),
    .A1(net6856),
    .A2(net7159));
 sg13g2_nand2_1 _18627_ (.Y(_03203_),
    .A(net2495),
    .B(net6855));
 sg13g2_o21ai_1 _18628_ (.B1(_03203_),
    .Y(_01905_),
    .A1(net6855),
    .A2(net7456));
 sg13g2_nand2_1 _18629_ (.Y(_03204_),
    .A(net4334),
    .B(net6855));
 sg13g2_o21ai_1 _18630_ (.B1(_03204_),
    .Y(_01906_),
    .A1(net6855),
    .A2(net7614));
 sg13g2_nand2_1 _18631_ (.Y(_03205_),
    .A(net3866),
    .B(net6857));
 sg13g2_o21ai_1 _18632_ (.B1(_03205_),
    .Y(_01907_),
    .A1(net6857),
    .A2(net7139));
 sg13g2_nand2_1 _18633_ (.Y(_03206_),
    .A(net3005),
    .B(net6857));
 sg13g2_o21ai_1 _18634_ (.B1(_03206_),
    .Y(_01908_),
    .A1(net6857),
    .A2(net7433));
 sg13g2_nand2_1 _18635_ (.Y(_03207_),
    .A(net2756),
    .B(net6857));
 sg13g2_o21ai_1 _18636_ (.B1(_03207_),
    .Y(_01909_),
    .A1(net6857),
    .A2(net7593));
 sg13g2_nand2_1 _18637_ (.Y(_03208_),
    .A(net3594),
    .B(net6859));
 sg13g2_o21ai_1 _18638_ (.B1(_03208_),
    .Y(_01910_),
    .A1(net6859),
    .A2(net7139));
 sg13g2_nand2_1 _18639_ (.Y(_03209_),
    .A(net2500),
    .B(net6859));
 sg13g2_o21ai_1 _18640_ (.B1(_03209_),
    .Y(_01911_),
    .A1(net6859),
    .A2(net7432));
 sg13g2_nand2_1 _18641_ (.Y(_03210_),
    .A(net4132),
    .B(net6859));
 sg13g2_o21ai_1 _18642_ (.B1(_03210_),
    .Y(_01912_),
    .A1(net6859),
    .A2(net7593));
 sg13g2_nand2_1 _18643_ (.Y(_03211_),
    .A(net2713),
    .B(net6861));
 sg13g2_o21ai_1 _18644_ (.B1(_03211_),
    .Y(_01913_),
    .A1(net6861),
    .A2(net7138));
 sg13g2_nand2_1 _18645_ (.Y(_03212_),
    .A(net3963),
    .B(net6861));
 sg13g2_o21ai_1 _18646_ (.B1(_03212_),
    .Y(_01914_),
    .A1(net6861),
    .A2(net7433));
 sg13g2_nand2_1 _18647_ (.Y(_03213_),
    .A(net2736),
    .B(net6861));
 sg13g2_o21ai_1 _18648_ (.B1(_03213_),
    .Y(_01915_),
    .A1(net6861),
    .A2(net7593));
 sg13g2_nand2_1 _18649_ (.Y(_03214_),
    .A(net3144),
    .B(net6863));
 sg13g2_o21ai_1 _18650_ (.B1(_03214_),
    .Y(_01916_),
    .A1(net6863),
    .A2(net7139));
 sg13g2_nand2_1 _18651_ (.Y(_03215_),
    .A(net2978),
    .B(net6863));
 sg13g2_o21ai_1 _18652_ (.B1(_03215_),
    .Y(_01917_),
    .A1(net6864),
    .A2(net7432));
 sg13g2_nand2_1 _18653_ (.Y(_03216_),
    .A(net2711),
    .B(net6863));
 sg13g2_o21ai_1 _18654_ (.B1(_03216_),
    .Y(_01918_),
    .A1(net6863),
    .A2(net7593));
 sg13g2_nand2_1 _18655_ (.Y(_03217_),
    .A(net2709),
    .B(net6865));
 sg13g2_o21ai_1 _18656_ (.B1(_03217_),
    .Y(_01919_),
    .A1(net6865),
    .A2(net7138));
 sg13g2_nand2_1 _18657_ (.Y(_03218_),
    .A(net2541),
    .B(net6865));
 sg13g2_o21ai_1 _18658_ (.B1(_03218_),
    .Y(_01920_),
    .A1(net6865),
    .A2(net7432));
 sg13g2_nand2_1 _18659_ (.Y(_03219_),
    .A(net2741),
    .B(net6866));
 sg13g2_o21ai_1 _18660_ (.B1(_03219_),
    .Y(_01921_),
    .A1(net6866),
    .A2(net7592));
 sg13g2_nand2_1 _18661_ (.Y(_03220_),
    .A(net3377),
    .B(net6869));
 sg13g2_o21ai_1 _18662_ (.B1(_03220_),
    .Y(_01922_),
    .A1(net6869),
    .A2(net7138));
 sg13g2_nand2_1 _18663_ (.Y(_03221_),
    .A(net3624),
    .B(net6869));
 sg13g2_o21ai_1 _18664_ (.B1(_03221_),
    .Y(_01923_),
    .A1(net6869),
    .A2(net7432));
 sg13g2_nand2_1 _18665_ (.Y(_03222_),
    .A(net3642),
    .B(net6870));
 sg13g2_o21ai_1 _18666_ (.B1(_03222_),
    .Y(_01924_),
    .A1(net6870),
    .A2(net7592));
 sg13g2_nand2_1 _18667_ (.Y(_03223_),
    .A(net2591),
    .B(net6871));
 sg13g2_o21ai_1 _18668_ (.B1(_03223_),
    .Y(_01925_),
    .A1(net6871),
    .A2(net7138));
 sg13g2_nand2_1 _18669_ (.Y(_03224_),
    .A(net3273),
    .B(net6871));
 sg13g2_o21ai_1 _18670_ (.B1(_03224_),
    .Y(_01926_),
    .A1(net6871),
    .A2(net7433));
 sg13g2_nand2_1 _18671_ (.Y(_03225_),
    .A(net3292),
    .B(net6872));
 sg13g2_o21ai_1 _18672_ (.B1(_03225_),
    .Y(_01927_),
    .A1(net6872),
    .A2(net7592));
 sg13g2_nor2_1 _18673_ (.A(net4278),
    .B(net6922),
    .Y(_03226_));
 sg13g2_a21oi_1 _18674_ (.A1(net6922),
    .A2(net7140),
    .Y(_01928_),
    .B1(_03226_));
 sg13g2_nor2_1 _18675_ (.A(net3894),
    .B(net6922),
    .Y(_03227_));
 sg13g2_a21oi_1 _18676_ (.A1(net6922),
    .A2(net7434),
    .Y(_01929_),
    .B1(_03227_));
 sg13g2_nor2_1 _18677_ (.A(net4121),
    .B(net6923),
    .Y(_03228_));
 sg13g2_a21oi_1 _18678_ (.A1(net6923),
    .A2(net7595),
    .Y(_01930_),
    .B1(_03228_));
 sg13g2_nand2_1 _18679_ (.Y(_03229_),
    .A(net2695),
    .B(net6924));
 sg13g2_o21ai_1 _18680_ (.B1(_03229_),
    .Y(_01931_),
    .A1(net6924),
    .A2(net7164));
 sg13g2_nand2_1 _18681_ (.Y(_03230_),
    .A(net3062),
    .B(net6924));
 sg13g2_o21ai_1 _18682_ (.B1(_03230_),
    .Y(_01932_),
    .A1(net6924),
    .A2(net7458));
 sg13g2_nand2_1 _18683_ (.Y(_03231_),
    .A(net3257),
    .B(net6924));
 sg13g2_o21ai_1 _18684_ (.B1(_03231_),
    .Y(_01933_),
    .A1(net6924),
    .A2(net7619));
 sg13g2_nand2_1 _18685_ (.Y(_03232_),
    .A(net3540),
    .B(net6926));
 sg13g2_o21ai_1 _18686_ (.B1(_03232_),
    .Y(_01934_),
    .A1(net6927),
    .A2(net7151));
 sg13g2_nand2_1 _18687_ (.Y(_03233_),
    .A(net2994),
    .B(net6926));
 sg13g2_o21ai_1 _18688_ (.B1(_03233_),
    .Y(_01935_),
    .A1(net6926),
    .A2(net7444));
 sg13g2_nand2_1 _18689_ (.Y(_03234_),
    .A(net3493),
    .B(net6926));
 sg13g2_o21ai_1 _18690_ (.B1(_03234_),
    .Y(_01936_),
    .A1(net6927),
    .A2(net7604));
 sg13g2_nand2_1 _18691_ (.Y(_03235_),
    .A(net3946),
    .B(net6521));
 sg13g2_o21ai_1 _18692_ (.B1(_03235_),
    .Y(_01937_),
    .A1(net6521),
    .A2(net7167));
 sg13g2_nand2_1 _18693_ (.Y(_03236_),
    .A(net2914),
    .B(net6520));
 sg13g2_o21ai_1 _18694_ (.B1(_03236_),
    .Y(_01938_),
    .A1(net6520),
    .A2(net7465));
 sg13g2_nand2_1 _18695_ (.Y(_03237_),
    .A(net2520),
    .B(net6520));
 sg13g2_o21ai_1 _18696_ (.B1(_03237_),
    .Y(_01939_),
    .A1(net6520),
    .A2(net7624));
 sg13g2_nand2_1 _18697_ (.Y(_03238_),
    .A(net2565),
    .B(net6929));
 sg13g2_o21ai_1 _18698_ (.B1(_03238_),
    .Y(_01940_),
    .A1(net6929),
    .A2(net7184));
 sg13g2_nand2_1 _18699_ (.Y(_03239_),
    .A(net3803),
    .B(net6928));
 sg13g2_o21ai_1 _18700_ (.B1(_03239_),
    .Y(_01941_),
    .A1(net6928),
    .A2(net7481));
 sg13g2_nand2_1 _18701_ (.Y(_03240_),
    .A(net3296),
    .B(net6928));
 sg13g2_o21ai_1 _18702_ (.B1(_03240_),
    .Y(_01942_),
    .A1(net6928),
    .A2(net7637));
 sg13g2_nand2_1 _18703_ (.Y(_03241_),
    .A(net3611),
    .B(net6524));
 sg13g2_o21ai_1 _18704_ (.B1(_03241_),
    .Y(_01943_),
    .A1(net6524),
    .A2(net7182));
 sg13g2_nand2_1 _18705_ (.Y(_03242_),
    .A(net3848),
    .B(net6524));
 sg13g2_o21ai_1 _18706_ (.B1(_03242_),
    .Y(_01944_),
    .A1(net6524),
    .A2(net7479));
 sg13g2_nand2_1 _18707_ (.Y(_03243_),
    .A(net4545),
    .B(net6524));
 sg13g2_o21ai_1 _18708_ (.B1(_03243_),
    .Y(_01945_),
    .A1(net6524),
    .A2(net7638));
 sg13g2_nor2_1 _18709_ (.A(net4118),
    .B(net6526),
    .Y(_03244_));
 sg13g2_a21oi_1 _18710_ (.A1(net6526),
    .A2(net7124),
    .Y(_01946_),
    .B1(_03244_));
 sg13g2_nor2_1 _18711_ (.A(net4208),
    .B(net6527),
    .Y(_03245_));
 sg13g2_a21oi_1 _18712_ (.A1(net6527),
    .A2(net7419),
    .Y(_01947_),
    .B1(_03245_));
 sg13g2_nor2_1 _18713_ (.A(net4645),
    .B(net6527),
    .Y(_03246_));
 sg13g2_a21oi_1 _18714_ (.A1(net6527),
    .A2(net7578),
    .Y(_01948_),
    .B1(_03246_));
 sg13g2_nor2_1 _18715_ (.A(net4831),
    .B(net6704),
    .Y(_03247_));
 sg13g2_a21oi_1 _18716_ (.A1(net6704),
    .A2(net7118),
    .Y(_01949_),
    .B1(_03247_));
 sg13g2_nor2_1 _18717_ (.A(net4513),
    .B(net6704),
    .Y(_03248_));
 sg13g2_a21oi_1 _18718_ (.A1(net6704),
    .A2(net7414),
    .Y(_01950_),
    .B1(_03248_));
 sg13g2_nor2_1 _18719_ (.A(net4751),
    .B(net6704),
    .Y(_03249_));
 sg13g2_a21oi_1 _18720_ (.A1(net6704),
    .A2(net7573),
    .Y(_01951_),
    .B1(_03249_));
 sg13g2_nand2_1 _18721_ (.Y(_03250_),
    .A(net3222),
    .B(net6706));
 sg13g2_o21ai_1 _18722_ (.B1(_03250_),
    .Y(_01952_),
    .A1(net6706),
    .A2(net7125));
 sg13g2_nand2_1 _18723_ (.Y(_03251_),
    .A(net2544),
    .B(net6706));
 sg13g2_o21ai_1 _18724_ (.B1(_03251_),
    .Y(_01953_),
    .A1(net6706),
    .A2(net7417));
 sg13g2_nand2_1 _18725_ (.Y(_03252_),
    .A(net2518),
    .B(net6706));
 sg13g2_o21ai_1 _18726_ (.B1(_03252_),
    .Y(_01954_),
    .A1(net6706),
    .A2(net7579));
 sg13g2_nor2_1 _18727_ (.A(net4460),
    .B(net6709),
    .Y(_03253_));
 sg13g2_a21oi_1 _18728_ (.A1(net6708),
    .A2(net7157),
    .Y(_01955_),
    .B1(_03253_));
 sg13g2_nor2_1 _18729_ (.A(net4265),
    .B(net6709),
    .Y(_03254_));
 sg13g2_a21oi_1 _18730_ (.A1(net6709),
    .A2(net7454),
    .Y(_01956_),
    .B1(_03254_));
 sg13g2_nor2_1 _18731_ (.A(net4310),
    .B(net6708),
    .Y(_03255_));
 sg13g2_a21oi_1 _18732_ (.A1(net6708),
    .A2(net7615),
    .Y(_01957_),
    .B1(_03255_));
 sg13g2_nand2_1 _18733_ (.Y(_03256_),
    .A(net2727),
    .B(net6710));
 sg13g2_o21ai_1 _18734_ (.B1(_03256_),
    .Y(_01958_),
    .A1(net6710),
    .A2(net7171));
 sg13g2_nand2_1 _18735_ (.Y(_03257_),
    .A(net3391),
    .B(net6711));
 sg13g2_o21ai_1 _18736_ (.B1(_03257_),
    .Y(_01959_),
    .A1(net6711),
    .A2(net7467));
 sg13g2_nand2_1 _18737_ (.Y(_03258_),
    .A(net4268),
    .B(net6710));
 sg13g2_o21ai_1 _18738_ (.B1(_03258_),
    .Y(_01960_),
    .A1(net6710),
    .A2(net7626));
 sg13g2_nand2_1 _18739_ (.Y(_03259_),
    .A(net4097),
    .B(net6712));
 sg13g2_o21ai_1 _18740_ (.B1(_03259_),
    .Y(_01961_),
    .A1(net6712),
    .A2(net7175));
 sg13g2_nand2_1 _18741_ (.Y(_03260_),
    .A(net2747),
    .B(net6713));
 sg13g2_o21ai_1 _18742_ (.B1(_03260_),
    .Y(_01962_),
    .A1(net6713),
    .A2(net7471));
 sg13g2_nand2_1 _18743_ (.Y(_03261_),
    .A(net3962),
    .B(net6712));
 sg13g2_o21ai_1 _18744_ (.B1(_03261_),
    .Y(_01963_),
    .A1(net6712),
    .A2(net7627));
 sg13g2_nor2_1 _18745_ (.A(net4333),
    .B(net7061),
    .Y(_03262_));
 sg13g2_a21oi_1 _18746_ (.A1(net7061),
    .A2(net7129),
    .Y(_01964_),
    .B1(_03262_));
 sg13g2_nor2_1 _18747_ (.A(net4659),
    .B(net7061),
    .Y(_03263_));
 sg13g2_a21oi_1 _18748_ (.A1(net7061),
    .A2(net7424),
    .Y(_01965_),
    .B1(_03263_));
 sg13g2_nor2_1 _18749_ (.A(net4806),
    .B(net7061),
    .Y(_03264_));
 sg13g2_a21oi_1 _18750_ (.A1(net7061),
    .A2(net7583),
    .Y(_01966_),
    .B1(_03264_));
 sg13g2_nor2_1 _18751_ (.A(net4139),
    .B(net7063),
    .Y(_03265_));
 sg13g2_a21oi_1 _18752_ (.A1(net7063),
    .A2(net7130),
    .Y(_01967_),
    .B1(_03265_));
 sg13g2_nor2_1 _18753_ (.A(net4081),
    .B(net7063),
    .Y(_03266_));
 sg13g2_a21oi_1 _18754_ (.A1(net7063),
    .A2(net7425),
    .Y(_01968_),
    .B1(_03266_));
 sg13g2_nor2_1 _18755_ (.A(net4149),
    .B(net7063),
    .Y(_03267_));
 sg13g2_a21oi_1 _18756_ (.A1(net7063),
    .A2(net7584),
    .Y(_01969_),
    .B1(_03267_));
 sg13g2_nand2_1 _18757_ (.Y(_03268_),
    .A(net3204),
    .B(net7068));
 sg13g2_o21ai_1 _18758_ (.B1(_03268_),
    .Y(_01970_),
    .A1(net7068),
    .A2(net7132));
 sg13g2_nand2_1 _18759_ (.Y(_03269_),
    .A(net2688),
    .B(net7069));
 sg13g2_o21ai_1 _18760_ (.B1(_03269_),
    .Y(_01971_),
    .A1(net7069),
    .A2(net7441));
 sg13g2_nand2_1 _18761_ (.Y(_03270_),
    .A(net3512),
    .B(net7068));
 sg13g2_o21ai_1 _18762_ (.B1(_03270_),
    .Y(_01972_),
    .A1(net7068),
    .A2(net7587));
 sg13g2_nand2_1 _18763_ (.Y(_03271_),
    .A(net2639),
    .B(net7070));
 sg13g2_o21ai_1 _18764_ (.B1(_03271_),
    .Y(_01973_),
    .A1(net7070),
    .A2(net7132));
 sg13g2_nand2_1 _18765_ (.Y(_03272_),
    .A(net2439),
    .B(net7071));
 sg13g2_o21ai_1 _18766_ (.B1(_03272_),
    .Y(_01974_),
    .A1(net7070),
    .A2(net7439));
 sg13g2_nand2_1 _18767_ (.Y(_03273_),
    .A(net3236),
    .B(net7070));
 sg13g2_o21ai_1 _18768_ (.B1(_03273_),
    .Y(_01975_),
    .A1(net7071),
    .A2(net7588));
 sg13g2_nand2_1 _18769_ (.Y(_03274_),
    .A(net3012),
    .B(net6725));
 sg13g2_o21ai_1 _18770_ (.B1(_03274_),
    .Y(_01976_),
    .A1(net6724),
    .A2(net7148));
 sg13g2_nand2_1 _18771_ (.Y(_03275_),
    .A(net2478),
    .B(net6724));
 sg13g2_o21ai_1 _18772_ (.B1(_03275_),
    .Y(_01977_),
    .A1(net6724),
    .A2(net7443));
 sg13g2_nand2_1 _18773_ (.Y(_03276_),
    .A(net3547),
    .B(net6724));
 sg13g2_o21ai_1 _18774_ (.B1(_03276_),
    .Y(_01978_),
    .A1(net6725),
    .A2(net7601));
 sg13g2_nand2_1 _18775_ (.Y(_03277_),
    .A(net3880),
    .B(net7087));
 sg13g2_o21ai_1 _18776_ (.B1(_03277_),
    .Y(_01979_),
    .A1(net7087),
    .A2(net7168));
 sg13g2_nand2_1 _18777_ (.Y(_03278_),
    .A(net3241),
    .B(net7086));
 sg13g2_o21ai_1 _18778_ (.B1(_03278_),
    .Y(_01980_),
    .A1(net7086),
    .A2(net7466));
 sg13g2_nand2_1 _18779_ (.Y(_03279_),
    .A(net3248),
    .B(net7086));
 sg13g2_o21ai_1 _18780_ (.B1(_03279_),
    .Y(_01981_),
    .A1(net7086),
    .A2(net7623));
 sg13g2_nand2_1 _18781_ (.Y(_03280_),
    .A(net2918),
    .B(net7089));
 sg13g2_o21ai_1 _18782_ (.B1(_03280_),
    .Y(_01982_),
    .A1(net7089),
    .A2(net7168));
 sg13g2_nand2_1 _18783_ (.Y(_03281_),
    .A(net3080),
    .B(net7089));
 sg13g2_o21ai_1 _18784_ (.B1(_03281_),
    .Y(_01983_),
    .A1(net7089),
    .A2(net7463));
 sg13g2_nand2_1 _18785_ (.Y(_03282_),
    .A(net3345),
    .B(net7088));
 sg13g2_o21ai_1 _18786_ (.B1(_03282_),
    .Y(_01984_),
    .A1(net7088),
    .A2(net7623));
 sg13g2_nor2_1 _18787_ (.A(net4402),
    .B(net6726),
    .Y(_03283_));
 sg13g2_a21oi_1 _18788_ (.A1(net6726),
    .A2(net7145),
    .Y(_01985_),
    .B1(_03283_));
 sg13g2_nor2_1 _18789_ (.A(net4611),
    .B(net6727),
    .Y(_03284_));
 sg13g2_a21oi_1 _18790_ (.A1(net6727),
    .A2(net7438),
    .Y(_01986_),
    .B1(_03284_));
 sg13g2_nor2_1 _18791_ (.A(net4737),
    .B(net6726),
    .Y(_03285_));
 sg13g2_a21oi_1 _18792_ (.A1(net6726),
    .A2(net7600),
    .Y(_01987_),
    .B1(_03285_));
 sg13g2_nor2_1 _18793_ (.A(net4084),
    .B(net7090),
    .Y(_03286_));
 sg13g2_a21oi_1 _18794_ (.A1(net7090),
    .A2(net7150),
    .Y(_01988_),
    .B1(_03286_));
 sg13g2_nor2_1 _18795_ (.A(net4825),
    .B(net7091),
    .Y(_03287_));
 sg13g2_a21oi_1 _18796_ (.A1(net7091),
    .A2(net7445),
    .Y(_01989_),
    .B1(_03287_));
 sg13g2_nor2_1 _18797_ (.A(net3701),
    .B(net7090),
    .Y(_03288_));
 sg13g2_a21oi_1 _18798_ (.A1(net7090),
    .A2(net7603),
    .Y(_01990_),
    .B1(_03288_));
 sg13g2_nand2_1 _18799_ (.Y(_03289_),
    .A(net4091),
    .B(net6912));
 sg13g2_o21ai_1 _18800_ (.B1(_03289_),
    .Y(_01991_),
    .A1(net6912),
    .A2(net7163));
 sg13g2_nand2_1 _18801_ (.Y(_03290_),
    .A(net3002),
    .B(net6912));
 sg13g2_o21ai_1 _18802_ (.B1(_03290_),
    .Y(_01992_),
    .A1(net6912),
    .A2(net7460));
 sg13g2_nand2_1 _18803_ (.Y(_03291_),
    .A(net3753),
    .B(net6912));
 sg13g2_o21ai_1 _18804_ (.B1(_03291_),
    .Y(_01993_),
    .A1(net6912),
    .A2(net7617));
 sg13g2_nand2_1 _18805_ (.Y(_03292_),
    .A(net3131),
    .B(net6916));
 sg13g2_o21ai_1 _18806_ (.B1(_03292_),
    .Y(_01994_),
    .A1(net6916),
    .A2(net7163));
 sg13g2_nand2_1 _18807_ (.Y(_03293_),
    .A(net3135),
    .B(net6916));
 sg13g2_o21ai_1 _18808_ (.B1(_03293_),
    .Y(_01995_),
    .A1(net6916),
    .A2(net7460));
 sg13g2_nand2_1 _18809_ (.Y(_03294_),
    .A(net3443),
    .B(net6916));
 sg13g2_o21ai_1 _18810_ (.B1(_03294_),
    .Y(_01996_),
    .A1(net6916),
    .A2(net7617));
 sg13g2_nand2_1 _18811_ (.Y(_03295_),
    .A(net2698),
    .B(net6918));
 sg13g2_o21ai_1 _18812_ (.B1(_03295_),
    .Y(_01997_),
    .A1(net6918),
    .A2(net7165));
 sg13g2_nand2_1 _18813_ (.Y(_03296_),
    .A(net3544),
    .B(net6918));
 sg13g2_o21ai_1 _18814_ (.B1(_03296_),
    .Y(_01998_),
    .A1(net6918),
    .A2(net7461));
 sg13g2_nand2_1 _18815_ (.Y(_03297_),
    .A(net3412),
    .B(net6918));
 sg13g2_o21ai_1 _18816_ (.B1(_03297_),
    .Y(_01999_),
    .A1(net6918),
    .A2(net7616));
 sg13g2_nand2_1 _18817_ (.Y(_03298_),
    .A(net3950),
    .B(net6920));
 sg13g2_o21ai_1 _18818_ (.B1(_03298_),
    .Y(_02000_),
    .A1(net6920),
    .A2(net7163));
 sg13g2_nand2_1 _18819_ (.Y(_03299_),
    .A(net3455),
    .B(net6920));
 sg13g2_o21ai_1 _18820_ (.B1(_03299_),
    .Y(_02001_),
    .A1(net6920),
    .A2(net7460));
 sg13g2_nand2_1 _18821_ (.Y(_03300_),
    .A(net3099),
    .B(net6920));
 sg13g2_o21ai_1 _18822_ (.B1(_03300_),
    .Y(_02002_),
    .A1(net6920),
    .A2(net7616));
 sg13g2_nand2_1 _18823_ (.Y(_03301_),
    .A(net2477),
    .B(net6517));
 sg13g2_o21ai_1 _18824_ (.B1(_03301_),
    .Y(_02003_),
    .A1(net6517),
    .A2(net7163));
 sg13g2_nand2_1 _18825_ (.Y(_03302_),
    .A(net2630),
    .B(net6516));
 sg13g2_o21ai_1 _18826_ (.B1(_03302_),
    .Y(_02004_),
    .A1(net6516),
    .A2(net7458));
 sg13g2_nand2_1 _18827_ (.Y(_03303_),
    .A(net4317),
    .B(net6516));
 sg13g2_o21ai_1 _18828_ (.B1(_03303_),
    .Y(_02005_),
    .A1(net6516),
    .A2(net7618));
 sg13g2_nand2_1 _18829_ (.Y(_03304_),
    .A(net3603),
    .B(net6519));
 sg13g2_o21ai_1 _18830_ (.B1(_03304_),
    .Y(_02006_),
    .A1(net6519),
    .A2(net7163));
 sg13g2_nand2_1 _18831_ (.Y(_03305_),
    .A(net3746),
    .B(net6518));
 sg13g2_o21ai_1 _18832_ (.B1(_03305_),
    .Y(_02007_),
    .A1(net6518),
    .A2(net7458));
 sg13g2_nand2_1 _18833_ (.Y(_03306_),
    .A(net2685),
    .B(net6518));
 sg13g2_o21ai_1 _18834_ (.B1(_03306_),
    .Y(_02008_),
    .A1(net6518),
    .A2(net7618));
 sg13g2_nand2_1 _18835_ (.Y(_03307_),
    .A(net4013),
    .B(net6523));
 sg13g2_o21ai_1 _18836_ (.B1(_03307_),
    .Y(_02009_),
    .A1(net6523),
    .A2(net7163));
 sg13g2_nand2_1 _18837_ (.Y(_03308_),
    .A(net2673),
    .B(net6522));
 sg13g2_o21ai_1 _18838_ (.B1(_03308_),
    .Y(_02010_),
    .A1(net6522),
    .A2(net7458));
 sg13g2_nand2_1 _18839_ (.Y(_03309_),
    .A(net3582),
    .B(net6522));
 sg13g2_o21ai_1 _18840_ (.B1(_03309_),
    .Y(_02011_),
    .A1(net6522),
    .A2(net7618));
 sg13g2_nand2_1 _18841_ (.Y(_03310_),
    .A(net2606),
    .B(net6703));
 sg13g2_o21ai_1 _18842_ (.B1(_03310_),
    .Y(_02012_),
    .A1(net6703),
    .A2(net7163));
 sg13g2_nand2_1 _18843_ (.Y(_03311_),
    .A(net4294),
    .B(net6702));
 sg13g2_o21ai_1 _18844_ (.B1(_03311_),
    .Y(_02013_),
    .A1(net6702),
    .A2(net7458));
 sg13g2_nand2_1 _18845_ (.Y(_03312_),
    .A(net2619),
    .B(net6702));
 sg13g2_o21ai_1 _18846_ (.B1(_03312_),
    .Y(_02014_),
    .A1(net6702),
    .A2(net7618));
 sg13g2_nand2_1 _18847_ (.Y(_03313_),
    .A(net2486),
    .B(net7053));
 sg13g2_o21ai_1 _18848_ (.B1(_03313_),
    .Y(_02015_),
    .A1(net7054),
    .A2(net7151));
 sg13g2_nand2_1 _18849_ (.Y(_03314_),
    .A(net4231),
    .B(net7053));
 sg13g2_o21ai_1 _18850_ (.B1(_03314_),
    .Y(_02016_),
    .A1(net7053),
    .A2(net7444));
 sg13g2_nand2_1 _18851_ (.Y(_03315_),
    .A(net2555),
    .B(net7053));
 sg13g2_o21ai_1 _18852_ (.B1(_03315_),
    .Y(_02017_),
    .A1(net7054),
    .A2(net7604));
 sg13g2_nor2_1 _18853_ (.A(net4133),
    .B(net7055),
    .Y(_03316_));
 sg13g2_a21oi_1 _18854_ (.A1(net7055),
    .A2(net7150),
    .Y(_02018_),
    .B1(_03316_));
 sg13g2_nor2_1 _18855_ (.A(net4316),
    .B(net7055),
    .Y(_03317_));
 sg13g2_a21oi_1 _18856_ (.A1(net7056),
    .A2(net7445),
    .Y(_02019_),
    .B1(_03317_));
 sg13g2_nor2_1 _18857_ (.A(net4753),
    .B(net7055),
    .Y(_03318_));
 sg13g2_a21oi_1 _18858_ (.A1(net7055),
    .A2(net7603),
    .Y(_02020_),
    .B1(_03318_));
 sg13g2_nand2_1 _18859_ (.Y(_03319_),
    .A(net3645),
    .B(net7058));
 sg13g2_o21ai_1 _18860_ (.B1(_03319_),
    .Y(_02021_),
    .A1(net7058),
    .A2(net7163));
 sg13g2_nand2_1 _18861_ (.Y(_03320_),
    .A(net3243),
    .B(net7057));
 sg13g2_o21ai_1 _18862_ (.B1(_03320_),
    .Y(_02022_),
    .A1(net7057),
    .A2(net7444));
 sg13g2_nand2_1 _18863_ (.Y(_03321_),
    .A(net2609),
    .B(net7057));
 sg13g2_o21ai_1 _18864_ (.B1(_03321_),
    .Y(_02023_),
    .A1(net7057),
    .A2(net7604));
 sg13g2_nand2_1 _18865_ (.Y(_03322_),
    .A(net2474),
    .B(net7059));
 sg13g2_o21ai_1 _18866_ (.B1(_03322_),
    .Y(_02024_),
    .A1(net7059),
    .A2(net7151));
 sg13g2_nand2_1 _18867_ (.Y(_03323_),
    .A(net2981),
    .B(net7060));
 sg13g2_o21ai_1 _18868_ (.B1(_03323_),
    .Y(_02025_),
    .A1(net7060),
    .A2(net7444));
 sg13g2_nand2_1 _18869_ (.Y(_03324_),
    .A(net3163),
    .B(net7059));
 sg13g2_o21ai_1 _18870_ (.B1(_03324_),
    .Y(_02026_),
    .A1(net7059),
    .A2(net7604));
 sg13g2_nand2_1 _18871_ (.Y(_03325_),
    .A(net3636),
    .B(net6714));
 sg13g2_o21ai_1 _18872_ (.B1(_03325_),
    .Y(_02027_),
    .A1(net6714),
    .A2(net7169));
 sg13g2_nand2_1 _18873_ (.Y(_03326_),
    .A(net3198),
    .B(net6715));
 sg13g2_o21ai_1 _18874_ (.B1(_03326_),
    .Y(_02028_),
    .A1(net6715),
    .A2(net7464));
 sg13g2_nand2_1 _18875_ (.Y(_03327_),
    .A(net2548),
    .B(net6714));
 sg13g2_o21ai_1 _18876_ (.B1(_03327_),
    .Y(_02029_),
    .A1(net6714),
    .A2(net7621));
 sg13g2_nand2_1 _18877_ (.Y(_03328_),
    .A(net3961),
    .B(net6716));
 sg13g2_o21ai_1 _18878_ (.B1(_03328_),
    .Y(_02030_),
    .A1(net6716),
    .A2(net7169));
 sg13g2_nand2_1 _18879_ (.Y(_03329_),
    .A(net4088),
    .B(net6717));
 sg13g2_o21ai_1 _18880_ (.B1(_03329_),
    .Y(_02031_),
    .A1(net6717),
    .A2(net7464));
 sg13g2_nand2_1 _18881_ (.Y(_03330_),
    .A(net2979),
    .B(net6716));
 sg13g2_o21ai_1 _18882_ (.B1(_03330_),
    .Y(_02032_),
    .A1(net6716),
    .A2(net7621));
 sg13g2_nand2_1 _18883_ (.Y(_03331_),
    .A(net3185),
    .B(net6718));
 sg13g2_o21ai_1 _18884_ (.B1(_03331_),
    .Y(_02033_),
    .A1(net6718),
    .A2(net7169));
 sg13g2_nand2_1 _18885_ (.Y(_03332_),
    .A(net2902),
    .B(net6719));
 sg13g2_o21ai_1 _18886_ (.B1(_03332_),
    .Y(_02034_),
    .A1(net6719),
    .A2(net7464));
 sg13g2_nand2_1 _18887_ (.Y(_03333_),
    .A(net2682),
    .B(net6718));
 sg13g2_o21ai_1 _18888_ (.B1(_03333_),
    .Y(_02035_),
    .A1(net6718),
    .A2(net7620));
 sg13g2_nand2_1 _18889_ (.Y(_03334_),
    .A(net2888),
    .B(net6720));
 sg13g2_o21ai_1 _18890_ (.B1(_03334_),
    .Y(_02036_),
    .A1(net6720),
    .A2(net7169));
 sg13g2_nand2_1 _18891_ (.Y(_03335_),
    .A(net4290),
    .B(net6721));
 sg13g2_o21ai_1 _18892_ (.B1(_03335_),
    .Y(_02037_),
    .A1(net6721),
    .A2(net7464));
 sg13g2_nand2_1 _18893_ (.Y(_03336_),
    .A(net3195),
    .B(net6720));
 sg13g2_o21ai_1 _18894_ (.B1(_03336_),
    .Y(_02038_),
    .A1(net6720),
    .A2(net7620));
 sg13g2_nand2_1 _18895_ (.Y(_03337_),
    .A(net2626),
    .B(net6723));
 sg13g2_o21ai_1 _18896_ (.B1(_03337_),
    .Y(_02039_),
    .A1(net6723),
    .A2(net7167));
 sg13g2_nand2_1 _18897_ (.Y(_03338_),
    .A(net2554),
    .B(net6722));
 sg13g2_o21ai_1 _18898_ (.B1(_03338_),
    .Y(_02040_),
    .A1(net6722),
    .A2(net7465));
 sg13g2_nand2_1 _18899_ (.Y(_03339_),
    .A(net2538),
    .B(net6722));
 sg13g2_o21ai_1 _18900_ (.B1(_03339_),
    .Y(_02041_),
    .A1(net6722),
    .A2(net7624));
 sg13g2_nand2_1 _18901_ (.Y(_03340_),
    .A(net3925),
    .B(net6501));
 sg13g2_o21ai_1 _18902_ (.B1(_03340_),
    .Y(_02042_),
    .A1(net6501),
    .A2(net7166));
 sg13g2_nand2_1 _18903_ (.Y(_03341_),
    .A(net2483),
    .B(net6500));
 sg13g2_o21ai_1 _18904_ (.B1(_03341_),
    .Y(_02043_),
    .A1(net6500),
    .A2(net7465));
 sg13g2_nand2_1 _18905_ (.Y(_03342_),
    .A(net3397),
    .B(net6500));
 sg13g2_o21ai_1 _18906_ (.B1(_03342_),
    .Y(_02044_),
    .A1(net6500),
    .A2(net7624));
 sg13g2_nand2_1 _18907_ (.Y(_03343_),
    .A(net4108),
    .B(net6531));
 sg13g2_o21ai_1 _18908_ (.B1(_03343_),
    .Y(_02045_),
    .A1(net6531),
    .A2(net7166));
 sg13g2_nand2_1 _18909_ (.Y(_03344_),
    .A(net3094),
    .B(net6530));
 sg13g2_o21ai_1 _18910_ (.B1(_03344_),
    .Y(_02046_),
    .A1(net6530),
    .A2(net7465));
 sg13g2_nand2_1 _18911_ (.Y(_03345_),
    .A(net3318),
    .B(net6530));
 sg13g2_o21ai_1 _18912_ (.B1(_03345_),
    .Y(_02047_),
    .A1(net6530),
    .A2(net7624));
 sg13g2_nor2_1 _18913_ (.A(net4330),
    .B(net7046),
    .Y(_03346_));
 sg13g2_a21oi_1 _18914_ (.A1(net7046),
    .A2(net7150),
    .Y(_02048_),
    .B1(_03346_));
 sg13g2_nor2_1 _18915_ (.A(net4455),
    .B(net7046),
    .Y(_03347_));
 sg13g2_a21oi_1 _18916_ (.A1(net7047),
    .A2(net7446),
    .Y(_02049_),
    .B1(_03347_));
 sg13g2_nor2_1 _18917_ (.A(net4707),
    .B(net7046),
    .Y(_03348_));
 sg13g2_a21oi_1 _18918_ (.A1(net7046),
    .A2(net7603),
    .Y(_02050_),
    .B1(_03348_));
 sg13g2_nand2_1 _18919_ (.Y(_03349_),
    .A(net2468),
    .B(net6529));
 sg13g2_o21ai_1 _18920_ (.B1(_03349_),
    .Y(_02051_),
    .A1(net6529),
    .A2(net7166));
 sg13g2_nand2_1 _18921_ (.Y(_03350_),
    .A(net3055),
    .B(net6528));
 sg13g2_o21ai_1 _18922_ (.B1(_03350_),
    .Y(_02052_),
    .A1(net6528),
    .A2(net7478));
 sg13g2_nand2_1 _18923_ (.Y(_03351_),
    .A(net2459),
    .B(net6528));
 sg13g2_o21ai_1 _18924_ (.B1(_03351_),
    .Y(_02053_),
    .A1(net6528),
    .A2(net7621));
 sg13g2_nand2_1 _18925_ (.Y(_03352_),
    .A(net3253),
    .B(net6503));
 sg13g2_o21ai_1 _18926_ (.B1(_03352_),
    .Y(_02054_),
    .A1(net6503),
    .A2(net7166));
 sg13g2_nand2_1 _18927_ (.Y(_03353_),
    .A(net2765),
    .B(net6502));
 sg13g2_o21ai_1 _18928_ (.B1(_03353_),
    .Y(_02055_),
    .A1(net6502),
    .A2(net7478));
 sg13g2_nand2_1 _18929_ (.Y(_03354_),
    .A(net3609),
    .B(net6502));
 sg13g2_o21ai_1 _18930_ (.B1(_03354_),
    .Y(_02056_),
    .A1(net6502),
    .A2(net7621));
 sg13g2_nand2_1 _18931_ (.Y(_03355_),
    .A(net3912),
    .B(net6533));
 sg13g2_o21ai_1 _18932_ (.B1(_03355_),
    .Y(_02057_),
    .A1(net6533),
    .A2(net7166));
 sg13g2_nand2_1 _18933_ (.Y(_03356_),
    .A(net3472),
    .B(net6532));
 sg13g2_o21ai_1 _18934_ (.B1(_03356_),
    .Y(_02058_),
    .A1(net6532),
    .A2(net7478));
 sg13g2_nand2_1 _18935_ (.Y(_03357_),
    .A(net3759),
    .B(net6532));
 sg13g2_o21ai_1 _18936_ (.B1(_03357_),
    .Y(_02059_),
    .A1(net6532),
    .A2(net7620));
 sg13g2_nand2_1 _18937_ (.Y(_03358_),
    .A(net2646),
    .B(net6537));
 sg13g2_o21ai_1 _18938_ (.B1(_03358_),
    .Y(_02060_),
    .A1(net6537),
    .A2(net7166));
 sg13g2_nand2_1 _18939_ (.Y(_03359_),
    .A(net2753),
    .B(net6536));
 sg13g2_o21ai_1 _18940_ (.B1(_03359_),
    .Y(_02061_),
    .A1(net6536),
    .A2(net7477));
 sg13g2_nand2_1 _18941_ (.Y(_03360_),
    .A(net2745),
    .B(net6536));
 sg13g2_o21ai_1 _18942_ (.B1(_03360_),
    .Y(_02062_),
    .A1(net6536),
    .A2(net7620));
 sg13g2_nand2_1 _18943_ (.Y(_03361_),
    .A(net2553),
    .B(net6538));
 sg13g2_o21ai_1 _18944_ (.B1(_03361_),
    .Y(_02063_),
    .A1(net6538),
    .A2(net7167));
 sg13g2_nand2_1 _18945_ (.Y(_03362_),
    .A(net3001),
    .B(net6538));
 sg13g2_o21ai_1 _18946_ (.B1(_03362_),
    .Y(_02064_),
    .A1(net6538),
    .A2(net7480));
 sg13g2_nand2_1 _18947_ (.Y(_03363_),
    .A(net2484),
    .B(net6538));
 sg13g2_o21ai_1 _18948_ (.B1(_03363_),
    .Y(_02065_),
    .A1(net6538),
    .A2(net7624));
 sg13g2_nand2_1 _18949_ (.Y(_03364_),
    .A(net3471),
    .B(net6700));
 sg13g2_o21ai_1 _18950_ (.B1(_03364_),
    .Y(_02066_),
    .A1(net6700),
    .A2(net7167));
 sg13g2_nand2_1 _18951_ (.Y(_03365_),
    .A(net3562),
    .B(net6700));
 sg13g2_o21ai_1 _18952_ (.B1(_03365_),
    .Y(_02067_),
    .A1(net6700),
    .A2(net7480));
 sg13g2_nand2_1 _18953_ (.Y(_03366_),
    .A(net2998),
    .B(net6700));
 sg13g2_o21ai_1 _18954_ (.B1(_03366_),
    .Y(_02068_),
    .A1(net6700),
    .A2(net7624));
 sg13g2_nand2_1 _18955_ (.Y(_03367_),
    .A(net3999),
    .B(net6534));
 sg13g2_o21ai_1 _18956_ (.B1(_03367_),
    .Y(_02069_),
    .A1(net6534),
    .A2(net7166));
 sg13g2_nand2_1 _18957_ (.Y(_03368_),
    .A(net4384),
    .B(net6534));
 sg13g2_o21ai_1 _18958_ (.B1(_03368_),
    .Y(_02070_),
    .A1(net6534),
    .A2(net7480));
 sg13g2_nand2_1 _18959_ (.Y(_03369_),
    .A(net2650),
    .B(net6534));
 sg13g2_o21ai_1 _18960_ (.B1(_03369_),
    .Y(_02071_),
    .A1(net6534),
    .A2(net7624));
 sg13g2_nand2_1 _18961_ (.Y(_03370_),
    .A(net3324),
    .B(net6504));
 sg13g2_o21ai_1 _18962_ (.B1(_03370_),
    .Y(_02072_),
    .A1(net6504),
    .A2(net7166));
 sg13g2_nand2_1 _18963_ (.Y(_03371_),
    .A(net3794),
    .B(net6504));
 sg13g2_o21ai_1 _18964_ (.B1(_03371_),
    .Y(_02073_),
    .A1(net6504),
    .A2(net7480));
 sg13g2_nand2_1 _18965_ (.Y(_03372_),
    .A(net2653),
    .B(net6504));
 sg13g2_o21ai_1 _18966_ (.B1(_03372_),
    .Y(_02074_),
    .A1(net6504),
    .A2(net7624));
 sg13g2_nand2_1 _18967_ (.Y(_03373_),
    .A(net2687),
    .B(net6915));
 sg13g2_o21ai_1 _18968_ (.B1(_03373_),
    .Y(_02075_),
    .A1(net6915),
    .A2(net7184));
 sg13g2_nand2_1 _18969_ (.Y(_03374_),
    .A(net2924),
    .B(net6914));
 sg13g2_o21ai_1 _18970_ (.B1(_03374_),
    .Y(_02076_),
    .A1(net6914),
    .A2(net7481));
 sg13g2_nand2_1 _18971_ (.Y(_03375_),
    .A(net2628),
    .B(net6914));
 sg13g2_o21ai_1 _18972_ (.B1(_03375_),
    .Y(_02077_),
    .A1(net6914),
    .A2(net7637));
 sg13g2_nor2_1 _18973_ (.A(net4162),
    .B(net6542),
    .Y(_03376_));
 sg13g2_a21oi_1 _18974_ (.A1(net6542),
    .A2(net7149),
    .Y(_02078_),
    .B1(_03376_));
 sg13g2_nor2_1 _18975_ (.A(net3855),
    .B(net6542),
    .Y(_03377_));
 sg13g2_a21oi_1 _18976_ (.A1(net6542),
    .A2(net7444),
    .Y(_02079_),
    .B1(_03377_));
 sg13g2_nor2_1 _18977_ (.A(net4743),
    .B(net6542),
    .Y(_03378_));
 sg13g2_a21oi_1 _18978_ (.A1(net6542),
    .A2(net7603),
    .Y(_02080_),
    .B1(_03378_));
 sg13g2_nand2_1 _18979_ (.Y(_03379_),
    .A(net3574),
    .B(net6931));
 sg13g2_o21ai_1 _18980_ (.B1(_03379_),
    .Y(_02081_),
    .A1(net6931),
    .A2(net7184));
 sg13g2_nand2_1 _18981_ (.Y(_03380_),
    .A(net4419),
    .B(net6930));
 sg13g2_o21ai_1 _18982_ (.B1(_03380_),
    .Y(_02082_),
    .A1(net6930),
    .A2(net7481));
 sg13g2_nand2_1 _18983_ (.Y(_03381_),
    .A(net3581),
    .B(net6930));
 sg13g2_o21ai_1 _18984_ (.B1(_03381_),
    .Y(_02083_),
    .A1(net6930),
    .A2(net7637));
 sg13g2_nand2_1 _18985_ (.Y(_03382_),
    .A(net2828),
    .B(net6933));
 sg13g2_o21ai_1 _18986_ (.B1(_03382_),
    .Y(_02084_),
    .A1(net6933),
    .A2(net7184));
 sg13g2_nand2_1 _18987_ (.Y(_03383_),
    .A(net2552),
    .B(net6932));
 sg13g2_o21ai_1 _18988_ (.B1(_03383_),
    .Y(_02085_),
    .A1(net6932),
    .A2(net7481));
 sg13g2_nand2_1 _18989_ (.Y(_03384_),
    .A(net3552),
    .B(net6932));
 sg13g2_o21ai_1 _18990_ (.B1(_03384_),
    .Y(_02086_),
    .A1(net6932),
    .A2(net7637));
 sg13g2_nand2_1 _18991_ (.Y(_03385_),
    .A(net4082),
    .B(net6934));
 sg13g2_o21ai_1 _18992_ (.B1(_03385_),
    .Y(_02087_),
    .A1(net6934),
    .A2(net7183));
 sg13g2_nand2_1 _18993_ (.Y(_03386_),
    .A(net2652),
    .B(net6934));
 sg13g2_o21ai_1 _18994_ (.B1(_03386_),
    .Y(_02088_),
    .A1(net6934),
    .A2(net7477));
 sg13g2_nand2_1 _18995_ (.Y(_03387_),
    .A(net3838),
    .B(net6934));
 sg13g2_o21ai_1 _18996_ (.B1(_03387_),
    .Y(_02089_),
    .A1(net6934),
    .A2(net7636));
 sg13g2_nand2_1 _18997_ (.Y(_03388_),
    .A(net4257),
    .B(net6936));
 sg13g2_o21ai_1 _18998_ (.B1(_03388_),
    .Y(_02090_),
    .A1(net6936),
    .A2(net7183));
 sg13g2_nand2_1 _18999_ (.Y(_03389_),
    .A(net4170),
    .B(net6936));
 sg13g2_o21ai_1 _19000_ (.B1(_03389_),
    .Y(_02091_),
    .A1(net6936),
    .A2(net7477));
 sg13g2_nand2_1 _19001_ (.Y(_03390_),
    .A(net3277),
    .B(net6936));
 sg13g2_o21ai_1 _19002_ (.B1(_03390_),
    .Y(_02092_),
    .A1(net6936),
    .A2(net7637));
 sg13g2_nand2_1 _19003_ (.Y(_03391_),
    .A(net4044),
    .B(net6938));
 sg13g2_o21ai_1 _19004_ (.B1(_03391_),
    .Y(_02093_),
    .A1(net6938),
    .A2(net7183));
 sg13g2_nand2_1 _19005_ (.Y(_03392_),
    .A(net3006),
    .B(net6938));
 sg13g2_o21ai_1 _19006_ (.B1(_03392_),
    .Y(_02094_),
    .A1(net6938),
    .A2(net7477));
 sg13g2_nand2_1 _19007_ (.Y(_03393_),
    .A(net3489),
    .B(net6938));
 sg13g2_o21ai_1 _19008_ (.B1(_03393_),
    .Y(_02095_),
    .A1(net6938),
    .A2(net7637));
 sg13g2_nand2_1 _19009_ (.Y(_03394_),
    .A(net2465),
    .B(net6940));
 sg13g2_o21ai_1 _19010_ (.B1(_03394_),
    .Y(_02096_),
    .A1(net6940),
    .A2(net7183));
 sg13g2_nand2_1 _19011_ (.Y(_03395_),
    .A(net3671),
    .B(net6940));
 sg13g2_o21ai_1 _19012_ (.B1(_03395_),
    .Y(_02097_),
    .A1(net6940),
    .A2(net7480));
 sg13g2_nand2_1 _19013_ (.Y(_03396_),
    .A(net2543),
    .B(net6940));
 sg13g2_o21ai_1 _19014_ (.B1(_03396_),
    .Y(_02098_),
    .A1(net6940),
    .A2(net7637));
 sg13g2_nand2_1 _19015_ (.Y(_03397_),
    .A(net2900),
    .B(net6550));
 sg13g2_o21ai_1 _19016_ (.B1(_03397_),
    .Y(_02099_),
    .A1(net6550),
    .A2(net7182));
 sg13g2_nand2_1 _19017_ (.Y(_03398_),
    .A(net2545),
    .B(net6550));
 sg13g2_o21ai_1 _19018_ (.B1(_03398_),
    .Y(_02100_),
    .A1(net6550),
    .A2(net7479));
 sg13g2_nand2_1 _19019_ (.Y(_03399_),
    .A(net2480),
    .B(net6550));
 sg13g2_o21ai_1 _19020_ (.B1(_03399_),
    .Y(_02101_),
    .A1(net6550),
    .A2(net7636));
 sg13g2_nand2_1 _19021_ (.Y(_03400_),
    .A(net3587),
    .B(net6552));
 sg13g2_o21ai_1 _19022_ (.B1(_03400_),
    .Y(_02102_),
    .A1(net6552),
    .A2(net7182));
 sg13g2_nand2_1 _19023_ (.Y(_03401_),
    .A(net2733),
    .B(net6552));
 sg13g2_o21ai_1 _19024_ (.B1(_03401_),
    .Y(_02103_),
    .A1(net6552),
    .A2(net7479));
 sg13g2_nand2_1 _19025_ (.Y(_03402_),
    .A(net3758),
    .B(net6552));
 sg13g2_o21ai_1 _19026_ (.B1(_03402_),
    .Y(_02104_),
    .A1(net6552),
    .A2(net7638));
 sg13g2_nand2_1 _19027_ (.Y(_03403_),
    .A(net4370),
    .B(net6554));
 sg13g2_o21ai_1 _19028_ (.B1(_03403_),
    .Y(_02105_),
    .A1(net6554),
    .A2(net7182));
 sg13g2_nand2_1 _19029_ (.Y(_03404_),
    .A(net3368),
    .B(net6554));
 sg13g2_o21ai_1 _19030_ (.B1(_03404_),
    .Y(_02106_),
    .A1(net6554),
    .A2(net7479));
 sg13g2_nand2_1 _19031_ (.Y(_03405_),
    .A(net3004),
    .B(net6554));
 sg13g2_o21ai_1 _19032_ (.B1(_03405_),
    .Y(_02107_),
    .A1(net6554),
    .A2(net7636));
 sg13g2_nor2_1 _19033_ (.A(net4087),
    .B(net6558),
    .Y(_03406_));
 sg13g2_a21oi_1 _19034_ (.A1(net6558),
    .A2(net7149),
    .Y(_02108_),
    .B1(_03406_));
 sg13g2_nor2_1 _19035_ (.A(net4263),
    .B(net6558),
    .Y(_03407_));
 sg13g2_a21oi_1 _19036_ (.A1(net6558),
    .A2(net7444),
    .Y(_02109_),
    .B1(_03407_));
 sg13g2_nor2_1 _19037_ (.A(net4423),
    .B(net6558),
    .Y(_03408_));
 sg13g2_a21oi_1 _19038_ (.A1(net6558),
    .A2(net7601),
    .Y(_02110_),
    .B1(_03408_));
 sg13g2_nand2_1 _19039_ (.Y(_03409_),
    .A(net3196),
    .B(net6945));
 sg13g2_o21ai_1 _19040_ (.B1(_03409_),
    .Y(_02111_),
    .A1(net6945),
    .A2(net7183));
 sg13g2_nand2_1 _19041_ (.Y(_03410_),
    .A(net3445),
    .B(net6944));
 sg13g2_o21ai_1 _19042_ (.B1(_03410_),
    .Y(_02112_),
    .A1(net6944),
    .A2(net7481));
 sg13g2_nand2_1 _19043_ (.Y(_03411_),
    .A(net4184),
    .B(net6944));
 sg13g2_o21ai_1 _19044_ (.B1(_03411_),
    .Y(_02113_),
    .A1(net6944),
    .A2(net7638));
 sg13g2_nand2_1 _19045_ (.Y(_03412_),
    .A(net2922),
    .B(net6947));
 sg13g2_o21ai_1 _19046_ (.B1(_03412_),
    .Y(_02114_),
    .A1(net6947),
    .A2(net7183));
 sg13g2_nand2_1 _19047_ (.Y(_03413_),
    .A(net2781),
    .B(net6946));
 sg13g2_o21ai_1 _19048_ (.B1(_03413_),
    .Y(_02115_),
    .A1(net6946),
    .A2(net7480));
 sg13g2_nand2_1 _19049_ (.Y(_03414_),
    .A(net3687),
    .B(net6946));
 sg13g2_o21ai_1 _19050_ (.B1(_03414_),
    .Y(_02116_),
    .A1(net6946),
    .A2(net7638));
 sg13g2_nand2_1 _19051_ (.Y(_03415_),
    .A(net3791),
    .B(net6949));
 sg13g2_o21ai_1 _19052_ (.B1(_03415_),
    .Y(_02117_),
    .A1(net6949),
    .A2(net7183));
 sg13g2_nand2_1 _19053_ (.Y(_03416_),
    .A(net3618),
    .B(net6948));
 sg13g2_o21ai_1 _19054_ (.B1(_03416_),
    .Y(_02118_),
    .A1(net6948),
    .A2(net7480));
 sg13g2_nand2_1 _19055_ (.Y(_03417_),
    .A(net2802),
    .B(net6948));
 sg13g2_o21ai_1 _19056_ (.B1(_03417_),
    .Y(_02119_),
    .A1(net6948),
    .A2(net7638));
 sg13g2_nand2_1 _19057_ (.Y(_03418_),
    .A(net3520),
    .B(net6951));
 sg13g2_o21ai_1 _19058_ (.B1(_03418_),
    .Y(_02120_),
    .A1(net6951),
    .A2(net7183));
 sg13g2_nand2_1 _19059_ (.Y(_03419_),
    .A(net3857),
    .B(net6950));
 sg13g2_o21ai_1 _19060_ (.B1(_03419_),
    .Y(_02121_),
    .A1(net6950),
    .A2(net7480));
 sg13g2_nand2_1 _19061_ (.Y(_03420_),
    .A(net3413),
    .B(net6950));
 sg13g2_o21ai_1 _19062_ (.B1(_03420_),
    .Y(_02122_),
    .A1(net6950),
    .A2(net7637));
 sg13g2_nor2_1 _19063_ (.A(net4681),
    .B(net6564),
    .Y(_03421_));
 sg13g2_a21oi_1 _19064_ (.A1(net6564),
    .A2(net7118),
    .Y(_02123_),
    .B1(_03421_));
 sg13g2_nor2_1 _19065_ (.A(net4629),
    .B(net6564),
    .Y(_03422_));
 sg13g2_a21oi_1 _19066_ (.A1(net6564),
    .A2(net7413),
    .Y(_02124_),
    .B1(_03422_));
 sg13g2_nor2_1 _19067_ (.A(net4762),
    .B(net6564),
    .Y(_03423_));
 sg13g2_a21oi_1 _19068_ (.A1(net6564),
    .A2(net7573),
    .Y(_02125_),
    .B1(_03423_));
 sg13g2_nor2_1 _19069_ (.A(net4124),
    .B(net6568),
    .Y(_03424_));
 sg13g2_a21oi_1 _19070_ (.A1(net6568),
    .A2(net7118),
    .Y(_02126_),
    .B1(_03424_));
 sg13g2_nor2_1 _19071_ (.A(net4723),
    .B(net6568),
    .Y(_03425_));
 sg13g2_a21oi_1 _19072_ (.A1(net6568),
    .A2(net7413),
    .Y(_02127_),
    .B1(_03425_));
 sg13g2_nor2_1 _19073_ (.A(net4644),
    .B(net6568),
    .Y(_03426_));
 sg13g2_a21oi_1 _19074_ (.A1(net6568),
    .A2(net7573),
    .Y(_02128_),
    .B1(_03426_));
 sg13g2_nor2_1 _19075_ (.A(net4225),
    .B(net6570),
    .Y(_03427_));
 sg13g2_a21oi_1 _19076_ (.A1(net6570),
    .A2(net7118),
    .Y(_02129_),
    .B1(_03427_));
 sg13g2_nor2_1 _19077_ (.A(net4812),
    .B(net6570),
    .Y(_03428_));
 sg13g2_a21oi_1 _19078_ (.A1(net6570),
    .A2(net7413),
    .Y(_02130_),
    .B1(_03428_));
 sg13g2_nor2_1 _19079_ (.A(net4643),
    .B(net6570),
    .Y(_03429_));
 sg13g2_a21oi_1 _19080_ (.A1(net6570),
    .A2(net7573),
    .Y(_02131_),
    .B1(_03429_));
 sg13g2_nor2_1 _19081_ (.A(net4790),
    .B(net6574),
    .Y(_03430_));
 sg13g2_a21oi_1 _19082_ (.A1(net6574),
    .A2(net7118),
    .Y(_02132_),
    .B1(_03430_));
 sg13g2_nor2_1 _19083_ (.A(net4510),
    .B(net6574),
    .Y(_03431_));
 sg13g2_a21oi_1 _19084_ (.A1(net6574),
    .A2(net7413),
    .Y(_02133_),
    .B1(_03431_));
 sg13g2_nor2_1 _19085_ (.A(net3875),
    .B(net6574),
    .Y(_03432_));
 sg13g2_a21oi_1 _19086_ (.A1(net6574),
    .A2(net7573),
    .Y(_02134_),
    .B1(_03432_));
 sg13g2_nor2_1 _19087_ (.A(net4365),
    .B(net6576),
    .Y(_03433_));
 sg13g2_a21oi_1 _19088_ (.A1(net6577),
    .A2(net7124),
    .Y(_02135_),
    .B1(_03433_));
 sg13g2_nor2_1 _19089_ (.A(net3783),
    .B(net6576),
    .Y(_03434_));
 sg13g2_a21oi_1 _19090_ (.A1(net6576),
    .A2(net7419),
    .Y(_02136_),
    .B1(_03434_));
 sg13g2_nor2_1 _19091_ (.A(net4688),
    .B(net6577),
    .Y(_03435_));
 sg13g2_a21oi_1 _19092_ (.A1(net6577),
    .A2(net7578),
    .Y(_02137_),
    .B1(_03435_));
 sg13g2_nor2_1 _19093_ (.A(net4010),
    .B(net6674),
    .Y(_03436_));
 sg13g2_a21oi_1 _19094_ (.A1(net6674),
    .A2(net7149),
    .Y(_02138_),
    .B1(_03436_));
 sg13g2_nor2_1 _19095_ (.A(net4255),
    .B(net6674),
    .Y(_03437_));
 sg13g2_a21oi_1 _19096_ (.A1(net6674),
    .A2(net7444),
    .Y(_02139_),
    .B1(_03437_));
 sg13g2_nor2_1 _19097_ (.A(net4433),
    .B(net6674),
    .Y(_03438_));
 sg13g2_a21oi_1 _19098_ (.A1(net6674),
    .A2(net7601),
    .Y(_02140_),
    .B1(_03438_));
 sg13g2_nor2_1 _19099_ (.A(net4653),
    .B(net6678),
    .Y(_03439_));
 sg13g2_a21oi_1 _19100_ (.A1(net6678),
    .A2(net7124),
    .Y(_02141_),
    .B1(_03439_));
 sg13g2_nor2_1 _19101_ (.A(net4622),
    .B(net6679),
    .Y(_03440_));
 sg13g2_a21oi_1 _19102_ (.A1(net6679),
    .A2(net7419),
    .Y(_02142_),
    .B1(_03440_));
 sg13g2_nor2_1 _19103_ (.A(net4837),
    .B(net6679),
    .Y(_03441_));
 sg13g2_a21oi_1 _19104_ (.A1(net6679),
    .A2(net7578),
    .Y(_02143_),
    .B1(_03441_));
 sg13g2_nand2_1 _19105_ (.Y(_03442_),
    .A(net2919),
    .B(net6682));
 sg13g2_o21ai_1 _19106_ (.B1(_03442_),
    .Y(_02144_),
    .A1(net6682),
    .A2(net7124));
 sg13g2_nand2_1 _19107_ (.Y(_03443_),
    .A(net2572),
    .B(net6683));
 sg13g2_o21ai_1 _19108_ (.B1(_03443_),
    .Y(_02145_),
    .A1(net6683),
    .A2(net7419));
 sg13g2_nand2_1 _19109_ (.Y(_03444_),
    .A(net3075),
    .B(net6683));
 sg13g2_o21ai_1 _19110_ (.B1(_03444_),
    .Y(_02146_),
    .A1(net6683),
    .A2(net7578));
 sg13g2_nor2_1 _19111_ (.A(net4481),
    .B(net6684),
    .Y(_03445_));
 sg13g2_a21oi_1 _19112_ (.A1(net6684),
    .A2(net7124),
    .Y(_02147_),
    .B1(_03445_));
 sg13g2_nor2_1 _19113_ (.A(net4319),
    .B(net6684),
    .Y(_03446_));
 sg13g2_a21oi_1 _19114_ (.A1(net6684),
    .A2(net7413),
    .Y(_02148_),
    .B1(_03446_));
 sg13g2_nor2_1 _19115_ (.A(net4218),
    .B(net6684),
    .Y(_03447_));
 sg13g2_a21oi_1 _19116_ (.A1(net6684),
    .A2(net7574),
    .Y(_02149_),
    .B1(_03447_));
 sg13g2_nor2_1 _19117_ (.A(net4807),
    .B(net6686),
    .Y(_03448_));
 sg13g2_a21oi_1 _19118_ (.A1(net6686),
    .A2(net7124),
    .Y(_02150_),
    .B1(_03448_));
 sg13g2_nor2_1 _19119_ (.A(net4764),
    .B(net6686),
    .Y(_03449_));
 sg13g2_a21oi_1 _19120_ (.A1(net6686),
    .A2(net7418),
    .Y(_02151_),
    .B1(_03449_));
 sg13g2_nor2_1 _19121_ (.A(net4578),
    .B(net6686),
    .Y(_03450_));
 sg13g2_a21oi_1 _19122_ (.A1(net6686),
    .A2(net7577),
    .Y(_02152_),
    .B1(_03450_));
 sg13g2_nor2_1 _19123_ (.A(net4612),
    .B(net6688),
    .Y(_03451_));
 sg13g2_a21oi_1 _19124_ (.A1(net6688),
    .A2(net7124),
    .Y(_02153_),
    .B1(_03451_));
 sg13g2_nor2_1 _19125_ (.A(net4818),
    .B(net6688),
    .Y(_03452_));
 sg13g2_a21oi_1 _19126_ (.A1(net6688),
    .A2(net7418),
    .Y(_02154_),
    .B1(_03452_));
 sg13g2_nor2_1 _19127_ (.A(net4725),
    .B(net6688),
    .Y(_03453_));
 sg13g2_a21oi_1 _19128_ (.A1(net6688),
    .A2(net7577),
    .Y(_02155_),
    .B1(_03453_));
 sg13g2_nor2_1 _19129_ (.A(net4844),
    .B(net6690),
    .Y(_03454_));
 sg13g2_a21oi_1 _19130_ (.A1(net6690),
    .A2(net7124),
    .Y(_02156_),
    .B1(_03454_));
 sg13g2_nor2_1 _19131_ (.A(net3952),
    .B(net6690),
    .Y(_03455_));
 sg13g2_a21oi_1 _19132_ (.A1(net6690),
    .A2(net7418),
    .Y(_02157_),
    .B1(_03455_));
 sg13g2_nor2_1 _19133_ (.A(net4769),
    .B(net6690),
    .Y(_03456_));
 sg13g2_a21oi_1 _19134_ (.A1(net6690),
    .A2(net7577),
    .Y(_02158_),
    .B1(_03456_));
 sg13g2_nor2_1 _19135_ (.A(net4832),
    .B(net6692),
    .Y(_03457_));
 sg13g2_a21oi_1 _19136_ (.A1(net6692),
    .A2(net7118),
    .Y(_02159_),
    .B1(_03457_));
 sg13g2_nor2_1 _19137_ (.A(net4680),
    .B(net6692),
    .Y(_03458_));
 sg13g2_a21oi_1 _19138_ (.A1(net6692),
    .A2(net7414),
    .Y(_02160_),
    .B1(_03458_));
 sg13g2_nor2_1 _19139_ (.A(net4656),
    .B(net6692),
    .Y(_03459_));
 sg13g2_a21oi_1 _19140_ (.A1(net6692),
    .A2(net7573),
    .Y(_02161_),
    .B1(_03459_));
 sg13g2_nor2_1 _19141_ (.A(net4672),
    .B(net6694),
    .Y(_03460_));
 sg13g2_a21oi_1 _19142_ (.A1(net6694),
    .A2(net7118),
    .Y(_02162_),
    .B1(_03460_));
 sg13g2_nor2_1 _19143_ (.A(net4106),
    .B(net6694),
    .Y(_03461_));
 sg13g2_a21oi_1 _19144_ (.A1(net6694),
    .A2(net7414),
    .Y(_02163_),
    .B1(_03461_));
 sg13g2_nor2_1 _19145_ (.A(net4779),
    .B(net6694),
    .Y(_03462_));
 sg13g2_a21oi_1 _19146_ (.A1(net6694),
    .A2(net7573),
    .Y(_02164_),
    .B1(_03462_));
 sg13g2_nor2_1 _19147_ (.A(net4810),
    .B(net6696),
    .Y(_03463_));
 sg13g2_a21oi_1 _19148_ (.A1(net6696),
    .A2(net7118),
    .Y(_02165_),
    .B1(_03463_));
 sg13g2_nor2_1 _19149_ (.A(net3760),
    .B(net6696),
    .Y(_03464_));
 sg13g2_a21oi_1 _19150_ (.A1(net6696),
    .A2(net7414),
    .Y(_02166_),
    .B1(_03464_));
 sg13g2_nor2_1 _19151_ (.A(net4266),
    .B(net6696),
    .Y(_03465_));
 sg13g2_a21oi_1 _19152_ (.A1(net6696),
    .A2(net7573),
    .Y(_02167_),
    .B1(_03465_));
 sg13g2_nand2_1 _19153_ (.Y(_03466_),
    .A(net3220),
    .B(net7044));
 sg13g2_o21ai_1 _19154_ (.B1(_03466_),
    .Y(_02168_),
    .A1(net7044),
    .A2(net7149));
 sg13g2_nand2_1 _19155_ (.Y(_03467_),
    .A(net4228),
    .B(net7045));
 sg13g2_o21ai_1 _19156_ (.B1(_03467_),
    .Y(_02169_),
    .A1(net7045),
    .A2(net7444));
 sg13g2_nand2_1 _19157_ (.Y(_03468_),
    .A(net3191),
    .B(net7044));
 sg13g2_o21ai_1 _19158_ (.B1(_03468_),
    .Y(_02170_),
    .A1(net7044),
    .A2(net7603));
 sg13g2_nor2_1 _19159_ (.A(net4525),
    .B(net6699),
    .Y(_03469_));
 sg13g2_a21oi_1 _19160_ (.A1(net6699),
    .A2(net7123),
    .Y(_02171_),
    .B1(_03469_));
 sg13g2_nor2_1 _19161_ (.A(net3710),
    .B(net6698),
    .Y(_03470_));
 sg13g2_a21oi_1 _19162_ (.A1(net6698),
    .A2(net7418),
    .Y(_02172_),
    .B1(_03470_));
 sg13g2_nor2_1 _19163_ (.A(net4791),
    .B(net6698),
    .Y(_03471_));
 sg13g2_a21oi_1 _19164_ (.A1(net6698),
    .A2(net7577),
    .Y(_02173_),
    .B1(_03471_));
 sg13g2_nor2_1 _19165_ (.A(net4529),
    .B(net6729),
    .Y(_03472_));
 sg13g2_a21oi_1 _19166_ (.A1(net6729),
    .A2(net7123),
    .Y(_02174_),
    .B1(_03472_));
 sg13g2_nor2_1 _19167_ (.A(net4173),
    .B(net6728),
    .Y(_03473_));
 sg13g2_a21oi_1 _19168_ (.A1(net6728),
    .A2(net7418),
    .Y(_02175_),
    .B1(_03473_));
 sg13g2_nor2_1 _19169_ (.A(net3879),
    .B(net6728),
    .Y(_03474_));
 sg13g2_a21oi_1 _19170_ (.A1(net6728),
    .A2(net7577),
    .Y(_02176_),
    .B1(_03474_));
 sg13g2_nor2_1 _19171_ (.A(net4727),
    .B(net6731),
    .Y(_03475_));
 sg13g2_a21oi_1 _19172_ (.A1(net6731),
    .A2(net7123),
    .Y(_02177_),
    .B1(_03475_));
 sg13g2_nor2_1 _19173_ (.A(net4846),
    .B(net6730),
    .Y(_03476_));
 sg13g2_a21oi_1 _19174_ (.A1(net6730),
    .A2(net7418),
    .Y(_02178_),
    .B1(_03476_));
 sg13g2_nor2_1 _19175_ (.A(net4704),
    .B(net6730),
    .Y(_03477_));
 sg13g2_a21oi_1 _19176_ (.A1(net6730),
    .A2(net7577),
    .Y(_02179_),
    .B1(_03477_));
 sg13g2_nor2_1 _19177_ (.A(net4454),
    .B(net6507),
    .Y(_03478_));
 sg13g2_a21oi_1 _19178_ (.A1(net6507),
    .A2(net7123),
    .Y(_02180_),
    .B1(_03478_));
 sg13g2_nor2_1 _19179_ (.A(net4020),
    .B(net6506),
    .Y(_03479_));
 sg13g2_a21oi_1 _19180_ (.A1(net6506),
    .A2(net7417),
    .Y(_02181_),
    .B1(_03479_));
 sg13g2_nor2_1 _19181_ (.A(net4401),
    .B(net6506),
    .Y(_03480_));
 sg13g2_a21oi_1 _19182_ (.A1(net6506),
    .A2(net7577),
    .Y(_02182_),
    .B1(_03480_));
 sg13g2_nor2_1 _19183_ (.A(net4788),
    .B(net6508),
    .Y(_03481_));
 sg13g2_a21oi_1 _19184_ (.A1(net6509),
    .A2(net7126),
    .Y(_02183_),
    .B1(_03481_));
 sg13g2_nor2_1 _19185_ (.A(net4528),
    .B(net6508),
    .Y(_03482_));
 sg13g2_a21oi_1 _19186_ (.A1(net6508),
    .A2(net7421),
    .Y(_02184_),
    .B1(_03482_));
 sg13g2_nor2_1 _19187_ (.A(net3795),
    .B(net6508),
    .Y(_03483_));
 sg13g2_a21oi_1 _19188_ (.A1(net6508),
    .A2(net7579),
    .Y(_02185_),
    .B1(_03483_));
 sg13g2_nand2_1 _19189_ (.Y(_03484_),
    .A(net3888),
    .B(net6540));
 sg13g2_o21ai_1 _19190_ (.B1(_03484_),
    .Y(_02186_),
    .A1(net6541),
    .A2(net7125));
 sg13g2_nand2_1 _19191_ (.Y(_03485_),
    .A(net3429),
    .B(net6540));
 sg13g2_o21ai_1 _19192_ (.B1(_03485_),
    .Y(_02187_),
    .A1(net6540),
    .A2(net7420));
 sg13g2_nand2_1 _19193_ (.Y(_03486_),
    .A(net2675),
    .B(net6540));
 sg13g2_o21ai_1 _19194_ (.B1(_03486_),
    .Y(_02188_),
    .A1(net6540),
    .A2(net7579));
 sg13g2_nand2_1 _19195_ (.Y(_03487_),
    .A(net3339),
    .B(net6544));
 sg13g2_o21ai_1 _19196_ (.B1(_03487_),
    .Y(_02189_),
    .A1(net6545),
    .A2(net7125));
 sg13g2_nand2_1 _19197_ (.Y(_03488_),
    .A(net2894),
    .B(net6544));
 sg13g2_o21ai_1 _19198_ (.B1(_03488_),
    .Y(_02190_),
    .A1(net6544),
    .A2(net7420));
 sg13g2_nand2_1 _19199_ (.Y(_03489_),
    .A(net3150),
    .B(net6544));
 sg13g2_o21ai_1 _19200_ (.B1(_03489_),
    .Y(_02191_),
    .A1(net6544),
    .A2(net7579));
 sg13g2_nand2_1 _19201_ (.Y(_03490_),
    .A(net2752),
    .B(net6546));
 sg13g2_o21ai_1 _19202_ (.B1(_03490_),
    .Y(_02192_),
    .A1(net6547),
    .A2(net7125));
 sg13g2_nand2_1 _19203_ (.Y(_03491_),
    .A(net2578),
    .B(net6546));
 sg13g2_o21ai_1 _19204_ (.B1(_03491_),
    .Y(_02193_),
    .A1(net6546),
    .A2(net7420));
 sg13g2_nand2_1 _19205_ (.Y(_03492_),
    .A(net2712),
    .B(net6546));
 sg13g2_o21ai_1 _19206_ (.B1(_03492_),
    .Y(_02194_),
    .A1(net6546),
    .A2(net7579));
 sg13g2_nor2_1 _19207_ (.A(net4639),
    .B(net6549),
    .Y(_03493_));
 sg13g2_a21oi_1 _19208_ (.A1(net6548),
    .A2(net7126),
    .Y(_02195_),
    .B1(_03493_));
 sg13g2_nor2_1 _19209_ (.A(net4487),
    .B(net6548),
    .Y(_03494_));
 sg13g2_a21oi_1 _19210_ (.A1(net6548),
    .A2(net7417),
    .Y(_02196_),
    .B1(_03494_));
 sg13g2_nor2_1 _19211_ (.A(net4229),
    .B(net6548),
    .Y(_03495_));
 sg13g2_a21oi_1 _19212_ (.A1(net6548),
    .A2(net7579),
    .Y(_02197_),
    .B1(_03495_));
 sg13g2_nor2_1 _19213_ (.A(net4177),
    .B(net6943),
    .Y(_03496_));
 sg13g2_a21oi_1 _19214_ (.A1(net6943),
    .A2(net7149),
    .Y(_02198_),
    .B1(_03496_));
 sg13g2_nor2_1 _19215_ (.A(net4336),
    .B(net6942),
    .Y(_03497_));
 sg13g2_a21oi_1 _19216_ (.A1(net6942),
    .A2(net7445),
    .Y(_02199_),
    .B1(_03497_));
 sg13g2_nor2_1 _19217_ (.A(net3935),
    .B(net6942),
    .Y(_03498_));
 sg13g2_a21oi_1 _19218_ (.A1(net6942),
    .A2(net7599),
    .Y(_02200_),
    .B1(_03498_));
 sg13g2_nand2_1 _19219_ (.Y(_03499_),
    .A(net2642),
    .B(net6556));
 sg13g2_o21ai_1 _19220_ (.B1(_03499_),
    .Y(_02201_),
    .A1(net6556),
    .A2(net7126));
 sg13g2_nand2_1 _19221_ (.Y(_03500_),
    .A(net3505),
    .B(net6556));
 sg13g2_o21ai_1 _19222_ (.B1(_03500_),
    .Y(_02202_),
    .A1(net6556),
    .A2(net7417));
 sg13g2_nand2_1 _19223_ (.Y(_03501_),
    .A(net4071),
    .B(net6556));
 sg13g2_o21ai_1 _19224_ (.B1(_03501_),
    .Y(_02203_),
    .A1(net6556),
    .A2(net7579));
 sg13g2_nand2_1 _19225_ (.Y(_03502_),
    .A(net2725),
    .B(net6561));
 sg13g2_o21ai_1 _19226_ (.B1(_03502_),
    .Y(_02204_),
    .A1(net6561),
    .A2(net7125));
 sg13g2_nand2_1 _19227_ (.Y(_03503_),
    .A(net3509),
    .B(net6560));
 sg13g2_o21ai_1 _19228_ (.B1(_03503_),
    .Y(_02205_),
    .A1(net6560),
    .A2(net7417));
 sg13g2_nand2_1 _19229_ (.Y(_03504_),
    .A(net2949),
    .B(net6560));
 sg13g2_o21ai_1 _19230_ (.B1(_03504_),
    .Y(_02206_),
    .A1(net6560),
    .A2(net7579));
 sg13g2_nand2_1 _19231_ (.Y(_03505_),
    .A(net3678),
    .B(net6562));
 sg13g2_o21ai_1 _19232_ (.B1(_03505_),
    .Y(_02207_),
    .A1(net6562),
    .A2(net7123));
 sg13g2_nand2_1 _19233_ (.Y(_03506_),
    .A(net3151),
    .B(net6563));
 sg13g2_o21ai_1 _19234_ (.B1(_03506_),
    .Y(_02208_),
    .A1(net6563),
    .A2(net7417));
 sg13g2_nand2_1 _19235_ (.Y(_03507_),
    .A(net3022),
    .B(net6563));
 sg13g2_o21ai_1 _19236_ (.B1(_03507_),
    .Y(_02209_),
    .A1(net6563),
    .A2(net7580));
 sg13g2_nand2_1 _19237_ (.Y(_03508_),
    .A(net4461),
    .B(net6566));
 sg13g2_o21ai_1 _19238_ (.B1(_03508_),
    .Y(_02210_),
    .A1(net6566),
    .A2(net7123));
 sg13g2_nand2_1 _19239_ (.Y(_03509_),
    .A(net3393),
    .B(net6567));
 sg13g2_o21ai_1 _19240_ (.B1(_03509_),
    .Y(_02211_),
    .A1(net6567),
    .A2(net7417));
 sg13g2_nand2_1 _19241_ (.Y(_03510_),
    .A(net2443),
    .B(net6567));
 sg13g2_o21ai_1 _19242_ (.B1(_03510_),
    .Y(_02212_),
    .A1(net6567),
    .A2(net7580));
 sg13g2_nand2_1 _19243_ (.Y(_03511_),
    .A(net3668),
    .B(net6572));
 sg13g2_o21ai_1 _19244_ (.B1(_03511_),
    .Y(_02213_),
    .A1(net6572),
    .A2(net7123));
 sg13g2_nand2_1 _19245_ (.Y(_03512_),
    .A(net3597),
    .B(net6572));
 sg13g2_o21ai_1 _19246_ (.B1(_03512_),
    .Y(_02214_),
    .A1(net6572),
    .A2(net7418));
 sg13g2_nand2_1 _19247_ (.Y(_03513_),
    .A(net3419),
    .B(net6572));
 sg13g2_o21ai_1 _19248_ (.B1(_03513_),
    .Y(_02215_),
    .A1(net6572),
    .A2(net7580));
 sg13g2_nand2_1 _19249_ (.Y(_03514_),
    .A(net3330),
    .B(net6676));
 sg13g2_o21ai_1 _19250_ (.B1(_03514_),
    .Y(_02216_),
    .A1(net6676),
    .A2(net7123));
 sg13g2_nand2_1 _19251_ (.Y(_03515_),
    .A(net2482),
    .B(net6677));
 sg13g2_o21ai_1 _19252_ (.B1(_03515_),
    .Y(_02217_),
    .A1(net6677),
    .A2(net7417));
 sg13g2_nand2_1 _19253_ (.Y(_03516_),
    .A(net2968),
    .B(net6677));
 sg13g2_o21ai_1 _19254_ (.B1(_03516_),
    .Y(_02218_),
    .A1(net6677),
    .A2(net7577));
 sg13g2_nor2_1 _19255_ (.A(net4468),
    .B(net6681),
    .Y(_03517_));
 sg13g2_a21oi_1 _19256_ (.A1(net6680),
    .A2(net7157),
    .Y(_02219_),
    .B1(_03517_));
 sg13g2_nor2_1 _19257_ (.A(net3814),
    .B(net6681),
    .Y(_03518_));
 sg13g2_a21oi_1 _19258_ (.A1(net6681),
    .A2(net7454),
    .Y(_02220_),
    .B1(_03518_));
 sg13g2_nor2_1 _19259_ (.A(net4804),
    .B(net6680),
    .Y(_03519_));
 sg13g2_a21oi_1 _19260_ (.A1(net6680),
    .A2(net7612),
    .Y(_02221_),
    .B1(_03519_));
 sg13g2_nor2_1 _19261_ (.A(net4352),
    .B(net6733),
    .Y(_03520_));
 sg13g2_a21oi_1 _19262_ (.A1(net6732),
    .A2(net7157),
    .Y(_02222_),
    .B1(_03520_));
 sg13g2_nor2_1 _19263_ (.A(net4344),
    .B(net6733),
    .Y(_03521_));
 sg13g2_a21oi_1 _19264_ (.A1(net6733),
    .A2(net7454),
    .Y(_02223_),
    .B1(_03521_));
 sg13g2_nor2_1 _19265_ (.A(net4532),
    .B(net6732),
    .Y(_03522_));
 sg13g2_a21oi_1 _19266_ (.A1(net6732),
    .A2(net7612),
    .Y(_02224_),
    .B1(_03522_));
 sg13g2_nor2_1 _19267_ (.A(net4801),
    .B(net6579),
    .Y(_03523_));
 sg13g2_a21oi_1 _19268_ (.A1(net6578),
    .A2(net7157),
    .Y(_02225_),
    .B1(_03523_));
 sg13g2_nor2_1 _19269_ (.A(net4828),
    .B(net6579),
    .Y(_03524_));
 sg13g2_a21oi_1 _19270_ (.A1(net6579),
    .A2(net7454),
    .Y(_02226_),
    .B1(_03524_));
 sg13g2_nor2_1 _19271_ (.A(net4752),
    .B(net6578),
    .Y(_03525_));
 sg13g2_a21oi_1 _19272_ (.A1(net6578),
    .A2(net7612),
    .Y(_02227_),
    .B1(_03525_));
 sg13g2_nor2_1 _19273_ (.A(net4034),
    .B(net6954),
    .Y(_03526_));
 sg13g2_a21oi_1 _19274_ (.A1(net6954),
    .A2(net7150),
    .Y(_02228_),
    .B1(_03526_));
 sg13g2_nor2_1 _19275_ (.A(net4726),
    .B(net6955),
    .Y(_03527_));
 sg13g2_a21oi_1 _19276_ (.A1(net6955),
    .A2(net7445),
    .Y(_02229_),
    .B1(_03527_));
 sg13g2_nor2_1 _19277_ (.A(net4168),
    .B(net6954),
    .Y(_03528_));
 sg13g2_a21oi_1 _19278_ (.A1(net6954),
    .A2(net7603),
    .Y(_02230_),
    .B1(_03528_));
 sg13g2_nor2_1 _19279_ (.A(net4376),
    .B(net6580),
    .Y(_03529_));
 sg13g2_a21oi_1 _19280_ (.A1(net6580),
    .A2(net7158),
    .Y(_02231_),
    .B1(_03529_));
 sg13g2_nor2_1 _19281_ (.A(net4165),
    .B(net6580),
    .Y(_03530_));
 sg13g2_a21oi_1 _19282_ (.A1(net6580),
    .A2(net7455),
    .Y(_02232_),
    .B1(_03530_));
 sg13g2_nor2_1 _19283_ (.A(net4780),
    .B(net6580),
    .Y(_03531_));
 sg13g2_a21oi_1 _19284_ (.A1(net6580),
    .A2(net7612),
    .Y(_02233_),
    .B1(_03531_));
 sg13g2_nand2_1 _19285_ (.Y(_03532_),
    .A(net4379),
    .B(net6583));
 sg13g2_o21ai_1 _19286_ (.B1(_03532_),
    .Y(_02234_),
    .A1(net6583),
    .A2(net7158));
 sg13g2_nand2_1 _19287_ (.Y(_03533_),
    .A(net3676),
    .B(net6582));
 sg13g2_o21ai_1 _19288_ (.B1(_03533_),
    .Y(_02235_),
    .A1(net6583),
    .A2(net7455));
 sg13g2_nand2_1 _19289_ (.Y(_03534_),
    .A(net2851),
    .B(net6583));
 sg13g2_o21ai_1 _19290_ (.B1(_03534_),
    .Y(_02236_),
    .A1(net6582),
    .A2(net7612));
 sg13g2_nand2_1 _19291_ (.Y(_03535_),
    .A(net2664),
    .B(net6585));
 sg13g2_o21ai_1 _19292_ (.B1(_03535_),
    .Y(_02237_),
    .A1(net6585),
    .A2(net7158));
 sg13g2_nand2_1 _19293_ (.Y(_03536_),
    .A(net3911),
    .B(net6585));
 sg13g2_o21ai_1 _19294_ (.B1(_03536_),
    .Y(_02238_),
    .A1(net6585),
    .A2(net7455));
 sg13g2_nand2_1 _19295_ (.Y(_03537_),
    .A(net3929),
    .B(net6584));
 sg13g2_o21ai_1 _19296_ (.B1(_03537_),
    .Y(_02239_),
    .A1(net6584),
    .A2(net7612));
 sg13g2_nand2_1 _19297_ (.Y(_03538_),
    .A(net3066),
    .B(net6587));
 sg13g2_o21ai_1 _19298_ (.B1(_03538_),
    .Y(_02240_),
    .A1(net6587),
    .A2(net7158));
 sg13g2_nand2_1 _19299_ (.Y(_03539_),
    .A(net4062),
    .B(net6586));
 sg13g2_o21ai_1 _19300_ (.B1(_03539_),
    .Y(_02241_),
    .A1(net6586),
    .A2(net7455));
 sg13g2_nand2_1 _19301_ (.Y(_03540_),
    .A(net3314),
    .B(net6587));
 sg13g2_o21ai_1 _19302_ (.B1(_03540_),
    .Y(_02242_),
    .A1(net6586),
    .A2(net7612));
 sg13g2_nor2_1 _19303_ (.A(net4464),
    .B(net6590),
    .Y(_03541_));
 sg13g2_a21oi_1 _19304_ (.A1(net6590),
    .A2(net7171),
    .Y(_02243_),
    .B1(_03541_));
 sg13g2_nor2_1 _19305_ (.A(net4428),
    .B(net6591),
    .Y(_03542_));
 sg13g2_a21oi_1 _19306_ (.A1(net6591),
    .A2(net7467),
    .Y(_02244_),
    .B1(_03542_));
 sg13g2_nor2_1 _19307_ (.A(net4843),
    .B(net6590),
    .Y(_03543_));
 sg13g2_a21oi_1 _19308_ (.A1(net6590),
    .A2(net7626),
    .Y(_02245_),
    .B1(_03543_));
 sg13g2_nand2_1 _19309_ (.Y(_03544_),
    .A(net4603),
    .B(net6592));
 sg13g2_o21ai_1 _19310_ (.B1(_03544_),
    .Y(_02246_),
    .A1(net6592),
    .A2(net7171));
 sg13g2_nand2_1 _19311_ (.Y(_03545_),
    .A(net3549),
    .B(net6593));
 sg13g2_o21ai_1 _19312_ (.B1(_03545_),
    .Y(_02247_),
    .A1(net6593),
    .A2(net7467));
 sg13g2_nand2_1 _19313_ (.Y(_03546_),
    .A(net3970),
    .B(net6592));
 sg13g2_o21ai_1 _19314_ (.B1(_03546_),
    .Y(_02248_),
    .A1(net6592),
    .A2(net7626));
 sg13g2_nand2_1 _19315_ (.Y(_03547_),
    .A(net3464),
    .B(net6596));
 sg13g2_o21ai_1 _19316_ (.B1(_03547_),
    .Y(_02249_),
    .A1(net6596),
    .A2(net7171));
 sg13g2_nand2_1 _19317_ (.Y(_03548_),
    .A(net4009),
    .B(net6596));
 sg13g2_o21ai_1 _19318_ (.B1(_03548_),
    .Y(_02250_),
    .A1(net6597),
    .A2(net7467));
 sg13g2_nand2_1 _19319_ (.Y(_03549_),
    .A(net3380),
    .B(net6596));
 sg13g2_o21ai_1 _19320_ (.B1(_03549_),
    .Y(_02251_),
    .A1(net6596),
    .A2(net7626));
 sg13g2_nand2_1 _19321_ (.Y(_03550_),
    .A(net3650),
    .B(net6598));
 sg13g2_o21ai_1 _19322_ (.B1(_03550_),
    .Y(_02252_),
    .A1(net6598),
    .A2(net7171));
 sg13g2_nand2_1 _19323_ (.Y(_03551_),
    .A(net3596),
    .B(net6599));
 sg13g2_o21ai_1 _19324_ (.B1(_03551_),
    .Y(_02253_),
    .A1(net6599),
    .A2(net7467));
 sg13g2_nand2_1 _19325_ (.Y(_03552_),
    .A(net3096),
    .B(net6598));
 sg13g2_o21ai_1 _19326_ (.B1(_03552_),
    .Y(_02254_),
    .A1(net6598),
    .A2(net7626));
 sg13g2_nand2_1 _19327_ (.Y(_03553_),
    .A(net2878),
    .B(net6602));
 sg13g2_o21ai_1 _19328_ (.B1(_03553_),
    .Y(_02255_),
    .A1(net6602),
    .A2(net7171));
 sg13g2_nand2_1 _19329_ (.Y(_03554_),
    .A(net3152),
    .B(net6603));
 sg13g2_o21ai_1 _19330_ (.B1(_03554_),
    .Y(_02256_),
    .A1(net6603),
    .A2(net7467));
 sg13g2_nand2_1 _19331_ (.Y(_03555_),
    .A(net2842),
    .B(net6602));
 sg13g2_o21ai_1 _19332_ (.B1(_03555_),
    .Y(_02257_),
    .A1(net6602),
    .A2(net7612));
 sg13g2_nor2_1 _19333_ (.A(net4230),
    .B(net6959),
    .Y(_03556_));
 sg13g2_a21oi_1 _19334_ (.A1(net6959),
    .A2(net7149),
    .Y(_02258_),
    .B1(_03556_));
 sg13g2_nor2_1 _19335_ (.A(net4711),
    .B(net6959),
    .Y(_03557_));
 sg13g2_a21oi_1 _19336_ (.A1(net6959),
    .A2(net7445),
    .Y(_02259_),
    .B1(_03557_));
 sg13g2_nor2_1 _19337_ (.A(net3981),
    .B(net6958),
    .Y(_03558_));
 sg13g2_a21oi_1 _19338_ (.A1(net6958),
    .A2(net7603),
    .Y(_02260_),
    .B1(_03558_));
 sg13g2_nand2_1 _19339_ (.Y(_03559_),
    .A(net3829),
    .B(net6606));
 sg13g2_o21ai_1 _19340_ (.B1(_03559_),
    .Y(_02261_),
    .A1(net6606),
    .A2(net7171));
 sg13g2_nand2_1 _19341_ (.Y(_03560_),
    .A(net4248),
    .B(net6607));
 sg13g2_o21ai_1 _19342_ (.B1(_03560_),
    .Y(_02262_),
    .A1(net6607),
    .A2(net7467));
 sg13g2_nand2_1 _19343_ (.Y(_03561_),
    .A(net3323),
    .B(net6606));
 sg13g2_o21ai_1 _19344_ (.B1(_03561_),
    .Y(_02263_),
    .A1(net6606),
    .A2(net7626));
 sg13g2_nand2_1 _19345_ (.Y(_03562_),
    .A(net3598),
    .B(net6608));
 sg13g2_o21ai_1 _19346_ (.B1(_03562_),
    .Y(_02264_),
    .A1(net6608),
    .A2(net7171));
 sg13g2_nand2_1 _19347_ (.Y(_03563_),
    .A(net3048),
    .B(net6609));
 sg13g2_o21ai_1 _19348_ (.B1(_03563_),
    .Y(_02265_),
    .A1(net6609),
    .A2(net7467));
 sg13g2_nand2_1 _19349_ (.Y(_03564_),
    .A(net2694),
    .B(net6608));
 sg13g2_o21ai_1 _19350_ (.B1(_03564_),
    .Y(_02266_),
    .A1(net6608),
    .A2(net7626));
 sg13g2_nand2_1 _19351_ (.Y(_03565_),
    .A(net2917),
    .B(net6612));
 sg13g2_o21ai_1 _19352_ (.B1(_03565_),
    .Y(_02267_),
    .A1(net6612),
    .A2(net7178));
 sg13g2_nand2_1 _19353_ (.Y(_03566_),
    .A(net3319),
    .B(net6613));
 sg13g2_o21ai_1 _19354_ (.B1(_03566_),
    .Y(_02268_),
    .A1(net6613),
    .A2(net7473));
 sg13g2_nand2_1 _19355_ (.Y(_03567_),
    .A(net3287),
    .B(net6612));
 sg13g2_o21ai_1 _19356_ (.B1(_03567_),
    .Y(_02269_),
    .A1(net6612),
    .A2(net7633));
 sg13g2_nand2_1 _19357_ (.Y(_03568_),
    .A(net3306),
    .B(net6614));
 sg13g2_o21ai_1 _19358_ (.B1(_03568_),
    .Y(_02270_),
    .A1(net6614),
    .A2(net7178));
 sg13g2_nand2_1 _19359_ (.Y(_03569_),
    .A(net2728),
    .B(net6615));
 sg13g2_o21ai_1 _19360_ (.B1(_03569_),
    .Y(_02271_),
    .A1(net6615),
    .A2(net7473));
 sg13g2_nand2_1 _19361_ (.Y(_03570_),
    .A(net3208),
    .B(net6614));
 sg13g2_o21ai_1 _19362_ (.B1(_03570_),
    .Y(_02272_),
    .A1(net6614),
    .A2(net7633));
 sg13g2_nand2_1 _19363_ (.Y(_03571_),
    .A(net3283),
    .B(net6616));
 sg13g2_o21ai_1 _19364_ (.B1(_03571_),
    .Y(_02273_),
    .A1(net6616),
    .A2(net7179));
 sg13g2_nand2_1 _19365_ (.Y(_03572_),
    .A(net3978),
    .B(net6617));
 sg13g2_o21ai_1 _19366_ (.B1(_03572_),
    .Y(_02274_),
    .A1(net6617),
    .A2(net7473));
 sg13g2_nand2_1 _19367_ (.Y(_03573_),
    .A(net3213),
    .B(net6616));
 sg13g2_o21ai_1 _19368_ (.B1(_03573_),
    .Y(_02275_),
    .A1(net6616),
    .A2(net7633));
 sg13g2_nand2_1 _19369_ (.Y(_03574_),
    .A(net3663),
    .B(net6618));
 sg13g2_o21ai_1 _19370_ (.B1(_03574_),
    .Y(_02276_),
    .A1(net6618),
    .A2(net7179));
 sg13g2_nand2_1 _19371_ (.Y(_03575_),
    .A(net3998),
    .B(net6619));
 sg13g2_o21ai_1 _19372_ (.B1(_03575_),
    .Y(_02277_),
    .A1(net6619),
    .A2(net7473));
 sg13g2_nand2_1 _19373_ (.Y(_03576_),
    .A(net3519),
    .B(net6618));
 sg13g2_o21ai_1 _19374_ (.B1(_03576_),
    .Y(_02278_),
    .A1(net6618),
    .A2(net7633));
 sg13g2_nand2_1 _19375_ (.Y(_03577_),
    .A(net2505),
    .B(net6620));
 sg13g2_o21ai_1 _19376_ (.B1(_03577_),
    .Y(_02279_),
    .A1(net6621),
    .A2(net7175));
 sg13g2_nand2_1 _19377_ (.Y(_03578_),
    .A(net3224),
    .B(net6620));
 sg13g2_o21ai_1 _19378_ (.B1(_03578_),
    .Y(_02280_),
    .A1(net6621),
    .A2(net7471));
 sg13g2_nand2_1 _19379_ (.Y(_03579_),
    .A(net3388),
    .B(net6620));
 sg13g2_o21ai_1 _19380_ (.B1(_03579_),
    .Y(_02281_),
    .A1(net6620),
    .A2(net7627));
 sg13g2_nand2_1 _19381_ (.Y(_03580_),
    .A(net3773),
    .B(net6664));
 sg13g2_o21ai_1 _19382_ (.B1(_03580_),
    .Y(_02282_),
    .A1(net6664),
    .A2(net7175));
 sg13g2_nand2_1 _19383_ (.Y(_03581_),
    .A(net2907),
    .B(net6665));
 sg13g2_o21ai_1 _19384_ (.B1(_03581_),
    .Y(_02283_),
    .A1(net6665),
    .A2(net7471));
 sg13g2_nand2_1 _19385_ (.Y(_03582_),
    .A(net2681),
    .B(net6664));
 sg13g2_o21ai_1 _19386_ (.B1(_03582_),
    .Y(_02284_),
    .A1(net6664),
    .A2(net7627));
 sg13g2_nand2_1 _19387_ (.Y(_03583_),
    .A(net3994),
    .B(net6666));
 sg13g2_o21ai_1 _19388_ (.B1(_03583_),
    .Y(_02285_),
    .A1(net6666),
    .A2(net7175));
 sg13g2_nand2_1 _19389_ (.Y(_03584_),
    .A(net4418),
    .B(net6667));
 sg13g2_o21ai_1 _19390_ (.B1(_03584_),
    .Y(_02286_),
    .A1(net6667),
    .A2(net7471));
 sg13g2_nand2_1 _19391_ (.Y(_03585_),
    .A(net3098),
    .B(net6666));
 sg13g2_o21ai_1 _19392_ (.B1(_03585_),
    .Y(_02287_),
    .A1(net6666),
    .A2(net7626));
 sg13g2_nand2_1 _19393_ (.Y(_03586_),
    .A(net2631),
    .B(net6669));
 sg13g2_o21ai_1 _19394_ (.B1(_03586_),
    .Y(_02288_),
    .A1(net6669),
    .A2(net7149));
 sg13g2_nand2_1 _19395_ (.Y(_03587_),
    .A(net3212),
    .B(net6668));
 sg13g2_o21ai_1 _19396_ (.B1(_03587_),
    .Y(_02289_),
    .A1(net6668),
    .A2(net7445));
 sg13g2_nand2_1 _19397_ (.Y(_03588_),
    .A(net2462),
    .B(net6668));
 sg13g2_o21ai_1 _19398_ (.B1(_03588_),
    .Y(_02290_),
    .A1(net6668),
    .A2(net7603));
 sg13g2_nand2_1 _19399_ (.Y(_03589_),
    .A(net2580),
    .B(net6670));
 sg13g2_o21ai_1 _19400_ (.B1(_03589_),
    .Y(_02291_),
    .A1(net6670),
    .A2(net7173));
 sg13g2_nand2_1 _19401_ (.Y(_03590_),
    .A(net3028),
    .B(net6670));
 sg13g2_o21ai_1 _19402_ (.B1(_03590_),
    .Y(_02292_),
    .A1(net6670),
    .A2(net7469));
 sg13g2_nand2_1 _19403_ (.Y(_03591_),
    .A(net3010),
    .B(net6671));
 sg13g2_o21ai_1 _19404_ (.B1(_03591_),
    .Y(_02293_),
    .A1(net6671),
    .A2(net7629));
 sg13g2_nand2_1 _19405_ (.Y(_03592_),
    .A(net3886),
    .B(net6672));
 sg13g2_o21ai_1 _19406_ (.B1(_03592_),
    .Y(_02294_),
    .A1(net6672),
    .A2(net7173));
 sg13g2_nand2_1 _19407_ (.Y(_03593_),
    .A(net3781),
    .B(net6672));
 sg13g2_o21ai_1 _19408_ (.B1(_03593_),
    .Y(_02295_),
    .A1(net6672),
    .A2(net7469));
 sg13g2_nand2_1 _19409_ (.Y(_03594_),
    .A(net3285),
    .B(net6673));
 sg13g2_o21ai_1 _19410_ (.B1(_03594_),
    .Y(_02296_),
    .A1(net6673),
    .A2(net7629));
 sg13g2_nand2_1 _19411_ (.Y(_03595_),
    .A(net4247),
    .B(net6734));
 sg13g2_o21ai_1 _19412_ (.B1(_03595_),
    .Y(_02297_),
    .A1(net6734),
    .A2(net7173));
 sg13g2_nand2_1 _19413_ (.Y(_03596_),
    .A(net3165),
    .B(net6734));
 sg13g2_o21ai_1 _19414_ (.B1(_03596_),
    .Y(_02298_),
    .A1(net6734),
    .A2(net7470));
 sg13g2_nand2_1 _19415_ (.Y(_03597_),
    .A(net3739),
    .B(net6735));
 sg13g2_o21ai_1 _19416_ (.B1(_03597_),
    .Y(_02299_),
    .A1(net6735),
    .A2(net7629));
 sg13g2_nand2_1 _19417_ (.Y(_03598_),
    .A(net4007),
    .B(net6588));
 sg13g2_o21ai_1 _19418_ (.B1(_03598_),
    .Y(_02300_),
    .A1(net6588),
    .A2(net7173));
 sg13g2_nand2_1 _19419_ (.Y(_03599_),
    .A(net3824),
    .B(net6588));
 sg13g2_o21ai_1 _19420_ (.B1(_03599_),
    .Y(_02301_),
    .A1(net6588),
    .A2(net7469));
 sg13g2_nand2_1 _19421_ (.Y(_03600_),
    .A(net4579),
    .B(net6589));
 sg13g2_o21ai_1 _19422_ (.B1(_03600_),
    .Y(_02302_),
    .A1(net6589),
    .A2(net7629));
 sg13g2_nand2_1 _19423_ (.Y(_03601_),
    .A(net3401),
    .B(net6595));
 sg13g2_o21ai_1 _19424_ (.B1(_03601_),
    .Y(_02303_),
    .A1(net6595),
    .A2(net7172));
 sg13g2_nand2_1 _19425_ (.Y(_03602_),
    .A(net3447),
    .B(net6594));
 sg13g2_o21ai_1 _19426_ (.B1(_03602_),
    .Y(_02304_),
    .A1(net6594),
    .A2(net7468));
 sg13g2_nand2_1 _19427_ (.Y(_03603_),
    .A(net3115),
    .B(net6594));
 sg13g2_o21ai_1 _19428_ (.B1(_03603_),
    .Y(_02305_),
    .A1(net6594),
    .A2(net7627));
 sg13g2_nand2_1 _19429_ (.Y(_03604_),
    .A(net3786),
    .B(net6601));
 sg13g2_o21ai_1 _19430_ (.B1(_03604_),
    .Y(_02306_),
    .A1(net6601),
    .A2(net7172));
 sg13g2_nand2_1 _19431_ (.Y(_03605_),
    .A(net4373),
    .B(net6600));
 sg13g2_o21ai_1 _19432_ (.B1(_03605_),
    .Y(_02307_),
    .A1(net6600),
    .A2(net7468));
 sg13g2_nand2_1 _19433_ (.Y(_03606_),
    .A(net2454),
    .B(net6600));
 sg13g2_o21ai_1 _19434_ (.B1(_03606_),
    .Y(_02308_),
    .A1(net6600),
    .A2(net7627));
 sg13g2_nand2_1 _19435_ (.Y(_03607_),
    .A(net4243),
    .B(net6605));
 sg13g2_o21ai_1 _19436_ (.B1(_03607_),
    .Y(_02309_),
    .A1(net6605),
    .A2(net7172));
 sg13g2_nand2_1 _19437_ (.Y(_03608_),
    .A(net3654),
    .B(net6604));
 sg13g2_o21ai_1 _19438_ (.B1(_03608_),
    .Y(_02310_),
    .A1(net6604),
    .A2(net7468));
 sg13g2_nand2_1 _19439_ (.Y(_03609_),
    .A(net2967),
    .B(net6604));
 sg13g2_o21ai_1 _19440_ (.B1(_03609_),
    .Y(_02311_),
    .A1(net6604),
    .A2(net7627));
 sg13g2_nor2_1 _19441_ (.A(net4759),
    .B(net6611),
    .Y(_03610_));
 sg13g2_a21oi_1 _19442_ (.A1(net6610),
    .A2(net7172),
    .Y(_02312_),
    .B1(_03610_));
 sg13g2_nor2_1 _19443_ (.A(net4755),
    .B(net6611),
    .Y(_03611_));
 sg13g2_a21oi_1 _19444_ (.A1(net6610),
    .A2(net7468),
    .Y(_02313_),
    .B1(_03611_));
 sg13g2_nor2_1 _19445_ (.A(net4596),
    .B(net6610),
    .Y(_03612_));
 sg13g2_a21oi_1 _19446_ (.A1(net6610),
    .A2(net7627),
    .Y(_02314_),
    .B1(_03612_));
 sg13g2_nor2_1 _19447_ (.A(net4800),
    .B(net6960),
    .Y(_03613_));
 sg13g2_a21oi_1 _19448_ (.A1(net6960),
    .A2(net7129),
    .Y(_02315_),
    .B1(_03613_));
 sg13g2_nor2_1 _19449_ (.A(net4028),
    .B(net6960),
    .Y(_03614_));
 sg13g2_a21oi_1 _19450_ (.A1(net6960),
    .A2(net7424),
    .Y(_02316_),
    .B1(_03614_));
 sg13g2_nor2_1 _19451_ (.A(net3666),
    .B(net6961),
    .Y(_03615_));
 sg13g2_a21oi_1 _19452_ (.A1(net6961),
    .A2(net7583),
    .Y(_02317_),
    .B1(_03615_));
 sg13g2_nor2_1 _19453_ (.A(net3756),
    .B(net6962),
    .Y(_03616_));
 sg13g2_a21oi_1 _19454_ (.A1(net6962),
    .A2(net7147),
    .Y(_02318_),
    .B1(_03616_));
 sg13g2_nor2_1 _19455_ (.A(net4037),
    .B(net6962),
    .Y(_03617_));
 sg13g2_a21oi_1 _19456_ (.A1(net6962),
    .A2(net7442),
    .Y(_02319_),
    .B1(_03617_));
 sg13g2_nor2_1 _19457_ (.A(net4568),
    .B(net6962),
    .Y(_03618_));
 sg13g2_a21oi_1 _19458_ (.A1(net6962),
    .A2(net7606),
    .Y(_02320_),
    .B1(_03618_));
 sg13g2_nor2_1 _19459_ (.A(net4538),
    .B(net6956),
    .Y(_03619_));
 sg13g2_a21oi_1 _19460_ (.A1(net6956),
    .A2(net7129),
    .Y(_02321_),
    .B1(_03619_));
 sg13g2_nor2_1 _19461_ (.A(net4750),
    .B(net6957),
    .Y(_03620_));
 sg13g2_a21oi_1 _19462_ (.A1(net6957),
    .A2(net7424),
    .Y(_02322_),
    .B1(_03620_));
 sg13g2_nor2_1 _19463_ (.A(net4614),
    .B(net6956),
    .Y(_03621_));
 sg13g2_a21oi_1 _19464_ (.A1(net6956),
    .A2(net7583),
    .Y(_02323_),
    .B1(_03621_));
 sg13g2_nor2_1 _19465_ (.A(net4295),
    .B(net6952),
    .Y(_03622_));
 sg13g2_a21oi_1 _19466_ (.A1(net6952),
    .A2(net7129),
    .Y(_02324_),
    .B1(_03622_));
 sg13g2_nor2_1 _19467_ (.A(net3652),
    .B(net6953),
    .Y(_03623_));
 sg13g2_a21oi_1 _19468_ (.A1(net6953),
    .A2(net7424),
    .Y(_02325_),
    .B1(_03623_));
 sg13g2_nor2_1 _19469_ (.A(net4279),
    .B(net6952),
    .Y(_03624_));
 sg13g2_a21oi_1 _19470_ (.A1(net6952),
    .A2(net7583),
    .Y(_02326_),
    .B1(_03624_));
 sg13g2_nor2_1 _19471_ (.A(net4561),
    .B(net6510),
    .Y(_03625_));
 sg13g2_a21oi_1 _19472_ (.A1(net6510),
    .A2(net7130),
    .Y(_02327_),
    .B1(_03625_));
 sg13g2_nor2_1 _19473_ (.A(net4437),
    .B(net6510),
    .Y(_03626_));
 sg13g2_a21oi_1 _19474_ (.A1(net6510),
    .A2(net7425),
    .Y(_02328_),
    .B1(_03626_));
 sg13g2_nor2_1 _19475_ (.A(net4051),
    .B(net6511),
    .Y(_03627_));
 sg13g2_a21oi_1 _19476_ (.A1(net6511),
    .A2(net7584),
    .Y(_02329_),
    .B1(_03627_));
 sg13g2_nor2_1 _19477_ (.A(net4049),
    .B(net6513),
    .Y(_03628_));
 sg13g2_a21oi_1 _19478_ (.A1(net6513),
    .A2(net7130),
    .Y(_02330_),
    .B1(_03628_));
 sg13g2_nor2_1 _19479_ (.A(net3990),
    .B(net6512),
    .Y(_03629_));
 sg13g2_a21oi_1 _19480_ (.A1(net6512),
    .A2(net7425),
    .Y(_02331_),
    .B1(_03629_));
 sg13g2_nor2_1 _19481_ (.A(net4125),
    .B(net6513),
    .Y(_03630_));
 sg13g2_a21oi_1 _19482_ (.A1(net6513),
    .A2(net7584),
    .Y(_02332_),
    .B1(_03630_));
 sg13g2_nor2_1 _19483_ (.A(net3936),
    .B(net6514),
    .Y(_03631_));
 sg13g2_a21oi_1 _19484_ (.A1(net6514),
    .A2(net7130),
    .Y(_02333_),
    .B1(_03631_));
 sg13g2_nor2_1 _19485_ (.A(net4761),
    .B(net6514),
    .Y(_03632_));
 sg13g2_a21oi_1 _19486_ (.A1(net6514),
    .A2(net7425),
    .Y(_02334_),
    .B1(_03632_));
 sg13g2_nor2_1 _19487_ (.A(net4371),
    .B(net6515),
    .Y(_03633_));
 sg13g2_a21oi_1 _19488_ (.A1(net6515),
    .A2(net7584),
    .Y(_02335_),
    .B1(_03633_));
 sg13g2_nor2_1 _19489_ (.A(net4296),
    .B(net6623),
    .Y(_03634_));
 sg13g2_a21oi_1 _19490_ (.A1(net6622),
    .A2(net7130),
    .Y(_02336_),
    .B1(_03634_));
 sg13g2_nor2_1 _19491_ (.A(net4138),
    .B(net6622),
    .Y(_03635_));
 sg13g2_a21oi_1 _19492_ (.A1(net6622),
    .A2(net7425),
    .Y(_02337_),
    .B1(_03635_));
 sg13g2_nor2_1 _19493_ (.A(net4142),
    .B(net6622),
    .Y(_03636_));
 sg13g2_a21oi_1 _19494_ (.A1(net6623),
    .A2(net7584),
    .Y(_02338_),
    .B1(_03636_));
 sg13g2_nor2_1 _19495_ (.A(net4794),
    .B(net6964),
    .Y(_03637_));
 sg13g2_a21oi_1 _19496_ (.A1(net6964),
    .A2(net7130),
    .Y(_02339_),
    .B1(_03637_));
 sg13g2_nor2_1 _19497_ (.A(net3904),
    .B(net6964),
    .Y(_03638_));
 sg13g2_a21oi_1 _19498_ (.A1(net6964),
    .A2(net7425),
    .Y(_02340_),
    .B1(_03638_));
 sg13g2_nor2_1 _19499_ (.A(net4763),
    .B(net6964),
    .Y(_03639_));
 sg13g2_a21oi_1 _19500_ (.A1(net6964),
    .A2(net7584),
    .Y(_02341_),
    .B1(_03639_));
 sg13g2_nor2_1 _19501_ (.A(net4696),
    .B(net6966),
    .Y(_03640_));
 sg13g2_a21oi_1 _19502_ (.A1(net6966),
    .A2(net7130),
    .Y(_02342_),
    .B1(_03640_));
 sg13g2_nor2_1 _19503_ (.A(net4235),
    .B(net6966),
    .Y(_03641_));
 sg13g2_a21oi_1 _19504_ (.A1(net6966),
    .A2(net7425),
    .Y(_02343_),
    .B1(_03641_));
 sg13g2_nor2_1 _19505_ (.A(net4453),
    .B(net6966),
    .Y(_03642_));
 sg13g2_a21oi_1 _19506_ (.A1(net6966),
    .A2(net7584),
    .Y(_02344_),
    .B1(_03642_));
 sg13g2_nor2_1 _19507_ (.A(net4412),
    .B(net6968),
    .Y(_03643_));
 sg13g2_a21oi_1 _19508_ (.A1(net6968),
    .A2(net7130),
    .Y(_02345_),
    .B1(_03643_));
 sg13g2_nor2_1 _19509_ (.A(net4708),
    .B(net6968),
    .Y(_03644_));
 sg13g2_a21oi_1 _19510_ (.A1(net6968),
    .A2(net7425),
    .Y(_02346_),
    .B1(_03644_));
 sg13g2_nor2_1 _19511_ (.A(net4583),
    .B(net6968),
    .Y(_03645_));
 sg13g2_a21oi_1 _19512_ (.A1(net6968),
    .A2(net7584),
    .Y(_02347_),
    .B1(_03645_));
 sg13g2_nand2_1 _19513_ (.Y(_03646_),
    .A(net2496),
    .B(net6970));
 sg13g2_o21ai_1 _19514_ (.B1(_03646_),
    .Y(_02348_),
    .A1(net6970),
    .A2(net7146));
 sg13g2_nand2_1 _19515_ (.Y(_03647_),
    .A(net2837),
    .B(net6970));
 sg13g2_o21ai_1 _19516_ (.B1(_03647_),
    .Y(_02349_),
    .A1(net6970),
    .A2(net7442));
 sg13g2_nand2_1 _19517_ (.Y(_03648_),
    .A(net3215),
    .B(net6970));
 sg13g2_o21ai_1 _19518_ (.B1(_03648_),
    .Y(_02350_),
    .A1(net6970),
    .A2(net7606));
 sg13g2_nor2_1 _19519_ (.A(net3949),
    .B(net6972),
    .Y(_03649_));
 sg13g2_a21oi_1 _19520_ (.A1(net6972),
    .A2(net7129),
    .Y(_02351_),
    .B1(_03649_));
 sg13g2_nor2_1 _19521_ (.A(net3890),
    .B(net6972),
    .Y(_03650_));
 sg13g2_a21oi_1 _19522_ (.A1(net6972),
    .A2(net7424),
    .Y(_02352_),
    .B1(_03650_));
 sg13g2_nor2_1 _19523_ (.A(net4729),
    .B(net6973),
    .Y(_03651_));
 sg13g2_a21oi_1 _19524_ (.A1(net6973),
    .A2(net7583),
    .Y(_02353_),
    .B1(_03651_));
 sg13g2_nor2_1 _19525_ (.A(net4793),
    .B(net6974),
    .Y(_03652_));
 sg13g2_a21oi_1 _19526_ (.A1(net6974),
    .A2(net7129),
    .Y(_02354_),
    .B1(_03652_));
 sg13g2_nor2_1 _19527_ (.A(net4260),
    .B(net6974),
    .Y(_03653_));
 sg13g2_a21oi_1 _19528_ (.A1(net6974),
    .A2(net7424),
    .Y(_02355_),
    .B1(_03653_));
 sg13g2_nor2_1 _19529_ (.A(net4524),
    .B(net6975),
    .Y(_03654_));
 sg13g2_a21oi_1 _19530_ (.A1(net6975),
    .A2(net7583),
    .Y(_02356_),
    .B1(_03654_));
 sg13g2_nor2_1 _19531_ (.A(net3948),
    .B(net6976),
    .Y(_03655_));
 sg13g2_a21oi_1 _19532_ (.A1(net6976),
    .A2(net7129),
    .Y(_02357_),
    .B1(_03655_));
 sg13g2_nor2_1 _19533_ (.A(net4171),
    .B(net6976),
    .Y(_03656_));
 sg13g2_a21oi_1 _19534_ (.A1(net6976),
    .A2(net7424),
    .Y(_02358_),
    .B1(_03656_));
 sg13g2_nor2_1 _19535_ (.A(net4702),
    .B(net6977),
    .Y(_03657_));
 sg13g2_a21oi_1 _19536_ (.A1(net6977),
    .A2(net7583),
    .Y(_02359_),
    .B1(_03657_));
 sg13g2_nor2_1 _19537_ (.A(net4555),
    .B(net6978),
    .Y(_03658_));
 sg13g2_a21oi_1 _19538_ (.A1(net6978),
    .A2(net7129),
    .Y(_02360_),
    .B1(_03658_));
 sg13g2_nor2_1 _19539_ (.A(net4205),
    .B(net6978),
    .Y(_03659_));
 sg13g2_a21oi_1 _19540_ (.A1(net6978),
    .A2(net7424),
    .Y(_02361_),
    .B1(_03659_));
 sg13g2_nor2_1 _19541_ (.A(net4777),
    .B(net6979),
    .Y(_03660_));
 sg13g2_a21oi_1 _19542_ (.A1(net6979),
    .A2(net7583),
    .Y(_02362_),
    .B1(_03660_));
 sg13g2_nor2_1 _19543_ (.A(net4190),
    .B(net6980),
    .Y(_03661_));
 sg13g2_a21oi_1 _19544_ (.A1(net6980),
    .A2(net7132),
    .Y(_02363_),
    .B1(_03661_));
 sg13g2_nor2_1 _19545_ (.A(net3627),
    .B(net6980),
    .Y(_03662_));
 sg13g2_a21oi_1 _19546_ (.A1(net6980),
    .A2(net7439),
    .Y(_02364_),
    .B1(_03662_));
 sg13g2_nor2_1 _19547_ (.A(net4459),
    .B(net6981),
    .Y(_03663_));
 sg13g2_a21oi_1 _19548_ (.A1(net6981),
    .A2(net7587),
    .Y(_02365_),
    .B1(_03663_));
 sg13g2_nor2_1 _19549_ (.A(net4465),
    .B(net6982),
    .Y(_03664_));
 sg13g2_a21oi_1 _19550_ (.A1(net6982),
    .A2(net7132),
    .Y(_02366_),
    .B1(_03664_));
 sg13g2_nor2_1 _19551_ (.A(net3809),
    .B(net6983),
    .Y(_03665_));
 sg13g2_a21oi_1 _19552_ (.A1(net6982),
    .A2(net7439),
    .Y(_02367_),
    .B1(_03665_));
 sg13g2_nor2_1 _19553_ (.A(net4677),
    .B(net6982),
    .Y(_03666_));
 sg13g2_a21oi_1 _19554_ (.A1(net6983),
    .A2(net7587),
    .Y(_02368_),
    .B1(_03666_));
 sg13g2_nor2_1 _19555_ (.A(net4569),
    .B(net6984),
    .Y(_03667_));
 sg13g2_a21oi_1 _19556_ (.A1(net6984),
    .A2(net7132),
    .Y(_02369_),
    .B1(_03667_));
 sg13g2_nor2_1 _19557_ (.A(net4830),
    .B(net6985),
    .Y(_03668_));
 sg13g2_a21oi_1 _19558_ (.A1(net6985),
    .A2(net7439),
    .Y(_02370_),
    .B1(_03668_));
 sg13g2_nor2_1 _19559_ (.A(net4222),
    .B(net6984),
    .Y(_03669_));
 sg13g2_a21oi_1 _19560_ (.A1(net6984),
    .A2(net7587),
    .Y(_02371_),
    .B1(_03669_));
 sg13g2_nand2_1 _19561_ (.Y(_03670_),
    .A(net2971),
    .B(net6986));
 sg13g2_o21ai_1 _19562_ (.B1(_03670_),
    .Y(_02372_),
    .A1(net6986),
    .A2(net7132));
 sg13g2_nand2_1 _19563_ (.Y(_03671_),
    .A(net2452),
    .B(net6987));
 sg13g2_o21ai_1 _19564_ (.B1(_03671_),
    .Y(_02373_),
    .A1(net6986),
    .A2(net7439));
 sg13g2_nand2_1 _19565_ (.Y(_03672_),
    .A(net3527),
    .B(net6986));
 sg13g2_o21ai_1 _19566_ (.B1(_03672_),
    .Y(_02374_),
    .A1(net6987),
    .A2(net7587));
 sg13g2_nand2_1 _19567_ (.Y(_03673_),
    .A(net3568),
    .B(net6988));
 sg13g2_o21ai_1 _19568_ (.B1(_03673_),
    .Y(_02375_),
    .A1(net6988),
    .A2(net7146));
 sg13g2_nand2_1 _19569_ (.Y(_03674_),
    .A(net3774),
    .B(net6989));
 sg13g2_o21ai_1 _19570_ (.B1(_03674_),
    .Y(_02376_),
    .A1(net6989),
    .A2(net7441));
 sg13g2_nand2_1 _19571_ (.Y(_03675_),
    .A(net3526),
    .B(net6988));
 sg13g2_o21ai_1 _19572_ (.B1(_03675_),
    .Y(_02377_),
    .A1(net6988),
    .A2(net7587));
 sg13g2_nand2_1 _19573_ (.Y(_03676_),
    .A(net4206),
    .B(net6991));
 sg13g2_o21ai_1 _19574_ (.B1(_03676_),
    .Y(_02378_),
    .A1(net6991),
    .A2(net7146));
 sg13g2_nand2_1 _19575_ (.Y(_03677_),
    .A(net3024),
    .B(net6991));
 sg13g2_o21ai_1 _19576_ (.B1(_03677_),
    .Y(_02379_),
    .A1(net6991),
    .A2(net7442));
 sg13g2_nand2_1 _19577_ (.Y(_03678_),
    .A(net3020),
    .B(net6990));
 sg13g2_o21ai_1 _19578_ (.B1(_03678_),
    .Y(_02380_),
    .A1(net6990),
    .A2(net7599));
 sg13g2_nand2_1 _19579_ (.Y(_03679_),
    .A(net3513),
    .B(net6992));
 sg13g2_o21ai_1 _19580_ (.B1(_03679_),
    .Y(_02381_),
    .A1(net6993),
    .A2(net7145));
 sg13g2_nand2_1 _19581_ (.Y(_03680_),
    .A(net3974),
    .B(net6993));
 sg13g2_o21ai_1 _19582_ (.B1(_03680_),
    .Y(_02382_),
    .A1(net6992),
    .A2(net7441));
 sg13g2_nand2_1 _19583_ (.Y(_03681_),
    .A(net3465),
    .B(net6992));
 sg13g2_o21ai_1 _19584_ (.B1(_03681_),
    .Y(_02383_),
    .A1(net6992),
    .A2(net7589));
 sg13g2_nand2_1 _19585_ (.Y(_03682_),
    .A(net3499),
    .B(net6994));
 sg13g2_o21ai_1 _19586_ (.B1(_03682_),
    .Y(_02384_),
    .A1(net6994),
    .A2(net7132));
 sg13g2_nand2_1 _19587_ (.Y(_03683_),
    .A(net3507),
    .B(net6995));
 sg13g2_o21ai_1 _19588_ (.B1(_03683_),
    .Y(_02385_),
    .A1(net6995),
    .A2(net7441));
 sg13g2_nand2_1 _19589_ (.Y(_03684_),
    .A(net2913),
    .B(net6994));
 sg13g2_o21ai_1 _19590_ (.B1(_03684_),
    .Y(_02386_),
    .A1(net6994),
    .A2(net7587));
 sg13g2_nand2_1 _19591_ (.Y(_03685_),
    .A(net3181),
    .B(net6624));
 sg13g2_o21ai_1 _19592_ (.B1(_03685_),
    .Y(_02387_),
    .A1(net6624),
    .A2(net7146));
 sg13g2_nand2_1 _19593_ (.Y(_03686_),
    .A(net2862),
    .B(net6625));
 sg13g2_o21ai_1 _19594_ (.B1(_03686_),
    .Y(_02388_),
    .A1(net6625),
    .A2(net7440));
 sg13g2_nand2_1 _19595_ (.Y(_03687_),
    .A(net2699),
    .B(net6624));
 sg13g2_o21ai_1 _19596_ (.B1(_03687_),
    .Y(_02389_),
    .A1(net6624),
    .A2(net7599));
 sg13g2_nand2_1 _19597_ (.Y(_03688_),
    .A(net3134),
    .B(net6626));
 sg13g2_o21ai_1 _19598_ (.B1(_03688_),
    .Y(_02390_),
    .A1(net6626),
    .A2(net7146));
 sg13g2_nand2_1 _19599_ (.Y(_03689_),
    .A(net4012),
    .B(net6627));
 sg13g2_o21ai_1 _19600_ (.B1(_03689_),
    .Y(_02391_),
    .A1(net6627),
    .A2(net7440));
 sg13g2_nand2_1 _19601_ (.Y(_03690_),
    .A(net2821),
    .B(net6626));
 sg13g2_o21ai_1 _19602_ (.B1(_03690_),
    .Y(_02392_),
    .A1(net6626),
    .A2(net7599));
 sg13g2_nand2_1 _19603_ (.Y(_03691_),
    .A(net2786),
    .B(net6628));
 sg13g2_o21ai_1 _19604_ (.B1(_03691_),
    .Y(_02393_),
    .A1(net6628),
    .A2(net7146));
 sg13g2_nand2_1 _19605_ (.Y(_03692_),
    .A(net3089),
    .B(net6629));
 sg13g2_o21ai_1 _19606_ (.B1(_03692_),
    .Y(_02394_),
    .A1(net6629),
    .A2(net7440));
 sg13g2_nand2_1 _19607_ (.Y(_03693_),
    .A(net3889),
    .B(net6628));
 sg13g2_o21ai_1 _19608_ (.B1(_03693_),
    .Y(_02395_),
    .A1(net6628),
    .A2(net7599));
 sg13g2_nand2_1 _19609_ (.Y(_03694_),
    .A(net3301),
    .B(net6630));
 sg13g2_o21ai_1 _19610_ (.B1(_03694_),
    .Y(_02396_),
    .A1(net6630),
    .A2(net7146));
 sg13g2_nand2_1 _19611_ (.Y(_03695_),
    .A(net3737),
    .B(net6631));
 sg13g2_o21ai_1 _19612_ (.B1(_03695_),
    .Y(_02397_),
    .A1(net6631),
    .A2(net7440));
 sg13g2_nand2_1 _19613_ (.Y(_03696_),
    .A(net2874),
    .B(net6630));
 sg13g2_o21ai_1 _19614_ (.B1(_03696_),
    .Y(_02398_),
    .A1(net6630),
    .A2(net7599));
 sg13g2_nand2_1 _19615_ (.Y(_03697_),
    .A(net4366),
    .B(net6996));
 sg13g2_o21ai_1 _19616_ (.B1(_03697_),
    .Y(_02399_),
    .A1(net6996),
    .A2(net7133));
 sg13g2_nand2_1 _19617_ (.Y(_03698_),
    .A(net3579),
    .B(net6996));
 sg13g2_o21ai_1 _19618_ (.B1(_03698_),
    .Y(_02400_),
    .A1(net6996),
    .A2(net7439));
 sg13g2_nand2_1 _19619_ (.Y(_03699_),
    .A(net3344),
    .B(net6997));
 sg13g2_o21ai_1 _19620_ (.B1(_03699_),
    .Y(_02401_),
    .A1(net6997),
    .A2(net7588));
 sg13g2_nand2_1 _19621_ (.Y(_03700_),
    .A(net3619),
    .B(net6998));
 sg13g2_o21ai_1 _19622_ (.B1(_03700_),
    .Y(_02402_),
    .A1(net6998),
    .A2(net7133));
 sg13g2_nand2_1 _19623_ (.Y(_03701_),
    .A(net2481),
    .B(net6998));
 sg13g2_o21ai_1 _19624_ (.B1(_03701_),
    .Y(_02403_),
    .A1(net6998),
    .A2(net7439));
 sg13g2_nand2_1 _19625_ (.Y(_03702_),
    .A(net3564),
    .B(net6999));
 sg13g2_o21ai_1 _19626_ (.B1(_03702_),
    .Y(_02404_),
    .A1(net6999),
    .A2(net7588));
 sg13g2_nand2_1 _19627_ (.Y(_03703_),
    .A(net2841),
    .B(net7000));
 sg13g2_o21ai_1 _19628_ (.B1(_03703_),
    .Y(_02405_),
    .A1(net7000),
    .A2(net7132));
 sg13g2_nand2_1 _19629_ (.Y(_03704_),
    .A(net3040),
    .B(net7001));
 sg13g2_o21ai_1 _19630_ (.B1(_03704_),
    .Y(_02406_),
    .A1(net7000),
    .A2(net7439));
 sg13g2_nand2_1 _19631_ (.Y(_03705_),
    .A(net3357),
    .B(net7000));
 sg13g2_o21ai_1 _19632_ (.B1(_03705_),
    .Y(_02407_),
    .A1(net7001),
    .A2(net7587));
 sg13g2_nor2_1 _19633_ (.A(net4631),
    .B(net7002),
    .Y(_03706_));
 sg13g2_a21oi_1 _19634_ (.A1(net7003),
    .A2(net7146),
    .Y(_02408_),
    .B1(_03706_));
 sg13g2_nor2_1 _19635_ (.A(net4686),
    .B(net7002),
    .Y(_03707_));
 sg13g2_a21oi_1 _19636_ (.A1(net7002),
    .A2(net7442),
    .Y(_02409_),
    .B1(_03707_));
 sg13g2_nor2_1 _19637_ (.A(net3463),
    .B(net7002),
    .Y(_03708_));
 sg13g2_a21oi_1 _19638_ (.A1(net7002),
    .A2(net7599),
    .Y(_02410_),
    .B1(_03708_));
 sg13g2_nor2_1 _19639_ (.A(net4796),
    .B(net7004),
    .Y(_03709_));
 sg13g2_a21oi_1 _19640_ (.A1(net7005),
    .A2(net7148),
    .Y(_02411_),
    .B1(_03709_));
 sg13g2_nor2_1 _19641_ (.A(net4634),
    .B(net7004),
    .Y(_03710_));
 sg13g2_a21oi_1 _19642_ (.A1(net7005),
    .A2(net7443),
    .Y(_02412_),
    .B1(_03710_));
 sg13g2_nor2_1 _19643_ (.A(net4176),
    .B(net7004),
    .Y(_03711_));
 sg13g2_a21oi_1 _19644_ (.A1(net7004),
    .A2(net7601),
    .Y(_02413_),
    .B1(_03711_));
 sg13g2_nor2_1 _19645_ (.A(net4613),
    .B(net7007),
    .Y(_03712_));
 sg13g2_a21oi_1 _19646_ (.A1(net7006),
    .A2(net7148),
    .Y(_02414_),
    .B1(_03712_));
 sg13g2_nor2_1 _19647_ (.A(net4714),
    .B(net7006),
    .Y(_03713_));
 sg13g2_a21oi_1 _19648_ (.A1(net7007),
    .A2(net7443),
    .Y(_02415_),
    .B1(_03713_));
 sg13g2_nor2_1 _19649_ (.A(net4808),
    .B(net7006),
    .Y(_03714_));
 sg13g2_a21oi_1 _19650_ (.A1(net7006),
    .A2(net7601),
    .Y(_02416_),
    .B1(_03714_));
 sg13g2_nor2_1 _19651_ (.A(net4717),
    .B(net7009),
    .Y(_03715_));
 sg13g2_a21oi_1 _19652_ (.A1(net7009),
    .A2(net7148),
    .Y(_02417_),
    .B1(_03715_));
 sg13g2_nor2_1 _19653_ (.A(net4079),
    .B(net7008),
    .Y(_03716_));
 sg13g2_a21oi_1 _19654_ (.A1(net7008),
    .A2(net7443),
    .Y(_02418_),
    .B1(_03716_));
 sg13g2_nor2_1 _19655_ (.A(net4400),
    .B(net7008),
    .Y(_03717_));
 sg13g2_a21oi_1 _19656_ (.A1(net7008),
    .A2(net7601),
    .Y(_02419_),
    .B1(_03717_));
 sg13g2_nand2_1 _19657_ (.Y(_03718_),
    .A(net3305),
    .B(net6633));
 sg13g2_o21ai_1 _19658_ (.B1(_03718_),
    .Y(_02420_),
    .A1(net6633),
    .A2(net7148));
 sg13g2_nand2_1 _19659_ (.Y(_03719_),
    .A(net3027),
    .B(net6632));
 sg13g2_o21ai_1 _19660_ (.B1(_03719_),
    .Y(_02421_),
    .A1(net6632),
    .A2(net7443));
 sg13g2_nand2_1 _19661_ (.Y(_03720_),
    .A(net2847),
    .B(net6632));
 sg13g2_o21ai_1 _19662_ (.B1(_03720_),
    .Y(_02422_),
    .A1(net6632),
    .A2(net7601));
 sg13g2_nand2_1 _19663_ (.Y(_03721_),
    .A(net2526),
    .B(net6634));
 sg13g2_o21ai_1 _19664_ (.B1(_03721_),
    .Y(_02423_),
    .A1(net6634),
    .A2(net7152));
 sg13g2_nand2_1 _19665_ (.Y(_03722_),
    .A(net2511),
    .B(net6635));
 sg13g2_o21ai_1 _19666_ (.B1(_03722_),
    .Y(_02424_),
    .A1(net6634),
    .A2(net7443));
 sg13g2_nand2_1 _19667_ (.Y(_03723_),
    .A(net3026),
    .B(net6635));
 sg13g2_o21ai_1 _19668_ (.B1(_03723_),
    .Y(_02425_),
    .A1(net6634),
    .A2(net7602));
 sg13g2_nand2_1 _19669_ (.Y(_03724_),
    .A(net3118),
    .B(net6636));
 sg13g2_o21ai_1 _19670_ (.B1(_03724_),
    .Y(_02426_),
    .A1(net6636),
    .A2(net7148));
 sg13g2_nand2_1 _19671_ (.Y(_03725_),
    .A(net2932),
    .B(net6636));
 sg13g2_o21ai_1 _19672_ (.B1(_03725_),
    .Y(_02427_),
    .A1(net6636),
    .A2(net7443));
 sg13g2_nand2_1 _19673_ (.Y(_03726_),
    .A(net3556),
    .B(net6637));
 sg13g2_o21ai_1 _19674_ (.B1(_03726_),
    .Y(_02428_),
    .A1(net6637),
    .A2(net7602));
 sg13g2_nand2_1 _19675_ (.Y(_03727_),
    .A(net3270),
    .B(net6638));
 sg13g2_o21ai_1 _19676_ (.B1(_03727_),
    .Y(_02429_),
    .A1(net6638),
    .A2(net7148));
 sg13g2_nand2_1 _19677_ (.Y(_03728_),
    .A(net2714),
    .B(net6638));
 sg13g2_o21ai_1 _19678_ (.B1(_03728_),
    .Y(_02430_),
    .A1(net6638),
    .A2(net7446));
 sg13g2_nand2_1 _19679_ (.Y(_03729_),
    .A(net3173),
    .B(net6639));
 sg13g2_o21ai_1 _19680_ (.B1(_03729_),
    .Y(_02431_),
    .A1(net6639),
    .A2(net7602));
 sg13g2_nand2_1 _19681_ (.Y(_03730_),
    .A(net2990),
    .B(net6640));
 sg13g2_o21ai_1 _19682_ (.B1(_03730_),
    .Y(_02432_),
    .A1(net6640),
    .A2(net7148));
 sg13g2_nand2_1 _19683_ (.Y(_03731_),
    .A(net3769),
    .B(net6640));
 sg13g2_o21ai_1 _19684_ (.B1(_03731_),
    .Y(_02433_),
    .A1(net6640),
    .A2(net7446));
 sg13g2_nand2_1 _19685_ (.Y(_03732_),
    .A(net3983),
    .B(net6641));
 sg13g2_o21ai_1 _19686_ (.B1(_03732_),
    .Y(_02434_),
    .A1(net6641),
    .A2(net7602));
 sg13g2_nand2_1 _19687_ (.Y(_03733_),
    .A(net2502),
    .B(net6643));
 sg13g2_o21ai_1 _19688_ (.B1(_03733_),
    .Y(_02435_),
    .A1(net6642),
    .A2(net7143));
 sg13g2_nand2_1 _19689_ (.Y(_03734_),
    .A(net2442),
    .B(net6642));
 sg13g2_o21ai_1 _19690_ (.B1(_03734_),
    .Y(_02436_),
    .A1(net6642),
    .A2(net7443));
 sg13g2_nand2_1 _19691_ (.Y(_03735_),
    .A(net3039),
    .B(net6642));
 sg13g2_o21ai_1 _19692_ (.B1(_03735_),
    .Y(_02437_),
    .A1(net6643),
    .A2(net7601));
 sg13g2_nand2_1 _19693_ (.Y(_03736_),
    .A(net3188),
    .B(net7010));
 sg13g2_o21ai_1 _19694_ (.B1(_03736_),
    .Y(_02438_),
    .A1(net7010),
    .A2(net7164));
 sg13g2_nand2_1 _19695_ (.Y(_03737_),
    .A(net3083),
    .B(net7010));
 sg13g2_o21ai_1 _19696_ (.B1(_03737_),
    .Y(_02439_),
    .A1(net7010),
    .A2(net7458));
 sg13g2_nand2_1 _19697_ (.Y(_03738_),
    .A(net2943),
    .B(net7010));
 sg13g2_o21ai_1 _19698_ (.B1(_03738_),
    .Y(_02440_),
    .A1(net7010),
    .A2(net7619));
 sg13g2_nand2_1 _19699_ (.Y(_03739_),
    .A(net4099),
    .B(net6644));
 sg13g2_o21ai_1 _19700_ (.B1(_03739_),
    .Y(_02441_),
    .A1(net6644),
    .A2(net7165));
 sg13g2_nand2_1 _19701_ (.Y(_03740_),
    .A(net3819),
    .B(net6645));
 sg13g2_o21ai_1 _19702_ (.B1(_03740_),
    .Y(_02442_),
    .A1(net6645),
    .A2(net7461));
 sg13g2_nand2_1 _19703_ (.Y(_03741_),
    .A(net4202),
    .B(net6644));
 sg13g2_o21ai_1 _19704_ (.B1(_03741_),
    .Y(_02443_),
    .A1(net6644),
    .A2(net7616));
 sg13g2_nand2_1 _19705_ (.Y(_03742_),
    .A(net3363),
    .B(net6646));
 sg13g2_o21ai_1 _19706_ (.B1(_03742_),
    .Y(_02444_),
    .A1(net6646),
    .A2(net7165));
 sg13g2_nand2_1 _19707_ (.Y(_03743_),
    .A(net2622),
    .B(net6647));
 sg13g2_o21ai_1 _19708_ (.B1(_03743_),
    .Y(_02445_),
    .A1(net6647),
    .A2(net7461));
 sg13g2_nand2_1 _19709_ (.Y(_03744_),
    .A(net2799),
    .B(net6646));
 sg13g2_o21ai_1 _19710_ (.B1(_03744_),
    .Y(_02446_),
    .A1(net6646),
    .A2(net7616));
 sg13g2_nand2_1 _19711_ (.Y(_03745_),
    .A(net2872),
    .B(net6649));
 sg13g2_o21ai_1 _19712_ (.B1(_03745_),
    .Y(_02447_),
    .A1(net6649),
    .A2(net7143));
 sg13g2_nand2_1 _19713_ (.Y(_03746_),
    .A(net3504),
    .B(net6648));
 sg13g2_o21ai_1 _19714_ (.B1(_03746_),
    .Y(_02448_),
    .A1(net6648),
    .A2(net7437));
 sg13g2_nand2_1 _19715_ (.Y(_03747_),
    .A(net3927),
    .B(net6648));
 sg13g2_o21ai_1 _19716_ (.B1(_03747_),
    .Y(_02449_),
    .A1(net6648),
    .A2(net7597));
 sg13g2_nand2_1 _19717_ (.Y(_03748_),
    .A(net4628),
    .B(net6651));
 sg13g2_o21ai_1 _19718_ (.B1(_03748_),
    .Y(_02450_),
    .A1(net6651),
    .A2(net7143));
 sg13g2_nand2_1 _19719_ (.Y(_03749_),
    .A(net2776),
    .B(net6650));
 sg13g2_o21ai_1 _19720_ (.B1(_03749_),
    .Y(_02451_),
    .A1(net6650),
    .A2(net7437));
 sg13g2_nand2_1 _19721_ (.Y(_03750_),
    .A(net3023),
    .B(net6650));
 sg13g2_o21ai_1 _19722_ (.B1(_03750_),
    .Y(_02452_),
    .A1(net6650),
    .A2(net7597));
 sg13g2_nand2_1 _19723_ (.Y(_03751_),
    .A(net3156),
    .B(net6652));
 sg13g2_o21ai_1 _19724_ (.B1(_03751_),
    .Y(_02453_),
    .A1(net6652),
    .A2(net7143));
 sg13g2_nand2_1 _19725_ (.Y(_03752_),
    .A(net2624),
    .B(net6653));
 sg13g2_o21ai_1 _19726_ (.B1(_03752_),
    .Y(_02454_),
    .A1(net6652),
    .A2(net7436));
 sg13g2_nand2_1 _19727_ (.Y(_03753_),
    .A(net3078),
    .B(net6652));
 sg13g2_o21ai_1 _19728_ (.B1(_03753_),
    .Y(_02455_),
    .A1(net6652),
    .A2(net7597));
 sg13g2_nand2_1 _19729_ (.Y(_03754_),
    .A(net3541),
    .B(net6655));
 sg13g2_o21ai_1 _19730_ (.B1(_03754_),
    .Y(_02456_),
    .A1(net6654),
    .A2(net7142));
 sg13g2_nand2_1 _19731_ (.Y(_03755_),
    .A(net3744),
    .B(net6654));
 sg13g2_o21ai_1 _19732_ (.B1(_03755_),
    .Y(_02457_),
    .A1(net6654),
    .A2(net7437));
 sg13g2_nand2_1 _19733_ (.Y(_03756_),
    .A(net2577),
    .B(net6654));
 sg13g2_o21ai_1 _19734_ (.B1(_03756_),
    .Y(_02458_),
    .A1(net6654),
    .A2(net7597));
 sg13g2_nand2_1 _19735_ (.Y(_03757_),
    .A(net3259),
    .B(net7013));
 sg13g2_o21ai_1 _19736_ (.B1(_03757_),
    .Y(_02459_),
    .A1(net7013),
    .A2(net7168));
 sg13g2_nand2_1 _19737_ (.Y(_03758_),
    .A(net3074),
    .B(net7013));
 sg13g2_o21ai_1 _19738_ (.B1(_03758_),
    .Y(_02460_),
    .A1(net7013),
    .A2(net7465));
 sg13g2_nand2_1 _19739_ (.Y(_03759_),
    .A(net3320),
    .B(net7012));
 sg13g2_o21ai_1 _19740_ (.B1(_03759_),
    .Y(_02461_),
    .A1(net7012),
    .A2(net7623));
 sg13g2_nand2_1 _19741_ (.Y(_03760_),
    .A(net3583),
    .B(net7015));
 sg13g2_o21ai_1 _19742_ (.B1(_03760_),
    .Y(_02462_),
    .A1(net7015),
    .A2(net7168));
 sg13g2_nand2_1 _19743_ (.Y(_03761_),
    .A(net2534),
    .B(net7015));
 sg13g2_o21ai_1 _19744_ (.B1(_03761_),
    .Y(_02463_),
    .A1(net7015),
    .A2(net7465));
 sg13g2_nand2_1 _19745_ (.Y(_03762_),
    .A(net2689),
    .B(net7014));
 sg13g2_o21ai_1 _19746_ (.B1(_03762_),
    .Y(_02464_),
    .A1(net7014),
    .A2(net7623));
 sg13g2_nand2_1 _19747_ (.Y(_03763_),
    .A(net3514),
    .B(net7017));
 sg13g2_o21ai_1 _19748_ (.B1(_03763_),
    .Y(_02465_),
    .A1(net7017),
    .A2(net7168));
 sg13g2_nand2_1 _19749_ (.Y(_03764_),
    .A(net3805),
    .B(net7016));
 sg13g2_o21ai_1 _19750_ (.B1(_03764_),
    .Y(_02466_),
    .A1(net7016),
    .A2(net7465));
 sg13g2_nand2_1 _19751_ (.Y(_03765_),
    .A(net3728),
    .B(net7016));
 sg13g2_o21ai_1 _19752_ (.B1(_03765_),
    .Y(_02467_),
    .A1(net7016),
    .A2(net7623));
 sg13g2_nand2_1 _19753_ (.Y(_03766_),
    .A(net2466),
    .B(net7018));
 sg13g2_o21ai_1 _19754_ (.B1(_03766_),
    .Y(_02468_),
    .A1(net7018),
    .A2(net7164));
 sg13g2_nand2_1 _19755_ (.Y(_03767_),
    .A(net3909),
    .B(net7018));
 sg13g2_o21ai_1 _19756_ (.B1(_03767_),
    .Y(_02469_),
    .A1(net7018),
    .A2(net7458));
 sg13g2_nand2_1 _19757_ (.Y(_03768_),
    .A(net3484),
    .B(net7018));
 sg13g2_o21ai_1 _19758_ (.B1(_03768_),
    .Y(_02470_),
    .A1(net7018),
    .A2(net7619));
 sg13g2_nand2_1 _19759_ (.Y(_03769_),
    .A(net2540),
    .B(net7020));
 sg13g2_o21ai_1 _19760_ (.B1(_03769_),
    .Y(_02471_),
    .A1(net7020),
    .A2(net7169));
 sg13g2_nand2_1 _19761_ (.Y(_03770_),
    .A(net2570),
    .B(net7021));
 sg13g2_o21ai_1 _19762_ (.B1(_03770_),
    .Y(_02472_),
    .A1(net7021),
    .A2(net7462));
 sg13g2_nand2_1 _19763_ (.Y(_03771_),
    .A(net2683),
    .B(net7020));
 sg13g2_o21ai_1 _19764_ (.B1(_03771_),
    .Y(_02473_),
    .A1(net7020),
    .A2(net7617));
 sg13g2_nand2_1 _19765_ (.Y(_03772_),
    .A(net2598),
    .B(net7022));
 sg13g2_o21ai_1 _19766_ (.B1(_03772_),
    .Y(_02474_),
    .A1(net7022),
    .A2(net7169));
 sg13g2_nand2_1 _19767_ (.Y(_03773_),
    .A(net3106),
    .B(net7023));
 sg13g2_o21ai_1 _19768_ (.B1(_03773_),
    .Y(_02475_),
    .A1(net7023),
    .A2(net7462));
 sg13g2_nand2_1 _19769_ (.Y(_03774_),
    .A(net3531),
    .B(net7022));
 sg13g2_o21ai_1 _19770_ (.B1(_03774_),
    .Y(_02476_),
    .A1(net7022),
    .A2(net7617));
 sg13g2_nand2_1 _19771_ (.Y(_03775_),
    .A(net3137),
    .B(net7025));
 sg13g2_o21ai_1 _19772_ (.B1(_03775_),
    .Y(_02477_),
    .A1(net7024),
    .A2(net7169));
 sg13g2_nand2_1 _19773_ (.Y(_03776_),
    .A(net3362),
    .B(net7025));
 sg13g2_o21ai_1 _19774_ (.B1(_03776_),
    .Y(_02478_),
    .A1(net7025),
    .A2(net7462));
 sg13g2_nand2_1 _19775_ (.Y(_03777_),
    .A(net2716),
    .B(net7024));
 sg13g2_o21ai_1 _19776_ (.B1(_03777_),
    .Y(_02479_),
    .A1(net7024),
    .A2(net7622));
 sg13g2_nand2_1 _19777_ (.Y(_03778_),
    .A(net2915),
    .B(net7026));
 sg13g2_o21ai_1 _19778_ (.B1(_03778_),
    .Y(_02480_),
    .A1(net7026),
    .A2(net7169));
 sg13g2_nand2_1 _19779_ (.Y(_03779_),
    .A(net2953),
    .B(net7027));
 sg13g2_o21ai_1 _19780_ (.B1(_03779_),
    .Y(_02481_),
    .A1(net7027),
    .A2(net7462));
 sg13g2_nand2_1 _19781_ (.Y(_03780_),
    .A(net2593),
    .B(net7026));
 sg13g2_o21ai_1 _19782_ (.B1(_03780_),
    .Y(_02482_),
    .A1(net7026),
    .A2(net7622));
 sg13g2_nand2_1 _19783_ (.Y(_03781_),
    .A(net2560),
    .B(net6656));
 sg13g2_o21ai_1 _19784_ (.B1(_03781_),
    .Y(_02483_),
    .A1(net6656),
    .A2(net7164));
 sg13g2_nand2_1 _19785_ (.Y(_03782_),
    .A(net2750),
    .B(net6657));
 sg13g2_o21ai_1 _19786_ (.B1(_03782_),
    .Y(_02484_),
    .A1(net6656),
    .A2(net7459));
 sg13g2_nand2_1 _19787_ (.Y(_03783_),
    .A(net4436),
    .B(net6657));
 sg13g2_o21ai_1 _19788_ (.B1(_03783_),
    .Y(_02485_),
    .A1(net6657),
    .A2(net7618));
 sg13g2_nand2_1 _19789_ (.Y(_03784_),
    .A(net3452),
    .B(net6658));
 sg13g2_o21ai_1 _19790_ (.B1(_03784_),
    .Y(_02486_),
    .A1(net6658),
    .A2(net7164));
 sg13g2_nand2_1 _19791_ (.Y(_03785_),
    .A(net3180),
    .B(net6659));
 sg13g2_o21ai_1 _19792_ (.B1(_03785_),
    .Y(_02487_),
    .A1(net6658),
    .A2(net7459));
 sg13g2_nand2_1 _19793_ (.Y(_03786_),
    .A(net3337),
    .B(net6659));
 sg13g2_o21ai_1 _19794_ (.B1(_03786_),
    .Y(_02488_),
    .A1(net6659),
    .A2(net7618));
 sg13g2_nand2_1 _19795_ (.Y(_03787_),
    .A(net3887),
    .B(net6660));
 sg13g2_o21ai_1 _19796_ (.B1(_03787_),
    .Y(_02489_),
    .A1(net6660),
    .A2(net7164));
 sg13g2_nand2_1 _19797_ (.Y(_03788_),
    .A(net3575),
    .B(net6661));
 sg13g2_o21ai_1 _19798_ (.B1(_03788_),
    .Y(_02490_),
    .A1(net6661),
    .A2(net7459));
 sg13g2_nand2_1 _19799_ (.Y(_03789_),
    .A(net2843),
    .B(net6660));
 sg13g2_o21ai_1 _19800_ (.B1(_03789_),
    .Y(_02491_),
    .A1(net6661),
    .A2(net7618));
 sg13g2_nand2_1 _19801_ (.Y(_03790_),
    .A(net3145),
    .B(net6662));
 sg13g2_o21ai_1 _19802_ (.B1(_03790_),
    .Y(_02492_),
    .A1(net6662),
    .A2(net7164));
 sg13g2_nand2_1 _19803_ (.Y(_03791_),
    .A(net3242),
    .B(net6663));
 sg13g2_o21ai_1 _19804_ (.B1(_03791_),
    .Y(_02493_),
    .A1(net6662),
    .A2(net7459));
 sg13g2_nand2_1 _19805_ (.Y(_03792_),
    .A(net3223),
    .B(net6663));
 sg13g2_o21ai_1 _19806_ (.B1(_03792_),
    .Y(_02494_),
    .A1(net6663),
    .A2(net7618));
 sg13g2_nand2_1 _19807_ (.Y(_03793_),
    .A(net2579),
    .B(net7029));
 sg13g2_o21ai_1 _19808_ (.B1(_03793_),
    .Y(_02495_),
    .A1(net7029),
    .A2(net7168));
 sg13g2_nand2_1 _19809_ (.Y(_03794_),
    .A(net3130),
    .B(net7029));
 sg13g2_o21ai_1 _19810_ (.B1(_03794_),
    .Y(_02496_),
    .A1(net7029),
    .A2(net7463));
 sg13g2_nand2_1 _19811_ (.Y(_03795_),
    .A(net3046),
    .B(net7028));
 sg13g2_o21ai_1 _19812_ (.B1(_03795_),
    .Y(_02497_),
    .A1(net7028),
    .A2(net7623));
 sg13g2_nand2_1 _19813_ (.Y(_03796_),
    .A(net2531),
    .B(net7030));
 sg13g2_o21ai_1 _19814_ (.B1(_03796_),
    .Y(_02498_),
    .A1(net7030),
    .A2(net7164));
 sg13g2_nand2_1 _19815_ (.Y(_03797_),
    .A(net3454),
    .B(net7030));
 sg13g2_o21ai_1 _19816_ (.B1(_03797_),
    .Y(_02499_),
    .A1(net7030),
    .A2(net7458));
 sg13g2_nand2_1 _19817_ (.Y(_03798_),
    .A(net3939),
    .B(net7030));
 sg13g2_o21ai_1 _19818_ (.B1(_03798_),
    .Y(_02500_),
    .A1(net7030),
    .A2(net7619));
 sg13g2_nand2_1 _19819_ (.Y(_03799_),
    .A(net2798),
    .B(net7033));
 sg13g2_o21ai_1 _19820_ (.B1(_03799_),
    .Y(_02501_),
    .A1(net7033),
    .A2(net7168));
 sg13g2_nand2_1 _19821_ (.Y(_03800_),
    .A(net3717),
    .B(net7032));
 sg13g2_o21ai_1 _19822_ (.B1(_03800_),
    .Y(_02502_),
    .A1(net7032),
    .A2(net7463));
 sg13g2_nand2_1 _19823_ (.Y(_03801_),
    .A(net3167),
    .B(net7032));
 sg13g2_o21ai_1 _19824_ (.B1(_03801_),
    .Y(_02503_),
    .A1(net7032),
    .A2(net7623));
 sg13g2_nand2_1 _19825_ (.Y(_03802_),
    .A(net2746),
    .B(net7035));
 sg13g2_o21ai_1 _19826_ (.B1(_03802_),
    .Y(_02504_),
    .A1(net7035),
    .A2(net7168));
 sg13g2_nand2_1 _19827_ (.Y(_03803_),
    .A(net2897),
    .B(net7034));
 sg13g2_o21ai_1 _19828_ (.B1(_03803_),
    .Y(_02505_),
    .A1(net7034),
    .A2(net7463));
 sg13g2_nand2_1 _19829_ (.Y(_03804_),
    .A(net3085),
    .B(net7035));
 sg13g2_o21ai_1 _19830_ (.B1(_03804_),
    .Y(_02506_),
    .A1(net7034),
    .A2(net7623));
 sg13g2_nand2_1 _19831_ (.Y(_03805_),
    .A(net3340),
    .B(net7037));
 sg13g2_o21ai_1 _19832_ (.B1(_03805_),
    .Y(_02507_),
    .A1(net7037),
    .A2(net7147));
 sg13g2_nand2_1 _19833_ (.Y(_03806_),
    .A(net2846),
    .B(net7037));
 sg13g2_o21ai_1 _19834_ (.B1(_03806_),
    .Y(_02508_),
    .A1(net7037),
    .A2(net7447));
 sg13g2_nand2_1 _19835_ (.Y(_03807_),
    .A(net2984),
    .B(net7036));
 sg13g2_o21ai_1 _19836_ (.B1(_03807_),
    .Y(_02509_),
    .A1(net7036),
    .A2(net7600));
 sg13g2_nand2_1 _19837_ (.Y(_03808_),
    .A(net2724),
    .B(net7038));
 sg13g2_o21ai_1 _19838_ (.B1(_03808_),
    .Y(_02510_),
    .A1(net7038),
    .A2(net7147));
 sg13g2_nand2_1 _19839_ (.Y(_03809_),
    .A(net4499),
    .B(net7039));
 sg13g2_o21ai_1 _19840_ (.B1(_03809_),
    .Y(_02511_),
    .A1(net7039),
    .A2(net7438));
 sg13g2_nand2_1 _19841_ (.Y(_03810_),
    .A(net2754),
    .B(net7038));
 sg13g2_o21ai_1 _19842_ (.B1(_03810_),
    .Y(_02512_),
    .A1(net7038),
    .A2(net7600));
 sg13g2_nand2_1 _19843_ (.Y(_03811_),
    .A(net3297),
    .B(net7040));
 sg13g2_o21ai_1 _19844_ (.B1(_03811_),
    .Y(_02513_),
    .A1(net7040),
    .A2(net7145));
 sg13g2_nand2_1 _19845_ (.Y(_03812_),
    .A(net3375),
    .B(net7041));
 sg13g2_o21ai_1 _19846_ (.B1(_03812_),
    .Y(_02514_),
    .A1(net7040),
    .A2(net7438));
 sg13g2_nand2_1 _19847_ (.Y(_03813_),
    .A(net3109),
    .B(net7040));
 sg13g2_o21ai_1 _19848_ (.B1(_03813_),
    .Y(_02515_),
    .A1(net7040),
    .A2(net7600));
 sg13g2_nand2_1 _19849_ (.Y(_03814_),
    .A(net2453),
    .B(net7110));
 sg13g2_o21ai_1 _19850_ (.B1(_03814_),
    .Y(_02516_),
    .A1(net7110),
    .A2(net7145));
 sg13g2_nand2_1 _19851_ (.Y(_03815_),
    .A(net3602),
    .B(net7110));
 sg13g2_o21ai_1 _19852_ (.B1(_03815_),
    .Y(_02517_),
    .A1(net7110),
    .A2(net7438));
 sg13g2_nand2_1 _19853_ (.Y(_03816_),
    .A(net3260),
    .B(net7110));
 sg13g2_o21ai_1 _19854_ (.B1(_03816_),
    .Y(_02518_),
    .A1(net7110),
    .A2(net7600));
 sg13g2_nand2_1 _19855_ (.Y(_03817_),
    .A(net3743),
    .B(net7105));
 sg13g2_o21ai_1 _19856_ (.B1(_03817_),
    .Y(_02519_),
    .A1(net7105),
    .A2(net7145));
 sg13g2_nand2_1 _19857_ (.Y(_03818_),
    .A(net3571),
    .B(net7106));
 sg13g2_o21ai_1 _19858_ (.B1(_03818_),
    .Y(_02520_),
    .A1(net7105),
    .A2(net7438));
 sg13g2_nand2_1 _19859_ (.Y(_03819_),
    .A(net3761),
    .B(net7105));
 sg13g2_o21ai_1 _19860_ (.B1(_03819_),
    .Y(_02521_),
    .A1(net7105),
    .A2(net7600));
 sg13g2_nand2_1 _19861_ (.Y(_03820_),
    .A(net3325),
    .B(net7112));
 sg13g2_o21ai_1 _19862_ (.B1(_03820_),
    .Y(_02522_),
    .A1(net7112),
    .A2(net7145));
 sg13g2_nand2_1 _19863_ (.Y(_03821_),
    .A(net3674),
    .B(net7112));
 sg13g2_o21ai_1 _19864_ (.B1(_03821_),
    .Y(_02523_),
    .A1(net7112),
    .A2(net7438));
 sg13g2_nand2_1 _19865_ (.Y(_03822_),
    .A(net2999),
    .B(net7112));
 sg13g2_o21ai_1 _19866_ (.B1(_03822_),
    .Y(_02524_),
    .A1(net7112),
    .A2(net7600));
 sg13g2_nand2_1 _19867_ (.Y(_03823_),
    .A(net3479),
    .B(net7108));
 sg13g2_o21ai_1 _19868_ (.B1(_03823_),
    .Y(_02525_),
    .A1(net7108),
    .A2(net7145));
 sg13g2_nand2_1 _19869_ (.Y(_03824_),
    .A(net4188),
    .B(net7108));
 sg13g2_o21ai_1 _19870_ (.B1(_03824_),
    .Y(_02526_),
    .A1(net7108),
    .A2(net7438));
 sg13g2_nand2_1 _19871_ (.Y(_03825_),
    .A(net3272),
    .B(net7108));
 sg13g2_o21ai_1 _19872_ (.B1(_03825_),
    .Y(_02527_),
    .A1(net7108),
    .A2(net7600));
 sg13g2_dfrbp_1 _19873_ (.CLK(\clknet_leaf_40_top1.acquisition_clk ),
    .RESET_B(net904),
    .D(_00074_),
    .Q_N(_09905_),
    .Q(\top1.memory1.mem2[197][0] ));
 sg13g2_dfrbp_1 _19874_ (.CLK(\clknet_leaf_38_top1.acquisition_clk ),
    .RESET_B(net1304),
    .D(_00075_),
    .Q_N(_09904_),
    .Q(\top1.memory1.mem2[197][1] ));
 sg13g2_dfrbp_1 _19875_ (.CLK(\clknet_leaf_41_top1.acquisition_clk ),
    .RESET_B(net1303),
    .D(_00076_),
    .Q_N(_09903_),
    .Q(\top1.memory1.mem2[197][2] ));
 sg13g2_dfrbp_1 _19876_ (.CLK(\clknet_leaf_96_top1.acquisition_clk ),
    .RESET_B(net1302),
    .D(_00077_),
    .Q_N(_09902_),
    .Q(\top1.memory1.mem2[195][0] ));
 sg13g2_dfrbp_1 _19877_ (.CLK(\clknet_leaf_96_top1.acquisition_clk ),
    .RESET_B(net1301),
    .D(_00078_),
    .Q_N(_09901_),
    .Q(\top1.memory1.mem2[195][1] ));
 sg13g2_dfrbp_1 _19878_ (.CLK(\clknet_leaf_97_top1.acquisition_clk ),
    .RESET_B(net1300),
    .D(_00079_),
    .Q_N(_09900_),
    .Q(\top1.memory1.mem2[195][2] ));
 sg13g2_dfrbp_1 _19879_ (.CLK(\clknet_leaf_99_top1.acquisition_clk ),
    .RESET_B(net1299),
    .D(_00080_),
    .Q_N(_09899_),
    .Q(\top1.memory1.mem2[198][0] ));
 sg13g2_dfrbp_1 _19880_ (.CLK(\clknet_leaf_41_top1.acquisition_clk ),
    .RESET_B(net1298),
    .D(_00081_),
    .Q_N(_09898_),
    .Q(\top1.memory1.mem2[198][1] ));
 sg13g2_dfrbp_1 _19881_ (.CLK(\clknet_leaf_99_top1.acquisition_clk ),
    .RESET_B(net1297),
    .D(_00082_),
    .Q_N(_09897_),
    .Q(\top1.memory1.mem2[198][2] ));
 sg13g2_dfrbp_1 _19882_ (.CLK(\clknet_leaf_40_top1.acquisition_clk ),
    .RESET_B(net1296),
    .D(_00083_),
    .Q_N(_09896_),
    .Q(\top1.memory1.mem2[196][0] ));
 sg13g2_dfrbp_1 _19883_ (.CLK(\clknet_leaf_38_top1.acquisition_clk ),
    .RESET_B(net1295),
    .D(_00084_),
    .Q_N(_09895_),
    .Q(\top1.memory1.mem2[196][1] ));
 sg13g2_dfrbp_1 _19884_ (.CLK(\clknet_leaf_38_top1.acquisition_clk ),
    .RESET_B(net1294),
    .D(_00085_),
    .Q_N(_09894_),
    .Q(\top1.memory1.mem2[196][2] ));
 sg13g2_dfrbp_1 _19885_ (.CLK(\clknet_leaf_211_top1.acquisition_clk ),
    .RESET_B(net1293),
    .D(_00086_),
    .Q_N(_09893_),
    .Q(\top1.memory1.mem2[122][0] ));
 sg13g2_dfrbp_1 _19886_ (.CLK(\clknet_leaf_211_top1.acquisition_clk ),
    .RESET_B(net1292),
    .D(_00087_),
    .Q_N(_09892_),
    .Q(\top1.memory1.mem2[122][1] ));
 sg13g2_dfrbp_1 _19887_ (.CLK(\clknet_leaf_209_top1.acquisition_clk ),
    .RESET_B(net1291),
    .D(_00088_),
    .Q_N(_09891_),
    .Q(\top1.memory1.mem2[122][2] ));
 sg13g2_dfrbp_1 _19888_ (.CLK(\clknet_leaf_252_top1.acquisition_clk ),
    .RESET_B(net1290),
    .D(_00089_),
    .Q_N(_09890_),
    .Q(\top1.memory1.mem2[97][0] ));
 sg13g2_dfrbp_1 _19889_ (.CLK(\clknet_leaf_251_top1.acquisition_clk ),
    .RESET_B(net1289),
    .D(_00090_),
    .Q_N(_09889_),
    .Q(\top1.memory1.mem2[97][1] ));
 sg13g2_dfrbp_1 _19890_ (.CLK(\clknet_leaf_250_top1.acquisition_clk ),
    .RESET_B(net1288),
    .D(_00091_),
    .Q_N(_09888_),
    .Q(\top1.memory1.mem2[97][2] ));
 sg13g2_dfrbp_1 _19891_ (.CLK(\clknet_leaf_293_top1.acquisition_clk ),
    .RESET_B(net1287),
    .D(_00092_),
    .Q_N(_09887_),
    .Q(\top1.memory1.mem2[82][0] ));
 sg13g2_dfrbp_1 _19892_ (.CLK(\clknet_leaf_296_top1.acquisition_clk ),
    .RESET_B(net1286),
    .D(_00093_),
    .Q_N(_09886_),
    .Q(\top1.memory1.mem2[82][1] ));
 sg13g2_dfrbp_1 _19893_ (.CLK(\clknet_leaf_295_top1.acquisition_clk ),
    .RESET_B(net1285),
    .D(_00094_),
    .Q_N(_09885_),
    .Q(\top1.memory1.mem2[82][2] ));
 sg13g2_dfrbp_1 _19894_ (.CLK(\clknet_leaf_294_top1.acquisition_clk ),
    .RESET_B(net1284),
    .D(_00095_),
    .Q_N(_09884_),
    .Q(\top1.memory1.mem2[81][0] ));
 sg13g2_dfrbp_1 _19895_ (.CLK(\clknet_leaf_296_top1.acquisition_clk ),
    .RESET_B(net1283),
    .D(_00096_),
    .Q_N(_09883_),
    .Q(\top1.memory1.mem2[81][1] ));
 sg13g2_dfrbp_1 _19896_ (.CLK(\clknet_leaf_295_top1.acquisition_clk ),
    .RESET_B(net1282),
    .D(_00097_),
    .Q_N(_09882_),
    .Q(\top1.memory1.mem2[81][2] ));
 sg13g2_dfrbp_1 _19897_ (.CLK(\clknet_leaf_88_top1.acquisition_clk ),
    .RESET_B(net1281),
    .D(_00098_),
    .Q_N(_09881_),
    .Q(\top1.memory1.mem2[1][0] ));
 sg13g2_dfrbp_1 _19898_ (.CLK(\clknet_leaf_85_top1.acquisition_clk ),
    .RESET_B(net1280),
    .D(_00099_),
    .Q_N(_09880_),
    .Q(\top1.memory1.mem2[1][1] ));
 sg13g2_dfrbp_1 _19899_ (.CLK(\clknet_leaf_91_top1.acquisition_clk ),
    .RESET_B(net1279),
    .D(_00100_),
    .Q_N(_09879_),
    .Q(\top1.memory1.mem2[1][2] ));
 sg13g2_dfrbp_1 _19900_ (.CLK(\clknet_leaf_40_top1.acquisition_clk ),
    .RESET_B(net1278),
    .D(_00101_),
    .Q_N(_09878_),
    .Q(\top1.memory1.mem2[199][0] ));
 sg13g2_dfrbp_1 _19901_ (.CLK(\clknet_leaf_41_top1.acquisition_clk ),
    .RESET_B(net1277),
    .D(_00102_),
    .Q_N(_09877_),
    .Q(\top1.memory1.mem2[199][1] ));
 sg13g2_dfrbp_1 _19902_ (.CLK(\clknet_leaf_41_top1.acquisition_clk ),
    .RESET_B(net1276),
    .D(_00103_),
    .Q_N(_09876_),
    .Q(\top1.memory1.mem2[199][2] ));
 sg13g2_dfrbp_1 _19903_ (.CLK(\clknet_leaf_117_top1.acquisition_clk ),
    .RESET_B(net1275),
    .D(_00104_),
    .Q_N(_09875_),
    .Q(\top1.memory1.mem2[189][0] ));
 sg13g2_dfrbp_1 _19904_ (.CLK(\clknet_leaf_118_top1.acquisition_clk ),
    .RESET_B(net1274),
    .D(_00105_),
    .Q_N(_09874_),
    .Q(\top1.memory1.mem2[189][1] ));
 sg13g2_dfrbp_1 _19905_ (.CLK(\clknet_leaf_115_top1.acquisition_clk ),
    .RESET_B(net1273),
    .D(_00106_),
    .Q_N(_09873_),
    .Q(\top1.memory1.mem2[189][2] ));
 sg13g2_dfrbp_1 _19906_ (.CLK(\clknet_leaf_135_top1.acquisition_clk ),
    .RESET_B(net1272),
    .D(_00107_),
    .Q_N(_09872_),
    .Q(\top1.memory1.mem2[179][0] ));
 sg13g2_dfrbp_1 _19907_ (.CLK(\clknet_leaf_129_top1.acquisition_clk ),
    .RESET_B(net1271),
    .D(_00108_),
    .Q_N(_09871_),
    .Q(\top1.memory1.mem2[179][1] ));
 sg13g2_dfrbp_1 _19908_ (.CLK(\clknet_leaf_130_top1.acquisition_clk ),
    .RESET_B(net1270),
    .D(_00109_),
    .Q_N(_09870_),
    .Q(\top1.memory1.mem2[179][2] ));
 sg13g2_dfrbp_1 _19909_ (.CLK(\clknet_leaf_105_top1.acquisition_clk ),
    .RESET_B(net1269),
    .D(_00110_),
    .Q_N(_09869_),
    .Q(\top1.memory1.mem2[169][0] ));
 sg13g2_dfrbp_1 _19910_ (.CLK(\clknet_leaf_106_top1.acquisition_clk ),
    .RESET_B(net1268),
    .D(_00111_),
    .Q_N(_09868_),
    .Q(\top1.memory1.mem2[169][1] ));
 sg13g2_dfrbp_1 _19911_ (.CLK(\clknet_leaf_107_top1.acquisition_clk ),
    .RESET_B(net1267),
    .D(_00112_),
    .Q_N(_09867_),
    .Q(\top1.memory1.mem2[169][2] ));
 sg13g2_dfrbp_1 _19912_ (.CLK(\clknet_leaf_117_top1.acquisition_clk ),
    .RESET_B(net1266),
    .D(_00113_),
    .Q_N(_09866_),
    .Q(\top1.memory1.mem2[36][0] ));
 sg13g2_dfrbp_1 _19913_ (.CLK(\clknet_leaf_133_top1.acquisition_clk ),
    .RESET_B(net1265),
    .D(_00114_),
    .Q_N(_09865_),
    .Q(\top1.memory1.mem2[36][1] ));
 sg13g2_dfrbp_1 _19914_ (.CLK(\clknet_leaf_131_top1.acquisition_clk ),
    .RESET_B(net1264),
    .D(_00115_),
    .Q_N(_09864_),
    .Q(\top1.memory1.mem2[36][2] ));
 sg13g2_dfrbp_1 _19915_ (.CLK(\clknet_leaf_73_top1.acquisition_clk ),
    .RESET_B(net1263),
    .D(_00116_),
    .Q_N(_09863_),
    .Q(\top1.memory1.mem2[159][0] ));
 sg13g2_dfrbp_1 _19916_ (.CLK(\clknet_leaf_73_top1.acquisition_clk ),
    .RESET_B(net1262),
    .D(_00117_),
    .Q_N(_09862_),
    .Q(\top1.memory1.mem2[159][1] ));
 sg13g2_dfrbp_1 _19917_ (.CLK(\clknet_leaf_81_top1.acquisition_clk ),
    .RESET_B(net1261),
    .D(_00118_),
    .Q_N(_09861_),
    .Q(\top1.memory1.mem2[159][2] ));
 sg13g2_dfrbp_1 _19918_ (.CLK(\clknet_leaf_178_top1.acquisition_clk ),
    .RESET_B(net1260),
    .D(_00119_),
    .Q_N(_09860_),
    .Q(\top1.memory1.mem2[35][0] ));
 sg13g2_dfrbp_1 _19919_ (.CLK(\clknet_leaf_177_top1.acquisition_clk ),
    .RESET_B(net1259),
    .D(_00120_),
    .Q_N(_09859_),
    .Q(\top1.memory1.mem2[35][1] ));
 sg13g2_dfrbp_1 _19920_ (.CLK(\clknet_leaf_175_top1.acquisition_clk ),
    .RESET_B(net1258),
    .D(_00121_),
    .Q_N(_09858_),
    .Q(\top1.memory1.mem2[35][2] ));
 sg13g2_dfrbp_1 _19921_ (.CLK(\clknet_leaf_43_top1.acquisition_clk ),
    .RESET_B(net1257),
    .D(_00122_),
    .Q_N(_09857_),
    .Q(\top1.memory1.mem2[149][0] ));
 sg13g2_dfrbp_1 _19922_ (.CLK(\clknet_leaf_77_top1.acquisition_clk ),
    .RESET_B(net1256),
    .D(_00123_),
    .Q_N(_09856_),
    .Q(\top1.memory1.mem2[149][1] ));
 sg13g2_dfrbp_1 _19923_ (.CLK(\clknet_leaf_97_top1.acquisition_clk ),
    .RESET_B(net1255),
    .D(_00124_),
    .Q_N(_09855_),
    .Q(\top1.memory1.mem2[149][2] ));
 sg13g2_dfrbp_1 _19924_ (.CLK(\clknet_leaf_178_top1.acquisition_clk ),
    .RESET_B(net1254),
    .D(_00125_),
    .Q_N(_09854_),
    .Q(\top1.memory1.mem2[34][0] ));
 sg13g2_dfrbp_1 _19925_ (.CLK(\clknet_leaf_179_top1.acquisition_clk ),
    .RESET_B(net1253),
    .D(_00126_),
    .Q_N(_09853_),
    .Q(\top1.memory1.mem2[34][1] ));
 sg13g2_dfrbp_1 _19926_ (.CLK(\clknet_leaf_176_top1.acquisition_clk ),
    .RESET_B(net1252),
    .D(_00127_),
    .Q_N(_09852_),
    .Q(\top1.memory1.mem2[34][2] ));
 sg13g2_dfrbp_1 _19927_ (.CLK(\clknet_leaf_69_top1.acquisition_clk ),
    .RESET_B(net1251),
    .D(_00128_),
    .Q_N(_09851_),
    .Q(\top1.memory1.mem2[139][0] ));
 sg13g2_dfrbp_1 _19928_ (.CLK(\clknet_leaf_69_top1.acquisition_clk ),
    .RESET_B(net1250),
    .D(_00129_),
    .Q_N(_09850_),
    .Q(\top1.memory1.mem2[139][1] ));
 sg13g2_dfrbp_1 _19929_ (.CLK(\clknet_leaf_68_top1.acquisition_clk ),
    .RESET_B(net1249),
    .D(_00130_),
    .Q_N(_09849_),
    .Q(\top1.memory1.mem2[139][2] ));
 sg13g2_dfrbp_1 _19930_ (.CLK(\clknet_leaf_178_top1.acquisition_clk ),
    .RESET_B(net1248),
    .D(_00131_),
    .Q_N(_09848_),
    .Q(\top1.memory1.mem2[33][0] ));
 sg13g2_dfrbp_1 _19931_ (.CLK(\clknet_leaf_179_top1.acquisition_clk ),
    .RESET_B(net1247),
    .D(_00132_),
    .Q_N(_09847_),
    .Q(\top1.memory1.mem2[33][1] ));
 sg13g2_dfrbp_1 _19932_ (.CLK(\clknet_leaf_175_top1.acquisition_clk ),
    .RESET_B(net1246),
    .D(_00133_),
    .Q_N(_09846_),
    .Q(\top1.memory1.mem2[33][2] ));
 sg13g2_dfrbp_1 _19933_ (.CLK(\clknet_leaf_65_top1.acquisition_clk ),
    .RESET_B(net1245),
    .D(_00134_),
    .Q_N(_09845_),
    .Q(\top1.memory1.mem2[129][0] ));
 sg13g2_dfrbp_1 _19934_ (.CLK(\clknet_leaf_64_top1.acquisition_clk ),
    .RESET_B(net1244),
    .D(_00135_),
    .Q_N(_09844_),
    .Q(\top1.memory1.mem2[129][1] ));
 sg13g2_dfrbp_1 _19935_ (.CLK(\clknet_leaf_64_top1.acquisition_clk ),
    .RESET_B(net1243),
    .D(_00136_),
    .Q_N(_09843_),
    .Q(\top1.memory1.mem2[129][2] ));
 sg13g2_dfrbp_1 _19936_ (.CLK(\clknet_leaf_178_top1.acquisition_clk ),
    .RESET_B(net1242),
    .D(_00137_),
    .Q_N(_09842_),
    .Q(\top1.memory1.mem2[32][0] ));
 sg13g2_dfrbp_1 _19937_ (.CLK(\clknet_leaf_179_top1.acquisition_clk ),
    .RESET_B(net1241),
    .D(_00138_),
    .Q_N(_09841_),
    .Q(\top1.memory1.mem2[32][1] ));
 sg13g2_dfrbp_1 _19938_ (.CLK(\clknet_leaf_175_top1.acquisition_clk ),
    .RESET_B(net1240),
    .D(_00139_),
    .Q_N(_09840_),
    .Q(\top1.memory1.mem2[32][2] ));
 sg13g2_dfrbp_1 _19939_ (.CLK(\clknet_leaf_222_top1.acquisition_clk ),
    .RESET_B(net1238),
    .D(_00140_),
    .Q_N(_09839_),
    .Q(\top1.memory1.mem2[119][0] ));
 sg13g2_dfrbp_1 _19940_ (.CLK(\clknet_leaf_213_top1.acquisition_clk ),
    .RESET_B(net1237),
    .D(_00141_),
    .Q_N(_09838_),
    .Q(\top1.memory1.mem2[119][1] ));
 sg13g2_dfrbp_1 _19941_ (.CLK(\clknet_leaf_223_top1.acquisition_clk ),
    .RESET_B(net1236),
    .D(_00142_),
    .Q_N(_09837_),
    .Q(\top1.memory1.mem2[119][2] ));
 sg13g2_dfrbp_1 _19942_ (.CLK(\clknet_leaf_122_top1.acquisition_clk ),
    .RESET_B(net1235),
    .D(_00143_),
    .Q_N(_09836_),
    .Q(\top1.memory1.mem2[31][0] ));
 sg13g2_dfrbp_1 _19943_ (.CLK(\clknet_leaf_92_top1.acquisition_clk ),
    .RESET_B(net1234),
    .D(_00144_),
    .Q_N(_09835_),
    .Q(\top1.memory1.mem2[31][1] ));
 sg13g2_dfrbp_1 _19944_ (.CLK(\clknet_leaf_88_top1.acquisition_clk ),
    .RESET_B(net1233),
    .D(_00145_),
    .Q_N(_09834_),
    .Q(\top1.memory1.mem2[31][2] ));
 sg13g2_dfrbp_1 _19945_ (.CLK(\clknet_leaf_226_top1.acquisition_clk ),
    .RESET_B(net1232),
    .D(_00146_),
    .Q_N(_09833_),
    .Q(\top1.memory1.mem2[109][0] ));
 sg13g2_dfrbp_1 _19946_ (.CLK(\clknet_leaf_234_top1.acquisition_clk ),
    .RESET_B(net1231),
    .D(_00147_),
    .Q_N(_09832_),
    .Q(\top1.memory1.mem2[109][1] ));
 sg13g2_dfrbp_1 _19947_ (.CLK(\clknet_leaf_225_top1.acquisition_clk ),
    .RESET_B(net1230),
    .D(_00148_),
    .Q_N(_09831_),
    .Q(\top1.memory1.mem2[109][2] ));
 sg13g2_dfrbp_1 _19948_ (.CLK(\clknet_leaf_122_top1.acquisition_clk ),
    .RESET_B(net1229),
    .D(_00149_),
    .Q_N(_09830_),
    .Q(\top1.memory1.mem2[30][0] ));
 sg13g2_dfrbp_1 _19949_ (.CLK(\clknet_leaf_88_top1.acquisition_clk ),
    .RESET_B(net1228),
    .D(_00150_),
    .Q_N(_09829_),
    .Q(\top1.memory1.mem2[30][1] ));
 sg13g2_dfrbp_1 _19950_ (.CLK(\clknet_leaf_88_top1.acquisition_clk ),
    .RESET_B(net1227),
    .D(_00151_),
    .Q_N(_09828_),
    .Q(\top1.memory1.mem2[30][2] ));
 sg13g2_dfrbp_1 _19951_ (.CLK(\clknet_leaf_251_top1.acquisition_clk ),
    .RESET_B(net1226),
    .D(_00152_),
    .Q_N(_09827_),
    .Q(\top1.memory1.mem2[99][0] ));
 sg13g2_dfrbp_1 _19952_ (.CLK(\clknet_leaf_251_top1.acquisition_clk ),
    .RESET_B(net1225),
    .D(_00153_),
    .Q_N(_09826_),
    .Q(\top1.memory1.mem2[99][1] ));
 sg13g2_dfrbp_1 _19953_ (.CLK(\clknet_leaf_251_top1.acquisition_clk ),
    .RESET_B(net1224),
    .D(_00154_),
    .Q_N(_09825_),
    .Q(\top1.memory1.mem2[99][2] ));
 sg13g2_dfrbp_1 _19954_ (.CLK(\clknet_leaf_87_top1.acquisition_clk ),
    .RESET_B(net1223),
    .D(_00155_),
    .Q_N(_09824_),
    .Q(\top1.memory1.mem2[2][0] ));
 sg13g2_dfrbp_1 _19955_ (.CLK(\clknet_leaf_89_top1.acquisition_clk ),
    .RESET_B(net1222),
    .D(_00156_),
    .Q_N(_09823_),
    .Q(\top1.memory1.mem2[2][1] ));
 sg13g2_dfrbp_1 _19956_ (.CLK(\clknet_leaf_91_top1.acquisition_clk ),
    .RESET_B(net1221),
    .D(_00157_),
    .Q_N(_09822_),
    .Q(\top1.memory1.mem2[2][2] ));
 sg13g2_dfrbp_1 _19957_ (.CLK(\clknet_leaf_9_top1.acquisition_clk ),
    .RESET_B(net1220),
    .D(_00158_),
    .Q_N(_09821_),
    .Q(\top1.memory1.mem2[89][0] ));
 sg13g2_dfrbp_1 _19958_ (.CLK(\clknet_leaf_292_top1.acquisition_clk ),
    .RESET_B(net1219),
    .D(_00159_),
    .Q_N(_09820_),
    .Q(\top1.memory1.mem2[89][1] ));
 sg13g2_dfrbp_1 _19959_ (.CLK(\clknet_leaf_28_top1.acquisition_clk ),
    .RESET_B(net1218),
    .D(_00160_),
    .Q_N(_09819_),
    .Q(\top1.memory1.mem2[89][2] ));
 sg13g2_dfrbp_1 _19960_ (.CLK(\clknet_leaf_124_top1.acquisition_clk ),
    .RESET_B(net1217),
    .D(_00161_),
    .Q_N(_09818_),
    .Q(\top1.memory1.mem2[28][0] ));
 sg13g2_dfrbp_1 _19961_ (.CLK(\clknet_leaf_88_top1.acquisition_clk ),
    .RESET_B(net1216),
    .D(_00162_),
    .Q_N(_09817_),
    .Q(\top1.memory1.mem2[28][1] ));
 sg13g2_dfrbp_1 _19962_ (.CLK(\clknet_leaf_88_top1.acquisition_clk ),
    .RESET_B(net1215),
    .D(_00163_),
    .Q_N(_09816_),
    .Q(\top1.memory1.mem2[28][2] ));
 sg13g2_dfrbp_1 _19963_ (.CLK(\clknet_leaf_3_top1.acquisition_clk ),
    .RESET_B(net1214),
    .D(_00164_),
    .Q_N(_09815_),
    .Q(\top1.memory1.mem2[79][0] ));
 sg13g2_dfrbp_1 _19964_ (.CLK(\clknet_leaf_2_top1.acquisition_clk ),
    .RESET_B(net1213),
    .D(_00165_),
    .Q_N(_09814_),
    .Q(\top1.memory1.mem2[79][1] ));
 sg13g2_dfrbp_1 _19965_ (.CLK(\clknet_leaf_3_top1.acquisition_clk ),
    .RESET_B(net1212),
    .D(_00166_),
    .Q_N(_09813_),
    .Q(\top1.memory1.mem2[79][2] ));
 sg13g2_dfrbp_1 _19966_ (.CLK(\clknet_leaf_126_top1.acquisition_clk ),
    .RESET_B(net1211),
    .D(_00167_),
    .Q_N(_09812_),
    .Q(\top1.memory1.mem2[27][0] ));
 sg13g2_dfrbp_1 _19967_ (.CLK(\clknet_leaf_126_top1.acquisition_clk ),
    .RESET_B(net1210),
    .D(_00168_),
    .Q_N(_09811_),
    .Q(\top1.memory1.mem2[27][1] ));
 sg13g2_dfrbp_1 _19968_ (.CLK(\clknet_leaf_122_top1.acquisition_clk ),
    .RESET_B(net1209),
    .D(_00169_),
    .Q_N(_09810_),
    .Q(\top1.memory1.mem2[27][2] ));
 sg13g2_dfrbp_1 _19969_ (.CLK(\clknet_leaf_87_top1.acquisition_clk ),
    .RESET_B(net1208),
    .D(_00170_),
    .Q_N(_09809_),
    .Q(\top1.memory1.mem2[3][0] ));
 sg13g2_dfrbp_1 _19970_ (.CLK(\clknet_leaf_89_top1.acquisition_clk ),
    .RESET_B(net1207),
    .D(_00171_),
    .Q_N(_09808_),
    .Q(\top1.memory1.mem2[3][1] ));
 sg13g2_dfrbp_1 _19971_ (.CLK(\clknet_leaf_91_top1.acquisition_clk ),
    .RESET_B(net1206),
    .D(_00172_),
    .Q_N(_09807_),
    .Q(\top1.memory1.mem2[3][2] ));
 sg13g2_dfrbp_1 _19972_ (.CLK(\clknet_leaf_141_top1.acquisition_clk ),
    .RESET_B(net1205),
    .D(_00173_),
    .Q_N(_09806_),
    .Q(\top1.memory1.mem2[45][0] ));
 sg13g2_dfrbp_1 _19973_ (.CLK(\clknet_leaf_142_top1.acquisition_clk ),
    .RESET_B(net1204),
    .D(_00174_),
    .Q_N(_09805_),
    .Q(\top1.memory1.mem2[45][1] ));
 sg13g2_dfrbp_1 _19974_ (.CLK(\clknet_leaf_132_top1.acquisition_clk ),
    .RESET_B(net1203),
    .D(_00175_),
    .Q_N(_09804_),
    .Q(\top1.memory1.mem2[45][2] ));
 sg13g2_dfrbp_1 _19975_ (.CLK(\clknet_leaf_293_top1.acquisition_clk ),
    .RESET_B(net1202),
    .D(_00176_),
    .Q_N(_09803_),
    .Q(\top1.memory1.mem2[80][0] ));
 sg13g2_dfrbp_1 _19976_ (.CLK(\clknet_leaf_296_top1.acquisition_clk ),
    .RESET_B(net1201),
    .D(_00177_),
    .Q_N(_09802_),
    .Q(\top1.memory1.mem2[80][1] ));
 sg13g2_dfrbp_1 _19977_ (.CLK(\clknet_leaf_295_top1.acquisition_clk ),
    .RESET_B(net1200),
    .D(_00178_),
    .Q_N(_09801_),
    .Q(\top1.memory1.mem2[80][2] ));
 sg13g2_dfrbp_1 _19978_ (.CLK(\clknet_leaf_101_top1.acquisition_clk ),
    .RESET_B(net1199),
    .D(_00179_),
    .Q_N(_09800_),
    .Q(\top1.memory1.mem2[7][0] ));
 sg13g2_dfrbp_1 _19979_ (.CLK(\clknet_leaf_92_top1.acquisition_clk ),
    .RESET_B(net1198),
    .D(_00180_),
    .Q_N(_09799_),
    .Q(\top1.memory1.mem2[7][1] ));
 sg13g2_dfrbp_1 _19980_ (.CLK(\clknet_leaf_93_top1.acquisition_clk ),
    .RESET_B(net1197),
    .D(_00181_),
    .Q_N(_09798_),
    .Q(\top1.memory1.mem2[7][2] ));
 sg13g2_dfrbp_1 _19981_ (.CLK(\clknet_leaf_3_top1.acquisition_clk ),
    .RESET_B(net1196),
    .D(_00182_),
    .Q_N(_09797_),
    .Q(\top1.memory1.mem2[78][0] ));
 sg13g2_dfrbp_1 _19982_ (.CLK(\clknet_leaf_2_top1.acquisition_clk ),
    .RESET_B(net1195),
    .D(_00183_),
    .Q_N(_09796_),
    .Q(\top1.memory1.mem2[78][1] ));
 sg13g2_dfrbp_1 _19983_ (.CLK(\clknet_leaf_4_top1.acquisition_clk ),
    .RESET_B(net1194),
    .D(_00184_),
    .Q_N(_09795_),
    .Q(\top1.memory1.mem2[78][2] ));
 sg13g2_dfrbp_1 _19984_ (.CLK(\clknet_leaf_3_top1.acquisition_clk ),
    .RESET_B(net1193),
    .D(_00185_),
    .Q_N(_09794_),
    .Q(\top1.memory1.mem2[77][0] ));
 sg13g2_dfrbp_1 _19985_ (.CLK(\clknet_leaf_0_top1.acquisition_clk ),
    .RESET_B(net1192),
    .D(_00186_),
    .Q_N(_09793_),
    .Q(\top1.memory1.mem2[77][1] ));
 sg13g2_dfrbp_1 _19986_ (.CLK(\clknet_leaf_4_top1.acquisition_clk ),
    .RESET_B(net1191),
    .D(_00187_),
    .Q_N(_09792_),
    .Q(\top1.memory1.mem2[77][2] ));
 sg13g2_dfrbp_1 _19987_ (.CLK(\clknet_leaf_3_top1.acquisition_clk ),
    .RESET_B(net1190),
    .D(_00188_),
    .Q_N(_09791_),
    .Q(\top1.memory1.mem2[76][0] ));
 sg13g2_dfrbp_1 _19988_ (.CLK(\clknet_leaf_3_top1.acquisition_clk ),
    .RESET_B(net1189),
    .D(_00189_),
    .Q_N(_09790_),
    .Q(\top1.memory1.mem2[76][1] ));
 sg13g2_dfrbp_1 _19989_ (.CLK(\clknet_leaf_3_top1.acquisition_clk ),
    .RESET_B(net1188),
    .D(_00190_),
    .Q_N(_09789_),
    .Q(\top1.memory1.mem2[76][2] ));
 sg13g2_dfrbp_1 _19990_ (.CLK(\clknet_leaf_297_top1.acquisition_clk ),
    .RESET_B(net1187),
    .D(_00191_),
    .Q_N(_09788_),
    .Q(\top1.memory1.mem2[75][0] ));
 sg13g2_dfrbp_1 _19991_ (.CLK(\clknet_leaf_298_top1.acquisition_clk ),
    .RESET_B(net1186),
    .D(_00192_),
    .Q_N(_09787_),
    .Q(\top1.memory1.mem2[75][1] ));
 sg13g2_dfrbp_1 _19992_ (.CLK(\clknet_leaf_292_top1.acquisition_clk ),
    .RESET_B(net1185),
    .D(_00193_),
    .Q_N(_09786_),
    .Q(\top1.memory1.mem2[75][2] ));
 sg13g2_dfrbp_1 _19993_ (.CLK(\clknet_leaf_298_top1.acquisition_clk ),
    .RESET_B(net1184),
    .D(_00194_),
    .Q_N(_09785_),
    .Q(\top1.memory1.mem2[74][0] ));
 sg13g2_dfrbp_1 _19994_ (.CLK(\clknet_leaf_298_top1.acquisition_clk ),
    .RESET_B(net1183),
    .D(_00195_),
    .Q_N(_09784_),
    .Q(\top1.memory1.mem2[74][1] ));
 sg13g2_dfrbp_1 _19995_ (.CLK(\clknet_leaf_298_top1.acquisition_clk ),
    .RESET_B(net1182),
    .D(_00196_),
    .Q_N(_09783_),
    .Q(\top1.memory1.mem2[74][2] ));
 sg13g2_dfrbp_1 _19996_ (.CLK(\clknet_leaf_298_top1.acquisition_clk ),
    .RESET_B(net1181),
    .D(_00197_),
    .Q_N(_09782_),
    .Q(\top1.memory1.mem2[73][0] ));
 sg13g2_dfrbp_1 _19997_ (.CLK(\clknet_leaf_6_top1.acquisition_clk ),
    .RESET_B(net1180),
    .D(_00198_),
    .Q_N(_09781_),
    .Q(\top1.memory1.mem2[73][1] ));
 sg13g2_dfrbp_1 _19998_ (.CLK(\clknet_leaf_6_top1.acquisition_clk ),
    .RESET_B(net1179),
    .D(_00199_),
    .Q_N(_09780_),
    .Q(\top1.memory1.mem2[73][2] ));
 sg13g2_dfrbp_1 _19999_ (.CLK(\clknet_leaf_298_top1.acquisition_clk ),
    .RESET_B(net1178),
    .D(_00200_),
    .Q_N(_09779_),
    .Q(\top1.memory1.mem2[72][0] ));
 sg13g2_dfrbp_1 _20000_ (.CLK(\clknet_leaf_1_top1.acquisition_clk ),
    .RESET_B(net1177),
    .D(_00201_),
    .Q_N(_09778_),
    .Q(\top1.memory1.mem2[72][1] ));
 sg13g2_dfrbp_1 _20001_ (.CLK(\clknet_leaf_6_top1.acquisition_clk ),
    .RESET_B(net1176),
    .D(_00202_),
    .Q_N(_09777_),
    .Q(\top1.memory1.mem2[72][2] ));
 sg13g2_dfrbp_1 _20002_ (.CLK(\clknet_leaf_6_top1.acquisition_clk ),
    .RESET_B(net1175),
    .D(_00203_),
    .Q_N(_09776_),
    .Q(\top1.memory1.mem2[71][0] ));
 sg13g2_dfrbp_1 _20003_ (.CLK(\clknet_leaf_8_top1.acquisition_clk ),
    .RESET_B(net1174),
    .D(_00204_),
    .Q_N(_09775_),
    .Q(\top1.memory1.mem2[71][1] ));
 sg13g2_dfrbp_1 _20004_ (.CLK(\clknet_leaf_7_top1.acquisition_clk ),
    .RESET_B(net1173),
    .D(_00205_),
    .Q_N(_09774_),
    .Q(\top1.memory1.mem2[71][2] ));
 sg13g2_dfrbp_1 _20005_ (.CLK(\clknet_leaf_252_top1.acquisition_clk ),
    .RESET_B(net1172),
    .D(_00206_),
    .Q_N(_09773_),
    .Q(\top1.memory1.mem2[96][0] ));
 sg13g2_dfrbp_1 _20006_ (.CLK(\clknet_leaf_252_top1.acquisition_clk ),
    .RESET_B(net1171),
    .D(_00207_),
    .Q_N(_09772_),
    .Q(\top1.memory1.mem2[96][1] ));
 sg13g2_dfrbp_1 _20007_ (.CLK(\clknet_leaf_250_top1.acquisition_clk ),
    .RESET_B(net1170),
    .D(_00208_),
    .Q_N(_09771_),
    .Q(\top1.memory1.mem2[96][2] ));
 sg13g2_dfrbp_1 _20008_ (.CLK(\clknet_leaf_292_top1.acquisition_clk ),
    .RESET_B(net1169),
    .D(_00209_),
    .Q_N(_09770_),
    .Q(\top1.memory1.mem2[70][0] ));
 sg13g2_dfrbp_1 _20009_ (.CLK(\clknet_leaf_8_top1.acquisition_clk ),
    .RESET_B(net1168),
    .D(_00210_),
    .Q_N(_09769_),
    .Q(\top1.memory1.mem2[70][1] ));
 sg13g2_dfrbp_1 _20010_ (.CLK(\clknet_leaf_7_top1.acquisition_clk ),
    .RESET_B(net1167),
    .D(_00211_),
    .Q_N(_09768_),
    .Q(\top1.memory1.mem2[70][2] ));
 sg13g2_dfrbp_1 _20011_ (.CLK(\clknet_leaf_285_top1.acquisition_clk ),
    .RESET_B(net1166),
    .D(_00212_),
    .Q_N(_09767_),
    .Q(\top1.memory1.mem2[95][0] ));
 sg13g2_dfrbp_1 _20012_ (.CLK(\clknet_leaf_286_top1.acquisition_clk ),
    .RESET_B(net1165),
    .D(_00213_),
    .Q_N(_09766_),
    .Q(\top1.memory1.mem2[95][1] ));
 sg13g2_dfrbp_1 _20013_ (.CLK(\clknet_leaf_291_top1.acquisition_clk ),
    .RESET_B(net1164),
    .D(_00214_),
    .Q_N(_09765_),
    .Q(\top1.memory1.mem2[95][2] ));
 sg13g2_dfrbp_1 _20014_ (.CLK(\clknet_leaf_101_top1.acquisition_clk ),
    .RESET_B(net1163),
    .D(_00215_),
    .Q_N(_09764_),
    .Q(\top1.memory1.mem2[6][0] ));
 sg13g2_dfrbp_1 _20015_ (.CLK(\clknet_leaf_93_top1.acquisition_clk ),
    .RESET_B(net1162),
    .D(_00216_),
    .Q_N(_09763_),
    .Q(\top1.memory1.mem2[6][1] ));
 sg13g2_dfrbp_1 _20016_ (.CLK(\clknet_leaf_94_top1.acquisition_clk ),
    .RESET_B(net1161),
    .D(_00217_),
    .Q_N(_09762_),
    .Q(\top1.memory1.mem2[6][2] ));
 sg13g2_dfrbp_1 _20017_ (.CLK(\clknet_leaf_211_top1.acquisition_clk ),
    .RESET_B(net1160),
    .D(_00218_),
    .Q_N(_09761_),
    .Q(\top1.memory1.mem2[121][0] ));
 sg13g2_dfrbp_1 _20018_ (.CLK(\clknet_leaf_194_top1.acquisition_clk ),
    .RESET_B(net1159),
    .D(_00219_),
    .Q_N(_09760_),
    .Q(\top1.memory1.mem2[121][1] ));
 sg13g2_dfrbp_1 _20019_ (.CLK(\clknet_leaf_209_top1.acquisition_clk ),
    .RESET_B(net1158),
    .D(_00220_),
    .Q_N(_09759_),
    .Q(\top1.memory1.mem2[121][2] ));
 sg13g2_dfrbp_1 _20020_ (.CLK(\clknet_leaf_211_top1.acquisition_clk ),
    .RESET_B(net1157),
    .D(_00221_),
    .Q_N(_09758_),
    .Q(\top1.memory1.mem2[120][0] ));
 sg13g2_dfrbp_1 _20021_ (.CLK(\clknet_leaf_194_top1.acquisition_clk ),
    .RESET_B(net1156),
    .D(_00222_),
    .Q_N(_09757_),
    .Q(\top1.memory1.mem2[120][1] ));
 sg13g2_dfrbp_1 _20022_ (.CLK(\clknet_leaf_196_top1.acquisition_clk ),
    .RESET_B(net1155),
    .D(_00223_),
    .Q_N(_09756_),
    .Q(\top1.memory1.mem2[120][2] ));
 sg13g2_dfrbp_1 _20023_ (.CLK(\clknet_leaf_86_top1.acquisition_clk ),
    .RESET_B(net1154),
    .D(_00224_),
    .Q_N(_09755_),
    .Q(\top1.memory1.mem2[11][0] ));
 sg13g2_dfrbp_1 _20024_ (.CLK(\clknet_leaf_85_top1.acquisition_clk ),
    .RESET_B(net1153),
    .D(_00225_),
    .Q_N(_09754_),
    .Q(\top1.memory1.mem2[11][1] ));
 sg13g2_dfrbp_1 _20025_ (.CLK(\clknet_leaf_90_top1.acquisition_clk ),
    .RESET_B(net1152),
    .D(_00226_),
    .Q_N(_09753_),
    .Q(\top1.memory1.mem2[11][2] ));
 sg13g2_dfrbp_1 _20026_ (.CLK(\clknet_leaf_222_top1.acquisition_clk ),
    .RESET_B(net1151),
    .D(_00227_),
    .Q_N(_09752_),
    .Q(\top1.memory1.mem2[118][0] ));
 sg13g2_dfrbp_1 _20027_ (.CLK(\clknet_leaf_228_top1.acquisition_clk ),
    .RESET_B(net1150),
    .D(_00228_),
    .Q_N(_09751_),
    .Q(\top1.memory1.mem2[118][1] ));
 sg13g2_dfrbp_1 _20028_ (.CLK(\clknet_leaf_222_top1.acquisition_clk ),
    .RESET_B(net1149),
    .D(_00229_),
    .Q_N(_09750_),
    .Q(\top1.memory1.mem2[118][2] ));
 sg13g2_dfrbp_1 _20029_ (.CLK(\clknet_leaf_222_top1.acquisition_clk ),
    .RESET_B(net1148),
    .D(_00230_),
    .Q_N(_09749_),
    .Q(\top1.memory1.mem2[117][0] ));
 sg13g2_dfrbp_1 _20030_ (.CLK(\clknet_leaf_228_top1.acquisition_clk ),
    .RESET_B(net1147),
    .D(_00231_),
    .Q_N(_09748_),
    .Q(\top1.memory1.mem2[117][1] ));
 sg13g2_dfrbp_1 _20031_ (.CLK(\clknet_leaf_223_top1.acquisition_clk ),
    .RESET_B(net1146),
    .D(_00232_),
    .Q_N(_09747_),
    .Q(\top1.memory1.mem2[117][2] ));
 sg13g2_dfrbp_1 _20032_ (.CLK(\clknet_leaf_96_top1.acquisition_clk ),
    .RESET_B(net1145),
    .D(_00233_),
    .Q_N(_09746_),
    .Q(\top1.memory1.mem2[194][0] ));
 sg13g2_dfrbp_1 _20033_ (.CLK(\clknet_leaf_96_top1.acquisition_clk ),
    .RESET_B(net1144),
    .D(_00234_),
    .Q_N(_09745_),
    .Q(\top1.memory1.mem2[194][1] ));
 sg13g2_dfrbp_1 _20034_ (.CLK(\clknet_leaf_95_top1.acquisition_clk ),
    .RESET_B(net1143),
    .D(_00235_),
    .Q_N(_09744_),
    .Q(\top1.memory1.mem2[194][2] ));
 sg13g2_dfrbp_1 _20035_ (.CLK(\clknet_leaf_95_top1.acquisition_clk ),
    .RESET_B(net1142),
    .D(_00236_),
    .Q_N(_09743_),
    .Q(\top1.memory1.mem2[193][0] ));
 sg13g2_dfrbp_1 _20036_ (.CLK(\clknet_leaf_98_top1.acquisition_clk ),
    .RESET_B(net1141),
    .D(_00237_),
    .Q_N(_09742_),
    .Q(\top1.memory1.mem2[193][1] ));
 sg13g2_dfrbp_1 _20037_ (.CLK(\clknet_leaf_95_top1.acquisition_clk ),
    .RESET_B(net1140),
    .D(_00238_),
    .Q_N(_09741_),
    .Q(\top1.memory1.mem2[193][2] ));
 sg13g2_dfrbp_1 _20038_ (.CLK(\clknet_leaf_96_top1.acquisition_clk ),
    .RESET_B(net1139),
    .D(_00239_),
    .Q_N(_09740_),
    .Q(\top1.memory1.mem2[192][0] ));
 sg13g2_dfrbp_1 _20039_ (.CLK(\clknet_leaf_96_top1.acquisition_clk ),
    .RESET_B(net1138),
    .D(_00240_),
    .Q_N(_09739_),
    .Q(\top1.memory1.mem2[192][1] ));
 sg13g2_dfrbp_1 _20040_ (.CLK(\clknet_leaf_95_top1.acquisition_clk ),
    .RESET_B(net1137),
    .D(_00241_),
    .Q_N(_09738_),
    .Q(\top1.memory1.mem2[192][2] ));
 sg13g2_dfrbp_1 _20041_ (.CLK(\clknet_leaf_117_top1.acquisition_clk ),
    .RESET_B(net1136),
    .D(_00242_),
    .Q_N(_09737_),
    .Q(\top1.memory1.mem2[191][0] ));
 sg13g2_dfrbp_1 _20042_ (.CLK(\clknet_leaf_134_top1.acquisition_clk ),
    .RESET_B(net1135),
    .D(_00243_),
    .Q_N(_09736_),
    .Q(\top1.memory1.mem2[191][1] ));
 sg13g2_dfrbp_1 _20043_ (.CLK(\clknet_leaf_115_top1.acquisition_clk ),
    .RESET_B(net1134),
    .D(_00244_),
    .Q_N(_09735_),
    .Q(\top1.memory1.mem2[191][2] ));
 sg13g2_dfrbp_1 _20044_ (.CLK(\clknet_leaf_117_top1.acquisition_clk ),
    .RESET_B(net1133),
    .D(_00245_),
    .Q_N(_09734_),
    .Q(\top1.memory1.mem2[190][0] ));
 sg13g2_dfrbp_1 _20045_ (.CLK(\clknet_leaf_135_top1.acquisition_clk ),
    .RESET_B(net1132),
    .D(_00246_),
    .Q_N(_09733_),
    .Q(\top1.memory1.mem2[190][1] ));
 sg13g2_dfrbp_1 _20046_ (.CLK(\clknet_leaf_114_top1.acquisition_clk ),
    .RESET_B(net1131),
    .D(_00247_),
    .Q_N(_09732_),
    .Q(\top1.memory1.mem2[190][2] ));
 sg13g2_dfrbp_1 _20047_ (.CLK(\clknet_leaf_120_top1.acquisition_clk ),
    .RESET_B(net1130),
    .D(_00248_),
    .Q_N(_09731_),
    .Q(\top1.memory1.mem2[18][0] ));
 sg13g2_dfrbp_1 _20048_ (.CLK(\clknet_leaf_128_top1.acquisition_clk ),
    .RESET_B(net1129),
    .D(_00249_),
    .Q_N(_09730_),
    .Q(\top1.memory1.mem2[18][1] ));
 sg13g2_dfrbp_1 _20049_ (.CLK(\clknet_leaf_128_top1.acquisition_clk ),
    .RESET_B(net1128),
    .D(_00250_),
    .Q_N(_09729_),
    .Q(\top1.memory1.mem2[18][2] ));
 sg13g2_dfrbp_1 _20050_ (.CLK(\clknet_leaf_117_top1.acquisition_clk ),
    .RESET_B(net1127),
    .D(_00251_),
    .Q_N(_09728_),
    .Q(\top1.memory1.mem2[188][0] ));
 sg13g2_dfrbp_1 _20051_ (.CLK(\clknet_leaf_119_top1.acquisition_clk ),
    .RESET_B(net1126),
    .D(_00252_),
    .Q_N(_09727_),
    .Q(\top1.memory1.mem2[188][1] ));
 sg13g2_dfrbp_1 _20052_ (.CLK(\clknet_leaf_115_top1.acquisition_clk ),
    .RESET_B(net1125),
    .D(_00253_),
    .Q_N(_09726_),
    .Q(\top1.memory1.mem2[188][2] ));
 sg13g2_dfrbp_1 _20053_ (.CLK(\clknet_leaf_118_top1.acquisition_clk ),
    .RESET_B(net1124),
    .D(_00254_),
    .Q_N(_09725_),
    .Q(\top1.memory1.mem2[187][0] ));
 sg13g2_dfrbp_1 _20054_ (.CLK(\clknet_leaf_134_top1.acquisition_clk ),
    .RESET_B(net1123),
    .D(_00255_),
    .Q_N(_09724_),
    .Q(\top1.memory1.mem2[187][1] ));
 sg13g2_dfrbp_1 _20055_ (.CLK(\clknet_leaf_128_top1.acquisition_clk ),
    .RESET_B(net1122),
    .D(_00256_),
    .Q_N(_09723_),
    .Q(\top1.memory1.mem2[187][2] ));
 sg13g2_dfrbp_1 _20056_ (.CLK(\clknet_leaf_118_top1.acquisition_clk ),
    .RESET_B(net1121),
    .D(_00257_),
    .Q_N(_09722_),
    .Q(\top1.memory1.mem2[186][0] ));
 sg13g2_dfrbp_1 _20057_ (.CLK(\clknet_leaf_119_top1.acquisition_clk ),
    .RESET_B(net1120),
    .D(_00258_),
    .Q_N(_09721_),
    .Q(\top1.memory1.mem2[186][1] ));
 sg13g2_dfrbp_1 _20058_ (.CLK(\clknet_leaf_128_top1.acquisition_clk ),
    .RESET_B(net1119),
    .D(_00259_),
    .Q_N(_09720_),
    .Q(\top1.memory1.mem2[186][2] ));
 sg13g2_dfrbp_1 _20059_ (.CLK(\clknet_leaf_120_top1.acquisition_clk ),
    .RESET_B(net1118),
    .D(_00260_),
    .Q_N(_09719_),
    .Q(\top1.memory1.mem2[185][0] ));
 sg13g2_dfrbp_1 _20060_ (.CLK(\clknet_leaf_119_top1.acquisition_clk ),
    .RESET_B(net1117),
    .D(_00261_),
    .Q_N(_09718_),
    .Q(\top1.memory1.mem2[185][1] ));
 sg13g2_dfrbp_1 _20061_ (.CLK(\clknet_leaf_127_top1.acquisition_clk ),
    .RESET_B(net1116),
    .D(_00262_),
    .Q_N(_09717_),
    .Q(\top1.memory1.mem2[185][2] ));
 sg13g2_dfrbp_1 _20062_ (.CLK(\clknet_leaf_120_top1.acquisition_clk ),
    .RESET_B(net1115),
    .D(_00263_),
    .Q_N(_09716_),
    .Q(\top1.memory1.mem2[184][0] ));
 sg13g2_dfrbp_1 _20063_ (.CLK(\clknet_leaf_123_top1.acquisition_clk ),
    .RESET_B(net1114),
    .D(_00264_),
    .Q_N(_09715_),
    .Q(\top1.memory1.mem2[184][1] ));
 sg13g2_dfrbp_1 _20064_ (.CLK(\clknet_leaf_128_top1.acquisition_clk ),
    .RESET_B(net1113),
    .D(_00265_),
    .Q_N(_09714_),
    .Q(\top1.memory1.mem2[184][2] ));
 sg13g2_dfrbp_1 _20065_ (.CLK(\clknet_leaf_114_top1.acquisition_clk ),
    .RESET_B(net1112),
    .D(_00266_),
    .Q_N(_09713_),
    .Q(\top1.memory1.mem2[183][0] ));
 sg13g2_dfrbp_1 _20066_ (.CLK(\clknet_leaf_114_top1.acquisition_clk ),
    .RESET_B(net1111),
    .D(_00267_),
    .Q_N(_09712_),
    .Q(\top1.memory1.mem2[183][1] ));
 sg13g2_dfrbp_1 _20067_ (.CLK(\clknet_leaf_177_top1.acquisition_clk ),
    .RESET_B(net1110),
    .D(_00268_),
    .Q_N(_09711_),
    .Q(\top1.memory1.mem2[183][2] ));
 sg13g2_dfrbp_1 _20068_ (.CLK(\clknet_leaf_114_top1.acquisition_clk ),
    .RESET_B(net1109),
    .D(_00269_),
    .Q_N(_09710_),
    .Q(\top1.memory1.mem2[182][0] ));
 sg13g2_dfrbp_1 _20069_ (.CLK(\clknet_leaf_114_top1.acquisition_clk ),
    .RESET_B(net1108),
    .D(_00270_),
    .Q_N(_09709_),
    .Q(\top1.memory1.mem2[182][1] ));
 sg13g2_dfrbp_1 _20070_ (.CLK(\clknet_leaf_177_top1.acquisition_clk ),
    .RESET_B(net1107),
    .D(_00271_),
    .Q_N(_09708_),
    .Q(\top1.memory1.mem2[182][2] ));
 sg13g2_dfrbp_1 _20071_ (.CLK(\clknet_leaf_115_top1.acquisition_clk ),
    .RESET_B(net1106),
    .D(_00272_),
    .Q_N(_09707_),
    .Q(\top1.memory1.mem2[181][0] ));
 sg13g2_dfrbp_1 _20072_ (.CLK(\clknet_leaf_115_top1.acquisition_clk ),
    .RESET_B(net1105),
    .D(_00273_),
    .Q_N(_09706_),
    .Q(\top1.memory1.mem2[181][1] ));
 sg13g2_dfrbp_1 _20073_ (.CLK(\clknet_leaf_181_top1.acquisition_clk ),
    .RESET_B(net1104),
    .D(_00274_),
    .Q_N(_09705_),
    .Q(\top1.memory1.mem2[181][2] ));
 sg13g2_dfrbp_1 _20074_ (.CLK(\clknet_leaf_113_top1.acquisition_clk ),
    .RESET_B(net1103),
    .D(_00275_),
    .Q_N(_09704_),
    .Q(\top1.memory1.mem2[180][0] ));
 sg13g2_dfrbp_1 _20075_ (.CLK(\clknet_leaf_113_top1.acquisition_clk ),
    .RESET_B(net1102),
    .D(_00276_),
    .Q_N(_09703_),
    .Q(\top1.memory1.mem2[180][1] ));
 sg13g2_dfrbp_1 _20076_ (.CLK(\clknet_leaf_177_top1.acquisition_clk ),
    .RESET_B(net1101),
    .D(_00277_),
    .Q_N(_09702_),
    .Q(\top1.memory1.mem2[180][2] ));
 sg13g2_dfrbp_1 _20077_ (.CLK(\clknet_leaf_120_top1.acquisition_clk ),
    .RESET_B(net1100),
    .D(_00278_),
    .Q_N(_09701_),
    .Q(\top1.memory1.mem2[17][0] ));
 sg13g2_dfrbp_1 _20078_ (.CLK(\clknet_leaf_123_top1.acquisition_clk ),
    .RESET_B(net1099),
    .D(_00279_),
    .Q_N(_09700_),
    .Q(\top1.memory1.mem2[17][1] ));
 sg13g2_dfrbp_1 _20079_ (.CLK(\clknet_leaf_128_top1.acquisition_clk ),
    .RESET_B(net1098),
    .D(_00280_),
    .Q_N(_09699_),
    .Q(\top1.memory1.mem2[17][2] ));
 sg13g2_dfrbp_1 _20080_ (.CLK(\clknet_leaf_134_top1.acquisition_clk ),
    .RESET_B(net1097),
    .D(_00281_),
    .Q_N(_09698_),
    .Q(\top1.memory1.mem2[178][0] ));
 sg13g2_dfrbp_1 _20081_ (.CLK(\clknet_leaf_129_top1.acquisition_clk ),
    .RESET_B(net1096),
    .D(_00282_),
    .Q_N(_09697_),
    .Q(\top1.memory1.mem2[178][1] ));
 sg13g2_dfrbp_1 _20082_ (.CLK(\clknet_leaf_130_top1.acquisition_clk ),
    .RESET_B(net1095),
    .D(_00283_),
    .Q_N(_09696_),
    .Q(\top1.memory1.mem2[178][2] ));
 sg13g2_dfrbp_1 _20083_ (.CLK(\clknet_leaf_134_top1.acquisition_clk ),
    .RESET_B(net1094),
    .D(_00284_),
    .Q_N(_09695_),
    .Q(\top1.memory1.mem2[177][0] ));
 sg13g2_dfrbp_1 _20084_ (.CLK(\clknet_leaf_129_top1.acquisition_clk ),
    .RESET_B(net1093),
    .D(_00285_),
    .Q_N(_09694_),
    .Q(\top1.memory1.mem2[177][1] ));
 sg13g2_dfrbp_1 _20085_ (.CLK(\clknet_leaf_131_top1.acquisition_clk ),
    .RESET_B(net1092),
    .D(_00286_),
    .Q_N(_09693_),
    .Q(\top1.memory1.mem2[177][2] ));
 sg13g2_dfrbp_1 _20086_ (.CLK(\clknet_leaf_134_top1.acquisition_clk ),
    .RESET_B(net1091),
    .D(_00287_),
    .Q_N(_09692_),
    .Q(\top1.memory1.mem2[176][0] ));
 sg13g2_dfrbp_1 _20087_ (.CLK(\clknet_leaf_129_top1.acquisition_clk ),
    .RESET_B(net1090),
    .D(_00288_),
    .Q_N(_09691_),
    .Q(\top1.memory1.mem2[176][1] ));
 sg13g2_dfrbp_1 _20088_ (.CLK(\clknet_leaf_130_top1.acquisition_clk ),
    .RESET_B(net1089),
    .D(_00289_),
    .Q_N(_09690_),
    .Q(\top1.memory1.mem2[176][2] ));
 sg13g2_dfrbp_1 _20089_ (.CLK(\clknet_leaf_37_top1.acquisition_clk ),
    .RESET_B(net1088),
    .D(_00290_),
    .Q_N(_09689_),
    .Q(\top1.memory1.mem2[175][0] ));
 sg13g2_dfrbp_1 _20090_ (.CLK(\clknet_leaf_263_top1.acquisition_clk ),
    .RESET_B(net1087),
    .D(_00291_),
    .Q_N(_09688_),
    .Q(\top1.memory1.mem2[175][1] ));
 sg13g2_dfrbp_1 _20091_ (.CLK(\clknet_leaf_259_top1.acquisition_clk ),
    .RESET_B(net1086),
    .D(_00292_),
    .Q_N(_09687_),
    .Q(\top1.memory1.mem2[175][2] ));
 sg13g2_dfrbp_1 _20092_ (.CLK(\clknet_leaf_260_top1.acquisition_clk ),
    .RESET_B(net1085),
    .D(_00293_),
    .Q_N(_09686_),
    .Q(\top1.memory1.mem2[174][0] ));
 sg13g2_dfrbp_1 _20093_ (.CLK(\clknet_leaf_263_top1.acquisition_clk ),
    .RESET_B(net1084),
    .D(_00294_),
    .Q_N(_09685_),
    .Q(\top1.memory1.mem2[174][1] ));
 sg13g2_dfrbp_1 _20094_ (.CLK(\clknet_leaf_264_top1.acquisition_clk ),
    .RESET_B(net1083),
    .D(_00295_),
    .Q_N(_09684_),
    .Q(\top1.memory1.mem2[174][2] ));
 sg13g2_dfrbp_1 _20095_ (.CLK(\clknet_leaf_260_top1.acquisition_clk ),
    .RESET_B(net1082),
    .D(_00296_),
    .Q_N(_09683_),
    .Q(\top1.memory1.mem2[173][0] ));
 sg13g2_dfrbp_1 _20096_ (.CLK(\clknet_leaf_264_top1.acquisition_clk ),
    .RESET_B(net1081),
    .D(_00297_),
    .Q_N(_09682_),
    .Q(\top1.memory1.mem2[173][1] ));
 sg13g2_dfrbp_1 _20097_ (.CLK(\clknet_leaf_264_top1.acquisition_clk ),
    .RESET_B(net1080),
    .D(_00298_),
    .Q_N(_09681_),
    .Q(\top1.memory1.mem2[173][2] ));
 sg13g2_dfrbp_1 _20098_ (.CLK(\clknet_leaf_261_top1.acquisition_clk ),
    .RESET_B(net1079),
    .D(_00299_),
    .Q_N(_09680_),
    .Q(\top1.memory1.mem2[172][0] ));
 sg13g2_dfrbp_1 _20099_ (.CLK(\clknet_leaf_264_top1.acquisition_clk ),
    .RESET_B(net1078),
    .D(_00300_),
    .Q_N(_09679_),
    .Q(\top1.memory1.mem2[172][1] ));
 sg13g2_dfrbp_1 _20100_ (.CLK(\clknet_leaf_261_top1.acquisition_clk ),
    .RESET_B(net1077),
    .D(_00301_),
    .Q_N(_09678_),
    .Q(\top1.memory1.mem2[172][2] ));
 sg13g2_dfrbp_1 _20101_ (.CLK(\clknet_leaf_107_top1.acquisition_clk ),
    .RESET_B(net1076),
    .D(_00302_),
    .Q_N(_09677_),
    .Q(\top1.memory1.mem2[171][0] ));
 sg13g2_dfrbp_1 _20102_ (.CLK(\clknet_leaf_183_top1.acquisition_clk ),
    .RESET_B(net1075),
    .D(_00303_),
    .Q_N(_09676_),
    .Q(\top1.memory1.mem2[171][1] ));
 sg13g2_dfrbp_1 _20103_ (.CLK(\clknet_leaf_109_top1.acquisition_clk ),
    .RESET_B(net1074),
    .D(_00304_),
    .Q_N(_09675_),
    .Q(\top1.memory1.mem2[171][2] ));
 sg13g2_dfrbp_1 _20104_ (.CLK(\clknet_leaf_107_top1.acquisition_clk ),
    .RESET_B(net1073),
    .D(_00305_),
    .Q_N(_09674_),
    .Q(\top1.memory1.mem2[170][0] ));
 sg13g2_dfrbp_1 _20105_ (.CLK(\clknet_leaf_183_top1.acquisition_clk ),
    .RESET_B(net1072),
    .D(_00306_),
    .Q_N(_09673_),
    .Q(\top1.memory1.mem2[170][1] ));
 sg13g2_dfrbp_1 _20106_ (.CLK(\clknet_leaf_110_top1.acquisition_clk ),
    .RESET_B(net1071),
    .D(_00307_),
    .Q_N(_09672_),
    .Q(\top1.memory1.mem2[170][2] ));
 sg13g2_dfrbp_1 _20107_ (.CLK(\clknet_leaf_119_top1.acquisition_clk ),
    .RESET_B(net1070),
    .D(_00308_),
    .Q_N(_09671_),
    .Q(\top1.memory1.mem2[16][0] ));
 sg13g2_dfrbp_1 _20108_ (.CLK(\clknet_leaf_122_top1.acquisition_clk ),
    .RESET_B(net1069),
    .D(_00309_),
    .Q_N(_09670_),
    .Q(\top1.memory1.mem2[16][1] ));
 sg13g2_dfrbp_1 _20109_ (.CLK(\clknet_leaf_123_top1.acquisition_clk ),
    .RESET_B(net1068),
    .D(_00310_),
    .Q_N(_09669_),
    .Q(\top1.memory1.mem2[16][2] ));
 sg13g2_dfrbp_1 _20110_ (.CLK(\clknet_leaf_105_top1.acquisition_clk ),
    .RESET_B(net1067),
    .D(_00311_),
    .Q_N(_09668_),
    .Q(\top1.memory1.mem2[168][0] ));
 sg13g2_dfrbp_1 _20111_ (.CLK(\clknet_leaf_106_top1.acquisition_clk ),
    .RESET_B(net1066),
    .D(_00312_),
    .Q_N(_09667_),
    .Q(\top1.memory1.mem2[168][1] ));
 sg13g2_dfrbp_1 _20112_ (.CLK(\clknet_leaf_107_top1.acquisition_clk ),
    .RESET_B(net1065),
    .D(_00313_),
    .Q_N(_09666_),
    .Q(\top1.memory1.mem2[168][2] ));
 sg13g2_dfrbp_1 _20113_ (.CLK(\clknet_leaf_101_top1.acquisition_clk ),
    .RESET_B(net1064),
    .D(_00314_),
    .Q_N(_09665_),
    .Q(\top1.memory1.mem2[167][0] ));
 sg13g2_dfrbp_1 _20114_ (.CLK(\clknet_leaf_102_top1.acquisition_clk ),
    .RESET_B(net1062),
    .D(_00315_),
    .Q_N(_09664_),
    .Q(\top1.memory1.mem2[167][1] ));
 sg13g2_dfrbp_1 _20115_ (.CLK(\clknet_leaf_111_top1.acquisition_clk ),
    .RESET_B(net1061),
    .D(_00316_),
    .Q_N(_09663_),
    .Q(\top1.memory1.mem2[167][2] ));
 sg13g2_dfrbp_1 _20116_ (.CLK(\clknet_leaf_101_top1.acquisition_clk ),
    .RESET_B(net1060),
    .D(_00317_),
    .Q_N(_09662_),
    .Q(\top1.memory1.mem2[166][0] ));
 sg13g2_dfrbp_1 _20117_ (.CLK(\clknet_leaf_102_top1.acquisition_clk ),
    .RESET_B(net1059),
    .D(_00318_),
    .Q_N(_09661_),
    .Q(\top1.memory1.mem2[166][1] ));
 sg13g2_dfrbp_1 _20118_ (.CLK(\clknet_leaf_111_top1.acquisition_clk ),
    .RESET_B(net1058),
    .D(_00319_),
    .Q_N(_09660_),
    .Q(\top1.memory1.mem2[166][2] ));
 sg13g2_dfrbp_1 _20119_ (.CLK(\clknet_leaf_101_top1.acquisition_clk ),
    .RESET_B(net1057),
    .D(_00320_),
    .Q_N(_09659_),
    .Q(\top1.memory1.mem2[165][0] ));
 sg13g2_dfrbp_1 _20120_ (.CLK(\clknet_leaf_102_top1.acquisition_clk ),
    .RESET_B(net1056),
    .D(_00321_),
    .Q_N(_09658_),
    .Q(\top1.memory1.mem2[165][1] ));
 sg13g2_dfrbp_1 _20121_ (.CLK(\clknet_leaf_101_top1.acquisition_clk ),
    .RESET_B(net1055),
    .D(_00322_),
    .Q_N(_09657_),
    .Q(\top1.memory1.mem2[165][2] ));
 sg13g2_dfrbp_1 _20122_ (.CLK(\clknet_leaf_93_top1.acquisition_clk ),
    .RESET_B(net1054),
    .D(_00323_),
    .Q_N(_09656_),
    .Q(\top1.memory1.mem2[164][0] ));
 sg13g2_dfrbp_1 _20123_ (.CLK(\clknet_leaf_102_top1.acquisition_clk ),
    .RESET_B(net1053),
    .D(_00324_),
    .Q_N(_09655_),
    .Q(\top1.memory1.mem2[164][1] ));
 sg13g2_dfrbp_1 _20124_ (.CLK(\clknet_leaf_101_top1.acquisition_clk ),
    .RESET_B(net1052),
    .D(_00325_),
    .Q_N(_09654_),
    .Q(\top1.memory1.mem2[164][2] ));
 sg13g2_dfrbp_1 _20125_ (.CLK(\clknet_leaf_104_top1.acquisition_clk ),
    .RESET_B(net1051),
    .D(_00326_),
    .Q_N(_09653_),
    .Q(\top1.memory1.mem2[163][0] ));
 sg13g2_dfrbp_1 _20126_ (.CLK(\clknet_leaf_37_top1.acquisition_clk ),
    .RESET_B(net1049),
    .D(_00327_),
    .Q_N(_09652_),
    .Q(\top1.memory1.mem2[163][1] ));
 sg13g2_dfrbp_1 _20127_ (.CLK(\clknet_leaf_103_top1.acquisition_clk ),
    .RESET_B(net1048),
    .D(_00328_),
    .Q_N(_09651_),
    .Q(\top1.memory1.mem2[163][2] ));
 sg13g2_dfrbp_1 _20128_ (.CLK(\clknet_leaf_104_top1.acquisition_clk ),
    .RESET_B(net1047),
    .D(_00329_),
    .Q_N(_09650_),
    .Q(\top1.memory1.mem2[162][0] ));
 sg13g2_dfrbp_1 _20129_ (.CLK(\clknet_leaf_105_top1.acquisition_clk ),
    .RESET_B(net1046),
    .D(_00330_),
    .Q_N(_09649_),
    .Q(\top1.memory1.mem2[162][1] ));
 sg13g2_dfrbp_1 _20130_ (.CLK(\clknet_leaf_99_top1.acquisition_clk ),
    .RESET_B(net1045),
    .D(_00331_),
    .Q_N(_09648_),
    .Q(\top1.memory1.mem2[162][2] ));
 sg13g2_dfrbp_1 _20131_ (.CLK(\clknet_leaf_104_top1.acquisition_clk ),
    .RESET_B(net1044),
    .D(_00332_),
    .Q_N(_09647_),
    .Q(\top1.memory1.mem2[161][0] ));
 sg13g2_dfrbp_1 _20132_ (.CLK(\clknet_leaf_38_top1.acquisition_clk ),
    .RESET_B(net1043),
    .D(_00333_),
    .Q_N(_09646_),
    .Q(\top1.memory1.mem2[161][1] ));
 sg13g2_dfrbp_1 _20133_ (.CLK(\clknet_leaf_103_top1.acquisition_clk ),
    .RESET_B(net1042),
    .D(_00334_),
    .Q_N(_09645_),
    .Q(\top1.memory1.mem2[161][2] ));
 sg13g2_dfrbp_1 _20134_ (.CLK(\clknet_leaf_104_top1.acquisition_clk ),
    .RESET_B(net1041),
    .D(_00335_),
    .Q_N(_09644_),
    .Q(\top1.memory1.mem2[160][0] ));
 sg13g2_dfrbp_1 _20135_ (.CLK(\clknet_leaf_38_top1.acquisition_clk ),
    .RESET_B(net1040),
    .D(_00336_),
    .Q_N(_09643_),
    .Q(\top1.memory1.mem2[160][1] ));
 sg13g2_dfrbp_1 _20136_ (.CLK(\clknet_leaf_103_top1.acquisition_clk ),
    .RESET_B(net1039),
    .D(_00337_),
    .Q_N(_09642_),
    .Q(\top1.memory1.mem2[160][2] ));
 sg13g2_dfrbp_1 _20137_ (.CLK(\clknet_leaf_84_top1.acquisition_clk ),
    .RESET_B(net1038),
    .D(_00338_),
    .Q_N(_09641_),
    .Q(\top1.memory1.mem2[15][0] ));
 sg13g2_dfrbp_1 _20138_ (.CLK(\clknet_leaf_83_top1.acquisition_clk ),
    .RESET_B(net1037),
    .D(_00339_),
    .Q_N(_09640_),
    .Q(\top1.memory1.mem2[15][1] ));
 sg13g2_dfrbp_1 _20139_ (.CLK(\clknet_leaf_82_top1.acquisition_clk ),
    .RESET_B(net1036),
    .D(_00340_),
    .Q_N(_09639_),
    .Q(\top1.memory1.mem2[15][2] ));
 sg13g2_dfrbp_1 _20140_ (.CLK(\clknet_leaf_73_top1.acquisition_clk ),
    .RESET_B(net1035),
    .D(_00341_),
    .Q_N(_09638_),
    .Q(\top1.memory1.mem2[158][0] ));
 sg13g2_dfrbp_1 _20141_ (.CLK(\clknet_leaf_73_top1.acquisition_clk ),
    .RESET_B(net1034),
    .D(_00342_),
    .Q_N(_09637_),
    .Q(\top1.memory1.mem2[158][1] ));
 sg13g2_dfrbp_1 _20142_ (.CLK(\clknet_leaf_72_top1.acquisition_clk ),
    .RESET_B(net1033),
    .D(_00343_),
    .Q_N(_09636_),
    .Q(\top1.memory1.mem2[158][2] ));
 sg13g2_dfrbp_1 _20143_ (.CLK(\clknet_leaf_71_top1.acquisition_clk ),
    .RESET_B(net1032),
    .D(_00344_),
    .Q_N(_09635_),
    .Q(\top1.memory1.mem2[157][0] ));
 sg13g2_dfrbp_1 _20144_ (.CLK(\clknet_leaf_72_top1.acquisition_clk ),
    .RESET_B(net1031),
    .D(_00345_),
    .Q_N(_09634_),
    .Q(\top1.memory1.mem2[157][1] ));
 sg13g2_dfrbp_1 _20145_ (.CLK(\clknet_leaf_81_top1.acquisition_clk ),
    .RESET_B(net1030),
    .D(_00346_),
    .Q_N(_09633_),
    .Q(\top1.memory1.mem2[157][2] ));
 sg13g2_dfrbp_1 _20146_ (.CLK(\clknet_leaf_71_top1.acquisition_clk ),
    .RESET_B(net1029),
    .D(_00347_),
    .Q_N(_09632_),
    .Q(\top1.memory1.mem2[156][0] ));
 sg13g2_dfrbp_1 _20147_ (.CLK(\clknet_leaf_73_top1.acquisition_clk ),
    .RESET_B(net1028),
    .D(_00348_),
    .Q_N(_09631_),
    .Q(\top1.memory1.mem2[156][1] ));
 sg13g2_dfrbp_1 _20148_ (.CLK(\clknet_leaf_72_top1.acquisition_clk ),
    .RESET_B(net1027),
    .D(_00349_),
    .Q_N(_09630_),
    .Q(\top1.memory1.mem2[156][2] ));
 sg13g2_dfrbp_1 _20149_ (.CLK(\clknet_leaf_79_top1.acquisition_clk ),
    .RESET_B(net1026),
    .D(_00350_),
    .Q_N(_09629_),
    .Q(\top1.memory1.mem2[155][0] ));
 sg13g2_dfrbp_1 _20150_ (.CLK(\clknet_leaf_80_top1.acquisition_clk ),
    .RESET_B(net1025),
    .D(_00351_),
    .Q_N(_09628_),
    .Q(\top1.memory1.mem2[155][1] ));
 sg13g2_dfrbp_1 _20151_ (.CLK(\clknet_leaf_97_top1.acquisition_clk ),
    .RESET_B(net1024),
    .D(_00352_),
    .Q_N(_09627_),
    .Q(\top1.memory1.mem2[155][2] ));
 sg13g2_dfrbp_1 _20152_ (.CLK(\clknet_leaf_80_top1.acquisition_clk ),
    .RESET_B(net1023),
    .D(_00353_),
    .Q_N(_09626_),
    .Q(\top1.memory1.mem2[154][0] ));
 sg13g2_dfrbp_1 _20153_ (.CLK(\clknet_leaf_81_top1.acquisition_clk ),
    .RESET_B(net1022),
    .D(_00354_),
    .Q_N(_09625_),
    .Q(\top1.memory1.mem2[154][1] ));
 sg13g2_dfrbp_1 _20154_ (.CLK(\clknet_leaf_77_top1.acquisition_clk ),
    .RESET_B(net1021),
    .D(_00355_),
    .Q_N(_09624_),
    .Q(\top1.memory1.mem2[154][2] ));
 sg13g2_dfrbp_1 _20155_ (.CLK(\clknet_leaf_82_top1.acquisition_clk ),
    .RESET_B(net1020),
    .D(_00356_),
    .Q_N(_09623_),
    .Q(\top1.memory1.mem2[153][0] ));
 sg13g2_dfrbp_1 _20156_ (.CLK(\clknet_leaf_78_top1.acquisition_clk ),
    .RESET_B(net1019),
    .D(_00357_),
    .Q_N(_09622_),
    .Q(\top1.memory1.mem2[153][1] ));
 sg13g2_dfrbp_1 _20157_ (.CLK(\clknet_leaf_96_top1.acquisition_clk ),
    .RESET_B(net1018),
    .D(_00358_),
    .Q_N(_09621_),
    .Q(\top1.memory1.mem2[153][2] ));
 sg13g2_dfrbp_1 _20158_ (.CLK(\clknet_leaf_82_top1.acquisition_clk ),
    .RESET_B(net1017),
    .D(_00359_),
    .Q_N(_09620_),
    .Q(\top1.memory1.mem2[152][0] ));
 sg13g2_dfrbp_1 _20159_ (.CLK(\clknet_leaf_82_top1.acquisition_clk ),
    .RESET_B(net1016),
    .D(_00360_),
    .Q_N(_09619_),
    .Q(\top1.memory1.mem2[152][1] ));
 sg13g2_dfrbp_1 _20160_ (.CLK(\clknet_leaf_77_top1.acquisition_clk ),
    .RESET_B(net1015),
    .D(_00361_),
    .Q_N(_09618_),
    .Q(\top1.memory1.mem2[152][2] ));
 sg13g2_dfrbp_1 _20161_ (.CLK(\clknet_leaf_43_top1.acquisition_clk ),
    .RESET_B(net1014),
    .D(_00362_),
    .Q_N(_09617_),
    .Q(\top1.memory1.mem2[151][0] ));
 sg13g2_dfrbp_1 _20162_ (.CLK(\clknet_leaf_58_top1.acquisition_clk ),
    .RESET_B(net1013),
    .D(_00363_),
    .Q_N(_09616_),
    .Q(\top1.memory1.mem2[151][1] ));
 sg13g2_dfrbp_1 _20163_ (.CLK(\clknet_leaf_42_top1.acquisition_clk ),
    .RESET_B(net1012),
    .D(_00364_),
    .Q_N(_09615_),
    .Q(\top1.memory1.mem2[151][2] ));
 sg13g2_dfrbp_1 _20164_ (.CLK(\clknet_leaf_43_top1.acquisition_clk ),
    .RESET_B(net1011),
    .D(_00365_),
    .Q_N(_09614_),
    .Q(\top1.memory1.mem2[150][0] ));
 sg13g2_dfrbp_1 _20165_ (.CLK(\clknet_leaf_42_top1.acquisition_clk ),
    .RESET_B(net1010),
    .D(_00366_),
    .Q_N(_09613_),
    .Q(\top1.memory1.mem2[150][1] ));
 sg13g2_dfrbp_1 _20166_ (.CLK(\clknet_leaf_42_top1.acquisition_clk ),
    .RESET_B(net1009),
    .D(_00367_),
    .Q_N(_09612_),
    .Q(\top1.memory1.mem2[150][2] ));
 sg13g2_dfrbp_1 _20167_ (.CLK(\clknet_leaf_83_top1.acquisition_clk ),
    .RESET_B(net1008),
    .D(_00368_),
    .Q_N(_09611_),
    .Q(\top1.memory1.mem2[14][0] ));
 sg13g2_dfrbp_1 _20168_ (.CLK(\clknet_leaf_83_top1.acquisition_clk ),
    .RESET_B(net1007),
    .D(_00369_),
    .Q_N(_09610_),
    .Q(\top1.memory1.mem2[14][1] ));
 sg13g2_dfrbp_1 _20169_ (.CLK(\clknet_leaf_83_top1.acquisition_clk ),
    .RESET_B(net1006),
    .D(_00370_),
    .Q_N(_09609_),
    .Q(\top1.memory1.mem2[14][2] ));
 sg13g2_dfrbp_1 _20170_ (.CLK(\clknet_leaf_97_top1.acquisition_clk ),
    .RESET_B(net1005),
    .D(_00371_),
    .Q_N(_09608_),
    .Q(\top1.memory1.mem2[148][0] ));
 sg13g2_dfrbp_1 _20171_ (.CLK(\clknet_leaf_77_top1.acquisition_clk ),
    .RESET_B(net1004),
    .D(_00372_),
    .Q_N(_09607_),
    .Q(\top1.memory1.mem2[148][1] ));
 sg13g2_dfrbp_1 _20172_ (.CLK(\clknet_leaf_42_top1.acquisition_clk ),
    .RESET_B(net1003),
    .D(_00373_),
    .Q_N(_09606_),
    .Q(\top1.memory1.mem2[148][2] ));
 sg13g2_dfrbp_1 _20173_ (.CLK(\clknet_leaf_75_top1.acquisition_clk ),
    .RESET_B(net1002),
    .D(_00374_),
    .Q_N(_09605_),
    .Q(\top1.memory1.mem2[147][0] ));
 sg13g2_dfrbp_1 _20174_ (.CLK(\clknet_leaf_76_top1.acquisition_clk ),
    .RESET_B(net1001),
    .D(_00375_),
    .Q_N(_09604_),
    .Q(\top1.memory1.mem2[147][1] ));
 sg13g2_dfrbp_1 _20175_ (.CLK(\clknet_leaf_78_top1.acquisition_clk ),
    .RESET_B(net1000),
    .D(_00376_),
    .Q_N(_09603_),
    .Q(\top1.memory1.mem2[147][2] ));
 sg13g2_dfrbp_1 _20176_ (.CLK(\clknet_leaf_75_top1.acquisition_clk ),
    .RESET_B(net999),
    .D(_00377_),
    .Q_N(_09602_),
    .Q(\top1.memory1.mem2[146][0] ));
 sg13g2_dfrbp_1 _20177_ (.CLK(\clknet_leaf_59_top1.acquisition_clk ),
    .RESET_B(net998),
    .D(_00378_),
    .Q_N(_09601_),
    .Q(\top1.memory1.mem2[146][1] ));
 sg13g2_dfrbp_1 _20178_ (.CLK(\clknet_leaf_77_top1.acquisition_clk ),
    .RESET_B(net997),
    .D(_00379_),
    .Q_N(_09600_),
    .Q(\top1.memory1.mem2[146][2] ));
 sg13g2_dfrbp_1 _20179_ (.CLK(\clknet_leaf_72_top1.acquisition_clk ),
    .RESET_B(net996),
    .D(_00380_),
    .Q_N(_09599_),
    .Q(\top1.memory1.mem2[145][0] ));
 sg13g2_dfrbp_1 _20180_ (.CLK(\clknet_leaf_59_top1.acquisition_clk ),
    .RESET_B(net995),
    .D(_00381_),
    .Q_N(_09598_),
    .Q(\top1.memory1.mem2[145][1] ));
 sg13g2_dfrbp_1 _20181_ (.CLK(\clknet_leaf_78_top1.acquisition_clk ),
    .RESET_B(net994),
    .D(_00382_),
    .Q_N(_09597_),
    .Q(\top1.memory1.mem2[145][2] ));
 sg13g2_dfrbp_1 _20182_ (.CLK(\clknet_leaf_72_top1.acquisition_clk ),
    .RESET_B(net993),
    .D(_00383_),
    .Q_N(_09596_),
    .Q(\top1.memory1.mem2[144][0] ));
 sg13g2_dfrbp_1 _20183_ (.CLK(\clknet_leaf_76_top1.acquisition_clk ),
    .RESET_B(net992),
    .D(_00384_),
    .Q_N(_09595_),
    .Q(\top1.memory1.mem2[144][1] ));
 sg13g2_dfrbp_1 _20184_ (.CLK(\clknet_leaf_77_top1.acquisition_clk ),
    .RESET_B(net991),
    .D(_00385_),
    .Q_N(_09594_),
    .Q(\top1.memory1.mem2[144][2] ));
 sg13g2_dfrbp_1 _20185_ (.CLK(\clknet_leaf_55_top1.acquisition_clk ),
    .RESET_B(net990),
    .D(_00386_),
    .Q_N(_09593_),
    .Q(\top1.memory1.mem2[143][0] ));
 sg13g2_dfrbp_1 _20186_ (.CLK(\clknet_leaf_62_top1.acquisition_clk ),
    .RESET_B(net989),
    .D(_00387_),
    .Q_N(_09592_),
    .Q(\top1.memory1.mem2[143][1] ));
 sg13g2_dfrbp_1 _20187_ (.CLK(\clknet_leaf_64_top1.acquisition_clk ),
    .RESET_B(net988),
    .D(_00388_),
    .Q_N(_09591_),
    .Q(\top1.memory1.mem2[143][2] ));
 sg13g2_dfrbp_1 _20188_ (.CLK(\clknet_leaf_62_top1.acquisition_clk ),
    .RESET_B(net987),
    .D(_00389_),
    .Q_N(_09590_),
    .Q(\top1.memory1.mem2[142][0] ));
 sg13g2_dfrbp_1 _20189_ (.CLK(\clknet_leaf_63_top1.acquisition_clk ),
    .RESET_B(net986),
    .D(_00390_),
    .Q_N(_09589_),
    .Q(\top1.memory1.mem2[142][1] ));
 sg13g2_dfrbp_1 _20190_ (.CLK(\clknet_leaf_63_top1.acquisition_clk ),
    .RESET_B(net985),
    .D(_00391_),
    .Q_N(_09588_),
    .Q(\top1.memory1.mem2[142][2] ));
 sg13g2_dfrbp_1 _20191_ (.CLK(\clknet_leaf_62_top1.acquisition_clk ),
    .RESET_B(net984),
    .D(_00392_),
    .Q_N(_09587_),
    .Q(\top1.memory1.mem2[141][0] ));
 sg13g2_dfrbp_1 _20192_ (.CLK(\clknet_leaf_62_top1.acquisition_clk ),
    .RESET_B(net983),
    .D(_00393_),
    .Q_N(_09586_),
    .Q(\top1.memory1.mem2[141][1] ));
 sg13g2_dfrbp_1 _20193_ (.CLK(\clknet_leaf_65_top1.acquisition_clk ),
    .RESET_B(net982),
    .D(_00394_),
    .Q_N(_09585_),
    .Q(\top1.memory1.mem2[141][2] ));
 sg13g2_dfrbp_1 _20194_ (.CLK(\clknet_leaf_55_top1.acquisition_clk ),
    .RESET_B(net981),
    .D(_00395_),
    .Q_N(_09584_),
    .Q(\top1.memory1.mem2[140][0] ));
 sg13g2_dfrbp_1 _20195_ (.CLK(\clknet_leaf_61_top1.acquisition_clk ),
    .RESET_B(net980),
    .D(_00396_),
    .Q_N(_09583_),
    .Q(\top1.memory1.mem2[140][1] ));
 sg13g2_dfrbp_1 _20196_ (.CLK(\clknet_leaf_63_top1.acquisition_clk ),
    .RESET_B(net979),
    .D(_00397_),
    .Q_N(_09582_),
    .Q(\top1.memory1.mem2[140][2] ));
 sg13g2_dfrbp_1 _20197_ (.CLK(\clknet_leaf_83_top1.acquisition_clk ),
    .RESET_B(net978),
    .D(_00398_),
    .Q_N(_09581_),
    .Q(\top1.memory1.mem2[13][0] ));
 sg13g2_dfrbp_1 _20198_ (.CLK(\clknet_leaf_83_top1.acquisition_clk ),
    .RESET_B(net977),
    .D(_00399_),
    .Q_N(_09580_),
    .Q(\top1.memory1.mem2[13][1] ));
 sg13g2_dfrbp_1 _20199_ (.CLK(\clknet_leaf_82_top1.acquisition_clk ),
    .RESET_B(net976),
    .D(_00400_),
    .Q_N(_09579_),
    .Q(\top1.memory1.mem2[13][2] ));
 sg13g2_dfrbp_1 _20200_ (.CLK(\clknet_leaf_74_top1.acquisition_clk ),
    .RESET_B(net975),
    .D(_00401_),
    .Q_N(_09578_),
    .Q(\top1.memory1.mem2[138][0] ));
 sg13g2_dfrbp_1 _20201_ (.CLK(\clknet_leaf_74_top1.acquisition_clk ),
    .RESET_B(net974),
    .D(_00402_),
    .Q_N(_09577_),
    .Q(\top1.memory1.mem2[138][1] ));
 sg13g2_dfrbp_1 _20202_ (.CLK(\clknet_leaf_60_top1.acquisition_clk ),
    .RESET_B(net973),
    .D(_00403_),
    .Q_N(_09576_),
    .Q(\top1.memory1.mem2[138][2] ));
 sg13g2_dfrbp_1 _20203_ (.CLK(\clknet_leaf_69_top1.acquisition_clk ),
    .RESET_B(net972),
    .D(_00404_),
    .Q_N(_09575_),
    .Q(\top1.memory1.mem2[137][0] ));
 sg13g2_dfrbp_1 _20204_ (.CLK(\clknet_leaf_69_top1.acquisition_clk ),
    .RESET_B(net971),
    .D(_00405_),
    .Q_N(_09574_),
    .Q(\top1.memory1.mem2[137][1] ));
 sg13g2_dfrbp_1 _20205_ (.CLK(\clknet_leaf_67_top1.acquisition_clk ),
    .RESET_B(net970),
    .D(_00406_),
    .Q_N(_09573_),
    .Q(\top1.memory1.mem2[137][2] ));
 sg13g2_dfrbp_1 _20206_ (.CLK(\clknet_leaf_74_top1.acquisition_clk ),
    .RESET_B(net969),
    .D(_00407_),
    .Q_N(_09572_),
    .Q(\top1.memory1.mem2[136][0] ));
 sg13g2_dfrbp_1 _20207_ (.CLK(\clknet_leaf_60_top1.acquisition_clk ),
    .RESET_B(net968),
    .D(_00408_),
    .Q_N(_09571_),
    .Q(\top1.memory1.mem2[136][1] ));
 sg13g2_dfrbp_1 _20208_ (.CLK(\clknet_leaf_60_top1.acquisition_clk ),
    .RESET_B(net967),
    .D(_00409_),
    .Q_N(_09570_),
    .Q(\top1.memory1.mem2[136][2] ));
 sg13g2_dfrbp_1 _20209_ (.CLK(\clknet_leaf_55_top1.acquisition_clk ),
    .RESET_B(net966),
    .D(_00410_),
    .Q_N(_09569_),
    .Q(\top1.memory1.mem2[135][0] ));
 sg13g2_dfrbp_1 _20210_ (.CLK(\clknet_leaf_61_top1.acquisition_clk ),
    .RESET_B(net965),
    .D(_00411_),
    .Q_N(_09568_),
    .Q(\top1.memory1.mem2[135][1] ));
 sg13g2_dfrbp_1 _20211_ (.CLK(\clknet_leaf_60_top1.acquisition_clk ),
    .RESET_B(net964),
    .D(_00412_),
    .Q_N(_09567_),
    .Q(\top1.memory1.mem2[135][2] ));
 sg13g2_dfrbp_1 _20212_ (.CLK(\clknet_leaf_222_top1.acquisition_clk ),
    .RESET_B(net963),
    .D(_00413_),
    .Q_N(_09566_),
    .Q(\top1.memory1.mem2[116][0] ));
 sg13g2_dfrbp_1 _20213_ (.CLK(\clknet_leaf_228_top1.acquisition_clk ),
    .RESET_B(net962),
    .D(_00414_),
    .Q_N(_09565_),
    .Q(\top1.memory1.mem2[116][1] ));
 sg13g2_dfrbp_1 _20214_ (.CLK(\clknet_leaf_223_top1.acquisition_clk ),
    .RESET_B(net961),
    .D(_00415_),
    .Q_N(_09564_),
    .Q(\top1.memory1.mem2[116][2] ));
 sg13g2_dfrbp_1 _20215_ (.CLK(\clknet_leaf_83_top1.acquisition_clk ),
    .RESET_B(net960),
    .D(_00416_),
    .Q_N(_09563_),
    .Q(\top1.memory1.mem2[12][0] ));
 sg13g2_dfrbp_1 _20216_ (.CLK(\clknet_leaf_83_top1.acquisition_clk ),
    .RESET_B(net959),
    .D(_00417_),
    .Q_N(_09562_),
    .Q(\top1.memory1.mem2[12][1] ));
 sg13g2_dfrbp_1 _20217_ (.CLK(\clknet_leaf_82_top1.acquisition_clk ),
    .RESET_B(net958),
    .D(_00418_),
    .Q_N(_09561_),
    .Q(\top1.memory1.mem2[12][2] ));
 sg13g2_dfrbp_1 _20218_ (.CLK(\clknet_leaf_212_top1.acquisition_clk ),
    .RESET_B(net957),
    .D(_00419_),
    .Q_N(_09560_),
    .Q(\top1.memory1.mem2[115][0] ));
 sg13g2_dfrbp_1 _20219_ (.CLK(\clknet_leaf_208_top1.acquisition_clk ),
    .RESET_B(net956),
    .D(_00420_),
    .Q_N(_09559_),
    .Q(\top1.memory1.mem2[115][1] ));
 sg13g2_dfrbp_1 _20220_ (.CLK(\clknet_leaf_200_top1.acquisition_clk ),
    .RESET_B(net955),
    .D(_00421_),
    .Q_N(_09558_),
    .Q(\top1.memory1.mem2[115][2] ));
 sg13g2_dfrbp_1 _20221_ (.CLK(\clknet_leaf_212_top1.acquisition_clk ),
    .RESET_B(net954),
    .D(_00422_),
    .Q_N(_09557_),
    .Q(\top1.memory1.mem2[114][0] ));
 sg13g2_dfrbp_1 _20222_ (.CLK(\clknet_leaf_210_top1.acquisition_clk ),
    .RESET_B(net953),
    .D(_00423_),
    .Q_N(_09556_),
    .Q(\top1.memory1.mem2[114][1] ));
 sg13g2_dfrbp_1 _20223_ (.CLK(\clknet_leaf_196_top1.acquisition_clk ),
    .RESET_B(net952),
    .D(_00424_),
    .Q_N(_09555_),
    .Q(\top1.memory1.mem2[114][2] ));
 sg13g2_dfrbp_1 _20224_ (.CLK(\clknet_leaf_65_top1.acquisition_clk ),
    .RESET_B(net951),
    .D(_00425_),
    .Q_N(_09554_),
    .Q(\top1.memory1.mem2[128][0] ));
 sg13g2_dfrbp_1 _20225_ (.CLK(\clknet_leaf_65_top1.acquisition_clk ),
    .RESET_B(net950),
    .D(_00426_),
    .Q_N(_09553_),
    .Q(\top1.memory1.mem2[128][1] ));
 sg13g2_dfrbp_1 _20226_ (.CLK(\clknet_leaf_65_top1.acquisition_clk ),
    .RESET_B(net949),
    .D(_00427_),
    .Q_N(_09552_),
    .Q(\top1.memory1.mem2[128][2] ));
 sg13g2_dfrbp_1 _20227_ (.CLK(\clknet_leaf_213_top1.acquisition_clk ),
    .RESET_B(net948),
    .D(_00428_),
    .Q_N(_09551_),
    .Q(\top1.memory1.mem2[113][0] ));
 sg13g2_dfrbp_1 _20228_ (.CLK(\clknet_leaf_210_top1.acquisition_clk ),
    .RESET_B(net947),
    .D(_00429_),
    .Q_N(_09550_),
    .Q(\top1.memory1.mem2[113][1] ));
 sg13g2_dfrbp_1 _20229_ (.CLK(\clknet_leaf_196_top1.acquisition_clk ),
    .RESET_B(net946),
    .D(_00430_),
    .Q_N(_09549_),
    .Q(\top1.memory1.mem2[113][2] ));
 sg13g2_dfrbp_1 _20230_ (.CLK(\clknet_leaf_213_top1.acquisition_clk ),
    .RESET_B(net945),
    .D(_00431_),
    .Q_N(_09548_),
    .Q(\top1.memory1.mem2[112][0] ));
 sg13g2_dfrbp_1 _20231_ (.CLK(\clknet_leaf_210_top1.acquisition_clk ),
    .RESET_B(net944),
    .D(_00432_),
    .Q_N(_09547_),
    .Q(\top1.memory1.mem2[112][1] ));
 sg13g2_dfrbp_1 _20232_ (.CLK(\clknet_leaf_200_top1.acquisition_clk ),
    .RESET_B(net943),
    .D(_00433_),
    .Q_N(_09546_),
    .Q(\top1.memory1.mem2[112][2] ));
 sg13g2_dfrbp_1 _20233_ (.CLK(\clknet_leaf_229_top1.acquisition_clk ),
    .RESET_B(net942),
    .D(_00434_),
    .Q_N(_09545_),
    .Q(\top1.memory1.mem2[127][0] ));
 sg13g2_dfrbp_1 _20234_ (.CLK(\clknet_leaf_227_top1.acquisition_clk ),
    .RESET_B(net941),
    .D(_00435_),
    .Q_N(_09544_),
    .Q(\top1.memory1.mem2[127][1] ));
 sg13g2_dfrbp_1 _20235_ (.CLK(\clknet_leaf_224_top1.acquisition_clk ),
    .RESET_B(net940),
    .D(_00436_),
    .Q_N(_09543_),
    .Q(\top1.memory1.mem2[127][2] ));
 sg13g2_dfrbp_1 _20236_ (.CLK(\clknet_leaf_226_top1.acquisition_clk ),
    .RESET_B(net939),
    .D(_00437_),
    .Q_N(_09542_),
    .Q(\top1.memory1.mem2[111][0] ));
 sg13g2_dfrbp_1 _20237_ (.CLK(\clknet_leaf_234_top1.acquisition_clk ),
    .RESET_B(net938),
    .D(_00438_),
    .Q_N(_09541_),
    .Q(\top1.memory1.mem2[111][1] ));
 sg13g2_dfrbp_1 _20238_ (.CLK(\clknet_leaf_229_top1.acquisition_clk ),
    .RESET_B(net937),
    .D(_00439_),
    .Q_N(_09540_),
    .Q(\top1.memory1.mem2[111][2] ));
 sg13g2_dfrbp_1 _20239_ (.CLK(\clknet_leaf_226_top1.acquisition_clk ),
    .RESET_B(net936),
    .D(_00440_),
    .Q_N(_09539_),
    .Q(\top1.memory1.mem2[110][0] ));
 sg13g2_dfrbp_1 _20240_ (.CLK(\clknet_leaf_234_top1.acquisition_clk ),
    .RESET_B(net934),
    .D(_00441_),
    .Q_N(_09538_),
    .Q(\top1.memory1.mem2[110][1] ));
 sg13g2_dfrbp_1 _20241_ (.CLK(\clknet_leaf_225_top1.acquisition_clk ),
    .RESET_B(net933),
    .D(_00442_),
    .Q_N(_09537_),
    .Q(\top1.memory1.mem2[110][2] ));
 sg13g2_dfrbp_1 _20242_ (.CLK(\clknet_leaf_229_top1.acquisition_clk ),
    .RESET_B(net932),
    .D(_00443_),
    .Q_N(_09536_),
    .Q(\top1.memory1.mem2[126][0] ));
 sg13g2_dfrbp_1 _20243_ (.CLK(\clknet_leaf_227_top1.acquisition_clk ),
    .RESET_B(net931),
    .D(_00444_),
    .Q_N(_09535_),
    .Q(\top1.memory1.mem2[126][1] ));
 sg13g2_dfrbp_1 _20244_ (.CLK(\clknet_leaf_224_top1.acquisition_clk ),
    .RESET_B(net930),
    .D(_00445_),
    .Q_N(_09534_),
    .Q(\top1.memory1.mem2[126][2] ));
 sg13g2_dfrbp_1 _20245_ (.CLK(\clknet_leaf_86_top1.acquisition_clk ),
    .RESET_B(net929),
    .D(_00446_),
    .Q_N(_09533_),
    .Q(\top1.memory1.mem2[10][0] ));
 sg13g2_dfrbp_1 _20246_ (.CLK(\clknet_leaf_85_top1.acquisition_clk ),
    .RESET_B(net928),
    .D(_00447_),
    .Q_N(_09532_),
    .Q(\top1.memory1.mem2[10][1] ));
 sg13g2_dfrbp_1 _20247_ (.CLK(\clknet_leaf_94_top1.acquisition_clk ),
    .RESET_B(net927),
    .D(_00448_),
    .Q_N(_09531_),
    .Q(\top1.memory1.mem2[10][2] ));
 sg13g2_dfrbp_1 _20248_ (.CLK(\clknet_leaf_226_top1.acquisition_clk ),
    .RESET_B(net926),
    .D(_00449_),
    .Q_N(_09530_),
    .Q(\top1.memory1.mem2[108][0] ));
 sg13g2_dfrbp_1 _20249_ (.CLK(\clknet_leaf_233_top1.acquisition_clk ),
    .RESET_B(net925),
    .D(_00450_),
    .Q_N(_09529_),
    .Q(\top1.memory1.mem2[108][1] ));
 sg13g2_dfrbp_1 _20250_ (.CLK(\clknet_leaf_225_top1.acquisition_clk ),
    .RESET_B(net924),
    .D(_00451_),
    .Q_N(_09528_),
    .Q(\top1.memory1.mem2[108][2] ));
 sg13g2_dfrbp_1 _20251_ (.CLK(\clknet_leaf_228_top1.acquisition_clk ),
    .RESET_B(net923),
    .D(_00452_),
    .Q_N(_09527_),
    .Q(\top1.memory1.mem2[125][0] ));
 sg13g2_dfrbp_1 _20252_ (.CLK(\clknet_leaf_227_top1.acquisition_clk ),
    .RESET_B(net922),
    .D(_00453_),
    .Q_N(_09526_),
    .Q(\top1.memory1.mem2[125][1] ));
 sg13g2_dfrbp_1 _20253_ (.CLK(\clknet_leaf_225_top1.acquisition_clk ),
    .RESET_B(net921),
    .D(_00454_),
    .Q_N(_09525_),
    .Q(\top1.memory1.mem2[125][2] ));
 sg13g2_dfrbp_1 _20254_ (.CLK(\clknet_leaf_211_top1.acquisition_clk ),
    .RESET_B(net920),
    .D(_00455_),
    .Q_N(_09524_),
    .Q(\top1.memory1.mem2[107][0] ));
 sg13g2_dfrbp_1 _20255_ (.CLK(\clknet_leaf_193_top1.acquisition_clk ),
    .RESET_B(net919),
    .D(_00456_),
    .Q_N(_09523_),
    .Q(\top1.memory1.mem2[107][1] ));
 sg13g2_dfrbp_1 _20256_ (.CLK(\clknet_leaf_229_top1.acquisition_clk ),
    .RESET_B(net918),
    .D(_00457_),
    .Q_N(_09522_),
    .Q(\top1.memory1.mem2[107][2] ));
 sg13g2_dfrbp_1 _20257_ (.CLK(\clknet_leaf_211_top1.acquisition_clk ),
    .RESET_B(net917),
    .D(_00458_),
    .Q_N(_09521_),
    .Q(\top1.memory1.mem2[106][0] ));
 sg13g2_dfrbp_1 _20258_ (.CLK(\clknet_leaf_193_top1.acquisition_clk ),
    .RESET_B(net916),
    .D(_00459_),
    .Q_N(_09520_),
    .Q(\top1.memory1.mem2[106][1] ));
 sg13g2_dfrbp_1 _20259_ (.CLK(\clknet_leaf_229_top1.acquisition_clk ),
    .RESET_B(net915),
    .D(_00460_),
    .Q_N(_09519_),
    .Q(\top1.memory1.mem2[106][2] ));
 sg13g2_dfrbp_1 _20260_ (.CLK(\clknet_leaf_229_top1.acquisition_clk ),
    .RESET_B(net914),
    .D(_00461_),
    .Q_N(_09518_),
    .Q(\top1.memory1.mem2[124][0] ));
 sg13g2_dfrbp_1 _20261_ (.CLK(\clknet_leaf_227_top1.acquisition_clk ),
    .RESET_B(net913),
    .D(_00462_),
    .Q_N(_09517_),
    .Q(\top1.memory1.mem2[124][1] ));
 sg13g2_dfrbp_1 _20262_ (.CLK(\clknet_leaf_224_top1.acquisition_clk ),
    .RESET_B(net912),
    .D(_00463_),
    .Q_N(_09516_),
    .Q(\top1.memory1.mem2[124][2] ));
 sg13g2_dfrbp_1 _20263_ (.CLK(\clknet_leaf_211_top1.acquisition_clk ),
    .RESET_B(net911),
    .D(_00464_),
    .Q_N(_09515_),
    .Q(\top1.memory1.mem2[105][0] ));
 sg13g2_dfrbp_1 _20264_ (.CLK(\clknet_leaf_252_top1.acquisition_clk ),
    .RESET_B(net910),
    .D(_00465_),
    .Q_N(_09514_),
    .Q(\top1.memory1.mem2[105][1] ));
 sg13g2_dfrbp_1 _20265_ (.CLK(\clknet_leaf_229_top1.acquisition_clk ),
    .RESET_B(net909),
    .D(_00466_),
    .Q_N(_09513_),
    .Q(\top1.memory1.mem2[105][2] ));
 sg13g2_dfrbp_1 _20266_ (.CLK(\clknet_leaf_230_top1.acquisition_clk ),
    .RESET_B(net908),
    .D(_00467_),
    .Q_N(_09512_),
    .Q(\top1.memory1.mem2[104][0] ));
 sg13g2_dfrbp_1 _20267_ (.CLK(\clknet_leaf_193_top1.acquisition_clk ),
    .RESET_B(net907),
    .D(_00468_),
    .Q_N(_09511_),
    .Q(\top1.memory1.mem2[104][1] ));
 sg13g2_dfrbp_1 _20268_ (.CLK(\clknet_leaf_229_top1.acquisition_clk ),
    .RESET_B(net906),
    .D(_00469_),
    .Q_N(_09510_),
    .Q(\top1.memory1.mem2[104][2] ));
 sg13g2_dfrbp_1 _20269_ (.CLK(\clknet_leaf_211_top1.acquisition_clk ),
    .RESET_B(net905),
    .D(_00470_),
    .Q_N(_09509_),
    .Q(\top1.memory1.mem2[123][0] ));
 sg13g2_dfrbp_1 _20270_ (.CLK(\clknet_leaf_194_top1.acquisition_clk ),
    .RESET_B(net903),
    .D(_00471_),
    .Q_N(_09508_),
    .Q(\top1.memory1.mem2[123][1] ));
 sg13g2_dfrbp_1 _20271_ (.CLK(\clknet_leaf_195_top1.acquisition_clk ),
    .RESET_B(net902),
    .D(_00472_),
    .Q_N(_09507_),
    .Q(\top1.memory1.mem2[123][2] ));
 sg13g2_dfrbp_1 _20272_ (.CLK(\clknet_leaf_236_top1.acquisition_clk ),
    .RESET_B(net901),
    .D(_00473_),
    .Q_N(_09506_),
    .Q(\top1.memory1.mem2[103][0] ));
 sg13g2_dfrbp_1 _20273_ (.CLK(\clknet_leaf_232_top1.acquisition_clk ),
    .RESET_B(net900),
    .D(_00474_),
    .Q_N(_09505_),
    .Q(\top1.memory1.mem2[103][1] ));
 sg13g2_dfrbp_1 _20274_ (.CLK(\clknet_leaf_236_top1.acquisition_clk ),
    .RESET_B(net899),
    .D(_00475_),
    .Q_N(_09504_),
    .Q(\top1.memory1.mem2[103][2] ));
 sg13g2_dfrbp_1 _20275_ (.CLK(\clknet_leaf_235_top1.acquisition_clk ),
    .RESET_B(net898),
    .D(_00476_),
    .Q_N(_09503_),
    .Q(\top1.memory1.mem2[102][0] ));
 sg13g2_dfrbp_1 _20276_ (.CLK(\clknet_leaf_232_top1.acquisition_clk ),
    .RESET_B(net897),
    .D(_00477_),
    .Q_N(_09502_),
    .Q(\top1.memory1.mem2[102][1] ));
 sg13g2_dfrbp_1 _20277_ (.CLK(\clknet_leaf_236_top1.acquisition_clk ),
    .RESET_B(net896),
    .D(_00478_),
    .Q_N(_09501_),
    .Q(\top1.memory1.mem2[102][2] ));
 sg13g2_dfrbp_1 _20278_ (.CLK(\clknet_leaf_235_top1.acquisition_clk ),
    .RESET_B(net895),
    .D(_00479_),
    .Q_N(_09500_),
    .Q(\top1.memory1.mem2[101][0] ));
 sg13g2_dfrbp_1 _20279_ (.CLK(\clknet_leaf_233_top1.acquisition_clk ),
    .RESET_B(net894),
    .D(_00480_),
    .Q_N(_09499_),
    .Q(\top1.memory1.mem2[101][1] ));
 sg13g2_dfrbp_1 _20280_ (.CLK(\clknet_leaf_236_top1.acquisition_clk ),
    .RESET_B(net893),
    .D(_00481_),
    .Q_N(_09498_),
    .Q(\top1.memory1.mem2[101][2] ));
 sg13g2_dfrbp_1 _20281_ (.CLK(\clknet_leaf_65_top1.acquisition_clk ),
    .RESET_B(net892),
    .D(_00482_),
    .Q_N(_09497_),
    .Q(\top1.memory1.mem2[130][0] ));
 sg13g2_dfrbp_1 _20282_ (.CLK(\clknet_leaf_66_top1.acquisition_clk ),
    .RESET_B(net891),
    .D(_00483_),
    .Q_N(_09496_),
    .Q(\top1.memory1.mem2[130][1] ));
 sg13g2_dfrbp_1 _20283_ (.CLK(\clknet_leaf_67_top1.acquisition_clk ),
    .RESET_B(net890),
    .D(_00484_),
    .Q_N(_09495_),
    .Q(\top1.memory1.mem2[130][2] ));
 sg13g2_dfrbp_1 _20284_ (.CLK(\clknet_leaf_236_top1.acquisition_clk ),
    .RESET_B(net889),
    .D(_00485_),
    .Q_N(_09494_),
    .Q(\top1.memory1.mem2[100][0] ));
 sg13g2_dfrbp_1 _20285_ (.CLK(\clknet_leaf_237_top1.acquisition_clk ),
    .RESET_B(net888),
    .D(_00486_),
    .Q_N(_09493_),
    .Q(\top1.memory1.mem2[100][1] ));
 sg13g2_dfrbp_1 _20286_ (.CLK(\clknet_leaf_236_top1.acquisition_clk ),
    .RESET_B(net887),
    .D(_00487_),
    .Q_N(_09492_),
    .Q(\top1.memory1.mem2[100][2] ));
 sg13g2_dfrbp_1 _20287_ (.CLK(\clknet_leaf_87_top1.acquisition_clk ),
    .RESET_B(net886),
    .D(_00488_),
    .Q_N(_09491_),
    .Q(\top1.memory1.mem2[0][0] ));
 sg13g2_dfrbp_1 _20288_ (.CLK(\clknet_leaf_89_top1.acquisition_clk ),
    .RESET_B(net885),
    .D(_00489_),
    .Q_N(_09490_),
    .Q(\top1.memory1.mem2[0][1] ));
 sg13g2_dfrbp_1 _20289_ (.CLK(\clknet_leaf_91_top1.acquisition_clk ),
    .RESET_B(net884),
    .D(_00490_),
    .Q_N(_09489_),
    .Q(\top1.memory1.mem2[0][2] ));
 sg13g2_dfrbp_1 _20290_ (.CLK(\clknet_leaf_64_top1.acquisition_clk ),
    .RESET_B(net883),
    .D(_00491_),
    .Q_N(_09488_),
    .Q(\top1.memory1.mem2[131][0] ));
 sg13g2_dfrbp_1 _20291_ (.CLK(\clknet_leaf_68_top1.acquisition_clk ),
    .RESET_B(net882),
    .D(_00492_),
    .Q_N(_09487_),
    .Q(\top1.memory1.mem2[131][1] ));
 sg13g2_dfrbp_1 _20292_ (.CLK(\clknet_leaf_67_top1.acquisition_clk ),
    .RESET_B(net881),
    .D(_00493_),
    .Q_N(_09486_),
    .Q(\top1.memory1.mem2[131][2] ));
 sg13g2_dfrbp_1 _20293_ (.CLK(\clknet_leaf_251_top1.acquisition_clk ),
    .RESET_B(net880),
    .D(_00494_),
    .Q_N(_09485_),
    .Q(\top1.memory1.mem2[98][0] ));
 sg13g2_dfrbp_1 _20294_ (.CLK(\clknet_leaf_251_top1.acquisition_clk ),
    .RESET_B(net879),
    .D(_00495_),
    .Q_N(_09484_),
    .Q(\top1.memory1.mem2[98][1] ));
 sg13g2_dfrbp_1 _20295_ (.CLK(\clknet_leaf_249_top1.acquisition_clk ),
    .RESET_B(net878),
    .D(_00496_),
    .Q_N(_09483_),
    .Q(\top1.memory1.mem2[98][2] ));
 sg13g2_dfrbp_1 _20296_ (.CLK(\clknet_leaf_6_top1.acquisition_clk ),
    .RESET_B(net877),
    .D(_00497_),
    .Q_N(_09482_),
    .Q(\top1.memory1.mem2[68][0] ));
 sg13g2_dfrbp_1 _20297_ (.CLK(\clknet_leaf_7_top1.acquisition_clk ),
    .RESET_B(net876),
    .D(_00498_),
    .Q_N(_09481_),
    .Q(\top1.memory1.mem2[68][1] ));
 sg13g2_dfrbp_1 _20298_ (.CLK(\clknet_leaf_7_top1.acquisition_clk ),
    .RESET_B(net875),
    .D(_00499_),
    .Q_N(_09480_),
    .Q(\top1.memory1.mem2[68][2] ));
 sg13g2_dfrbp_1 _20299_ (.CLK(\clknet_leaf_298_top1.acquisition_clk ),
    .RESET_B(net874),
    .D(_00500_),
    .Q_N(_09479_),
    .Q(\top1.memory1.mem2[67][0] ));
 sg13g2_dfrbp_1 _20300_ (.CLK(\clknet_leaf_1_top1.acquisition_clk ),
    .RESET_B(net873),
    .D(_00501_),
    .Q_N(_09478_),
    .Q(\top1.memory1.mem2[67][1] ));
 sg13g2_dfrbp_1 _20301_ (.CLK(\clknet_leaf_300_top1.acquisition_clk ),
    .RESET_B(net872),
    .D(_00502_),
    .Q_N(_09477_),
    .Q(\top1.memory1.mem2[67][2] ));
 sg13g2_dfrbp_1 _20302_ (.CLK(\clknet_leaf_285_top1.acquisition_clk ),
    .RESET_B(net871),
    .D(_00503_),
    .Q_N(_09476_),
    .Q(\top1.memory1.mem2[94][0] ));
 sg13g2_dfrbp_1 _20303_ (.CLK(\clknet_leaf_286_top1.acquisition_clk ),
    .RESET_B(net870),
    .D(_00504_),
    .Q_N(_09475_),
    .Q(\top1.memory1.mem2[94][1] ));
 sg13g2_dfrbp_1 _20304_ (.CLK(\clknet_leaf_289_top1.acquisition_clk ),
    .RESET_B(net869),
    .D(_00505_),
    .Q_N(_09474_),
    .Q(\top1.memory1.mem2[94][2] ));
 sg13g2_dfrbp_1 _20305_ (.CLK(\clknet_leaf_299_top1.acquisition_clk ),
    .RESET_B(net868),
    .D(_00506_),
    .Q_N(_09473_),
    .Q(\top1.memory1.mem2[66][0] ));
 sg13g2_dfrbp_1 _20306_ (.CLK(\clknet_leaf_0_top1.acquisition_clk ),
    .RESET_B(net867),
    .D(_00507_),
    .Q_N(_09472_),
    .Q(\top1.memory1.mem2[66][1] ));
 sg13g2_dfrbp_1 _20307_ (.CLK(\clknet_leaf_300_top1.acquisition_clk ),
    .RESET_B(net866),
    .D(_00508_),
    .Q_N(_09471_),
    .Q(\top1.memory1.mem2[66][2] ));
 sg13g2_dfrbp_1 _20308_ (.CLK(\clknet_leaf_299_top1.acquisition_clk ),
    .RESET_B(net865),
    .D(_00509_),
    .Q_N(_09470_),
    .Q(\top1.memory1.mem2[65][0] ));
 sg13g2_dfrbp_1 _20309_ (.CLK(\clknet_leaf_0_top1.acquisition_clk ),
    .RESET_B(net864),
    .D(_00510_),
    .Q_N(_09469_),
    .Q(\top1.memory1.mem2[65][1] ));
 sg13g2_dfrbp_1 _20310_ (.CLK(\clknet_leaf_300_top1.acquisition_clk ),
    .RESET_B(net863),
    .D(_00511_),
    .Q_N(_09468_),
    .Q(\top1.memory1.mem2[65][2] ));
 sg13g2_dfrbp_1 _20311_ (.CLK(\clknet_leaf_285_top1.acquisition_clk ),
    .RESET_B(net862),
    .D(_00512_),
    .Q_N(_09467_),
    .Q(\top1.memory1.mem2[93][0] ));
 sg13g2_dfrbp_1 _20312_ (.CLK(\clknet_leaf_286_top1.acquisition_clk ),
    .RESET_B(net861),
    .D(_00513_),
    .Q_N(_09466_),
    .Q(\top1.memory1.mem2[93][1] ));
 sg13g2_dfrbp_1 _20313_ (.CLK(\clknet_leaf_290_top1.acquisition_clk ),
    .RESET_B(net860),
    .D(_00514_),
    .Q_N(_09465_),
    .Q(\top1.memory1.mem2[93][2] ));
 sg13g2_dfrbp_1 _20314_ (.CLK(\clknet_leaf_299_top1.acquisition_clk ),
    .RESET_B(net859),
    .D(_00515_),
    .Q_N(_09464_),
    .Q(\top1.memory1.mem2[64][0] ));
 sg13g2_dfrbp_1 _20315_ (.CLK(\clknet_leaf_0_top1.acquisition_clk ),
    .RESET_B(net858),
    .D(_00516_),
    .Q_N(_09463_),
    .Q(\top1.memory1.mem2[64][1] ));
 sg13g2_dfrbp_1 _20316_ (.CLK(\clknet_leaf_299_top1.acquisition_clk ),
    .RESET_B(net857),
    .D(_00517_),
    .Q_N(_09462_),
    .Q(\top1.memory1.mem2[64][2] ));
 sg13g2_dfrbp_1 _20317_ (.CLK(\clknet_leaf_149_top1.acquisition_clk ),
    .RESET_B(net856),
    .D(_00518_),
    .Q_N(_09461_),
    .Q(\top1.memory1.mem2[63][0] ));
 sg13g2_dfrbp_1 _20318_ (.CLK(\clknet_leaf_146_top1.acquisition_clk ),
    .RESET_B(net855),
    .D(_00519_),
    .Q_N(_09460_),
    .Q(\top1.memory1.mem2[63][1] ));
 sg13g2_dfrbp_1 _20319_ (.CLK(\clknet_leaf_146_top1.acquisition_clk ),
    .RESET_B(net854),
    .D(_00520_),
    .Q_N(_09459_),
    .Q(\top1.memory1.mem2[63][2] ));
 sg13g2_dfrbp_1 _20320_ (.CLK(\clknet_leaf_285_top1.acquisition_clk ),
    .RESET_B(net853),
    .D(_00521_),
    .Q_N(_09458_),
    .Q(\top1.memory1.mem2[92][0] ));
 sg13g2_dfrbp_1 _20321_ (.CLK(\clknet_leaf_294_top1.acquisition_clk ),
    .RESET_B(net852),
    .D(_00522_),
    .Q_N(_09457_),
    .Q(\top1.memory1.mem2[92][1] ));
 sg13g2_dfrbp_1 _20322_ (.CLK(\clknet_leaf_289_top1.acquisition_clk ),
    .RESET_B(net851),
    .D(_00523_),
    .Q_N(_09456_),
    .Q(\top1.memory1.mem2[92][2] ));
 sg13g2_dfrbp_1 _20323_ (.CLK(\clknet_leaf_144_top1.acquisition_clk ),
    .RESET_B(net850),
    .D(_00524_),
    .Q_N(_09455_),
    .Q(\top1.memory1.mem2[62][0] ));
 sg13g2_dfrbp_1 _20324_ (.CLK(\clknet_leaf_145_top1.acquisition_clk ),
    .RESET_B(net849),
    .D(_00525_),
    .Q_N(_09454_),
    .Q(\top1.memory1.mem2[62][1] ));
 sg13g2_dfrbp_1 _20325_ (.CLK(\clknet_leaf_146_top1.acquisition_clk ),
    .RESET_B(net848),
    .D(_00526_),
    .Q_N(_09453_),
    .Q(\top1.memory1.mem2[62][2] ));
 sg13g2_dfrbp_1 _20326_ (.CLK(\clknet_leaf_139_top1.acquisition_clk ),
    .RESET_B(net847),
    .D(_00527_),
    .Q_N(_09452_),
    .Q(\top1.memory1.mem2[61][0] ));
 sg13g2_dfrbp_1 _20327_ (.CLK(\clknet_leaf_145_top1.acquisition_clk ),
    .RESET_B(net846),
    .D(_00528_),
    .Q_N(_09451_),
    .Q(\top1.memory1.mem2[61][1] ));
 sg13g2_dfrbp_1 _20328_ (.CLK(\clknet_leaf_144_top1.acquisition_clk ),
    .RESET_B(net845),
    .D(_00529_),
    .Q_N(_09450_),
    .Q(\top1.memory1.mem2[61][2] ));
 sg13g2_dfrbp_1 _20329_ (.CLK(\clknet_leaf_9_top1.acquisition_clk ),
    .RESET_B(net844),
    .D(_00530_),
    .Q_N(_09449_),
    .Q(\top1.memory1.mem2[91][0] ));
 sg13g2_dfrbp_1 _20330_ (.CLK(\clknet_leaf_293_top1.acquisition_clk ),
    .RESET_B(net843),
    .D(_00531_),
    .Q_N(_09448_),
    .Q(\top1.memory1.mem2[91][1] ));
 sg13g2_dfrbp_1 _20331_ (.CLK(\clknet_leaf_28_top1.acquisition_clk ),
    .RESET_B(net842),
    .D(_00532_),
    .Q_N(_09447_),
    .Q(\top1.memory1.mem2[91][2] ));
 sg13g2_dfrbp_1 _20332_ (.CLK(\clknet_leaf_140_top1.acquisition_clk ),
    .RESET_B(net841),
    .D(_00533_),
    .Q_N(_09446_),
    .Q(\top1.memory1.mem2[60][0] ));
 sg13g2_dfrbp_1 _20333_ (.CLK(\clknet_leaf_146_top1.acquisition_clk ),
    .RESET_B(net840),
    .D(_00534_),
    .Q_N(_09445_),
    .Q(\top1.memory1.mem2[60][1] ));
 sg13g2_dfrbp_1 _20334_ (.CLK(\clknet_leaf_144_top1.acquisition_clk ),
    .RESET_B(net839),
    .D(_00535_),
    .Q_N(_09444_),
    .Q(\top1.memory1.mem2[60][2] ));
 sg13g2_dfrbp_1 _20335_ (.CLK(\clknet_leaf_100_top1.acquisition_clk ),
    .RESET_B(net838),
    .D(_00536_),
    .Q_N(_09443_),
    .Q(\top1.memory1.mem2[5][0] ));
 sg13g2_dfrbp_1 _20336_ (.CLK(\clknet_leaf_93_top1.acquisition_clk ),
    .RESET_B(net837),
    .D(_00537_),
    .Q_N(_09442_),
    .Q(\top1.memory1.mem2[5][1] ));
 sg13g2_dfrbp_1 _20337_ (.CLK(\clknet_leaf_94_top1.acquisition_clk ),
    .RESET_B(net836),
    .D(_00538_),
    .Q_N(_09441_),
    .Q(\top1.memory1.mem2[5][2] ));
 sg13g2_dfrbp_1 _20338_ (.CLK(\clknet_leaf_290_top1.acquisition_clk ),
    .RESET_B(net835),
    .D(_00539_),
    .Q_N(_09440_),
    .Q(\top1.memory1.mem2[90][0] ));
 sg13g2_dfrbp_1 _20339_ (.CLK(\clknet_leaf_293_top1.acquisition_clk ),
    .RESET_B(net834),
    .D(_00540_),
    .Q_N(_09439_),
    .Q(\top1.memory1.mem2[90][1] ));
 sg13g2_dfrbp_1 _20340_ (.CLK(\clknet_leaf_9_top1.acquisition_clk ),
    .RESET_B(net833),
    .D(_00541_),
    .Q_N(_09438_),
    .Q(\top1.memory1.mem2[90][2] ));
 sg13g2_dfrbp_1 _20341_ (.CLK(\clknet_leaf_168_top1.acquisition_clk ),
    .RESET_B(net832),
    .D(_00542_),
    .Q_N(_09437_),
    .Q(\top1.memory1.mem2[58][0] ));
 sg13g2_dfrbp_1 _20342_ (.CLK(\clknet_leaf_173_top1.acquisition_clk ),
    .RESET_B(net831),
    .D(_00543_),
    .Q_N(_09436_),
    .Q(\top1.memory1.mem2[58][1] ));
 sg13g2_dfrbp_1 _20343_ (.CLK(\clknet_leaf_157_top1.acquisition_clk ),
    .RESET_B(net830),
    .D(_00544_),
    .Q_N(_09435_),
    .Q(\top1.memory1.mem2[58][2] ));
 sg13g2_dfrbp_1 _20344_ (.CLK(\clknet_leaf_173_top1.acquisition_clk ),
    .RESET_B(net829),
    .D(_00545_),
    .Q_N(_09434_),
    .Q(\top1.memory1.mem2[57][0] ));
 sg13g2_dfrbp_1 _20345_ (.CLK(\clknet_leaf_172_top1.acquisition_clk ),
    .RESET_B(net828),
    .D(_00546_),
    .Q_N(_09433_),
    .Q(\top1.memory1.mem2[57][1] ));
 sg13g2_dfrbp_1 _20346_ (.CLK(\clknet_leaf_157_top1.acquisition_clk ),
    .RESET_B(net827),
    .D(_00547_),
    .Q_N(_09432_),
    .Q(\top1.memory1.mem2[57][2] ));
 sg13g2_dfrbp_1 _20347_ (.CLK(\clknet_leaf_86_top1.acquisition_clk ),
    .RESET_B(net826),
    .D(_00548_),
    .Q_N(_09431_),
    .Q(\top1.memory1.mem2[8][0] ));
 sg13g2_dfrbp_1 _20348_ (.CLK(\clknet_leaf_85_top1.acquisition_clk ),
    .RESET_B(net825),
    .D(_00549_),
    .Q_N(_09430_),
    .Q(\top1.memory1.mem2[8][1] ));
 sg13g2_dfrbp_1 _20349_ (.CLK(\clknet_leaf_90_top1.acquisition_clk ),
    .RESET_B(net824),
    .D(_00550_),
    .Q_N(_09429_),
    .Q(\top1.memory1.mem2[8][2] ));
 sg13g2_dfrbp_1 _20350_ (.CLK(\clknet_leaf_172_top1.acquisition_clk ),
    .RESET_B(net823),
    .D(_00551_),
    .Q_N(_09428_),
    .Q(\top1.memory1.mem2[56][0] ));
 sg13g2_dfrbp_1 _20351_ (.CLK(\clknet_leaf_173_top1.acquisition_clk ),
    .RESET_B(net822),
    .D(_00552_),
    .Q_N(_09427_),
    .Q(\top1.memory1.mem2[56][1] ));
 sg13g2_dfrbp_1 _20352_ (.CLK(\clknet_leaf_157_top1.acquisition_clk ),
    .RESET_B(net821),
    .D(_00553_),
    .Q_N(_09426_),
    .Q(\top1.memory1.mem2[56][2] ));
 sg13g2_dfrbp_1 _20353_ (.CLK(\clknet_leaf_154_top1.acquisition_clk ),
    .RESET_B(net820),
    .D(_00554_),
    .Q_N(_09425_),
    .Q(\top1.memory1.mem2[55][0] ));
 sg13g2_dfrbp_1 _20354_ (.CLK(\clknet_leaf_154_top1.acquisition_clk ),
    .RESET_B(net819),
    .D(_00555_),
    .Q_N(_09424_),
    .Q(\top1.memory1.mem2[55][1] ));
 sg13g2_dfrbp_1 _20355_ (.CLK(\clknet_leaf_139_top1.acquisition_clk ),
    .RESET_B(net818),
    .D(_00556_),
    .Q_N(_09423_),
    .Q(\top1.memory1.mem2[55][2] ));
 sg13g2_dfrbp_1 _20356_ (.CLK(\clknet_leaf_8_top1.acquisition_clk ),
    .RESET_B(net817),
    .D(_00557_),
    .Q_N(_09422_),
    .Q(\top1.memory1.mem2[88][0] ));
 sg13g2_dfrbp_1 _20357_ (.CLK(\clknet_leaf_292_top1.acquisition_clk ),
    .RESET_B(net816),
    .D(_00558_),
    .Q_N(_09421_),
    .Q(\top1.memory1.mem2[88][1] ));
 sg13g2_dfrbp_1 _20358_ (.CLK(\clknet_leaf_9_top1.acquisition_clk ),
    .RESET_B(net815),
    .D(_00559_),
    .Q_N(_09420_),
    .Q(\top1.memory1.mem2[88][2] ));
 sg13g2_dfrbp_1 _20359_ (.CLK(\clknet_leaf_154_top1.acquisition_clk ),
    .RESET_B(net814),
    .D(_00560_),
    .Q_N(_09419_),
    .Q(\top1.memory1.mem2[54][0] ));
 sg13g2_dfrbp_1 _20360_ (.CLK(\clknet_leaf_154_top1.acquisition_clk ),
    .RESET_B(net813),
    .D(_00561_),
    .Q_N(_09418_),
    .Q(\top1.memory1.mem2[54][1] ));
 sg13g2_dfrbp_1 _20361_ (.CLK(\clknet_leaf_138_top1.acquisition_clk ),
    .RESET_B(net812),
    .D(_00562_),
    .Q_N(_09417_),
    .Q(\top1.memory1.mem2[54][2] ));
 sg13g2_dfrbp_1 _20362_ (.CLK(\clknet_leaf_154_top1.acquisition_clk ),
    .RESET_B(net811),
    .D(_00563_),
    .Q_N(_09416_),
    .Q(\top1.memory1.mem2[53][0] ));
 sg13g2_dfrbp_1 _20363_ (.CLK(\clknet_leaf_137_top1.acquisition_clk ),
    .RESET_B(net810),
    .D(_00564_),
    .Q_N(_09415_),
    .Q(\top1.memory1.mem2[53][1] ));
 sg13g2_dfrbp_1 _20364_ (.CLK(\clknet_leaf_138_top1.acquisition_clk ),
    .RESET_B(net809),
    .D(_00565_),
    .Q_N(_09414_),
    .Q(\top1.memory1.mem2[53][2] ));
 sg13g2_dfrbp_1 _20365_ (.CLK(\clknet_leaf_27_top1.acquisition_clk ),
    .RESET_B(net808),
    .D(_00566_),
    .Q_N(_09413_),
    .Q(\top1.memory1.mem2[87][0] ));
 sg13g2_dfrbp_1 _20366_ (.CLK(\clknet_leaf_32_top1.acquisition_clk ),
    .RESET_B(net807),
    .D(_00567_),
    .Q_N(_09412_),
    .Q(\top1.memory1.mem2[87][1] ));
 sg13g2_dfrbp_1 _20367_ (.CLK(\clknet_leaf_27_top1.acquisition_clk ),
    .RESET_B(net806),
    .D(_00568_),
    .Q_N(_09411_),
    .Q(\top1.memory1.mem2[87][2] ));
 sg13g2_dfrbp_1 _20368_ (.CLK(\clknet_leaf_139_top1.acquisition_clk ),
    .RESET_B(net805),
    .D(_00569_),
    .Q_N(_09410_),
    .Q(\top1.memory1.mem2[52][0] ));
 sg13g2_dfrbp_1 _20369_ (.CLK(\clknet_leaf_154_top1.acquisition_clk ),
    .RESET_B(net804),
    .D(_00570_),
    .Q_N(_09409_),
    .Q(\top1.memory1.mem2[52][1] ));
 sg13g2_dfrbp_1 _20370_ (.CLK(\clknet_leaf_139_top1.acquisition_clk ),
    .RESET_B(net803),
    .D(_00571_),
    .Q_N(_09408_),
    .Q(\top1.memory1.mem2[52][2] ));
 sg13g2_dfrbp_1 _20371_ (.CLK(\clknet_leaf_144_top1.acquisition_clk ),
    .RESET_B(net802),
    .D(_00572_),
    .Q_N(_09407_),
    .Q(\top1.memory1.mem2[51][0] ));
 sg13g2_dfrbp_1 _20372_ (.CLK(\clknet_leaf_141_top1.acquisition_clk ),
    .RESET_B(net801),
    .D(_00573_),
    .Q_N(_09406_),
    .Q(\top1.memory1.mem2[51][1] ));
 sg13g2_dfrbp_1 _20373_ (.CLK(\clknet_leaf_140_top1.acquisition_clk ),
    .RESET_B(net800),
    .D(_00574_),
    .Q_N(_09405_),
    .Q(\top1.memory1.mem2[51][2] ));
 sg13g2_dfrbp_1 _20374_ (.CLK(\clknet_leaf_27_top1.acquisition_clk ),
    .RESET_B(net799),
    .D(_00575_),
    .Q_N(_09404_),
    .Q(\top1.memory1.mem2[86][0] ));
 sg13g2_dfrbp_1 _20375_ (.CLK(\clknet_leaf_29_top1.acquisition_clk ),
    .RESET_B(net798),
    .D(_00576_),
    .Q_N(_09403_),
    .Q(\top1.memory1.mem2[86][1] ));
 sg13g2_dfrbp_1 _20376_ (.CLK(\clknet_leaf_27_top1.acquisition_clk ),
    .RESET_B(net797),
    .D(_00577_),
    .Q_N(_09402_),
    .Q(\top1.memory1.mem2[86][2] ));
 sg13g2_dfrbp_1 _20377_ (.CLK(\clknet_leaf_140_top1.acquisition_clk ),
    .RESET_B(net796),
    .D(_00578_),
    .Q_N(_09401_),
    .Q(\top1.memory1.mem2[50][0] ));
 sg13g2_dfrbp_1 _20378_ (.CLK(\clknet_leaf_143_top1.acquisition_clk ),
    .RESET_B(net795),
    .D(_00579_),
    .Q_N(_09400_),
    .Q(\top1.memory1.mem2[50][1] ));
 sg13g2_dfrbp_1 _20379_ (.CLK(\clknet_leaf_143_top1.acquisition_clk ),
    .RESET_B(net794),
    .D(_00580_),
    .Q_N(_09399_),
    .Q(\top1.memory1.mem2[50][2] ));
 sg13g2_dfrbp_1 _20380_ (.CLK(\clknet_leaf_100_top1.acquisition_clk ),
    .RESET_B(net793),
    .D(_00581_),
    .Q_N(_09398_),
    .Q(\top1.memory1.mem2[4][0] ));
 sg13g2_dfrbp_1 _20381_ (.CLK(\clknet_leaf_93_top1.acquisition_clk ),
    .RESET_B(net792),
    .D(_00582_),
    .Q_N(_09397_),
    .Q(\top1.memory1.mem2[4][1] ));
 sg13g2_dfrbp_1 _20382_ (.CLK(\clknet_leaf_94_top1.acquisition_clk ),
    .RESET_B(net791),
    .D(_00583_),
    .Q_N(_09396_),
    .Q(\top1.memory1.mem2[4][2] ));
 sg13g2_dfrbp_1 _20383_ (.CLK(\clknet_leaf_28_top1.acquisition_clk ),
    .RESET_B(net790),
    .D(_00584_),
    .Q_N(_09395_),
    .Q(\top1.memory1.mem2[85][0] ));
 sg13g2_dfrbp_1 _20384_ (.CLK(\clknet_leaf_29_top1.acquisition_clk ),
    .RESET_B(net789),
    .D(_00585_),
    .Q_N(_09394_),
    .Q(\top1.memory1.mem2[85][1] ));
 sg13g2_dfrbp_1 _20385_ (.CLK(\clknet_leaf_27_top1.acquisition_clk ),
    .RESET_B(net788),
    .D(_00586_),
    .Q_N(_09393_),
    .Q(\top1.memory1.mem2[85][2] ));
 sg13g2_dfrbp_1 _20386_ (.CLK(\clknet_leaf_141_top1.acquisition_clk ),
    .RESET_B(net787),
    .D(_00587_),
    .Q_N(_09392_),
    .Q(\top1.memory1.mem2[44][0] ));
 sg13g2_dfrbp_1 _20387_ (.CLK(\clknet_leaf_142_top1.acquisition_clk ),
    .RESET_B(net786),
    .D(_00588_),
    .Q_N(_09391_),
    .Q(\top1.memory1.mem2[44][1] ));
 sg13g2_dfrbp_1 _20388_ (.CLK(\clknet_leaf_132_top1.acquisition_clk ),
    .RESET_B(net785),
    .D(_00589_),
    .Q_N(_09390_),
    .Q(\top1.memory1.mem2[44][2] ));
 sg13g2_dfrbp_1 _20389_ (.CLK(\clknet_leaf_137_top1.acquisition_clk ),
    .RESET_B(net784),
    .D(_00590_),
    .Q_N(_09389_),
    .Q(\top1.memory1.mem2[43][0] ));
 sg13g2_dfrbp_1 _20390_ (.CLK(\clknet_leaf_154_top1.acquisition_clk ),
    .RESET_B(net783),
    .D(_00591_),
    .Q_N(_09388_),
    .Q(\top1.memory1.mem2[43][1] ));
 sg13g2_dfrbp_1 _20391_ (.CLK(\clknet_leaf_173_top1.acquisition_clk ),
    .RESET_B(net782),
    .D(_00592_),
    .Q_N(_09387_),
    .Q(\top1.memory1.mem2[43][2] ));
 sg13g2_dfrbp_1 _20392_ (.CLK(\clknet_leaf_138_top1.acquisition_clk ),
    .RESET_B(net781),
    .D(_00593_),
    .Q_N(_09386_),
    .Q(\top1.memory1.mem2[46][0] ));
 sg13g2_dfrbp_1 _20393_ (.CLK(\clknet_leaf_141_top1.acquisition_clk ),
    .RESET_B(net780),
    .D(_00594_),
    .Q_N(_09385_),
    .Q(\top1.memory1.mem2[46][1] ));
 sg13g2_dfrbp_1 _20394_ (.CLK(\clknet_leaf_132_top1.acquisition_clk ),
    .RESET_B(net779),
    .D(_00595_),
    .Q_N(_09384_),
    .Q(\top1.memory1.mem2[46][2] ));
 sg13g2_dfrbp_1 _20395_ (.CLK(\clknet_leaf_137_top1.acquisition_clk ),
    .RESET_B(net778),
    .D(_00596_),
    .Q_N(_09383_),
    .Q(\top1.memory1.mem2[42][0] ));
 sg13g2_dfrbp_1 _20396_ (.CLK(\clknet_leaf_155_top1.acquisition_clk ),
    .RESET_B(net777),
    .D(_00597_),
    .Q_N(_09382_),
    .Q(\top1.memory1.mem2[42][1] ));
 sg13g2_dfrbp_1 _20397_ (.CLK(\clknet_leaf_174_top1.acquisition_clk ),
    .RESET_B(net776),
    .D(_00598_),
    .Q_N(_09381_),
    .Q(\top1.memory1.mem2[42][2] ));
 sg13g2_dfrbp_1 _20398_ (.CLK(\clknet_leaf_116_top1.acquisition_clk ),
    .RESET_B(net775),
    .D(_00599_),
    .Q_N(_09380_),
    .Q(\top1.memory1.mem2[38][0] ));
 sg13g2_dfrbp_1 _20399_ (.CLK(\clknet_leaf_135_top1.acquisition_clk ),
    .RESET_B(net774),
    .D(_00600_),
    .Q_N(_09379_),
    .Q(\top1.memory1.mem2[38][1] ));
 sg13g2_dfrbp_1 _20400_ (.CLK(\clknet_leaf_131_top1.acquisition_clk ),
    .RESET_B(net773),
    .D(_00601_),
    .Q_N(_09378_),
    .Q(\top1.memory1.mem2[38][2] ));
 sg13g2_dfrbp_1 _20401_ (.CLK(\clknet_leaf_138_top1.acquisition_clk ),
    .RESET_B(net772),
    .D(_00602_),
    .Q_N(_09377_),
    .Q(\top1.memory1.mem2[40][0] ));
 sg13g2_dfrbp_1 _20402_ (.CLK(\clknet_leaf_137_top1.acquisition_clk ),
    .RESET_B(net771),
    .D(_00603_),
    .Q_N(_09376_),
    .Q(\top1.memory1.mem2[40][1] ));
 sg13g2_dfrbp_1 _20403_ (.CLK(\clknet_leaf_174_top1.acquisition_clk ),
    .RESET_B(net770),
    .D(_00604_),
    .Q_N(_09375_),
    .Q(\top1.memory1.mem2[40][2] ));
 sg13g2_dfrbp_1 _20404_ (.CLK(\clknet_leaf_7_top1.acquisition_clk ),
    .RESET_B(net769),
    .D(_00605_),
    .Q_N(_09374_),
    .Q(\top1.memory1.mem2[69][0] ));
 sg13g2_dfrbp_1 _20405_ (.CLK(\clknet_leaf_8_top1.acquisition_clk ),
    .RESET_B(net768),
    .D(_00606_),
    .Q_N(_09373_),
    .Q(\top1.memory1.mem2[69][1] ));
 sg13g2_dfrbp_1 _20406_ (.CLK(\clknet_leaf_7_top1.acquisition_clk ),
    .RESET_B(net767),
    .D(_00607_),
    .Q_N(_09372_),
    .Q(\top1.memory1.mem2[69][2] ));
 sg13g2_dfrbp_1 _20407_ (.CLK(\clknet_leaf_158_top1.acquisition_clk ),
    .RESET_B(net766),
    .D(_00608_),
    .Q_N(_09371_),
    .Q(\top1.memory1.mem2[59][0] ));
 sg13g2_dfrbp_1 _20408_ (.CLK(\clknet_leaf_173_top1.acquisition_clk ),
    .RESET_B(net765),
    .D(_00609_),
    .Q_N(_09370_),
    .Q(\top1.memory1.mem2[59][1] ));
 sg13g2_dfrbp_1 _20409_ (.CLK(\clknet_leaf_157_top1.acquisition_clk ),
    .RESET_B(net764),
    .D(_00610_),
    .Q_N(_09369_),
    .Q(\top1.memory1.mem2[59][2] ));
 sg13g2_dfrbp_1 _20410_ (.CLK(\clknet_leaf_126_top1.acquisition_clk ),
    .RESET_B(net763),
    .D(_00611_),
    .Q_N(_09368_),
    .Q(\top1.memory1.mem2[26][0] ));
 sg13g2_dfrbp_1 _20411_ (.CLK(\clknet_leaf_126_top1.acquisition_clk ),
    .RESET_B(net762),
    .D(_00612_),
    .Q_N(_09367_),
    .Q(\top1.memory1.mem2[26][1] ));
 sg13g2_dfrbp_1 _20412_ (.CLK(\clknet_leaf_124_top1.acquisition_clk ),
    .RESET_B(net761),
    .D(_00613_),
    .Q_N(_09366_),
    .Q(\top1.memory1.mem2[26][2] ));
 sg13g2_dfrbp_1 _20413_ (.CLK(\clknet_leaf_140_top1.acquisition_clk ),
    .RESET_B(net760),
    .D(_00614_),
    .Q_N(_09365_),
    .Q(\top1.memory1.mem2[49][0] ));
 sg13g2_dfrbp_1 _20414_ (.CLK(\clknet_leaf_141_top1.acquisition_clk ),
    .RESET_B(net759),
    .D(_00615_),
    .Q_N(_09364_),
    .Q(\top1.memory1.mem2[49][1] ));
 sg13g2_dfrbp_1 _20415_ (.CLK(\clknet_leaf_143_top1.acquisition_clk ),
    .RESET_B(net758),
    .D(_00616_),
    .Q_N(_09363_),
    .Q(\top1.memory1.mem2[49][2] ));
 sg13g2_dfrbp_1 _20416_ (.CLK(\clknet_leaf_175_top1.acquisition_clk ),
    .RESET_B(net757),
    .D(_00617_),
    .Q_N(_09362_),
    .Q(\top1.memory1.mem2[39][0] ));
 sg13g2_dfrbp_1 _20417_ (.CLK(\clknet_leaf_136_top1.acquisition_clk ),
    .RESET_B(net756),
    .D(_00618_),
    .Q_N(_09361_),
    .Q(\top1.memory1.mem2[39][1] ));
 sg13g2_dfrbp_1 _20418_ (.CLK(\clknet_leaf_131_top1.acquisition_clk ),
    .RESET_B(net755),
    .D(_00619_),
    .Q_N(_09360_),
    .Q(\top1.memory1.mem2[39][2] ));
 sg13g2_dfrbp_1 _20419_ (.CLK(\clknet_leaf_125_top1.acquisition_clk ),
    .RESET_B(net754),
    .D(_00620_),
    .Q_N(_09359_),
    .Q(\top1.memory1.mem2[25][0] ));
 sg13g2_dfrbp_1 _20420_ (.CLK(\clknet_leaf_126_top1.acquisition_clk ),
    .RESET_B(net753),
    .D(_00621_),
    .Q_N(_09358_),
    .Q(\top1.memory1.mem2[25][1] ));
 sg13g2_dfrbp_1 _20421_ (.CLK(\clknet_leaf_123_top1.acquisition_clk ),
    .RESET_B(net752),
    .D(_00622_),
    .Q_N(_09357_),
    .Q(\top1.memory1.mem2[25][2] ));
 sg13g2_dfrbp_1 _20422_ (.CLK(\clknet_leaf_124_top1.acquisition_clk ),
    .RESET_B(net751),
    .D(_00623_),
    .Q_N(_09356_),
    .Q(\top1.memory1.mem2[29][0] ));
 sg13g2_dfrbp_1 _20423_ (.CLK(\clknet_leaf_125_top1.acquisition_clk ),
    .RESET_B(net750),
    .D(_00624_),
    .Q_N(_09355_),
    .Q(\top1.memory1.mem2[29][1] ));
 sg13g2_dfrbp_1 _20424_ (.CLK(\clknet_leaf_87_top1.acquisition_clk ),
    .RESET_B(net749),
    .D(_00625_),
    .Q_N(_09354_),
    .Q(\top1.memory1.mem2[29][2] ));
 sg13g2_dfrbp_1 _20425_ (.CLK(\clknet_leaf_119_top1.acquisition_clk ),
    .RESET_B(net748),
    .D(_00626_),
    .Q_N(_09353_),
    .Q(\top1.memory1.mem2[19][0] ));
 sg13g2_dfrbp_1 _20426_ (.CLK(\clknet_leaf_123_top1.acquisition_clk ),
    .RESET_B(net747),
    .D(_00627_),
    .Q_N(_09352_),
    .Q(\top1.memory1.mem2[19][1] ));
 sg13g2_dfrbp_1 _20427_ (.CLK(\clknet_leaf_123_top1.acquisition_clk ),
    .RESET_B(net746),
    .D(_00628_),
    .Q_N(_09351_),
    .Q(\top1.memory1.mem2[19][2] ));
 sg13g2_dfrbp_1 _20428_ (.CLK(\clknet_leaf_126_top1.acquisition_clk ),
    .RESET_B(net745),
    .D(_00629_),
    .Q_N(_09350_),
    .Q(\top1.memory1.mem2[24][0] ));
 sg13g2_dfrbp_1 _20429_ (.CLK(\clknet_leaf_125_top1.acquisition_clk ),
    .RESET_B(net744),
    .D(_00630_),
    .Q_N(_09349_),
    .Q(\top1.memory1.mem2[24][1] ));
 sg13g2_dfrbp_1 _20430_ (.CLK(\clknet_leaf_125_top1.acquisition_clk ),
    .RESET_B(net743),
    .D(_00631_),
    .Q_N(_09348_),
    .Q(\top1.memory1.mem2[24][2] ));
 sg13g2_dfrbp_1 _20431_ (.CLK(\clknet_leaf_265_top1.acquisition_clk ),
    .RESET_B(net742),
    .D(_00632_),
    .Q_N(_09347_),
    .Q(\top1.memory1.mem1[9][0] ));
 sg13g2_dfrbp_1 _20432_ (.CLK(\clknet_leaf_265_top1.acquisition_clk ),
    .RESET_B(net741),
    .D(_00633_),
    .Q_N(_09346_),
    .Q(\top1.memory1.mem1[9][1] ));
 sg13g2_dfrbp_1 _20433_ (.CLK(\clknet_leaf_276_top1.acquisition_clk ),
    .RESET_B(net740),
    .D(_00634_),
    .Q_N(_09345_),
    .Q(\top1.memory1.mem1[9][2] ));
 sg13g2_dfrbp_1 _20434_ (.CLK(\clknet_leaf_121_top1.acquisition_clk ),
    .RESET_B(net739),
    .D(_00635_),
    .Q_N(_09344_),
    .Q(\top1.memory1.mem2[23][0] ));
 sg13g2_dfrbp_1 _20435_ (.CLK(\clknet_leaf_121_top1.acquisition_clk ),
    .RESET_B(net738),
    .D(_00636_),
    .Q_N(_09343_),
    .Q(\top1.memory1.mem2[23][1] ));
 sg13g2_dfrbp_1 _20436_ (.CLK(\clknet_leaf_122_top1.acquisition_clk ),
    .RESET_B(net737),
    .D(_00637_),
    .Q_N(_09342_),
    .Q(\top1.memory1.mem2[23][2] ));
 sg13g2_dfrbp_1 _20437_ (.CLK(\clknet_leaf_121_top1.acquisition_clk ),
    .RESET_B(net736),
    .D(_00638_),
    .Q_N(_09341_),
    .Q(\top1.memory1.mem2[22][0] ));
 sg13g2_dfrbp_1 _20438_ (.CLK(\clknet_leaf_120_top1.acquisition_clk ),
    .RESET_B(net735),
    .D(_00639_),
    .Q_N(_09340_),
    .Q(\top1.memory1.mem2[22][1] ));
 sg13g2_dfrbp_1 _20439_ (.CLK(\clknet_leaf_121_top1.acquisition_clk ),
    .RESET_B(net734),
    .D(_00640_),
    .Q_N(_09339_),
    .Q(\top1.memory1.mem2[22][2] ));
 sg13g2_dfrbp_1 _20440_ (.CLK(\clknet_leaf_121_top1.acquisition_clk ),
    .RESET_B(net733),
    .D(_00641_),
    .Q_N(_09338_),
    .Q(\top1.memory1.mem2[21][0] ));
 sg13g2_dfrbp_1 _20441_ (.CLK(\clknet_leaf_121_top1.acquisition_clk ),
    .RESET_B(net732),
    .D(_00642_),
    .Q_N(_09337_),
    .Q(\top1.memory1.mem2[21][1] ));
 sg13g2_dfrbp_1 _20442_ (.CLK(\clknet_leaf_122_top1.acquisition_clk ),
    .RESET_B(net731),
    .D(_00643_),
    .Q_N(_09336_),
    .Q(\top1.memory1.mem2[21][2] ));
 sg13g2_dfrbp_1 _20443_ (.CLK(\clknet_leaf_55_top1.acquisition_clk ),
    .RESET_B(net730),
    .D(_00644_),
    .Q_N(_09335_),
    .Q(\top1.memory1.mem2[134][0] ));
 sg13g2_dfrbp_1 _20444_ (.CLK(\clknet_leaf_62_top1.acquisition_clk ),
    .RESET_B(net729),
    .D(_00645_),
    .Q_N(_09334_),
    .Q(\top1.memory1.mem2[134][1] ));
 sg13g2_dfrbp_1 _20445_ (.CLK(\clknet_leaf_74_top1.acquisition_clk ),
    .RESET_B(net728),
    .D(_00646_),
    .Q_N(_09333_),
    .Q(\top1.memory1.mem2[134][2] ));
 sg13g2_dfrbp_1 _20446_ (.CLK(\clknet_leaf_55_top1.acquisition_clk ),
    .RESET_B(net727),
    .D(_00647_),
    .Q_N(_09332_),
    .Q(\top1.memory1.mem2[133][0] ));
 sg13g2_dfrbp_1 _20447_ (.CLK(\clknet_leaf_55_top1.acquisition_clk ),
    .RESET_B(net726),
    .D(_00648_),
    .Q_N(_09331_),
    .Q(\top1.memory1.mem2[133][1] ));
 sg13g2_dfrbp_1 _20448_ (.CLK(\clknet_leaf_61_top1.acquisition_clk ),
    .RESET_B(net725),
    .D(_00649_),
    .Q_N(_09330_),
    .Q(\top1.memory1.mem2[133][2] ));
 sg13g2_dfrbp_1 _20449_ (.CLK(\clknet_leaf_62_top1.acquisition_clk ),
    .RESET_B(net724),
    .D(_00650_),
    .Q_N(_09329_),
    .Q(\top1.memory1.mem2[132][0] ));
 sg13g2_dfrbp_1 _20450_ (.CLK(\clknet_leaf_61_top1.acquisition_clk ),
    .RESET_B(net723),
    .D(_00651_),
    .Q_N(_09328_),
    .Q(\top1.memory1.mem2[132][1] ));
 sg13g2_dfrbp_1 _20451_ (.CLK(\clknet_leaf_68_top1.acquisition_clk ),
    .RESET_B(net722),
    .D(_00652_),
    .Q_N(_09327_),
    .Q(\top1.memory1.mem2[132][2] ));
 sg13g2_dfrbp_1 _20452_ (.CLK(\clknet_leaf_28_top1.acquisition_clk ),
    .RESET_B(net721),
    .D(_00653_),
    .Q_N(_09326_),
    .Q(\top1.memory1.mem2[84][0] ));
 sg13g2_dfrbp_1 _20453_ (.CLK(\clknet_leaf_29_top1.acquisition_clk ),
    .RESET_B(net720),
    .D(_00654_),
    .Q_N(_09325_),
    .Q(\top1.memory1.mem2[84][1] ));
 sg13g2_dfrbp_1 _20454_ (.CLK(\clknet_leaf_28_top1.acquisition_clk ),
    .RESET_B(net719),
    .D(_00655_),
    .Q_N(_09324_),
    .Q(\top1.memory1.mem2[84][2] ));
 sg13g2_dfrbp_1 _20455_ (.CLK(\clknet_leaf_294_top1.acquisition_clk ),
    .RESET_B(net718),
    .D(_00656_),
    .Q_N(_09323_),
    .Q(\top1.memory1.mem2[83][0] ));
 sg13g2_dfrbp_1 _20456_ (.CLK(\clknet_leaf_295_top1.acquisition_clk ),
    .RESET_B(net717),
    .D(_00657_),
    .Q_N(_09322_),
    .Q(\top1.memory1.mem2[83][1] ));
 sg13g2_dfrbp_1 _20457_ (.CLK(\clknet_leaf_295_top1.acquisition_clk ),
    .RESET_B(net716),
    .D(_00658_),
    .Q_N(_09321_),
    .Q(\top1.memory1.mem2[83][2] ));
 sg13g2_dfrbp_1 _20458_ (.CLK(\clknet_leaf_141_top1.acquisition_clk ),
    .RESET_B(net715),
    .D(_00659_),
    .Q_N(_09320_),
    .Q(\top1.memory1.mem2[47][0] ));
 sg13g2_dfrbp_1 _20459_ (.CLK(\clknet_leaf_142_top1.acquisition_clk ),
    .RESET_B(net714),
    .D(_00660_),
    .Q_N(_09319_),
    .Q(\top1.memory1.mem2[47][1] ));
 sg13g2_dfrbp_1 _20460_ (.CLK(\clknet_leaf_132_top1.acquisition_clk ),
    .RESET_B(net713),
    .D(_00661_),
    .Q_N(_09318_),
    .Q(\top1.memory1.mem2[47][2] ));
 sg13g2_dfrbp_1 _20461_ (.CLK(\clknet_leaf_138_top1.acquisition_clk ),
    .RESET_B(net712),
    .D(_00662_),
    .Q_N(_09317_),
    .Q(\top1.memory1.mem2[41][0] ));
 sg13g2_dfrbp_1 _20462_ (.CLK(\clknet_leaf_137_top1.acquisition_clk ),
    .RESET_B(net711),
    .D(_00663_),
    .Q_N(_09316_),
    .Q(\top1.memory1.mem2[41][1] ));
 sg13g2_dfrbp_1 _20463_ (.CLK(\clknet_leaf_174_top1.acquisition_clk ),
    .RESET_B(net710),
    .D(_00664_),
    .Q_N(_09315_),
    .Q(\top1.memory1.mem2[41][2] ));
 sg13g2_dfrbp_1 _20464_ (.CLK(\clknet_leaf_140_top1.acquisition_clk ),
    .RESET_B(net709),
    .D(_00665_),
    .Q_N(_09314_),
    .Q(\top1.memory1.mem2[48][0] ));
 sg13g2_dfrbp_1 _20465_ (.CLK(\clknet_leaf_142_top1.acquisition_clk ),
    .RESET_B(net708),
    .D(_00666_),
    .Q_N(_09313_),
    .Q(\top1.memory1.mem2[48][1] ));
 sg13g2_dfrbp_1 _20466_ (.CLK(\clknet_leaf_143_top1.acquisition_clk ),
    .RESET_B(net707),
    .D(_00667_),
    .Q_N(_09312_),
    .Q(\top1.memory1.mem2[48][2] ));
 sg13g2_dfrbp_1 _20467_ (.CLK(\clknet_leaf_120_top1.acquisition_clk ),
    .RESET_B(net706),
    .D(_00668_),
    .Q_N(_09311_),
    .Q(\top1.memory1.mem2[20][0] ));
 sg13g2_dfrbp_1 _20468_ (.CLK(\clknet_leaf_120_top1.acquisition_clk ),
    .RESET_B(net705),
    .D(_00669_),
    .Q_N(_09310_),
    .Q(\top1.memory1.mem2[20][1] ));
 sg13g2_dfrbp_1 _20469_ (.CLK(\clknet_leaf_122_top1.acquisition_clk ),
    .RESET_B(net704),
    .D(_00670_),
    .Q_N(_09309_),
    .Q(\top1.memory1.mem2[20][2] ));
 sg13g2_dfrbp_1 _20470_ (.CLK(\clknet_leaf_137_top1.acquisition_clk ),
    .RESET_B(net703),
    .D(_00671_),
    .Q_N(_09308_),
    .Q(\top1.memory1.mem2[37][0] ));
 sg13g2_dfrbp_1 _20471_ (.CLK(\clknet_leaf_132_top1.acquisition_clk ),
    .RESET_B(net702),
    .D(_00672_),
    .Q_N(_09307_),
    .Q(\top1.memory1.mem2[37][1] ));
 sg13g2_dfrbp_1 _20472_ (.CLK(\clknet_leaf_131_top1.acquisition_clk ),
    .RESET_B(net701),
    .D(_00673_),
    .Q_N(_09306_),
    .Q(\top1.memory1.mem2[37][2] ));
 sg13g2_dfrbp_1 _20473_ (.CLK(\clknet_leaf_270_top1.acquisition_clk ),
    .RESET_B(net700),
    .D(_00674_),
    .Q_N(_09305_),
    .Q(\top1.memory1.mem1[92][0] ));
 sg13g2_dfrbp_1 _20474_ (.CLK(\clknet_leaf_283_top1.acquisition_clk ),
    .RESET_B(net699),
    .D(_00675_),
    .Q_N(_09304_),
    .Q(\top1.memory1.mem1[92][1] ));
 sg13g2_dfrbp_1 _20475_ (.CLK(\clknet_leaf_288_top1.acquisition_clk ),
    .RESET_B(net698),
    .D(_00676_),
    .Q_N(_09303_),
    .Q(\top1.memory1.mem1[92][2] ));
 sg13g2_dfrbp_1 _20476_ (.CLK(\clknet_leaf_270_top1.acquisition_clk ),
    .RESET_B(net697),
    .D(_00677_),
    .Q_N(_09302_),
    .Q(\top1.memory1.mem1[93][0] ));
 sg13g2_dfrbp_1 _20477_ (.CLK(\clknet_leaf_283_top1.acquisition_clk ),
    .RESET_B(net696),
    .D(_00678_),
    .Q_N(_09301_),
    .Q(\top1.memory1.mem1[93][1] ));
 sg13g2_dfrbp_1 _20478_ (.CLK(\clknet_leaf_288_top1.acquisition_clk ),
    .RESET_B(net695),
    .D(_00679_),
    .Q_N(_09300_),
    .Q(\top1.memory1.mem1[93][2] ));
 sg13g2_dfrbp_1 _20479_ (.CLK(\clknet_leaf_270_top1.acquisition_clk ),
    .RESET_B(net694),
    .D(_00680_),
    .Q_N(_09299_),
    .Q(\top1.memory1.mem1[94][0] ));
 sg13g2_dfrbp_1 _20480_ (.CLK(\clknet_leaf_283_top1.acquisition_clk ),
    .RESET_B(net693),
    .D(_00681_),
    .Q_N(_09298_),
    .Q(\top1.memory1.mem1[94][1] ));
 sg13g2_dfrbp_1 _20481_ (.CLK(\clknet_leaf_282_top1.acquisition_clk ),
    .RESET_B(net692),
    .D(_00682_),
    .Q_N(_09297_),
    .Q(\top1.memory1.mem1[94][2] ));
 sg13g2_dfrbp_1 _20482_ (.CLK(\clknet_leaf_271_top1.acquisition_clk ),
    .RESET_B(net691),
    .D(_00683_),
    .Q_N(_09296_),
    .Q(\top1.memory1.mem1[95][0] ));
 sg13g2_dfrbp_1 _20483_ (.CLK(\clknet_leaf_283_top1.acquisition_clk ),
    .RESET_B(net690),
    .D(_00684_),
    .Q_N(_09295_),
    .Q(\top1.memory1.mem1[95][1] ));
 sg13g2_dfrbp_1 _20484_ (.CLK(\clknet_leaf_282_top1.acquisition_clk ),
    .RESET_B(net689),
    .D(_00685_),
    .Q_N(_09294_),
    .Q(\top1.memory1.mem1[95][2] ));
 sg13g2_dfrbp_1 _20485_ (.CLK(\clknet_leaf_242_top1.acquisition_clk ),
    .RESET_B(net688),
    .D(_00686_),
    .Q_N(_09293_),
    .Q(\top1.memory1.mem1[169][0] ));
 sg13g2_dfrbp_1 _20486_ (.CLK(\clknet_leaf_242_top1.acquisition_clk ),
    .RESET_B(net687),
    .D(_00687_),
    .Q_N(_09292_),
    .Q(\top1.memory1.mem1[169][1] ));
 sg13g2_dfrbp_1 _20487_ (.CLK(\clknet_leaf_264_top1.acquisition_clk ),
    .RESET_B(net686),
    .D(_00688_),
    .Q_N(_09291_),
    .Q(\top1.memory1.mem1[169][2] ));
 sg13g2_dfrbp_1 _20488_ (.CLK(\clknet_leaf_268_top1.acquisition_clk ),
    .RESET_B(net685),
    .D(_00689_),
    .Q_N(_09290_),
    .Q(\top1.memory1.mem1[91][0] ));
 sg13g2_dfrbp_1 _20489_ (.CLK(\clknet_leaf_284_top1.acquisition_clk ),
    .RESET_B(net684),
    .D(_00690_),
    .Q_N(_09289_),
    .Q(\top1.memory1.mem1[91][1] ));
 sg13g2_dfrbp_1 _20490_ (.CLK(\clknet_leaf_288_top1.acquisition_clk ),
    .RESET_B(net683),
    .D(_00691_),
    .Q_N(_09288_),
    .Q(\top1.memory1.mem1[91][2] ));
 sg13g2_dfrbp_1 _20491_ (.CLK(\clknet_leaf_270_top1.acquisition_clk ),
    .RESET_B(net682),
    .D(_00692_),
    .Q_N(_09287_),
    .Q(\top1.memory1.mem1[90][0] ));
 sg13g2_dfrbp_1 _20492_ (.CLK(\clknet_leaf_284_top1.acquisition_clk ),
    .RESET_B(net681),
    .D(_00693_),
    .Q_N(_09286_),
    .Q(\top1.memory1.mem1[90][1] ));
 sg13g2_dfrbp_1 _20493_ (.CLK(\clknet_leaf_270_top1.acquisition_clk ),
    .RESET_B(net680),
    .D(_00694_),
    .Q_N(_09285_),
    .Q(\top1.memory1.mem1[90][2] ));
 sg13g2_dfrbp_1 _20494_ (.CLK(\clknet_leaf_22_top1.acquisition_clk ),
    .RESET_B(net679),
    .D(_00695_),
    .Q_N(_09284_),
    .Q(\top1.memory1.mem1[149][0] ));
 sg13g2_dfrbp_1 _20495_ (.CLK(\clknet_leaf_22_top1.acquisition_clk ),
    .RESET_B(net678),
    .D(_00696_),
    .Q_N(_09283_),
    .Q(\top1.memory1.mem1[149][1] ));
 sg13g2_dfrbp_1 _20496_ (.CLK(\clknet_leaf_24_top1.acquisition_clk ),
    .RESET_B(net677),
    .D(_00697_),
    .Q_N(_09282_),
    .Q(\top1.memory1.mem1[149][2] ));
 sg13g2_dfrbp_1 _20497_ (.CLK(\clknet_leaf_285_top1.acquisition_clk ),
    .RESET_B(net676),
    .D(_00698_),
    .Q_N(_09281_),
    .Q(\top1.memory1.mem1[82][0] ));
 sg13g2_dfrbp_1 _20498_ (.CLK(\clknet_leaf_289_top1.acquisition_clk ),
    .RESET_B(net675),
    .D(_00699_),
    .Q_N(_09280_),
    .Q(\top1.memory1.mem1[82][1] ));
 sg13g2_dfrbp_1 _20499_ (.CLK(\clknet_leaf_287_top1.acquisition_clk ),
    .RESET_B(net674),
    .D(_00700_),
    .Q_N(_09279_),
    .Q(\top1.memory1.mem1[82][2] ));
 sg13g2_dfrbp_1 _20500_ (.CLK(\clknet_leaf_286_top1.acquisition_clk ),
    .RESET_B(net673),
    .D(_00701_),
    .Q_N(_09278_),
    .Q(\top1.memory1.mem1[83][0] ));
 sg13g2_dfrbp_1 _20501_ (.CLK(\clknet_leaf_289_top1.acquisition_clk ),
    .RESET_B(net672),
    .D(_00702_),
    .Q_N(_09277_),
    .Q(\top1.memory1.mem1[83][1] ));
 sg13g2_dfrbp_1 _20502_ (.CLK(\clknet_leaf_287_top1.acquisition_clk ),
    .RESET_B(net671),
    .D(_00703_),
    .Q_N(_09276_),
    .Q(\top1.memory1.mem1[83][2] ));
 sg13g2_dfrbp_1 _20503_ (.CLK(\clknet_leaf_75_top1.acquisition_clk ),
    .RESET_B(net670),
    .D(_00704_),
    .Q_N(_09275_),
    .Q(\top1.memory1.mem1[159][0] ));
 sg13g2_dfrbp_1 _20504_ (.CLK(\clknet_leaf_73_top1.acquisition_clk ),
    .RESET_B(net669),
    .D(_00705_),
    .Q_N(_09274_),
    .Q(\top1.memory1.mem1[159][1] ));
 sg13g2_dfrbp_1 _20505_ (.CLK(\clknet_leaf_59_top1.acquisition_clk ),
    .RESET_B(net668),
    .D(_00706_),
    .Q_N(_09273_),
    .Q(\top1.memory1.mem1[159][2] ));
 sg13g2_dfrbp_1 _20506_ (.CLK(\clknet_leaf_268_top1.acquisition_clk ),
    .RESET_B(net667),
    .D(_00707_),
    .Q_N(_09272_),
    .Q(\top1.memory1.mem1[84][0] ));
 sg13g2_dfrbp_1 _20507_ (.CLK(\clknet_leaf_30_top1.acquisition_clk ),
    .RESET_B(net666),
    .D(_00708_),
    .Q_N(_09271_),
    .Q(\top1.memory1.mem1[84][1] ));
 sg13g2_dfrbp_1 _20508_ (.CLK(\clknet_leaf_289_top1.acquisition_clk ),
    .RESET_B(net665),
    .D(_00709_),
    .Q_N(_09270_),
    .Q(\top1.memory1.mem1[84][2] ));
 sg13g2_dfrbp_1 _20509_ (.CLK(\clknet_leaf_269_top1.acquisition_clk ),
    .RESET_B(net664),
    .D(_00710_),
    .Q_N(_09269_),
    .Q(\top1.memory1.mem1[85][0] ));
 sg13g2_dfrbp_1 _20510_ (.CLK(\clknet_leaf_29_top1.acquisition_clk ),
    .RESET_B(net663),
    .D(_00711_),
    .Q_N(_09268_),
    .Q(\top1.memory1.mem1[85][1] ));
 sg13g2_dfrbp_1 _20511_ (.CLK(\clknet_leaf_290_top1.acquisition_clk ),
    .RESET_B(net662),
    .D(_00712_),
    .Q_N(_09267_),
    .Q(\top1.memory1.mem1[85][2] ));
 sg13g2_dfrbp_1 _20512_ (.CLK(\clknet_leaf_269_top1.acquisition_clk ),
    .RESET_B(net661),
    .D(_00713_),
    .Q_N(_09266_),
    .Q(\top1.memory1.mem1[86][0] ));
 sg13g2_dfrbp_1 _20513_ (.CLK(\clknet_leaf_268_top1.acquisition_clk ),
    .RESET_B(net660),
    .D(_00714_),
    .Q_N(_09265_),
    .Q(\top1.memory1.mem1[86][1] ));
 sg13g2_dfrbp_1 _20514_ (.CLK(\clknet_leaf_290_top1.acquisition_clk ),
    .RESET_B(net659),
    .D(_00715_),
    .Q_N(_09264_),
    .Q(\top1.memory1.mem1[86][2] ));
 sg13g2_dfrbp_1 _20515_ (.CLK(\clknet_leaf_268_top1.acquisition_clk ),
    .RESET_B(net658),
    .D(_00716_),
    .Q_N(_09263_),
    .Q(\top1.memory1.mem1[87][0] ));
 sg13g2_dfrbp_1 _20516_ (.CLK(\clknet_leaf_30_top1.acquisition_clk ),
    .RESET_B(net657),
    .D(_00717_),
    .Q_N(_09262_),
    .Q(\top1.memory1.mem1[87][1] ));
 sg13g2_dfrbp_1 _20517_ (.CLK(\clknet_leaf_289_top1.acquisition_clk ),
    .RESET_B(net656),
    .D(_00718_),
    .Q_N(_09261_),
    .Q(\top1.memory1.mem1[87][2] ));
 sg13g2_dfrbp_1 _20518_ (.CLK(\clknet_leaf_269_top1.acquisition_clk ),
    .RESET_B(net655),
    .D(_00719_),
    .Q_N(_09260_),
    .Q(\top1.memory1.mem1[88][0] ));
 sg13g2_dfrbp_1 _20519_ (.CLK(\clknet_leaf_284_top1.acquisition_clk ),
    .RESET_B(net654),
    .D(_00720_),
    .Q_N(_09259_),
    .Q(\top1.memory1.mem1[88][1] ));
 sg13g2_dfrbp_1 _20520_ (.CLK(\clknet_leaf_290_top1.acquisition_clk ),
    .RESET_B(net653),
    .D(_00721_),
    .Q_N(_09258_),
    .Q(\top1.memory1.mem1[88][2] ));
 sg13g2_dfrbp_1 _20521_ (.CLK(\clknet_leaf_265_top1.acquisition_clk ),
    .RESET_B(net652),
    .D(_00722_),
    .Q_N(_09257_),
    .Q(\top1.memory1.mem1[8][0] ));
 sg13g2_dfrbp_1 _20522_ (.CLK(\clknet_leaf_265_top1.acquisition_clk ),
    .RESET_B(net651),
    .D(_00723_),
    .Q_N(_09256_),
    .Q(\top1.memory1.mem1[8][1] ));
 sg13g2_dfrbp_1 _20523_ (.CLK(\clknet_leaf_271_top1.acquisition_clk ),
    .RESET_B(net650),
    .D(_00724_),
    .Q_N(_09255_),
    .Q(\top1.memory1.mem1[8][2] ));
 sg13g2_dfrbp_1 _20524_ (.CLK(\clknet_leaf_218_top1.acquisition_clk ),
    .RESET_B(net649),
    .D(_00725_),
    .Q_N(_09254_),
    .Q(\top1.memory1.mem1[119][0] ));
 sg13g2_dfrbp_1 _20525_ (.CLK(\clknet_leaf_217_top1.acquisition_clk ),
    .RESET_B(net648),
    .D(_00726_),
    .Q_N(_09253_),
    .Q(\top1.memory1.mem1[119][1] ));
 sg13g2_dfrbp_1 _20526_ (.CLK(\clknet_leaf_219_top1.acquisition_clk ),
    .RESET_B(net647),
    .D(_00727_),
    .Q_N(_09252_),
    .Q(\top1.memory1.mem1[119][2] ));
 sg13g2_dfrbp_1 _20527_ (.CLK(\clknet_leaf_18_top1.acquisition_clk ),
    .RESET_B(net646),
    .D(_00728_),
    .Q_N(_09251_),
    .Q(\top1.memory1.mem1[129][0] ));
 sg13g2_dfrbp_1 _20528_ (.CLK(\clknet_leaf_51_top1.acquisition_clk ),
    .RESET_B(net645),
    .D(_00729_),
    .Q_N(_09250_),
    .Q(\top1.memory1.mem1[129][1] ));
 sg13g2_dfrbp_1 _20529_ (.CLK(\clknet_leaf_19_top1.acquisition_clk ),
    .RESET_B(net644),
    .D(_00730_),
    .Q_N(_09249_),
    .Q(\top1.memory1.mem1[129][2] ));
 sg13g2_dfrbp_1 _20530_ (.CLK(\clknet_leaf_54_top1.acquisition_clk ),
    .RESET_B(net643),
    .D(_00731_),
    .Q_N(_09248_),
    .Q(\top1.memory1.mem1[139][0] ));
 sg13g2_dfrbp_1 _20531_ (.CLK(\clknet_leaf_56_top1.acquisition_clk ),
    .RESET_B(net642),
    .D(_00732_),
    .Q_N(_09247_),
    .Q(\top1.memory1.mem1[139][1] ));
 sg13g2_dfrbp_1 _20532_ (.CLK(\clknet_leaf_50_top1.acquisition_clk ),
    .RESET_B(net641),
    .D(_00733_),
    .Q_N(_09246_),
    .Q(\top1.memory1.mem1[139][2] ));
 sg13g2_dfrbp_1 _20533_ (.CLK(\clknet_leaf_13_top1.acquisition_clk ),
    .RESET_B(net640),
    .D(_00734_),
    .Q_N(_09245_),
    .Q(\top1.memory1.mem1[76][0] ));
 sg13g2_dfrbp_1 _20534_ (.CLK(\clknet_leaf_13_top1.acquisition_clk ),
    .RESET_B(net639),
    .D(_00735_),
    .Q_N(_09244_),
    .Q(\top1.memory1.mem1[76][1] ));
 sg13g2_dfrbp_1 _20535_ (.CLK(\clknet_leaf_15_top1.acquisition_clk ),
    .RESET_B(net638),
    .D(_00736_),
    .Q_N(_09243_),
    .Q(\top1.memory1.mem1[76][2] ));
 sg13g2_dfrbp_1 _20536_ (.CLK(\clknet_leaf_4_top1.acquisition_clk ),
    .RESET_B(net637),
    .D(_00737_),
    .Q_N(_09242_),
    .Q(\top1.memory1.mem1[77][0] ));
 sg13g2_dfrbp_1 _20537_ (.CLK(\clknet_leaf_13_top1.acquisition_clk ),
    .RESET_B(net636),
    .D(_00738_),
    .Q_N(_09241_),
    .Q(\top1.memory1.mem1[77][1] ));
 sg13g2_dfrbp_1 _20538_ (.CLK(\clknet_leaf_15_top1.acquisition_clk ),
    .RESET_B(net635),
    .D(_00739_),
    .Q_N(_09240_),
    .Q(\top1.memory1.mem1[77][2] ));
 sg13g2_dfrbp_1 _20539_ (.CLK(\clknet_leaf_13_top1.acquisition_clk ),
    .RESET_B(net634),
    .D(_00740_),
    .Q_N(_09239_),
    .Q(\top1.memory1.mem1[78][0] ));
 sg13g2_dfrbp_1 _20540_ (.CLK(\clknet_leaf_13_top1.acquisition_clk ),
    .RESET_B(net633),
    .D(_00741_),
    .Q_N(_09238_),
    .Q(\top1.memory1.mem1[78][1] ));
 sg13g2_dfrbp_1 _20541_ (.CLK(\clknet_leaf_14_top1.acquisition_clk ),
    .RESET_B(net632),
    .D(_00742_),
    .Q_N(_09237_),
    .Q(\top1.memory1.mem1[78][2] ));
 sg13g2_dfrbp_1 _20542_ (.CLK(\clknet_leaf_261_top1.acquisition_clk ),
    .RESET_B(net631),
    .D(_00743_),
    .Q_N(_09236_),
    .Q(\top1.memory1.mem1[7][0] ));
 sg13g2_dfrbp_1 _20543_ (.CLK(\clknet_leaf_263_top1.acquisition_clk ),
    .RESET_B(net630),
    .D(_00744_),
    .Q_N(_09235_),
    .Q(\top1.memory1.mem1[7][1] ));
 sg13g2_dfrbp_1 _20544_ (.CLK(\clknet_leaf_266_top1.acquisition_clk ),
    .RESET_B(net629),
    .D(_00745_),
    .Q_N(_09234_),
    .Q(\top1.memory1.mem1[7][2] ));
 sg13g2_dfrbp_1 _20545_ (.CLK(\clknet_leaf_285_top1.acquisition_clk ),
    .RESET_B(net628),
    .D(_00746_),
    .Q_N(_09233_),
    .Q(\top1.memory1.mem1[80][0] ));
 sg13g2_dfrbp_1 _20546_ (.CLK(\clknet_leaf_286_top1.acquisition_clk ),
    .RESET_B(net627),
    .D(_00747_),
    .Q_N(_09232_),
    .Q(\top1.memory1.mem1[80][1] ));
 sg13g2_dfrbp_1 _20547_ (.CLK(\clknet_leaf_287_top1.acquisition_clk ),
    .RESET_B(net626),
    .D(_00748_),
    .Q_N(_09231_),
    .Q(\top1.memory1.mem1[80][2] ));
 sg13g2_dfrbp_1 _20548_ (.CLK(\clknet_leaf_286_top1.acquisition_clk ),
    .RESET_B(net625),
    .D(_00749_),
    .Q_N(_09230_),
    .Q(\top1.memory1.mem1[81][0] ));
 sg13g2_dfrbp_1 _20549_ (.CLK(\clknet_leaf_286_top1.acquisition_clk ),
    .RESET_B(net624),
    .D(_00750_),
    .Q_N(_09229_),
    .Q(\top1.memory1.mem1[81][1] ));
 sg13g2_dfrbp_1 _20550_ (.CLK(\clknet_leaf_287_top1.acquisition_clk ),
    .RESET_B(net623),
    .D(_00751_),
    .Q_N(_09228_),
    .Q(\top1.memory1.mem1[81][2] ));
 sg13g2_dfrbp_1 _20551_ (.CLK(\clknet_leaf_257_top1.acquisition_clk ),
    .RESET_B(net622),
    .D(_00752_),
    .Q_N(_09227_),
    .Q(\top1.memory1.mem1[29][0] ));
 sg13g2_dfrbp_1 _20552_ (.CLK(\clknet_leaf_256_top1.acquisition_clk ),
    .RESET_B(net621),
    .D(_00753_),
    .Q_N(_09226_),
    .Q(\top1.memory1.mem1[29][1] ));
 sg13g2_dfrbp_1 _20553_ (.CLK(\clknet_leaf_259_top1.acquisition_clk ),
    .RESET_B(net620),
    .D(_00754_),
    .Q_N(_09225_),
    .Q(\top1.memory1.mem1[29][2] ));
 sg13g2_dfrbp_1 _20554_ (.CLK(net7718),
    .RESET_B(net7725),
    .D(_00755_),
    .Q_N(_09224_),
    .Q(\top1.event_time[27] ));
 sg13g2_dfrbp_1 _20555_ (.CLK(net7718),
    .RESET_B(net7723),
    .D(_00756_),
    .Q_N(_09223_),
    .Q(\top1.event_time[28] ));
 sg13g2_dfrbp_1 _20556_ (.CLK(net7718),
    .RESET_B(net7723),
    .D(_00757_),
    .Q_N(_09222_),
    .Q(\top1.event_time[29] ));
 sg13g2_dfrbp_1 _20557_ (.CLK(net7718),
    .RESET_B(net7723),
    .D(_00758_),
    .Q_N(_09221_),
    .Q(\top1.event_time[30] ));
 sg13g2_dfrbp_1 _20558_ (.CLK(net7718),
    .RESET_B(net7723),
    .D(_00759_),
    .Q_N(_09220_),
    .Q(\top1.event_time[31] ));
 sg13g2_dfrbp_1 _20559_ (.CLK(\clknet_leaf_147_top1.acquisition_clk ),
    .RESET_B(net619),
    .D(_00760_),
    .Q_N(_09219_),
    .Q(\top1.memory1.mem1[39][0] ));
 sg13g2_dfrbp_1 _20560_ (.CLK(\clknet_leaf_147_top1.acquisition_clk ),
    .RESET_B(net618),
    .D(_00761_),
    .Q_N(_09218_),
    .Q(\top1.memory1.mem1[39][1] ));
 sg13g2_dfrbp_1 _20561_ (.CLK(\clknet_leaf_151_top1.acquisition_clk ),
    .RESET_B(net617),
    .D(_00762_),
    .Q_N(_09217_),
    .Q(\top1.memory1.mem1[39][2] ));
 sg13g2_dfrbp_1 _20562_ (.CLK(\clknet_leaf_148_top1.acquisition_clk ),
    .RESET_B(net616),
    .D(_00763_),
    .Q_N(_09216_),
    .Q(\top1.memory1.mem1[38][0] ));
 sg13g2_dfrbp_1 _20563_ (.CLK(\clknet_leaf_148_top1.acquisition_clk ),
    .RESET_B(net615),
    .D(_00764_),
    .Q_N(_09215_),
    .Q(\top1.memory1.mem1[38][1] ));
 sg13g2_dfrbp_1 _20564_ (.CLK(\clknet_leaf_151_top1.acquisition_clk ),
    .RESET_B(net614),
    .D(_00765_),
    .Q_N(_09214_),
    .Q(\top1.memory1.mem1[38][2] ));
 sg13g2_dfrbp_1 _20565_ (.CLK(\clknet_leaf_277_top1.acquisition_clk ),
    .RESET_B(net613),
    .D(_00766_),
    .Q_N(_09213_),
    .Q(\top1.memory1.mem1[3][0] ));
 sg13g2_dfrbp_1 _20566_ (.CLK(\clknet_leaf_280_top1.acquisition_clk ),
    .RESET_B(net612),
    .D(_00767_),
    .Q_N(_09212_),
    .Q(\top1.memory1.mem1[3][1] ));
 sg13g2_dfrbp_1 _20567_ (.CLK(\clknet_leaf_281_top1.acquisition_clk ),
    .RESET_B(net611),
    .D(_00768_),
    .Q_N(_09211_),
    .Q(\top1.memory1.mem1[3][2] ));
 sg13g2_dfrbp_1 _20568_ (.CLK(\clknet_leaf_149_top1.acquisition_clk ),
    .RESET_B(net610),
    .D(_00769_),
    .Q_N(_09210_),
    .Q(\top1.memory1.mem1[40][0] ));
 sg13g2_dfrbp_1 _20569_ (.CLK(\clknet_leaf_158_top1.acquisition_clk ),
    .RESET_B(net609),
    .D(_00770_),
    .Q_N(_09209_),
    .Q(\top1.memory1.mem1[40][1] ));
 sg13g2_dfrbp_1 _20570_ (.CLK(\clknet_leaf_159_top1.acquisition_clk ),
    .RESET_B(net608),
    .D(_00771_),
    .Q_N(_09208_),
    .Q(\top1.memory1.mem1[40][2] ));
 sg13g2_dfrbp_1 _20571_ (.CLK(\clknet_leaf_145_top1.acquisition_clk ),
    .RESET_B(net607),
    .D(_00772_),
    .Q_N(_09207_),
    .Q(\top1.memory1.mem1[41][0] ));
 sg13g2_dfrbp_1 _20572_ (.CLK(\clknet_leaf_158_top1.acquisition_clk ),
    .RESET_B(net606),
    .D(_00773_),
    .Q_N(_09206_),
    .Q(\top1.memory1.mem1[41][1] ));
 sg13g2_dfrbp_1 _20573_ (.CLK(\clknet_leaf_152_top1.acquisition_clk ),
    .RESET_B(net605),
    .D(_00774_),
    .Q_N(_09205_),
    .Q(\top1.memory1.mem1[41][2] ));
 sg13g2_dfrbp_1 _20574_ (.CLK(\clknet_leaf_149_top1.acquisition_clk ),
    .RESET_B(net604),
    .D(_00775_),
    .Q_N(_09204_),
    .Q(\top1.memory1.mem1[42][0] ));
 sg13g2_dfrbp_1 _20575_ (.CLK(\clknet_leaf_158_top1.acquisition_clk ),
    .RESET_B(net603),
    .D(_00776_),
    .Q_N(_09203_),
    .Q(\top1.memory1.mem1[42][1] ));
 sg13g2_dfrbp_1 _20576_ (.CLK(\clknet_leaf_152_top1.acquisition_clk ),
    .RESET_B(net602),
    .D(_00777_),
    .Q_N(_09202_),
    .Q(\top1.memory1.mem1[42][2] ));
 sg13g2_dfrbp_1 _20577_ (.CLK(\clknet_leaf_149_top1.acquisition_clk ),
    .RESET_B(net601),
    .D(_00778_),
    .Q_N(_09201_),
    .Q(\top1.memory1.mem1[43][0] ));
 sg13g2_dfrbp_1 _20578_ (.CLK(\clknet_leaf_158_top1.acquisition_clk ),
    .RESET_B(net600),
    .D(_00779_),
    .Q_N(_09200_),
    .Q(\top1.memory1.mem1[43][1] ));
 sg13g2_dfrbp_1 _20579_ (.CLK(\clknet_leaf_152_top1.acquisition_clk ),
    .RESET_B(net599),
    .D(_00780_),
    .Q_N(_09199_),
    .Q(\top1.memory1.mem1[43][2] ));
 sg13g2_dfrbp_1 _20580_ (.CLK(\clknet_leaf_161_top1.acquisition_clk ),
    .RESET_B(net598),
    .D(_00781_),
    .Q_N(_09198_),
    .Q(\top1.memory1.mem1[44][0] ));
 sg13g2_dfrbp_1 _20581_ (.CLK(\clknet_leaf_162_top1.acquisition_clk ),
    .RESET_B(net597),
    .D(_00782_),
    .Q_N(_09197_),
    .Q(\top1.memory1.mem1[44][1] ));
 sg13g2_dfrbp_1 _20582_ (.CLK(\clknet_leaf_162_top1.acquisition_clk ),
    .RESET_B(net596),
    .D(_00783_),
    .Q_N(_09196_),
    .Q(\top1.memory1.mem1[44][2] ));
 sg13g2_dfrbp_1 _20583_ (.CLK(\clknet_leaf_160_top1.acquisition_clk ),
    .RESET_B(net595),
    .D(_00784_),
    .Q_N(_09195_),
    .Q(\top1.memory1.mem1[45][0] ));
 sg13g2_dfrbp_1 _20584_ (.CLK(\clknet_leaf_162_top1.acquisition_clk ),
    .RESET_B(net594),
    .D(_00785_),
    .Q_N(_09194_),
    .Q(\top1.memory1.mem1[45][1] ));
 sg13g2_dfrbp_1 _20585_ (.CLK(\clknet_leaf_161_top1.acquisition_clk ),
    .RESET_B(net593),
    .D(_00786_),
    .Q_N(_09193_),
    .Q(\top1.memory1.mem1[45][2] ));
 sg13g2_dfrbp_1 _20586_ (.CLK(\clknet_leaf_161_top1.acquisition_clk ),
    .RESET_B(net592),
    .D(_00787_),
    .Q_N(_09192_),
    .Q(\top1.memory1.mem1[46][0] ));
 sg13g2_dfrbp_1 _20587_ (.CLK(\clknet_leaf_162_top1.acquisition_clk ),
    .RESET_B(net591),
    .D(_00788_),
    .Q_N(_09191_),
    .Q(\top1.memory1.mem1[46][1] ));
 sg13g2_dfrbp_1 _20588_ (.CLK(\clknet_leaf_159_top1.acquisition_clk ),
    .RESET_B(net590),
    .D(_00789_),
    .Q_N(_09190_),
    .Q(\top1.memory1.mem1[46][2] ));
 sg13g2_dfrbp_1 _20589_ (.CLK(\clknet_leaf_160_top1.acquisition_clk ),
    .RESET_B(net589),
    .D(_00790_),
    .Q_N(_09189_),
    .Q(\top1.memory1.mem1[47][0] ));
 sg13g2_dfrbp_1 _20590_ (.CLK(\clknet_leaf_162_top1.acquisition_clk ),
    .RESET_B(net588),
    .D(_00791_),
    .Q_N(_09188_),
    .Q(\top1.memory1.mem1[47][1] ));
 sg13g2_dfrbp_1 _20591_ (.CLK(\clknet_leaf_161_top1.acquisition_clk ),
    .RESET_B(net587),
    .D(_00792_),
    .Q_N(_09187_),
    .Q(\top1.memory1.mem1[47][2] ));
 sg13g2_dfrbp_1 _20592_ (.CLK(\clknet_leaf_165_top1.acquisition_clk ),
    .RESET_B(net586),
    .D(_00793_),
    .Q_N(_09186_),
    .Q(\top1.memory1.mem1[48][0] ));
 sg13g2_dfrbp_1 _20593_ (.CLK(\clknet_leaf_166_top1.acquisition_clk ),
    .RESET_B(net585),
    .D(_00794_),
    .Q_N(_09185_),
    .Q(\top1.memory1.mem1[48][1] ));
 sg13g2_dfrbp_1 _20594_ (.CLK(\clknet_leaf_163_top1.acquisition_clk ),
    .RESET_B(net584),
    .D(_00795_),
    .Q_N(_09184_),
    .Q(\top1.memory1.mem1[48][2] ));
 sg13g2_dfrbp_1 _20595_ (.CLK(\clknet_leaf_261_top1.acquisition_clk ),
    .RESET_B(net583),
    .D(_00796_),
    .Q_N(_09183_),
    .Q(\top1.memory1.mem1[4][0] ));
 sg13g2_dfrbp_1 _20596_ (.CLK(\clknet_leaf_263_top1.acquisition_clk ),
    .RESET_B(net582),
    .D(_00797_),
    .Q_N(_09182_),
    .Q(\top1.memory1.mem1[4][1] ));
 sg13g2_dfrbp_1 _20597_ (.CLK(\clknet_leaf_266_top1.acquisition_clk ),
    .RESET_B(net581),
    .D(_00798_),
    .Q_N(_09181_),
    .Q(\top1.memory1.mem1[4][2] ));
 sg13g2_dfrbp_1 _20598_ (.CLK(\clknet_leaf_166_top1.acquisition_clk ),
    .RESET_B(net580),
    .D(_00799_),
    .Q_N(_09180_),
    .Q(\top1.memory1.mem1[50][0] ));
 sg13g2_dfrbp_1 _20599_ (.CLK(\clknet_leaf_166_top1.acquisition_clk ),
    .RESET_B(net579),
    .D(_00800_),
    .Q_N(_09179_),
    .Q(\top1.memory1.mem1[50][1] ));
 sg13g2_dfrbp_1 _20600_ (.CLK(\clknet_leaf_164_top1.acquisition_clk ),
    .RESET_B(net578),
    .D(_00801_),
    .Q_N(_09178_),
    .Q(\top1.memory1.mem1[50][2] ));
 sg13g2_dfrbp_1 _20601_ (.CLK(\clknet_leaf_165_top1.acquisition_clk ),
    .RESET_B(net577),
    .D(_00802_),
    .Q_N(_09177_),
    .Q(\top1.memory1.mem1[51][0] ));
 sg13g2_dfrbp_1 _20602_ (.CLK(\clknet_leaf_165_top1.acquisition_clk ),
    .RESET_B(net576),
    .D(_00803_),
    .Q_N(_09176_),
    .Q(\top1.memory1.mem1[51][1] ));
 sg13g2_dfrbp_1 _20603_ (.CLK(\clknet_leaf_163_top1.acquisition_clk ),
    .RESET_B(net575),
    .D(_00804_),
    .Q_N(_09175_),
    .Q(\top1.memory1.mem1[51][2] ));
 sg13g2_dfrbp_1 _20604_ (.CLK(\clknet_leaf_166_top1.acquisition_clk ),
    .RESET_B(net574),
    .D(_00805_),
    .Q_N(_09174_),
    .Q(\top1.memory1.mem1[52][0] ));
 sg13g2_dfrbp_1 _20605_ (.CLK(\clknet_leaf_201_top1.acquisition_clk ),
    .RESET_B(net573),
    .D(_00806_),
    .Q_N(_09173_),
    .Q(\top1.memory1.mem1[52][1] ));
 sg13g2_dfrbp_1 _20606_ (.CLK(\clknet_leaf_199_top1.acquisition_clk ),
    .RESET_B(net572),
    .D(_00807_),
    .Q_N(_09172_),
    .Q(\top1.memory1.mem1[52][2] ));
 sg13g2_dfrbp_1 _20607_ (.CLK(\clknet_leaf_201_top1.acquisition_clk ),
    .RESET_B(net571),
    .D(_00808_),
    .Q_N(_09171_),
    .Q(\top1.memory1.mem1[53][0] ));
 sg13g2_dfrbp_1 _20608_ (.CLK(\clknet_leaf_201_top1.acquisition_clk ),
    .RESET_B(net570),
    .D(_00809_),
    .Q_N(_09170_),
    .Q(\top1.memory1.mem1[53][1] ));
 sg13g2_dfrbp_1 _20609_ (.CLK(\clknet_leaf_201_top1.acquisition_clk ),
    .RESET_B(net569),
    .D(_00810_),
    .Q_N(_09169_),
    .Q(\top1.memory1.mem1[53][2] ));
 sg13g2_dfrbp_1 _20610_ (.CLK(\clknet_leaf_166_top1.acquisition_clk ),
    .RESET_B(net568),
    .D(_00811_),
    .Q_N(_09168_),
    .Q(\top1.memory1.mem1[54][0] ));
 sg13g2_dfrbp_1 _20611_ (.CLK(\clknet_leaf_201_top1.acquisition_clk ),
    .RESET_B(net567),
    .D(_00812_),
    .Q_N(_09167_),
    .Q(\top1.memory1.mem1[54][1] ));
 sg13g2_dfrbp_1 _20612_ (.CLK(\clknet_leaf_201_top1.acquisition_clk ),
    .RESET_B(net566),
    .D(_00813_),
    .Q_N(_09166_),
    .Q(\top1.memory1.mem1[54][2] ));
 sg13g2_dfrbp_1 _20613_ (.CLK(\clknet_leaf_166_top1.acquisition_clk ),
    .RESET_B(net565),
    .D(_00814_),
    .Q_N(_09165_),
    .Q(\top1.memory1.mem1[55][0] ));
 sg13g2_dfrbp_1 _20614_ (.CLK(\clknet_leaf_201_top1.acquisition_clk ),
    .RESET_B(net564),
    .D(_00815_),
    .Q_N(_09164_),
    .Q(\top1.memory1.mem1[55][1] ));
 sg13g2_dfrbp_1 _20615_ (.CLK(\clknet_leaf_201_top1.acquisition_clk ),
    .RESET_B(net563),
    .D(_00816_),
    .Q_N(_09163_),
    .Q(\top1.memory1.mem1[55][2] ));
 sg13g2_dfrbp_1 _20616_ (.CLK(\clknet_leaf_167_top1.acquisition_clk ),
    .RESET_B(net562),
    .D(_00817_),
    .Q_N(_09162_),
    .Q(\top1.memory1.mem1[56][0] ));
 sg13g2_dfrbp_1 _20617_ (.CLK(\clknet_leaf_162_top1.acquisition_clk ),
    .RESET_B(net561),
    .D(_00818_),
    .Q_N(_09161_),
    .Q(\top1.memory1.mem1[56][1] ));
 sg13g2_dfrbp_1 _20618_ (.CLK(\clknet_leaf_172_top1.acquisition_clk ),
    .RESET_B(net560),
    .D(_00819_),
    .Q_N(_09160_),
    .Q(\top1.memory1.mem1[56][2] ));
 sg13g2_dfrbp_1 _20619_ (.CLK(\clknet_leaf_167_top1.acquisition_clk ),
    .RESET_B(net559),
    .D(_00820_),
    .Q_N(_09159_),
    .Q(\top1.memory1.mem1[57][0] ));
 sg13g2_dfrbp_1 _20620_ (.CLK(\clknet_leaf_163_top1.acquisition_clk ),
    .RESET_B(net558),
    .D(_00821_),
    .Q_N(_09158_),
    .Q(\top1.memory1.mem1[57][1] ));
 sg13g2_dfrbp_1 _20621_ (.CLK(\clknet_leaf_173_top1.acquisition_clk ),
    .RESET_B(net557),
    .D(_00822_),
    .Q_N(_09157_),
    .Q(\top1.memory1.mem1[57][2] ));
 sg13g2_dfrbp_1 _20622_ (.CLK(\clknet_leaf_167_top1.acquisition_clk ),
    .RESET_B(net556),
    .D(_00823_),
    .Q_N(_09156_),
    .Q(\top1.memory1.mem1[58][0] ));
 sg13g2_dfrbp_1 _20623_ (.CLK(\clknet_leaf_163_top1.acquisition_clk ),
    .RESET_B(net555),
    .D(_00824_),
    .Q_N(_09155_),
    .Q(\top1.memory1.mem1[58][1] ));
 sg13g2_dfrbp_1 _20624_ (.CLK(\clknet_leaf_168_top1.acquisition_clk ),
    .RESET_B(net554),
    .D(_00825_),
    .Q_N(_09154_),
    .Q(\top1.memory1.mem1[58][2] ));
 sg13g2_dfrbp_1 _20625_ (.CLK(\clknet_leaf_262_top1.acquisition_clk ),
    .RESET_B(net553),
    .D(_00826_),
    .Q_N(_09153_),
    .Q(\top1.memory1.mem1[5][0] ));
 sg13g2_dfrbp_1 _20626_ (.CLK(\clknet_leaf_263_top1.acquisition_clk ),
    .RESET_B(net552),
    .D(_00827_),
    .Q_N(_09152_),
    .Q(\top1.memory1.mem1[5][1] ));
 sg13g2_dfrbp_1 _20627_ (.CLK(\clknet_leaf_266_top1.acquisition_clk ),
    .RESET_B(net551),
    .D(_00828_),
    .Q_N(_09151_),
    .Q(\top1.memory1.mem1[5][2] ));
 sg13g2_dfrbp_1 _20628_ (.CLK(\clknet_leaf_204_top1.acquisition_clk ),
    .RESET_B(net550),
    .D(_00829_),
    .Q_N(_09150_),
    .Q(\top1.memory1.mem1[60][0] ));
 sg13g2_dfrbp_1 _20629_ (.CLK(\clknet_leaf_205_top1.acquisition_clk ),
    .RESET_B(net549),
    .D(_00830_),
    .Q_N(_09149_),
    .Q(\top1.memory1.mem1[60][1] ));
 sg13g2_dfrbp_1 _20630_ (.CLK(\clknet_leaf_200_top1.acquisition_clk ),
    .RESET_B(net548),
    .D(_00831_),
    .Q_N(_09148_),
    .Q(\top1.memory1.mem1[60][2] ));
 sg13g2_dfrbp_1 _20631_ (.CLK(\clknet_leaf_204_top1.acquisition_clk ),
    .RESET_B(net547),
    .D(_00832_),
    .Q_N(_09147_),
    .Q(\top1.memory1.mem1[61][0] ));
 sg13g2_dfrbp_1 _20632_ (.CLK(\clknet_leaf_205_top1.acquisition_clk ),
    .RESET_B(net546),
    .D(_00833_),
    .Q_N(_09146_),
    .Q(\top1.memory1.mem1[61][1] ));
 sg13g2_dfrbp_1 _20633_ (.CLK(\clknet_leaf_202_top1.acquisition_clk ),
    .RESET_B(net545),
    .D(_00834_),
    .Q_N(_09145_),
    .Q(\top1.memory1.mem1[61][2] ));
 sg13g2_dfrbp_1 _20634_ (.CLK(\clknet_leaf_204_top1.acquisition_clk ),
    .RESET_B(net544),
    .D(_00835_),
    .Q_N(_09144_),
    .Q(\top1.memory1.mem1[62][0] ));
 sg13g2_dfrbp_1 _20635_ (.CLK(\clknet_leaf_203_top1.acquisition_clk ),
    .RESET_B(net543),
    .D(_00836_),
    .Q_N(_09143_),
    .Q(\top1.memory1.mem1[62][1] ));
 sg13g2_dfrbp_1 _20636_ (.CLK(\clknet_leaf_202_top1.acquisition_clk ),
    .RESET_B(net542),
    .D(_00837_),
    .Q_N(_09142_),
    .Q(\top1.memory1.mem1[62][2] ));
 sg13g2_dfrbp_1 _20637_ (.CLK(\clknet_leaf_165_top1.acquisition_clk ),
    .RESET_B(net541),
    .D(_00838_),
    .Q_N(_09141_),
    .Q(\top1.memory1.mem1[49][0] ));
 sg13g2_dfrbp_1 _20638_ (.CLK(\clknet_leaf_163_top1.acquisition_clk ),
    .RESET_B(net540),
    .D(_00839_),
    .Q_N(_09140_),
    .Q(\top1.memory1.mem1[49][1] ));
 sg13g2_dfrbp_1 _20639_ (.CLK(\clknet_leaf_163_top1.acquisition_clk ),
    .RESET_B(net539),
    .D(_00840_),
    .Q_N(_09139_),
    .Q(\top1.memory1.mem1[49][2] ));
 sg13g2_dfrbp_1 _20640_ (.CLK(\clknet_leaf_32_top1.acquisition_clk ),
    .RESET_B(net538),
    .D(_00841_),
    .Q_N(_09138_),
    .Q(\top1.memory1.mem1[198][0] ));
 sg13g2_dfrbp_1 _20641_ (.CLK(\clknet_leaf_31_top1.acquisition_clk ),
    .RESET_B(net537),
    .D(_00842_),
    .Q_N(_09137_),
    .Q(\top1.memory1.mem1[198][1] ));
 sg13g2_dfrbp_1 _20642_ (.CLK(\clknet_leaf_32_top1.acquisition_clk ),
    .RESET_B(net536),
    .D(_00843_),
    .Q_N(_09136_),
    .Q(\top1.memory1.mem1[198][2] ));
 sg13g2_dfrbp_1 _20643_ (.CLK(\clknet_leaf_33_top1.acquisition_clk ),
    .RESET_B(net535),
    .D(_00844_),
    .Q_N(_09135_),
    .Q(\top1.memory1.mem1[197][0] ));
 sg13g2_dfrbp_1 _20644_ (.CLK(\clknet_leaf_34_top1.acquisition_clk ),
    .RESET_B(net534),
    .D(_00845_),
    .Q_N(_09134_),
    .Q(\top1.memory1.mem1[197][1] ));
 sg13g2_dfrbp_1 _20645_ (.CLK(\clknet_leaf_33_top1.acquisition_clk ),
    .RESET_B(net533),
    .D(_00846_),
    .Q_N(_09133_),
    .Q(\top1.memory1.mem1[197][2] ));
 sg13g2_dfrbp_1 _20646_ (.CLK(\clknet_leaf_205_top1.acquisition_clk ),
    .RESET_B(net532),
    .D(_00847_),
    .Q_N(_09132_),
    .Q(\top1.memory1.mem1[63][0] ));
 sg13g2_dfrbp_1 _20647_ (.CLK(\clknet_leaf_203_top1.acquisition_clk ),
    .RESET_B(net531),
    .D(_00848_),
    .Q_N(_09131_),
    .Q(\top1.memory1.mem1[63][1] ));
 sg13g2_dfrbp_1 _20648_ (.CLK(\clknet_leaf_202_top1.acquisition_clk ),
    .RESET_B(net530),
    .D(_00849_),
    .Q_N(_09130_),
    .Q(\top1.memory1.mem1[63][2] ));
 sg13g2_dfrbp_1 _20649_ (.CLK(\clknet_leaf_6_top1.acquisition_clk ),
    .RESET_B(net529),
    .D(_00850_),
    .Q_N(_09129_),
    .Q(\top1.memory1.mem1[64][0] ));
 sg13g2_dfrbp_1 _20650_ (.CLK(\clknet_leaf_1_top1.acquisition_clk ),
    .RESET_B(net528),
    .D(_00851_),
    .Q_N(_09128_),
    .Q(\top1.memory1.mem1[64][1] ));
 sg13g2_dfrbp_1 _20651_ (.CLK(\clknet_leaf_1_top1.acquisition_clk ),
    .RESET_B(net527),
    .D(_00852_),
    .Q_N(_09127_),
    .Q(\top1.memory1.mem1[64][2] ));
 sg13g2_dfrbp_1 _20652_ (.CLK(\clknet_leaf_5_top1.acquisition_clk ),
    .RESET_B(net526),
    .D(_00853_),
    .Q_N(_09126_),
    .Q(\top1.memory1.mem1[65][0] ));
 sg13g2_dfrbp_1 _20653_ (.CLK(\clknet_leaf_1_top1.acquisition_clk ),
    .RESET_B(net525),
    .D(_00854_),
    .Q_N(_09125_),
    .Q(\top1.memory1.mem1[65][1] ));
 sg13g2_dfrbp_1 _20654_ (.CLK(\clknet_leaf_5_top1.acquisition_clk ),
    .RESET_B(net524),
    .D(_00855_),
    .Q_N(_09124_),
    .Q(\top1.memory1.mem1[65][2] ));
 sg13g2_dfrbp_1 _20655_ (.CLK(\clknet_leaf_33_top1.acquisition_clk ),
    .RESET_B(net523),
    .D(_00856_),
    .Q_N(_09123_),
    .Q(\top1.memory1.mem1[196][0] ));
 sg13g2_dfrbp_1 _20656_ (.CLK(\clknet_leaf_30_top1.acquisition_clk ),
    .RESET_B(net522),
    .D(_00857_),
    .Q_N(_09122_),
    .Q(\top1.memory1.mem1[196][1] ));
 sg13g2_dfrbp_1 _20657_ (.CLK(\clknet_leaf_32_top1.acquisition_clk ),
    .RESET_B(net521),
    .D(_00858_),
    .Q_N(_09121_),
    .Q(\top1.memory1.mem1[196][2] ));
 sg13g2_dfrbp_1 _20658_ (.CLK(\clknet_leaf_167_top1.acquisition_clk ),
    .RESET_B(net520),
    .D(_00859_),
    .Q_N(_09120_),
    .Q(\top1.memory1.mem1[59][0] ));
 sg13g2_dfrbp_1 _20659_ (.CLK(\clknet_leaf_163_top1.acquisition_clk ),
    .RESET_B(net519),
    .D(_00860_),
    .Q_N(_09119_),
    .Q(\top1.memory1.mem1[59][1] ));
 sg13g2_dfrbp_1 _20660_ (.CLK(\clknet_leaf_172_top1.acquisition_clk ),
    .RESET_B(net518),
    .D(_00861_),
    .Q_N(_09118_),
    .Q(\top1.memory1.mem1[59][2] ));
 sg13g2_dfrbp_1 _20661_ (.CLK(\clknet_leaf_5_top1.acquisition_clk ),
    .RESET_B(net517),
    .D(_00862_),
    .Q_N(_09117_),
    .Q(\top1.memory1.mem1[66][0] ));
 sg13g2_dfrbp_1 _20662_ (.CLK(\clknet_leaf_6_top1.acquisition_clk ),
    .RESET_B(net516),
    .D(_00863_),
    .Q_N(_09116_),
    .Q(\top1.memory1.mem1[66][1] ));
 sg13g2_dfrbp_1 _20663_ (.CLK(\clknet_leaf_5_top1.acquisition_clk ),
    .RESET_B(net515),
    .D(_00864_),
    .Q_N(_09115_),
    .Q(\top1.memory1.mem1[66][2] ));
 sg13g2_dfrbp_1 _20664_ (.CLK(\clknet_leaf_35_top1.acquisition_clk ),
    .RESET_B(net514),
    .D(_00865_),
    .Q_N(_09114_),
    .Q(\top1.memory1.mem1[195][0] ));
 sg13g2_dfrbp_1 _20665_ (.CLK(\clknet_leaf_35_top1.acquisition_clk ),
    .RESET_B(net513),
    .D(_00866_),
    .Q_N(_09113_),
    .Q(\top1.memory1.mem1[195][1] ));
 sg13g2_dfrbp_1 _20666_ (.CLK(\clknet_leaf_35_top1.acquisition_clk ),
    .RESET_B(net512),
    .D(_00867_),
    .Q_N(_09112_),
    .Q(\top1.memory1.mem1[195][2] ));
 sg13g2_dfrbp_1 _20667_ (.CLK(\clknet_leaf_6_top1.acquisition_clk ),
    .RESET_B(net511),
    .D(_00868_),
    .Q_N(_09111_),
    .Q(\top1.memory1.mem1[67][0] ));
 sg13g2_dfrbp_1 _20668_ (.CLK(\clknet_leaf_1_top1.acquisition_clk ),
    .RESET_B(net510),
    .D(_00869_),
    .Q_N(_09110_),
    .Q(\top1.memory1.mem1[67][1] ));
 sg13g2_dfrbp_1 _20669_ (.CLK(\clknet_leaf_1_top1.acquisition_clk ),
    .RESET_B(net509),
    .D(_00870_),
    .Q_N(_09109_),
    .Q(\top1.memory1.mem1[67][2] ));
 sg13g2_dfrbp_1 _20670_ (.CLK(\clknet_leaf_26_top1.acquisition_clk ),
    .RESET_B(net508),
    .D(_00871_),
    .Q_N(_09108_),
    .Q(\top1.memory1.mem1[68][0] ));
 sg13g2_dfrbp_1 _20671_ (.CLK(\clknet_leaf_11_top1.acquisition_clk ),
    .RESET_B(net507),
    .D(_00872_),
    .Q_N(_09107_),
    .Q(\top1.memory1.mem1[68][1] ));
 sg13g2_dfrbp_1 _20672_ (.CLK(\clknet_leaf_21_top1.acquisition_clk ),
    .RESET_B(net506),
    .D(_00873_),
    .Q_N(_09106_),
    .Q(\top1.memory1.mem1[68][2] ));
 sg13g2_dfrbp_1 _20673_ (.CLK(\clknet_leaf_267_top1.acquisition_clk ),
    .RESET_B(net505),
    .D(_00874_),
    .Q_N(_09105_),
    .Q(\top1.memory1.mem1[194][0] ));
 sg13g2_dfrbp_1 _20674_ (.CLK(\clknet_leaf_31_top1.acquisition_clk ),
    .RESET_B(net504),
    .D(_00875_),
    .Q_N(_09104_),
    .Q(\top1.memory1.mem1[194][1] ));
 sg13g2_dfrbp_1 _20675_ (.CLK(\clknet_leaf_31_top1.acquisition_clk ),
    .RESET_B(net503),
    .D(_00876_),
    .Q_N(_09103_),
    .Q(\top1.memory1.mem1[194][2] ));
 sg13g2_dfrbp_1 _20676_ (.CLK(\clknet_leaf_21_top1.acquisition_clk ),
    .RESET_B(net502),
    .D(_00877_),
    .Q_N(_09102_),
    .Q(\top1.memory1.mem1[69][0] ));
 sg13g2_dfrbp_1 _20677_ (.CLK(\clknet_leaf_21_top1.acquisition_clk ),
    .RESET_B(net501),
    .D(_00878_),
    .Q_N(_09101_),
    .Q(\top1.memory1.mem1[69][1] ));
 sg13g2_dfrbp_1 _20678_ (.CLK(\clknet_leaf_21_top1.acquisition_clk ),
    .RESET_B(net500),
    .D(_00879_),
    .Q_N(_09100_),
    .Q(\top1.memory1.mem1[69][2] ));
 sg13g2_dfrbp_1 _20679_ (.CLK(\clknet_leaf_36_top1.acquisition_clk ),
    .RESET_B(net499),
    .D(_00880_),
    .Q_N(_09099_),
    .Q(\top1.memory1.mem1[6][0] ));
 sg13g2_dfrbp_1 _20680_ (.CLK(\clknet_leaf_266_top1.acquisition_clk ),
    .RESET_B(net498),
    .D(_00881_),
    .Q_N(_09098_),
    .Q(\top1.memory1.mem1[6][1] ));
 sg13g2_dfrbp_1 _20681_ (.CLK(\clknet_leaf_266_top1.acquisition_clk ),
    .RESET_B(net497),
    .D(_00882_),
    .Q_N(_09097_),
    .Q(\top1.memory1.mem1[6][2] ));
 sg13g2_dfrbp_1 _20682_ (.CLK(\clknet_leaf_36_top1.acquisition_clk ),
    .RESET_B(net496),
    .D(_00883_),
    .Q_N(_09096_),
    .Q(\top1.memory1.mem1[193][0] ));
 sg13g2_dfrbp_1 _20683_ (.CLK(\clknet_leaf_35_top1.acquisition_clk ),
    .RESET_B(net495),
    .D(_00884_),
    .Q_N(_09095_),
    .Q(\top1.memory1.mem1[193][1] ));
 sg13g2_dfrbp_1 _20684_ (.CLK(\clknet_leaf_36_top1.acquisition_clk ),
    .RESET_B(net494),
    .D(_00885_),
    .Q_N(_09094_),
    .Q(\top1.memory1.mem1[193][2] ));
 sg13g2_dfrbp_1 _20685_ (.CLK(\clknet_leaf_21_top1.acquisition_clk ),
    .RESET_B(net493),
    .D(_00886_),
    .Q_N(_09093_),
    .Q(\top1.memory1.mem1[70][0] ));
 sg13g2_dfrbp_1 _20686_ (.CLK(\clknet_leaf_10_top1.acquisition_clk ),
    .RESET_B(net492),
    .D(_00887_),
    .Q_N(_09092_),
    .Q(\top1.memory1.mem1[70][1] ));
 sg13g2_dfrbp_1 _20687_ (.CLK(\clknet_leaf_22_top1.acquisition_clk ),
    .RESET_B(net491),
    .D(_00888_),
    .Q_N(_09091_),
    .Q(\top1.memory1.mem1[70][2] ));
 sg13g2_dfrbp_1 _20688_ (.CLK(\clknet_leaf_11_top1.acquisition_clk ),
    .RESET_B(net490),
    .D(_00889_),
    .Q_N(_09090_),
    .Q(\top1.memory1.mem1[71][0] ));
 sg13g2_dfrbp_1 _20689_ (.CLK(\clknet_leaf_10_top1.acquisition_clk ),
    .RESET_B(net489),
    .D(_00890_),
    .Q_N(_09089_),
    .Q(\top1.memory1.mem1[71][1] ));
 sg13g2_dfrbp_1 _20690_ (.CLK(\clknet_leaf_22_top1.acquisition_clk ),
    .RESET_B(net488),
    .D(_00891_),
    .Q_N(_09088_),
    .Q(\top1.memory1.mem1[71][2] ));
 sg13g2_dfrbp_1 _20691_ (.CLK(\clknet_leaf_5_top1.acquisition_clk ),
    .RESET_B(net487),
    .D(_00892_),
    .Q_N(_09087_),
    .Q(\top1.memory1.mem1[72][0] ));
 sg13g2_dfrbp_1 _20692_ (.CLK(\clknet_leaf_12_top1.acquisition_clk ),
    .RESET_B(net486),
    .D(_00893_),
    .Q_N(_09086_),
    .Q(\top1.memory1.mem1[72][1] ));
 sg13g2_dfrbp_1 _20693_ (.CLK(\clknet_leaf_5_top1.acquisition_clk ),
    .RESET_B(net485),
    .D(_00894_),
    .Q_N(_09085_),
    .Q(\top1.memory1.mem1[72][2] ));
 sg13g2_dfrbp_1 _20694_ (.CLK(\clknet_leaf_262_top1.acquisition_clk ),
    .RESET_B(net484),
    .D(_00895_),
    .Q_N(_09084_),
    .Q(\top1.memory1.mem1[192][0] ));
 sg13g2_dfrbp_1 _20695_ (.CLK(\clknet_leaf_267_top1.acquisition_clk ),
    .RESET_B(net483),
    .D(_00896_),
    .Q_N(_09083_),
    .Q(\top1.memory1.mem1[192][1] ));
 sg13g2_dfrbp_1 _20696_ (.CLK(\clknet_leaf_36_top1.acquisition_clk ),
    .RESET_B(net482),
    .D(_00897_),
    .Q_N(_09082_),
    .Q(\top1.memory1.mem1[192][2] ));
 sg13g2_dfrbp_1 _20697_ (.CLK(\clknet_leaf_253_top1.acquisition_clk ),
    .RESET_B(net481),
    .D(_00898_),
    .Q_N(_09081_),
    .Q(\top1.memory1.mem1[191][0] ));
 sg13g2_dfrbp_1 _20698_ (.CLK(\clknet_leaf_191_top1.acquisition_clk ),
    .RESET_B(net480),
    .D(_00899_),
    .Q_N(_09080_),
    .Q(\top1.memory1.mem1[191][1] ));
 sg13g2_dfrbp_1 _20699_ (.CLK(\clknet_leaf_186_top1.acquisition_clk ),
    .RESET_B(net479),
    .D(_00900_),
    .Q_N(_09079_),
    .Q(\top1.memory1.mem1[191][2] ));
 sg13g2_dfrbp_1 _20700_ (.CLK(\clknet_leaf_253_top1.acquisition_clk ),
    .RESET_B(net478),
    .D(_00901_),
    .Q_N(_09078_),
    .Q(\top1.memory1.mem1[190][0] ));
 sg13g2_dfrbp_1 _20701_ (.CLK(\clknet_leaf_186_top1.acquisition_clk ),
    .RESET_B(net477),
    .D(_00902_),
    .Q_N(_09077_),
    .Q(\top1.memory1.mem1[190][1] ));
 sg13g2_dfrbp_1 _20702_ (.CLK(\clknet_leaf_186_top1.acquisition_clk ),
    .RESET_B(net476),
    .D(_00903_),
    .Q_N(_09076_),
    .Q(\top1.memory1.mem1[190][2] ));
 sg13g2_dfrbp_1 _20703_ (.CLK(\clknet_leaf_108_top1.acquisition_clk ),
    .RESET_B(net475),
    .D(_00904_),
    .Q_N(_09075_),
    .Q(\top1.memory1.mem1[18][0] ));
 sg13g2_dfrbp_1 _20704_ (.CLK(\clknet_leaf_182_top1.acquisition_clk ),
    .RESET_B(net474),
    .D(_00905_),
    .Q_N(_09074_),
    .Q(\top1.memory1.mem1[18][1] ));
 sg13g2_dfrbp_1 _20705_ (.CLK(\clknet_leaf_108_top1.acquisition_clk ),
    .RESET_B(net473),
    .D(_00906_),
    .Q_N(_09073_),
    .Q(\top1.memory1.mem1[18][2] ));
 sg13g2_dfrbp_1 _20706_ (.CLK(\clknet_leaf_14_top1.acquisition_clk ),
    .RESET_B(net472),
    .D(_00907_),
    .Q_N(_09072_),
    .Q(\top1.memory1.mem1[79][0] ));
 sg13g2_dfrbp_1 _20707_ (.CLK(\clknet_leaf_13_top1.acquisition_clk ),
    .RESET_B(net471),
    .D(_00908_),
    .Q_N(_09071_),
    .Q(\top1.memory1.mem1[79][1] ));
 sg13g2_dfrbp_1 _20708_ (.CLK(\clknet_leaf_15_top1.acquisition_clk ),
    .RESET_B(net470),
    .D(_00909_),
    .Q_N(_09070_),
    .Q(\top1.memory1.mem1[79][2] ));
 sg13g2_dfrbp_1 _20709_ (.CLK(\clknet_leaf_268_top1.acquisition_clk ),
    .RESET_B(net469),
    .D(_00910_),
    .Q_N(_09069_),
    .Q(\top1.memory1.mem1[89][0] ));
 sg13g2_dfrbp_1 _20710_ (.CLK(\clknet_leaf_283_top1.acquisition_clk ),
    .RESET_B(net468),
    .D(_00911_),
    .Q_N(_09068_),
    .Q(\top1.memory1.mem1[89][1] ));
 sg13g2_dfrbp_1 _20711_ (.CLK(\clknet_leaf_288_top1.acquisition_clk ),
    .RESET_B(net467),
    .D(_00912_),
    .Q_N(_09067_),
    .Q(\top1.memory1.mem1[89][2] ));
 sg13g2_dfrbp_1 _20712_ (.CLK(\clknet_leaf_253_top1.acquisition_clk ),
    .RESET_B(net466),
    .D(_00913_),
    .Q_N(_09066_),
    .Q(\top1.memory1.mem1[188][0] ));
 sg13g2_dfrbp_1 _20713_ (.CLK(\clknet_leaf_258_top1.acquisition_clk ),
    .RESET_B(net465),
    .D(_00914_),
    .Q_N(_09065_),
    .Q(\top1.memory1.mem1[188][1] ));
 sg13g2_dfrbp_1 _20714_ (.CLK(\clknet_leaf_186_top1.acquisition_clk ),
    .RESET_B(net464),
    .D(_00915_),
    .Q_N(_09064_),
    .Q(\top1.memory1.mem1[188][2] ));
 sg13g2_dfrbp_1 _20715_ (.CLK(\clknet_leaf_232_top1.acquisition_clk ),
    .RESET_B(net463),
    .D(_00916_),
    .Q_N(_09063_),
    .Q(\top1.memory1.mem1[187][0] ));
 sg13g2_dfrbp_1 _20716_ (.CLK(\clknet_leaf_249_top1.acquisition_clk ),
    .RESET_B(net462),
    .D(_00917_),
    .Q_N(_09062_),
    .Q(\top1.memory1.mem1[187][1] ));
 sg13g2_dfrbp_1 _20717_ (.CLK(\clknet_leaf_255_top1.acquisition_clk ),
    .RESET_B(net461),
    .D(_00918_),
    .Q_N(_09061_),
    .Q(\top1.memory1.mem1[187][2] ));
 sg13g2_dfrbp_1 _20718_ (.CLK(\clknet_leaf_243_top1.acquisition_clk ),
    .RESET_B(net460),
    .D(_00919_),
    .Q_N(_09060_),
    .Q(\top1.memory1.mem1[186][0] ));
 sg13g2_dfrbp_1 _20719_ (.CLK(\clknet_leaf_244_top1.acquisition_clk ),
    .RESET_B(net459),
    .D(_00920_),
    .Q_N(_09059_),
    .Q(\top1.memory1.mem1[186][1] ));
 sg13g2_dfrbp_1 _20720_ (.CLK(\clknet_leaf_248_top1.acquisition_clk ),
    .RESET_B(net458),
    .D(_00921_),
    .Q_N(_09058_),
    .Q(\top1.memory1.mem1[186][2] ));
 sg13g2_dfrbp_1 _20721_ (.CLK(\clknet_leaf_5_top1.acquisition_clk ),
    .RESET_B(net457),
    .D(_00922_),
    .Q_N(_09057_),
    .Q(\top1.memory1.mem1[73][0] ));
 sg13g2_dfrbp_1 _20722_ (.CLK(\clknet_leaf_12_top1.acquisition_clk ),
    .RESET_B(net456),
    .D(_00923_),
    .Q_N(_09056_),
    .Q(\top1.memory1.mem1[73][1] ));
 sg13g2_dfrbp_1 _20723_ (.CLK(\clknet_leaf_10_top1.acquisition_clk ),
    .RESET_B(net455),
    .D(_00924_),
    .Q_N(_09055_),
    .Q(\top1.memory1.mem1[73][2] ));
 sg13g2_dfrbp_1 _20724_ (.CLK(\clknet_leaf_243_top1.acquisition_clk ),
    .RESET_B(net454),
    .D(_00925_),
    .Q_N(_09054_),
    .Q(\top1.memory1.mem1[185][0] ));
 sg13g2_dfrbp_1 _20725_ (.CLK(\clknet_leaf_248_top1.acquisition_clk ),
    .RESET_B(net453),
    .D(_00926_),
    .Q_N(_09053_),
    .Q(\top1.memory1.mem1[185][1] ));
 sg13g2_dfrbp_1 _20726_ (.CLK(\clknet_leaf_254_top1.acquisition_clk ),
    .RESET_B(net452),
    .D(_00927_),
    .Q_N(_09052_),
    .Q(\top1.memory1.mem1[185][2] ));
 sg13g2_dfrbp_1 _20727_ (.CLK(\clknet_leaf_12_top1.acquisition_clk ),
    .RESET_B(net451),
    .D(_00928_),
    .Q_N(_09051_),
    .Q(\top1.memory1.mem1[74][0] ));
 sg13g2_dfrbp_1 _20728_ (.CLK(\clknet_leaf_12_top1.acquisition_clk ),
    .RESET_B(net450),
    .D(_00929_),
    .Q_N(_09050_),
    .Q(\top1.memory1.mem1[74][1] ));
 sg13g2_dfrbp_1 _20729_ (.CLK(\clknet_leaf_11_top1.acquisition_clk ),
    .RESET_B(net449),
    .D(_00930_),
    .Q_N(_09049_),
    .Q(\top1.memory1.mem1[74][2] ));
 sg13g2_dfrbp_1 _20730_ (.CLK(\clknet_leaf_12_top1.acquisition_clk ),
    .RESET_B(net448),
    .D(_00931_),
    .Q_N(_09048_),
    .Q(\top1.memory1.mem1[75][0] ));
 sg13g2_dfrbp_1 _20731_ (.CLK(\clknet_leaf_12_top1.acquisition_clk ),
    .RESET_B(net447),
    .D(_00932_),
    .Q_N(_09047_),
    .Q(\top1.memory1.mem1[75][1] ));
 sg13g2_dfrbp_1 _20732_ (.CLK(\clknet_leaf_12_top1.acquisition_clk ),
    .RESET_B(net446),
    .D(_00933_),
    .Q_N(_09046_),
    .Q(\top1.memory1.mem1[75][2] ));
 sg13g2_dfrbp_1 _20733_ (.CLK(\clknet_leaf_244_top1.acquisition_clk ),
    .RESET_B(net445),
    .D(_00934_),
    .Q_N(_09045_),
    .Q(\top1.memory1.mem1[184][0] ));
 sg13g2_dfrbp_1 _20734_ (.CLK(\clknet_leaf_244_top1.acquisition_clk ),
    .RESET_B(net444),
    .D(_00935_),
    .Q_N(_09044_),
    .Q(\top1.memory1.mem1[184][1] ));
 sg13g2_dfrbp_1 _20735_ (.CLK(\clknet_leaf_254_top1.acquisition_clk ),
    .RESET_B(net443),
    .D(_00936_),
    .Q_N(_09043_),
    .Q(\top1.memory1.mem1[184][2] ));
 sg13g2_dfrbp_1 _20736_ (.CLK(\clknet_leaf_238_top1.acquisition_clk ),
    .RESET_B(net442),
    .D(_00937_),
    .Q_N(_09042_),
    .Q(\top1.memory1.mem1[183][0] ));
 sg13g2_dfrbp_1 _20737_ (.CLK(\clknet_leaf_239_top1.acquisition_clk ),
    .RESET_B(net441),
    .D(_00938_),
    .Q_N(_09041_),
    .Q(\top1.memory1.mem1[183][1] ));
 sg13g2_dfrbp_1 _20738_ (.CLK(\clknet_leaf_232_top1.acquisition_clk ),
    .RESET_B(net440),
    .D(_00939_),
    .Q_N(_09040_),
    .Q(\top1.memory1.mem1[183][2] ));
 sg13g2_dfrbp_1 _20739_ (.CLK(\clknet_leaf_238_top1.acquisition_clk ),
    .RESET_B(net439),
    .D(_00940_),
    .Q_N(_09039_),
    .Q(\top1.memory1.mem1[182][0] ));
 sg13g2_dfrbp_1 _20740_ (.CLK(\clknet_leaf_238_top1.acquisition_clk ),
    .RESET_B(net438),
    .D(_00941_),
    .Q_N(_09038_),
    .Q(\top1.memory1.mem1[182][1] ));
 sg13g2_dfrbp_1 _20741_ (.CLK(\clknet_leaf_232_top1.acquisition_clk ),
    .RESET_B(net437),
    .D(_00942_),
    .Q_N(_09037_),
    .Q(\top1.memory1.mem1[182][2] ));
 sg13g2_dfrbp_1 _20742_ (.CLK(\clknet_leaf_238_top1.acquisition_clk ),
    .RESET_B(net436),
    .D(_00943_),
    .Q_N(_09036_),
    .Q(\top1.memory1.mem1[181][0] ));
 sg13g2_dfrbp_1 _20743_ (.CLK(\clknet_leaf_239_top1.acquisition_clk ),
    .RESET_B(net435),
    .D(_00944_),
    .Q_N(_09035_),
    .Q(\top1.memory1.mem1[181][1] ));
 sg13g2_dfrbp_1 _20744_ (.CLK(\clknet_leaf_237_top1.acquisition_clk ),
    .RESET_B(net434),
    .D(_00945_),
    .Q_N(_09034_),
    .Q(\top1.memory1.mem1[181][2] ));
 sg13g2_dfrbp_1 _20745_ (.CLK(\clknet_leaf_238_top1.acquisition_clk ),
    .RESET_B(net433),
    .D(_00946_),
    .Q_N(_09033_),
    .Q(\top1.memory1.mem1[180][0] ));
 sg13g2_dfrbp_1 _20746_ (.CLK(\clknet_leaf_239_top1.acquisition_clk ),
    .RESET_B(net432),
    .D(_00947_),
    .Q_N(_09032_),
    .Q(\top1.memory1.mem1[180][1] ));
 sg13g2_dfrbp_1 _20747_ (.CLK(\clknet_leaf_237_top1.acquisition_clk ),
    .RESET_B(net431),
    .D(_00948_),
    .Q_N(_09031_),
    .Q(\top1.memory1.mem1[180][2] ));
 sg13g2_dfrbp_1 _20748_ (.CLK(\clknet_leaf_109_top1.acquisition_clk ),
    .RESET_B(net430),
    .D(_00949_),
    .Q_N(_09030_),
    .Q(\top1.memory1.mem1[17][0] ));
 sg13g2_dfrbp_1 _20749_ (.CLK(\clknet_leaf_182_top1.acquisition_clk ),
    .RESET_B(net429),
    .D(_00950_),
    .Q_N(_09029_),
    .Q(\top1.memory1.mem1[17][1] ));
 sg13g2_dfrbp_1 _20750_ (.CLK(\clknet_leaf_108_top1.acquisition_clk ),
    .RESET_B(net428),
    .D(_00951_),
    .Q_N(_09028_),
    .Q(\top1.memory1.mem1[17][2] ));
 sg13g2_dfrbp_1 _20751_ (.CLK(\clknet_leaf_188_top1.acquisition_clk ),
    .RESET_B(net427),
    .D(_00952_),
    .Q_N(_09027_),
    .Q(\top1.memory1.mem1[99][0] ));
 sg13g2_dfrbp_1 _20752_ (.CLK(\clknet_leaf_179_top1.acquisition_clk ),
    .RESET_B(net426),
    .D(_00953_),
    .Q_N(_09026_),
    .Q(\top1.memory1.mem1[99][1] ));
 sg13g2_dfrbp_1 _20753_ (.CLK(\clknet_leaf_187_top1.acquisition_clk ),
    .RESET_B(net425),
    .D(_00954_),
    .Q_N(_09025_),
    .Q(\top1.memory1.mem1[99][2] ));
 sg13g2_dfrbp_1 _20754_ (.CLK(\clknet_leaf_252_top1.acquisition_clk ),
    .RESET_B(net424),
    .D(_00955_),
    .Q_N(_09024_),
    .Q(\top1.memory1.mem1[178][0] ));
 sg13g2_dfrbp_1 _20755_ (.CLK(\clknet_leaf_248_top1.acquisition_clk ),
    .RESET_B(net423),
    .D(_00956_),
    .Q_N(_09023_),
    .Q(\top1.memory1.mem1[178][1] ));
 sg13g2_dfrbp_1 _20756_ (.CLK(\clknet_leaf_190_top1.acquisition_clk ),
    .RESET_B(net422),
    .D(_00957_),
    .Q_N(_09022_),
    .Q(\top1.memory1.mem1[178][2] ));
 sg13g2_dfrbp_1 _20757_ (.CLK(\clknet_leaf_252_top1.acquisition_clk ),
    .RESET_B(net421),
    .D(_00958_),
    .Q_N(_09021_),
    .Q(\top1.memory1.mem1[177][0] ));
 sg13g2_dfrbp_1 _20758_ (.CLK(\clknet_leaf_248_top1.acquisition_clk ),
    .RESET_B(net420),
    .D(_00959_),
    .Q_N(_09020_),
    .Q(\top1.memory1.mem1[177][1] ));
 sg13g2_dfrbp_1 _20759_ (.CLK(\clknet_leaf_191_top1.acquisition_clk ),
    .RESET_B(net419),
    .D(_00960_),
    .Q_N(_09019_),
    .Q(\top1.memory1.mem1[177][2] ));
 sg13g2_dfrbp_1 _20760_ (.CLK(\clknet_leaf_198_top1.acquisition_clk ),
    .RESET_B(net418),
    .D(_00961_),
    .Q_N(_09018_),
    .Q(\top1.memory1.mem1[109][0] ));
 sg13g2_dfrbp_1 _20761_ (.CLK(\clknet_leaf_197_top1.acquisition_clk ),
    .RESET_B(net417),
    .D(_00962_),
    .Q_N(_09017_),
    .Q(\top1.memory1.mem1[109][1] ));
 sg13g2_dfrbp_1 _20762_ (.CLK(\clknet_leaf_195_top1.acquisition_clk ),
    .RESET_B(net416),
    .D(_00963_),
    .Q_N(_09016_),
    .Q(\top1.memory1.mem1[109][2] ));
 sg13g2_dfrbp_1 _20763_ (.CLK(\clknet_leaf_253_top1.acquisition_clk ),
    .RESET_B(net415),
    .D(_00964_),
    .Q_N(_09015_),
    .Q(\top1.memory1.mem1[176][0] ));
 sg13g2_dfrbp_1 _20764_ (.CLK(\clknet_leaf_248_top1.acquisition_clk ),
    .RESET_B(net414),
    .D(_00965_),
    .Q_N(_09014_),
    .Q(\top1.memory1.mem1[176][1] ));
 sg13g2_dfrbp_1 _20765_ (.CLK(\clknet_leaf_253_top1.acquisition_clk ),
    .RESET_B(net413),
    .D(_00966_),
    .Q_N(_09013_),
    .Q(\top1.memory1.mem1[176][2] ));
 sg13g2_dfrbp_1 _20766_ (.CLK(\clknet_leaf_241_top1.acquisition_clk ),
    .RESET_B(net412),
    .D(_00967_),
    .Q_N(_09012_),
    .Q(\top1.memory1.mem1[175][0] ));
 sg13g2_dfrbp_1 _20767_ (.CLK(\clknet_leaf_240_top1.acquisition_clk ),
    .RESET_B(net411),
    .D(_00968_),
    .Q_N(_09011_),
    .Q(\top1.memory1.mem1[175][1] ));
 sg13g2_dfrbp_1 _20768_ (.CLK(\clknet_leaf_246_top1.acquisition_clk ),
    .RESET_B(net410),
    .D(_00969_),
    .Q_N(_09010_),
    .Q(\top1.memory1.mem1[175][2] ));
 sg13g2_dfrbp_1 _20769_ (.CLK(\clknet_leaf_241_top1.acquisition_clk ),
    .RESET_B(net409),
    .D(_00970_),
    .Q_N(_09009_),
    .Q(\top1.memory1.mem1[174][0] ));
 sg13g2_dfrbp_1 _20770_ (.CLK(\clknet_leaf_240_top1.acquisition_clk ),
    .RESET_B(net408),
    .D(_00971_),
    .Q_N(_09008_),
    .Q(\top1.memory1.mem1[174][1] ));
 sg13g2_dfrbp_1 _20771_ (.CLK(\clknet_leaf_246_top1.acquisition_clk ),
    .RESET_B(net407),
    .D(_00972_),
    .Q_N(_09007_),
    .Q(\top1.memory1.mem1[174][2] ));
 sg13g2_dfrbp_1 _20772_ (.CLK(\clknet_leaf_241_top1.acquisition_clk ),
    .RESET_B(net406),
    .D(_00973_),
    .Q_N(_09006_),
    .Q(\top1.memory1.mem1[173][0] ));
 sg13g2_dfrbp_1 _20773_ (.CLK(\clknet_leaf_240_top1.acquisition_clk ),
    .RESET_B(net405),
    .D(_00974_),
    .Q_N(_09005_),
    .Q(\top1.memory1.mem1[173][1] ));
 sg13g2_dfrbp_1 _20774_ (.CLK(\clknet_leaf_246_top1.acquisition_clk ),
    .RESET_B(net404),
    .D(_00975_),
    .Q_N(_09004_),
    .Q(\top1.memory1.mem1[173][2] ));
 sg13g2_dfrbp_1 _20775_ (.CLK(\clknet_leaf_242_top1.acquisition_clk ),
    .RESET_B(net403),
    .D(_00976_),
    .Q_N(_09003_),
    .Q(\top1.memory1.mem1[172][0] ));
 sg13g2_dfrbp_1 _20776_ (.CLK(\clknet_leaf_240_top1.acquisition_clk ),
    .RESET_B(net402),
    .D(_00977_),
    .Q_N(_09002_),
    .Q(\top1.memory1.mem1[172][1] ));
 sg13g2_dfrbp_1 _20777_ (.CLK(\clknet_leaf_246_top1.acquisition_clk ),
    .RESET_B(net401),
    .D(_00978_),
    .Q_N(_09001_),
    .Q(\top1.memory1.mem1[172][2] ));
 sg13g2_dfrbp_1 _20778_ (.CLK(\clknet_leaf_245_top1.acquisition_clk ),
    .RESET_B(net400),
    .D(_00979_),
    .Q_N(_09000_),
    .Q(\top1.memory1.mem1[171][0] ));
 sg13g2_dfrbp_1 _20779_ (.CLK(\clknet_leaf_245_top1.acquisition_clk ),
    .RESET_B(net399),
    .D(_00980_),
    .Q_N(_08999_),
    .Q(\top1.memory1.mem1[171][1] ));
 sg13g2_dfrbp_1 _20780_ (.CLK(\clknet_leaf_255_top1.acquisition_clk ),
    .RESET_B(net398),
    .D(_00981_),
    .Q_N(_08998_),
    .Q(\top1.memory1.mem1[171][2] ));
 sg13g2_dfrbp_1 _20781_ (.CLK(\clknet_leaf_245_top1.acquisition_clk ),
    .RESET_B(net397),
    .D(_00982_),
    .Q_N(_08997_),
    .Q(\top1.memory1.mem1[170][0] ));
 sg13g2_dfrbp_1 _20782_ (.CLK(\clknet_leaf_242_top1.acquisition_clk ),
    .RESET_B(net396),
    .D(_00983_),
    .Q_N(_08996_),
    .Q(\top1.memory1.mem1[170][1] ));
 sg13g2_dfrbp_1 _20783_ (.CLK(\clknet_leaf_256_top1.acquisition_clk ),
    .RESET_B(net395),
    .D(_00984_),
    .Q_N(_08995_),
    .Q(\top1.memory1.mem1[170][2] ));
 sg13g2_dfrbp_1 _20784_ (.CLK(\clknet_leaf_108_top1.acquisition_clk ),
    .RESET_B(net394),
    .D(_00985_),
    .Q_N(_08994_),
    .Q(\top1.memory1.mem1[16][0] ));
 sg13g2_dfrbp_1 _20785_ (.CLK(\clknet_leaf_183_top1.acquisition_clk ),
    .RESET_B(net393),
    .D(_00986_),
    .Q_N(_08993_),
    .Q(\top1.memory1.mem1[16][1] ));
 sg13g2_dfrbp_1 _20786_ (.CLK(\clknet_leaf_109_top1.acquisition_clk ),
    .RESET_B(net392),
    .D(_00987_),
    .Q_N(_08992_),
    .Q(\top1.memory1.mem1[16][2] ));
 sg13g2_dfrbp_1 _20787_ (.CLK(\clknet_leaf_245_top1.acquisition_clk ),
    .RESET_B(net391),
    .D(_00988_),
    .Q_N(_08991_),
    .Q(\top1.memory1.mem1[168][0] ));
 sg13g2_dfrbp_1 _20788_ (.CLK(\clknet_leaf_245_top1.acquisition_clk ),
    .RESET_B(net390),
    .D(_00989_),
    .Q_N(_08990_),
    .Q(\top1.memory1.mem1[168][1] ));
 sg13g2_dfrbp_1 _20789_ (.CLK(\clknet_leaf_256_top1.acquisition_clk ),
    .RESET_B(net389),
    .D(_00990_),
    .Q_N(_08989_),
    .Q(\top1.memory1.mem1[168][2] ));
 sg13g2_dfrbp_1 _20790_ (.CLK(\clknet_leaf_239_top1.acquisition_clk ),
    .RESET_B(net388),
    .D(_00991_),
    .Q_N(_08988_),
    .Q(\top1.memory1.mem1[167][0] ));
 sg13g2_dfrbp_1 _20791_ (.CLK(\clknet_leaf_240_top1.acquisition_clk ),
    .RESET_B(net387),
    .D(_00992_),
    .Q_N(_08987_),
    .Q(\top1.memory1.mem1[167][1] ));
 sg13g2_dfrbp_1 _20792_ (.CLK(\clknet_leaf_255_top1.acquisition_clk ),
    .RESET_B(net386),
    .D(_00993_),
    .Q_N(_08986_),
    .Q(\top1.memory1.mem1[167][2] ));
 sg13g2_dfrbp_1 _20793_ (.CLK(\clknet_leaf_240_top1.acquisition_clk ),
    .RESET_B(net385),
    .D(_00994_),
    .Q_N(_08985_),
    .Q(\top1.memory1.mem1[166][0] ));
 sg13g2_dfrbp_1 _20794_ (.CLK(\clknet_leaf_239_top1.acquisition_clk ),
    .RESET_B(net384),
    .D(_00995_),
    .Q_N(_08984_),
    .Q(\top1.memory1.mem1[166][1] ));
 sg13g2_dfrbp_1 _20795_ (.CLK(\clknet_leaf_255_top1.acquisition_clk ),
    .RESET_B(net935),
    .D(_00996_),
    .Q_N(_09906_),
    .Q(\top1.memory1.mem1[166][2] ));
 sg13g2_dfrbp_1 _20796_ (.CLK(net6740),
    .RESET_B(net7734),
    .D(_00046_),
    .Q_N(_08983_),
    .Q(\top1.PISO_time ));
 sg13g2_dfrbp_1 _20797_ (.CLK(\clknet_leaf_17_top1.acquisition_clk ),
    .RESET_B(net383),
    .D(_00997_),
    .Q_N(_08982_),
    .Q(\top1.memory1.mem1[128][0] ));
 sg13g2_dfrbp_1 _20798_ (.CLK(\clknet_leaf_19_top1.acquisition_clk ),
    .RESET_B(net382),
    .D(_00998_),
    .Q_N(_08981_),
    .Q(\top1.memory1.mem1[128][1] ));
 sg13g2_dfrbp_1 _20799_ (.CLK(\clknet_leaf_19_top1.acquisition_clk ),
    .RESET_B(net381),
    .D(_00999_),
    .Q_N(_08980_),
    .Q(\top1.memory1.mem1[128][2] ));
 sg13g2_dfrbp_1 _20800_ (.CLK(\clknet_leaf_208_top1.acquisition_clk ),
    .RESET_B(net380),
    .D(_01000_),
    .Q_N(_08979_),
    .Q(\top1.memory1.mem1[127][0] ));
 sg13g2_dfrbp_1 _20801_ (.CLK(\clknet_leaf_207_top1.acquisition_clk ),
    .RESET_B(net379),
    .D(_01001_),
    .Q_N(_08978_),
    .Q(\top1.memory1.mem1[127][1] ));
 sg13g2_dfrbp_1 _20802_ (.CLK(\clknet_leaf_205_top1.acquisition_clk ),
    .RESET_B(net378),
    .D(_01002_),
    .Q_N(_08977_),
    .Q(\top1.memory1.mem1[127][2] ));
 sg13g2_dfrbp_1 _20803_ (.CLK(\clknet_leaf_208_top1.acquisition_clk ),
    .RESET_B(net377),
    .D(_01003_),
    .Q_N(_08976_),
    .Q(\top1.memory1.mem1[126][0] ));
 sg13g2_dfrbp_1 _20804_ (.CLK(\clknet_leaf_207_top1.acquisition_clk ),
    .RESET_B(net376),
    .D(_01004_),
    .Q_N(_08975_),
    .Q(\top1.memory1.mem1[126][1] ));
 sg13g2_dfrbp_1 _20805_ (.CLK(\clknet_leaf_204_top1.acquisition_clk ),
    .RESET_B(net375),
    .D(_01005_),
    .Q_N(_08974_),
    .Q(\top1.memory1.mem1[126][2] ));
 sg13g2_dfrbp_1 _20806_ (.CLK(\clknet_leaf_207_top1.acquisition_clk ),
    .RESET_B(net374),
    .D(_01006_),
    .Q_N(_08973_),
    .Q(\top1.memory1.mem1[125][0] ));
 sg13g2_dfrbp_1 _20807_ (.CLK(\clknet_leaf_215_top1.acquisition_clk ),
    .RESET_B(net373),
    .D(_01007_),
    .Q_N(_08972_),
    .Q(\top1.memory1.mem1[125][1] ));
 sg13g2_dfrbp_1 _20808_ (.CLK(\clknet_leaf_204_top1.acquisition_clk ),
    .RESET_B(net372),
    .D(_01008_),
    .Q_N(_08971_),
    .Q(\top1.memory1.mem1[125][2] ));
 sg13g2_dfrbp_1 _20809_ (.CLK(\clknet_leaf_257_top1.acquisition_clk ),
    .RESET_B(net371),
    .D(_01009_),
    .Q_N(_08970_),
    .Q(\top1.memory1.mem1[31][0] ));
 sg13g2_dfrbp_1 _20810_ (.CLK(\clknet_leaf_256_top1.acquisition_clk ),
    .RESET_B(net370),
    .D(_01010_),
    .Q_N(_08969_),
    .Q(\top1.memory1.mem1[31][1] ));
 sg13g2_dfrbp_1 _20811_ (.CLK(\clknet_leaf_260_top1.acquisition_clk ),
    .RESET_B(net369),
    .D(_01011_),
    .Q_N(_08968_),
    .Q(\top1.memory1.mem1[31][2] ));
 sg13g2_dfrbp_1 _20812_ (.CLK(net7720),
    .RESET_B(net7735),
    .D(_01012_),
    .Q_N(_08967_),
    .Q(\top1.event_time[10] ));
 sg13g2_dfrbp_1 _20813_ (.CLK(net7720),
    .RESET_B(net7735),
    .D(_01013_),
    .Q_N(_08966_),
    .Q(\top1.event_time[11] ));
 sg13g2_dfrbp_1 _20814_ (.CLK(net7720),
    .RESET_B(net7735),
    .D(_01014_),
    .Q_N(_08965_),
    .Q(\top1.event_time[12] ));
 sg13g2_dfrbp_1 _20815_ (.CLK(net7721),
    .RESET_B(net7729),
    .D(_01015_),
    .Q_N(_08964_),
    .Q(\top1.event_time[13] ));
 sg13g2_dfrbp_1 _20816_ (.CLK(net7721),
    .RESET_B(net7730),
    .D(_01016_),
    .Q_N(_08963_),
    .Q(\top1.event_time[14] ));
 sg13g2_dfrbp_1 _20817_ (.CLK(net7721),
    .RESET_B(net7729),
    .D(_01017_),
    .Q_N(_08962_),
    .Q(\top1.event_time[15] ));
 sg13g2_dfrbp_1 _20818_ (.CLK(net6744),
    .RESET_B(net368),
    .D(_01018_),
    .Q_N(_08961_),
    .Q(\top1.memory2.data_out[0] ));
 sg13g2_dfrbp_1 _20819_ (.CLK(net6744),
    .RESET_B(net367),
    .D(_01019_),
    .Q_N(_08960_),
    .Q(\top1.memory2.data_out[1] ));
 sg13g2_dfrbp_1 _20820_ (.CLK(net6744),
    .RESET_B(net366),
    .D(_01020_),
    .Q_N(_08959_),
    .Q(\top1.memory2.data_out[2] ));
 sg13g2_dfrbp_1 _20821_ (.CLK(net7719),
    .RESET_B(net7727),
    .D(_01021_),
    .Q_N(_08958_),
    .Q(\top1.event_time[16] ));
 sg13g2_dfrbp_1 _20822_ (.CLK(net7719),
    .RESET_B(net7726),
    .D(_01022_),
    .Q_N(_08957_),
    .Q(\top1.event_time[17] ));
 sg13g2_dfrbp_1 _20823_ (.CLK(net7719),
    .RESET_B(net7726),
    .D(_01023_),
    .Q_N(_08956_),
    .Q(\top1.event_time[18] ));
 sg13g2_dfrbp_1 _20824_ (.CLK(net7719),
    .RESET_B(net7726),
    .D(_01024_),
    .Q_N(_08955_),
    .Q(\top1.event_time[19] ));
 sg13g2_dfrbp_1 _20825_ (.CLK(net8),
    .RESET_B(net7726),
    .D(_01025_),
    .Q_N(_08954_),
    .Q(\top1.event_time[20] ));
 sg13g2_dfrbp_1 _20826_ (.CLK(net7719),
    .RESET_B(net7726),
    .D(_01026_),
    .Q_N(_09907_),
    .Q(\top1.event_time[21] ));
 sg13g2_dfrbp_1 _20827_ (.CLK(net7722),
    .RESET_B(net7732),
    .D(_00053_),
    .Q_N(_09908_),
    .Q(\top1.event_time[0] ));
 sg13g2_dfrbp_1 _20828_ (.CLK(net7722),
    .RESET_B(net7732),
    .D(_00054_),
    .Q_N(_09909_),
    .Q(\top1.event_time[1] ));
 sg13g2_dfrbp_1 _20829_ (.CLK(net7722),
    .RESET_B(net7732),
    .D(_00055_),
    .Q_N(_09910_),
    .Q(\top1.event_time[2] ));
 sg13g2_dfrbp_1 _20830_ (.CLK(net7722),
    .RESET_B(net7732),
    .D(_00056_),
    .Q_N(_09911_),
    .Q(\top1.event_time[3] ));
 sg13g2_dfrbp_1 _20831_ (.CLK(net7722),
    .RESET_B(net7732),
    .D(_00057_),
    .Q_N(_09912_),
    .Q(\top1.event_time[4] ));
 sg13g2_dfrbp_1 _20832_ (.CLK(net7720),
    .RESET_B(net7736),
    .D(_00058_),
    .Q_N(_09913_),
    .Q(\top1.event_time[5] ));
 sg13g2_dfrbp_1 _20833_ (.CLK(net7720),
    .RESET_B(net7736),
    .D(_00059_),
    .Q_N(_09914_),
    .Q(\top1.event_time[6] ));
 sg13g2_dfrbp_1 _20834_ (.CLK(net7720),
    .RESET_B(net7736),
    .D(_00060_),
    .Q_N(_09915_),
    .Q(\top1.event_time[7] ));
 sg13g2_dfrbp_1 _20835_ (.CLK(net7720),
    .RESET_B(net7736),
    .D(_00061_),
    .Q_N(_09916_),
    .Q(\top1.event_time[8] ));
 sg13g2_dfrbp_1 _20836_ (.CLK(net7720),
    .RESET_B(net7736),
    .D(_00062_),
    .Q_N(_09917_),
    .Q(\top1.event_time[9] ));
 sg13g2_dfrbp_1 _20837_ (.CLK(net6737),
    .RESET_B(net7731),
    .D(_00052_),
    .Q_N(_08953_),
    .Q(\top1.reg2.serial_out ));
 sg13g2_dfrbp_1 _20838_ (.CLK(\clknet_leaf_253_top1.acquisition_clk ),
    .RESET_B(net365),
    .D(_01027_),
    .Q_N(_08952_),
    .Q(\top1.memory1.mem1[189][0] ));
 sg13g2_dfrbp_1 _20839_ (.CLK(\clknet_leaf_254_top1.acquisition_clk ),
    .RESET_B(net364),
    .D(_01028_),
    .Q_N(_08951_),
    .Q(\top1.memory1.mem1[189][1] ));
 sg13g2_dfrbp_1 _20840_ (.CLK(\clknet_leaf_187_top1.acquisition_clk ),
    .RESET_B(net1050),
    .D(_01029_),
    .Q_N(_09918_),
    .Q(\top1.memory1.mem1[189][2] ));
 sg13g2_dfrbp_1 _20841_ (.CLK(net6739),
    .RESET_B(net7741),
    .D(_00049_),
    .Q_N(_08950_),
    .Q(\top1.PISO_ch1 ));
 sg13g2_dfrbp_1 _20842_ (.CLK(\clknet_leaf_148_top1.acquisition_clk ),
    .RESET_B(net363),
    .D(_01030_),
    .Q_N(_08949_),
    .Q(\top1.memory1.mem1[33][0] ));
 sg13g2_dfrbp_1 _20843_ (.CLK(\clknet_leaf_147_top1.acquisition_clk ),
    .RESET_B(net362),
    .D(_01031_),
    .Q_N(_08948_),
    .Q(\top1.memory1.mem1[33][1] ));
 sg13g2_dfrbp_1 _20844_ (.CLK(\clknet_leaf_152_top1.acquisition_clk ),
    .RESET_B(net361),
    .D(_01032_),
    .Q_N(_08947_),
    .Q(\top1.memory1.mem1[33][2] ));
 sg13g2_dfrbp_1 _20845_ (.CLK(\clknet_leaf_145_top1.acquisition_clk ),
    .RESET_B(net360),
    .D(_01033_),
    .Q_N(_08946_),
    .Q(\top1.memory1.mem1[34][0] ));
 sg13g2_dfrbp_1 _20846_ (.CLK(\clknet_leaf_147_top1.acquisition_clk ),
    .RESET_B(net359),
    .D(_01034_),
    .Q_N(_08945_),
    .Q(\top1.memory1.mem1[34][1] ));
 sg13g2_dfrbp_1 _20847_ (.CLK(\clknet_leaf_152_top1.acquisition_clk ),
    .RESET_B(net358),
    .D(_01035_),
    .Q_N(_08944_),
    .Q(\top1.memory1.mem1[34][2] ));
 sg13g2_dfrbp_1 _20848_ (.CLK(\clknet_leaf_108_top1.acquisition_clk ),
    .RESET_B(net357),
    .D(_01036_),
    .Q_N(_08943_),
    .Q(\top1.memory1.mem1[19][0] ));
 sg13g2_dfrbp_1 _20849_ (.CLK(\clknet_leaf_182_top1.acquisition_clk ),
    .RESET_B(net356),
    .D(_01037_),
    .Q_N(_08942_),
    .Q(\top1.memory1.mem1[19][1] ));
 sg13g2_dfrbp_1 _20850_ (.CLK(\clknet_leaf_108_top1.acquisition_clk ),
    .RESET_B(net355),
    .D(_01038_),
    .Q_N(_08941_),
    .Q(\top1.memory1.mem1[19][2] ));
 sg13g2_dfrbp_1 _20851_ (.CLK(\clknet_leaf_188_top1.acquisition_clk ),
    .RESET_B(net354),
    .D(_01039_),
    .Q_N(_08940_),
    .Q(\top1.memory1.mem1[98][0] ));
 sg13g2_dfrbp_1 _20852_ (.CLK(\clknet_leaf_180_top1.acquisition_clk ),
    .RESET_B(net353),
    .D(_01040_),
    .Q_N(_08939_),
    .Q(\top1.memory1.mem1[98][1] ));
 sg13g2_dfrbp_1 _20853_ (.CLK(\clknet_leaf_190_top1.acquisition_clk ),
    .RESET_B(net352),
    .D(_01041_),
    .Q_N(_08938_),
    .Q(\top1.memory1.mem1[98][2] ));
 sg13g2_dfrbp_1 _20854_ (.CLK(\clknet_leaf_277_top1.acquisition_clk ),
    .RESET_B(net351),
    .D(_01042_),
    .Q_N(_08937_),
    .Q(\top1.memory1.mem1[2][0] ));
 sg13g2_dfrbp_1 _20855_ (.CLK(\clknet_leaf_278_top1.acquisition_clk ),
    .RESET_B(net350),
    .D(_01043_),
    .Q_N(_08936_),
    .Q(\top1.memory1.mem1[2][1] ));
 sg13g2_dfrbp_1 _20856_ (.CLK(\clknet_leaf_281_top1.acquisition_clk ),
    .RESET_B(net349),
    .D(_01044_),
    .Q_N(_08935_),
    .Q(\top1.memory1.mem1[2][2] ));
 sg13g2_dfrbp_1 _20857_ (.CLK(\clknet_leaf_188_top1.acquisition_clk ),
    .RESET_B(net348),
    .D(_01045_),
    .Q_N(_08934_),
    .Q(\top1.memory1.mem1[97][0] ));
 sg13g2_dfrbp_1 _20858_ (.CLK(\clknet_leaf_179_top1.acquisition_clk ),
    .RESET_B(net347),
    .D(_01046_),
    .Q_N(_08933_),
    .Q(\top1.memory1.mem1[97][1] ));
 sg13g2_dfrbp_1 _20859_ (.CLK(\clknet_leaf_190_top1.acquisition_clk ),
    .RESET_B(net346),
    .D(_01047_),
    .Q_N(_08932_),
    .Q(\top1.memory1.mem1[97][2] ));
 sg13g2_dfrbp_1 _20860_ (.CLK(\clknet_leaf_188_top1.acquisition_clk ),
    .RESET_B(net345),
    .D(_01048_),
    .Q_N(_08931_),
    .Q(\top1.memory1.mem1[96][0] ));
 sg13g2_dfrbp_1 _20861_ (.CLK(\clknet_leaf_180_top1.acquisition_clk ),
    .RESET_B(net344),
    .D(_01049_),
    .Q_N(_08930_),
    .Q(\top1.memory1.mem1[96][1] ));
 sg13g2_dfrbp_1 _20862_ (.CLK(\clknet_leaf_189_top1.acquisition_clk ),
    .RESET_B(net343),
    .D(_01050_),
    .Q_N(_08929_),
    .Q(\top1.memory1.mem1[96][2] ));
 sg13g2_dfrbp_1 _20863_ (.CLK(\clknet_leaf_257_top1.acquisition_clk ),
    .RESET_B(net342),
    .D(_01051_),
    .Q_N(_08928_),
    .Q(\top1.memory1.mem1[28][0] ));
 sg13g2_dfrbp_1 _20864_ (.CLK(\clknet_leaf_256_top1.acquisition_clk ),
    .RESET_B(net341),
    .D(_01052_),
    .Q_N(_08927_),
    .Q(\top1.memory1.mem1[28][1] ));
 sg13g2_dfrbp_1 _20865_ (.CLK(\clknet_leaf_259_top1.acquisition_clk ),
    .RESET_B(net340),
    .D(_01053_),
    .Q_N(_08926_),
    .Q(\top1.memory1.mem1[28][2] ));
 sg13g2_dfrbp_1 _20866_ (.CLK(net6744),
    .RESET_B(net339),
    .D(_01054_),
    .Q_N(_08925_),
    .Q(\top1.memory1.data_out[0] ));
 sg13g2_dfrbp_1 _20867_ (.CLK(net6744),
    .RESET_B(net338),
    .D(_01055_),
    .Q_N(_08924_),
    .Q(\top1.memory1.data_out[1] ));
 sg13g2_dfrbp_1 _20868_ (.CLK(net6744),
    .RESET_B(net337),
    .D(_01056_),
    .Q_N(_08923_),
    .Q(\top1.memory1.data_out[2] ));
 sg13g2_dfrbp_1 _20869_ (.CLK(\clknet_leaf_145_top1.acquisition_clk ),
    .RESET_B(net336),
    .D(_01057_),
    .Q_N(_08922_),
    .Q(\top1.memory1.mem1[35][0] ));
 sg13g2_dfrbp_1 _20870_ (.CLK(\clknet_leaf_147_top1.acquisition_clk ),
    .RESET_B(net335),
    .D(_01058_),
    .Q_N(_08921_),
    .Q(\top1.memory1.mem1[35][1] ));
 sg13g2_dfrbp_1 _20871_ (.CLK(\clknet_leaf_150_top1.acquisition_clk ),
    .RESET_B(net334),
    .D(_01059_),
    .Q_N(_08920_),
    .Q(\top1.memory1.mem1[35][2] ));
 sg13g2_dfrbp_1 _20872_ (.CLK(\clknet_leaf_188_top1.acquisition_clk ),
    .RESET_B(net333),
    .D(_01060_),
    .Q_N(_08919_),
    .Q(\top1.memory1.mem1[102][0] ));
 sg13g2_dfrbp_1 _20873_ (.CLK(\clknet_leaf_194_top1.acquisition_clk ),
    .RESET_B(net332),
    .D(_01061_),
    .Q_N(_08918_),
    .Q(\top1.memory1.mem1[102][1] ));
 sg13g2_dfrbp_1 _20874_ (.CLK(\clknet_leaf_190_top1.acquisition_clk ),
    .RESET_B(net331),
    .D(_01062_),
    .Q_N(_08917_),
    .Q(\top1.memory1.mem1[102][2] ));
 sg13g2_dfrbp_1 _20875_ (.CLK(\clknet_leaf_188_top1.acquisition_clk ),
    .RESET_B(net330),
    .D(_01063_),
    .Q_N(_08916_),
    .Q(\top1.memory1.mem1[101][0] ));
 sg13g2_dfrbp_1 _20876_ (.CLK(\clknet_leaf_195_top1.acquisition_clk ),
    .RESET_B(net329),
    .D(_01064_),
    .Q_N(_08915_),
    .Q(\top1.memory1.mem1[101][1] ));
 sg13g2_dfrbp_1 _20877_ (.CLK(\clknet_leaf_192_top1.acquisition_clk ),
    .RESET_B(net328),
    .D(_01065_),
    .Q_N(_08914_),
    .Q(\top1.memory1.mem1[101][2] ));
 sg13g2_dfrbp_1 _20878_ (.CLK(\clknet_leaf_189_top1.acquisition_clk ),
    .RESET_B(net327),
    .D(_01066_),
    .Q_N(_08913_),
    .Q(\top1.memory1.mem1[100][0] ));
 sg13g2_dfrbp_1 _20879_ (.CLK(\clknet_leaf_192_top1.acquisition_clk ),
    .RESET_B(net326),
    .D(_01067_),
    .Q_N(_08912_),
    .Q(\top1.memory1.mem1[100][1] ));
 sg13g2_dfrbp_1 _20880_ (.CLK(\clknet_leaf_192_top1.acquisition_clk ),
    .RESET_B(net325),
    .D(_01068_),
    .Q_N(_08911_),
    .Q(\top1.memory1.mem1[100][2] ));
 sg13g2_dfrbp_1 _20881_ (.CLK(\clknet_leaf_277_top1.acquisition_clk ),
    .RESET_B(net324),
    .D(_01069_),
    .Q_N(_08910_),
    .Q(\top1.memory1.mem1[0][0] ));
 sg13g2_dfrbp_1 _20882_ (.CLK(\clknet_leaf_280_top1.acquisition_clk ),
    .RESET_B(net323),
    .D(_01070_),
    .Q_N(_08909_),
    .Q(\top1.memory1.mem1[0][1] ));
 sg13g2_dfrbp_1 _20883_ (.CLK(\clknet_leaf_281_top1.acquisition_clk ),
    .RESET_B(net322),
    .D(_01071_),
    .Q_N(_08908_),
    .Q(\top1.memory1.mem1[0][2] ));
 sg13g2_dfrbp_1 _20884_ (.CLK(\clknet_leaf_181_top1.acquisition_clk ),
    .RESET_B(net321),
    .D(_01072_),
    .Q_N(_08907_),
    .Q(\top1.memory1.mem1[27][0] ));
 sg13g2_dfrbp_1 _20885_ (.CLK(\clknet_leaf_181_top1.acquisition_clk ),
    .RESET_B(net320),
    .D(_01073_),
    .Q_N(_08906_),
    .Q(\top1.memory1.mem1[27][1] ));
 sg13g2_dfrbp_1 _20886_ (.CLK(\clknet_leaf_182_top1.acquisition_clk ),
    .RESET_B(net319),
    .D(_01074_),
    .Q_N(_08905_),
    .Q(\top1.memory1.mem1[27][2] ));
 sg13g2_dfrbp_1 _20887_ (.CLK(\clknet_leaf_182_top1.acquisition_clk ),
    .RESET_B(net318),
    .D(_01075_),
    .Q_N(_08904_),
    .Q(\top1.memory1.mem1[26][0] ));
 sg13g2_dfrbp_1 _20888_ (.CLK(\clknet_leaf_181_top1.acquisition_clk ),
    .RESET_B(net317),
    .D(_01076_),
    .Q_N(_08903_),
    .Q(\top1.memory1.mem1[26][1] ));
 sg13g2_dfrbp_1 _20889_ (.CLK(\clknet_leaf_108_top1.acquisition_clk ),
    .RESET_B(net316),
    .D(_01077_),
    .Q_N(_08902_),
    .Q(\top1.memory1.mem1[26][2] ));
 sg13g2_dfrbp_1 _20890_ (.CLK(\clknet_leaf_182_top1.acquisition_clk ),
    .RESET_B(net315),
    .D(_01078_),
    .Q_N(_08901_),
    .Q(\top1.memory1.mem1[25][0] ));
 sg13g2_dfrbp_1 _20891_ (.CLK(\clknet_leaf_181_top1.acquisition_clk ),
    .RESET_B(net314),
    .D(_01079_),
    .Q_N(_08900_),
    .Q(\top1.memory1.mem1[25][1] ));
 sg13g2_dfrbp_1 _20892_ (.CLK(\clknet_leaf_113_top1.acquisition_clk ),
    .RESET_B(net313),
    .D(_01080_),
    .Q_N(_08899_),
    .Q(\top1.memory1.mem1[25][2] ));
 sg13g2_dfrbp_1 _20893_ (.CLK(\clknet_leaf_40_top1.acquisition_clk ),
    .RESET_B(net7743),
    .D(_01081_),
    .Q_N(_08898_),
    .Q(\top1.mem_ctl.state_reg[0] ));
 sg13g2_dfrbp_1 _20894_ (.CLK(\clknet_leaf_40_top1.acquisition_clk ),
    .RESET_B(net7742),
    .D(_01082_),
    .Q_N(_08897_),
    .Q(\top1.mem_ctl.state_reg[1] ));
 sg13g2_dfrbp_1 _20895_ (.CLK(\clknet_leaf_171_top1.acquisition_clk ),
    .RESET_B(net312),
    .D(_01083_),
    .Q_N(_08896_),
    .Q(\top1.memory1.mem1[105][0] ));
 sg13g2_dfrbp_1 _20896_ (.CLK(\clknet_leaf_172_top1.acquisition_clk ),
    .RESET_B(net311),
    .D(_01084_),
    .Q_N(_08895_),
    .Q(\top1.memory1.mem1[105][1] ));
 sg13g2_dfrbp_1 _20897_ (.CLK(\clknet_leaf_169_top1.acquisition_clk ),
    .RESET_B(net310),
    .D(_01085_),
    .Q_N(_08894_),
    .Q(\top1.memory1.mem1[105][2] ));
 sg13g2_dfrbp_1 _20898_ (.CLK(\clknet_leaf_171_top1.acquisition_clk ),
    .RESET_B(net309),
    .D(_01086_),
    .Q_N(_08893_),
    .Q(\top1.memory1.mem1[106][0] ));
 sg13g2_dfrbp_1 _20899_ (.CLK(\clknet_leaf_171_top1.acquisition_clk ),
    .RESET_B(net308),
    .D(_01087_),
    .Q_N(_08892_),
    .Q(\top1.memory1.mem1[106][1] ));
 sg13g2_dfrbp_1 _20900_ (.CLK(\clknet_leaf_170_top1.acquisition_clk ),
    .RESET_B(net307),
    .D(_01088_),
    .Q_N(_08891_),
    .Q(\top1.memory1.mem1[106][2] ));
 sg13g2_dfrbp_1 _20901_ (.CLK(\clknet_leaf_198_top1.acquisition_clk ),
    .RESET_B(net306),
    .D(_01089_),
    .Q_N(_08890_),
    .Q(\top1.memory1.mem1[111][0] ));
 sg13g2_dfrbp_1 _20902_ (.CLK(\clknet_leaf_194_top1.acquisition_clk ),
    .RESET_B(net305),
    .D(_01090_),
    .Q_N(_08889_),
    .Q(\top1.memory1.mem1[111][1] ));
 sg13g2_dfrbp_1 _20903_ (.CLK(\clknet_leaf_195_top1.acquisition_clk ),
    .RESET_B(net304),
    .D(_01091_),
    .Q_N(_08888_),
    .Q(\top1.memory1.mem1[111][2] ));
 sg13g2_dfrbp_1 _20904_ (.CLK(\clknet_leaf_197_top1.acquisition_clk ),
    .RESET_B(net303),
    .D(_01092_),
    .Q_N(_08887_),
    .Q(\top1.memory1.mem1[110][0] ));
 sg13g2_dfrbp_1 _20905_ (.CLK(\clknet_leaf_195_top1.acquisition_clk ),
    .RESET_B(net302),
    .D(_01093_),
    .Q_N(_08886_),
    .Q(\top1.memory1.mem1[110][1] ));
 sg13g2_dfrbp_1 _20906_ (.CLK(\clknet_leaf_197_top1.acquisition_clk ),
    .RESET_B(net301),
    .D(_01094_),
    .Q_N(_08885_),
    .Q(\top1.memory1.mem1[110][2] ));
 sg13g2_dfrbp_1 _20907_ (.CLK(\clknet_leaf_274_top1.acquisition_clk ),
    .RESET_B(net300),
    .D(_01095_),
    .Q_N(_08884_),
    .Q(\top1.memory1.mem1[10][0] ));
 sg13g2_dfrbp_1 _20908_ (.CLK(\clknet_leaf_273_top1.acquisition_clk ),
    .RESET_B(net299),
    .D(_01096_),
    .Q_N(_08883_),
    .Q(\top1.memory1.mem1[10][1] ));
 sg13g2_dfrbp_1 _20909_ (.CLK(\clknet_leaf_282_top1.acquisition_clk ),
    .RESET_B(net298),
    .D(_01097_),
    .Q_N(_08882_),
    .Q(\top1.memory1.mem1[10][2] ));
 sg13g2_dfrbp_1 _20910_ (.CLK(\clknet_leaf_197_top1.acquisition_clk ),
    .RESET_B(net297),
    .D(_01098_),
    .Q_N(_08881_),
    .Q(\top1.memory1.mem1[108][0] ));
 sg13g2_dfrbp_1 _20911_ (.CLK(\clknet_leaf_195_top1.acquisition_clk ),
    .RESET_B(net296),
    .D(_01099_),
    .Q_N(_08880_),
    .Q(\top1.memory1.mem1[108][1] ));
 sg13g2_dfrbp_1 _20912_ (.CLK(\clknet_leaf_195_top1.acquisition_clk ),
    .RESET_B(net295),
    .D(_01100_),
    .Q_N(_08879_),
    .Q(\top1.memory1.mem1[108][2] ));
 sg13g2_dfrbp_1 _20913_ (.CLK(\clknet_leaf_171_top1.acquisition_clk ),
    .RESET_B(net294),
    .D(_01101_),
    .Q_N(_08878_),
    .Q(\top1.memory1.mem1[107][0] ));
 sg13g2_dfrbp_1 _20914_ (.CLK(\clknet_leaf_171_top1.acquisition_clk ),
    .RESET_B(net293),
    .D(_01102_),
    .Q_N(_08877_),
    .Q(\top1.memory1.mem1[107][1] ));
 sg13g2_dfrbp_1 _20915_ (.CLK(\clknet_leaf_170_top1.acquisition_clk ),
    .RESET_B(net292),
    .D(_01103_),
    .Q_N(_08876_),
    .Q(\top1.memory1.mem1[107][2] ));
 sg13g2_dfrbp_1 _20916_ (.CLK(\clknet_leaf_206_top1.acquisition_clk ),
    .RESET_B(net291),
    .D(_01104_),
    .Q_N(_08875_),
    .Q(\top1.memory1.mem1[112][0] ));
 sg13g2_dfrbp_1 _20917_ (.CLK(\clknet_leaf_217_top1.acquisition_clk ),
    .RESET_B(net290),
    .D(_01105_),
    .Q_N(_08874_),
    .Q(\top1.memory1.mem1[112][1] ));
 sg13g2_dfrbp_1 _20918_ (.CLK(\clknet_leaf_206_top1.acquisition_clk ),
    .RESET_B(net289),
    .D(_01106_),
    .Q_N(_08873_),
    .Q(\top1.memory1.mem1[112][2] ));
 sg13g2_dfrbp_1 _20919_ (.CLK(\clknet_leaf_205_top1.acquisition_clk ),
    .RESET_B(net288),
    .D(_01107_),
    .Q_N(_08872_),
    .Q(\top1.memory1.mem1[113][0] ));
 sg13g2_dfrbp_1 _20920_ (.CLK(\clknet_leaf_217_top1.acquisition_clk ),
    .RESET_B(net287),
    .D(_01108_),
    .Q_N(_08871_),
    .Q(\top1.memory1.mem1[113][1] ));
 sg13g2_dfrbp_1 _20921_ (.CLK(\clknet_leaf_205_top1.acquisition_clk ),
    .RESET_B(net286),
    .D(_01109_),
    .Q_N(_08870_),
    .Q(\top1.memory1.mem1[113][2] ));
 sg13g2_dfrbp_1 _20922_ (.CLK(\clknet_leaf_171_top1.acquisition_clk ),
    .RESET_B(net285),
    .D(_01110_),
    .Q_N(_08869_),
    .Q(\top1.memory1.mem1[104][0] ));
 sg13g2_dfrbp_1 _20923_ (.CLK(\clknet_leaf_171_top1.acquisition_clk ),
    .RESET_B(net284),
    .D(_01111_),
    .Q_N(_08868_),
    .Q(\top1.memory1.mem1[104][1] ));
 sg13g2_dfrbp_1 _20924_ (.CLK(\clknet_leaf_170_top1.acquisition_clk ),
    .RESET_B(net283),
    .D(_01112_),
    .Q_N(_08867_),
    .Q(\top1.memory1.mem1[104][2] ));
 sg13g2_dfrbp_1 _20925_ (.CLK(\clknet_leaf_198_top1.acquisition_clk ),
    .RESET_B(net282),
    .D(_01113_),
    .Q_N(_08866_),
    .Q(\top1.memory1.mem1[103][0] ));
 sg13g2_dfrbp_1 _20926_ (.CLK(\clknet_leaf_195_top1.acquisition_clk ),
    .RESET_B(net281),
    .D(_01114_),
    .Q_N(_08865_),
    .Q(\top1.memory1.mem1[103][1] ));
 sg13g2_dfrbp_1 _20927_ (.CLK(\clknet_leaf_192_top1.acquisition_clk ),
    .RESET_B(net280),
    .D(_01115_),
    .Q_N(_08864_),
    .Q(\top1.memory1.mem1[103][2] ));
 sg13g2_dfrbp_1 _20928_ (.CLK(\clknet_leaf_218_top1.acquisition_clk ),
    .RESET_B(net279),
    .D(_01116_),
    .Q_N(_08863_),
    .Q(\top1.memory1.mem1[122][0] ));
 sg13g2_dfrbp_1 _20929_ (.CLK(\clknet_leaf_221_top1.acquisition_clk ),
    .RESET_B(net278),
    .D(_01117_),
    .Q_N(_08862_),
    .Q(\top1.memory1.mem1[122][1] ));
 sg13g2_dfrbp_1 _20930_ (.CLK(\clknet_leaf_220_top1.acquisition_clk ),
    .RESET_B(net277),
    .D(_01118_),
    .Q_N(_08861_),
    .Q(\top1.memory1.mem1[122][2] ));
 sg13g2_dfrbp_1 _20931_ (.CLK(\clknet_leaf_214_top1.acquisition_clk ),
    .RESET_B(net276),
    .D(_01119_),
    .Q_N(_08860_),
    .Q(\top1.memory1.mem1[121][0] ));
 sg13g2_dfrbp_1 _20932_ (.CLK(\clknet_leaf_221_top1.acquisition_clk ),
    .RESET_B(net275),
    .D(_01120_),
    .Q_N(_08859_),
    .Q(\top1.memory1.mem1[121][1] ));
 sg13g2_dfrbp_1 _20933_ (.CLK(\clknet_leaf_220_top1.acquisition_clk ),
    .RESET_B(net274),
    .D(_01121_),
    .Q_N(_08858_),
    .Q(\top1.memory1.mem1[121][2] ));
 sg13g2_dfrbp_1 _20934_ (.CLK(\clknet_leaf_215_top1.acquisition_clk ),
    .RESET_B(net273),
    .D(_01122_),
    .Q_N(_08857_),
    .Q(\top1.memory1.mem1[120][0] ));
 sg13g2_dfrbp_1 _20935_ (.CLK(\clknet_leaf_221_top1.acquisition_clk ),
    .RESET_B(net272),
    .D(_01123_),
    .Q_N(_08856_),
    .Q(\top1.memory1.mem1[120][1] ));
 sg13g2_dfrbp_1 _20936_ (.CLK(\clknet_leaf_220_top1.acquisition_clk ),
    .RESET_B(net271),
    .D(_01124_),
    .Q_N(_08855_),
    .Q(\top1.memory1.mem1[120][2] ));
 sg13g2_dfrbp_1 _20937_ (.CLK(\clknet_leaf_265_top1.acquisition_clk ),
    .RESET_B(net270),
    .D(_01125_),
    .Q_N(_08854_),
    .Q(\top1.memory1.mem1[11][0] ));
 sg13g2_dfrbp_1 _20938_ (.CLK(\clknet_leaf_265_top1.acquisition_clk ),
    .RESET_B(net269),
    .D(_01126_),
    .Q_N(_08853_),
    .Q(\top1.memory1.mem1[11][1] ));
 sg13g2_dfrbp_1 _20939_ (.CLK(\clknet_leaf_276_top1.acquisition_clk ),
    .RESET_B(net268),
    .D(_01127_),
    .Q_N(_08852_),
    .Q(\top1.memory1.mem1[11][2] ));
 sg13g2_dfrbp_1 _20940_ (.CLK(\clknet_leaf_206_top1.acquisition_clk ),
    .RESET_B(net267),
    .D(_01128_),
    .Q_N(_08851_),
    .Q(\top1.memory1.mem1[114][0] ));
 sg13g2_dfrbp_1 _20941_ (.CLK(\clknet_leaf_216_top1.acquisition_clk ),
    .RESET_B(net266),
    .D(_01129_),
    .Q_N(_08850_),
    .Q(\top1.memory1.mem1[114][1] ));
 sg13g2_dfrbp_1 _20942_ (.CLK(\clknet_leaf_205_top1.acquisition_clk ),
    .RESET_B(net265),
    .D(_01130_),
    .Q_N(_08849_),
    .Q(\top1.memory1.mem1[114][2] ));
 sg13g2_dfrbp_1 _20943_ (.CLK(\clknet_leaf_240_top1.acquisition_clk ),
    .RESET_B(net264),
    .D(_01131_),
    .Q_N(_08848_),
    .Q(\top1.memory1.mem1[165][0] ));
 sg13g2_dfrbp_1 _20944_ (.CLK(\clknet_leaf_238_top1.acquisition_clk ),
    .RESET_B(net263),
    .D(_01132_),
    .Q_N(_08847_),
    .Q(\top1.memory1.mem1[165][1] ));
 sg13g2_dfrbp_1 _20945_ (.CLK(\clknet_leaf_255_top1.acquisition_clk ),
    .RESET_B(net262),
    .D(_01133_),
    .Q_N(_08846_),
    .Q(\top1.memory1.mem1[165][2] ));
 sg13g2_dfrbp_1 _20946_ (.CLK(\clknet_leaf_274_top1.acquisition_clk ),
    .RESET_B(net261),
    .D(_01134_),
    .Q_N(_08845_),
    .Q(\top1.memory1.mem1[162][0] ));
 sg13g2_dfrbp_1 _20947_ (.CLK(\clknet_leaf_279_top1.acquisition_clk ),
    .RESET_B(net260),
    .D(_01135_),
    .Q_N(_08844_),
    .Q(\top1.memory1.mem1[162][1] ));
 sg13g2_dfrbp_1 _20948_ (.CLK(\clknet_leaf_264_top1.acquisition_clk ),
    .RESET_B(net259),
    .D(_01136_),
    .Q_N(_08843_),
    .Q(\top1.memory1.mem1[162][2] ));
 sg13g2_dfrbp_1 _20949_ (.CLK(\clknet_leaf_274_top1.acquisition_clk ),
    .RESET_B(net258),
    .D(_01137_),
    .Q_N(_08842_),
    .Q(\top1.memory1.mem1[161][0] ));
 sg13g2_dfrbp_1 _20950_ (.CLK(\clknet_leaf_279_top1.acquisition_clk ),
    .RESET_B(net257),
    .D(_01138_),
    .Q_N(_08841_),
    .Q(\top1.memory1.mem1[161][1] ));
 sg13g2_dfrbp_1 _20951_ (.CLK(\clknet_leaf_274_top1.acquisition_clk ),
    .RESET_B(net256),
    .D(_01139_),
    .Q_N(_08840_),
    .Q(\top1.memory1.mem1[161][2] ));
 sg13g2_dfrbp_1 _20952_ (.CLK(net6742),
    .RESET_B(net7750),
    .D(_01140_),
    .Q_N(_09919_),
    .Q(\top1.fsm.sending_data ));
 sg13g2_dfrbp_1 _20953_ (.CLK(net7559),
    .RESET_B(net7746),
    .D(\top1.fsm.idx_final[0] ),
    .Q_N(_09920_),
    .Q(\top1.fsm.reg_idx_final[0] ));
 sg13g2_dfrbp_1 _20954_ (.CLK(net7560),
    .RESET_B(net7746),
    .D(\top1.fsm.idx_final[1] ),
    .Q_N(_09921_),
    .Q(\top1.fsm.reg_idx_final[1] ));
 sg13g2_dfrbp_1 _20955_ (.CLK(net7560),
    .RESET_B(net7745),
    .D(\top1.fsm.idx_final[2] ),
    .Q_N(_09922_),
    .Q(\top1.fsm.reg_idx_final[2] ));
 sg13g2_dfrbp_1 _20956_ (.CLK(net7559),
    .RESET_B(net7746),
    .D(\top1.fsm.idx_final[3] ),
    .Q_N(_09923_),
    .Q(\top1.fsm.reg_idx_final[3] ));
 sg13g2_dfrbp_1 _20957_ (.CLK(net7559),
    .RESET_B(net7745),
    .D(\top1.fsm.idx_final[4] ),
    .Q_N(_09924_),
    .Q(\top1.fsm.reg_idx_final[4] ));
 sg13g2_dfrbp_1 _20958_ (.CLK(net7559),
    .RESET_B(net7745),
    .D(\top1.fsm.idx_final[5] ),
    .Q_N(_09925_),
    .Q(\top1.fsm.reg_idx_final[5] ));
 sg13g2_dfrbp_1 _20959_ (.CLK(net7559),
    .RESET_B(net7745),
    .D(\top1.fsm.idx_final[6] ),
    .Q_N(_09926_),
    .Q(\top1.fsm.reg_idx_final[6] ));
 sg13g2_dfrbp_1 _20960_ (.CLK(net7559),
    .RESET_B(net7745),
    .D(\top1.fsm.idx_final[7] ),
    .Q_N(_08839_),
    .Q(\top1.fsm.reg_idx_final[7] ));
 sg13g2_dfrbp_1 _20961_ (.CLK(net6743),
    .RESET_B(net7741),
    .D(_01141_),
    .Q_N(_00065_),
    .Q(\top1.fsm.sending_pending ));
 sg13g2_dfrbp_1 _20962_ (.CLK(\clknet_leaf_274_top1.acquisition_clk ),
    .RESET_B(net255),
    .D(_01142_),
    .Q_N(_08838_),
    .Q(\top1.memory1.mem1[160][0] ));
 sg13g2_dfrbp_1 _20963_ (.CLK(\clknet_leaf_279_top1.acquisition_clk ),
    .RESET_B(net254),
    .D(_01143_),
    .Q_N(_08837_),
    .Q(\top1.memory1.mem1[160][1] ));
 sg13g2_dfrbp_1 _20964_ (.CLK(\clknet_leaf_275_top1.acquisition_clk ),
    .RESET_B(net253),
    .D(_01144_),
    .Q_N(_08836_),
    .Q(\top1.memory1.mem1[160][2] ));
 sg13g2_dfrbp_1 _20965_ (.CLK(net6739),
    .RESET_B(net7741),
    .D(_01145_),
    .Q_N(_08835_),
    .Q(\top1.fsm.signal_duration ));
 sg13g2_dfrbp_1 _20966_ (.CLK(net6739),
    .RESET_B(net7741),
    .D(_01146_),
    .Q_N(_00066_),
    .Q(\top1.fsm.re ));
 sg13g2_dfrbp_1 _20967_ (.CLK(\clknet_leaf_147_top1.acquisition_clk ),
    .RESET_B(net252),
    .D(_01147_),
    .Q_N(_08834_),
    .Q(\top1.memory1.mem1[37][0] ));
 sg13g2_dfrbp_1 _20968_ (.CLK(\clknet_leaf_148_top1.acquisition_clk ),
    .RESET_B(net251),
    .D(_01148_),
    .Q_N(_08833_),
    .Q(\top1.memory1.mem1[37][1] ));
 sg13g2_dfrbp_1 _20969_ (.CLK(\clknet_leaf_151_top1.acquisition_clk ),
    .RESET_B(net250),
    .D(_01149_),
    .Q_N(_08832_),
    .Q(\top1.memory1.mem1[37][2] ));
 sg13g2_dfrbp_1 _20970_ (.CLK(\clknet_leaf_240_top1.acquisition_clk ),
    .RESET_B(net249),
    .D(_01150_),
    .Q_N(_08831_),
    .Q(\top1.memory1.mem1[164][0] ));
 sg13g2_dfrbp_1 _20971_ (.CLK(\clknet_leaf_239_top1.acquisition_clk ),
    .RESET_B(net248),
    .D(_01151_),
    .Q_N(_08830_),
    .Q(\top1.memory1.mem1[164][1] ));
 sg13g2_dfrbp_1 _20972_ (.CLK(\clknet_leaf_255_top1.acquisition_clk ),
    .RESET_B(net1063),
    .D(_01152_),
    .Q_N(_09927_),
    .Q(\top1.memory1.mem1[164][2] ));
 sg13g2_dfrbp_1 _20973_ (.CLK(net6739),
    .RESET_B(net7734),
    .D(_00001_),
    .Q_N(_09928_),
    .Q(\top1.fsm.cpt[0] ));
 sg13g2_dfrbp_1 _20974_ (.CLK(net6739),
    .RESET_B(net7734),
    .D(_00002_),
    .Q_N(_09929_),
    .Q(\top1.fsm.cpt[1] ));
 sg13g2_dfrbp_1 _20975_ (.CLK(net6739),
    .RESET_B(net7734),
    .D(_00003_),
    .Q_N(_09930_),
    .Q(\top1.fsm.cpt[2] ));
 sg13g2_dfrbp_1 _20976_ (.CLK(net6739),
    .RESET_B(net7734),
    .D(_00004_),
    .Q_N(_09931_),
    .Q(\top1.fsm.cpt[3] ));
 sg13g2_dfrbp_1 _20977_ (.CLK(net6739),
    .RESET_B(net7734),
    .D(_00005_),
    .Q_N(_00064_),
    .Q(\top1.fsm.cpt[4] ));
 sg13g2_dfrbp_1 _20978_ (.CLK(\clknet_leaf_48_top1.acquisition_clk ),
    .RESET_B(net247),
    .D(_01153_),
    .Q_N(_08829_),
    .Q(\top1.memory1.mem1[132][0] ));
 sg13g2_dfrbp_1 _20979_ (.CLK(\clknet_leaf_56_top1.acquisition_clk ),
    .RESET_B(net246),
    .D(_01154_),
    .Q_N(_08828_),
    .Q(\top1.memory1.mem1[132][1] ));
 sg13g2_dfrbp_1 _20980_ (.CLK(\clknet_leaf_22_top1.acquisition_clk ),
    .RESET_B(net245),
    .D(_01155_),
    .Q_N(_08827_),
    .Q(\top1.memory1.mem1[132][2] ));
 sg13g2_dfrbp_1 _20981_ (.CLK(net6745),
    .RESET_B(net7747),
    .D(_01156_),
    .Q_N(_08826_),
    .Q(\top1.addr_out[0] ));
 sg13g2_dfrbp_1 _20982_ (.CLK(net6745),
    .RESET_B(net7749),
    .D(_01157_),
    .Q_N(_08825_),
    .Q(\top1.addr_out[1] ));
 sg13g2_dfrbp_1 _20983_ (.CLK(net6745),
    .RESET_B(net7747),
    .D(_01158_),
    .Q_N(_00073_),
    .Q(\top1.addr_out[2] ));
 sg13g2_dfrbp_1 _20984_ (.CLK(net6745),
    .RESET_B(net7747),
    .D(_01159_),
    .Q_N(_00072_),
    .Q(\top1.addr_out[3] ));
 sg13g2_dfrbp_1 _20985_ (.CLK(net6746),
    .RESET_B(net7743),
    .D(_01160_),
    .Q_N(_00071_),
    .Q(\top1.addr_out[4] ));
 sg13g2_dfrbp_1 _20986_ (.CLK(net6746),
    .RESET_B(net7743),
    .D(_01161_),
    .Q_N(_00070_),
    .Q(\top1.addr_out[5] ));
 sg13g2_dfrbp_1 _20987_ (.CLK(net6745),
    .RESET_B(net7746),
    .D(_01162_),
    .Q_N(_00069_),
    .Q(\top1.addr_out[6] ));
 sg13g2_dfrbp_1 _20988_ (.CLK(net6745),
    .RESET_B(net7746),
    .D(_01163_),
    .Q_N(_00068_),
    .Q(\top1.addr_out[7] ));
 sg13g2_dfrbp_1 _20989_ (.CLK(net6742),
    .RESET_B(net7741),
    .D(\top1.fsm.state_next[0] ),
    .Q_N(_09932_),
    .Q(\top1.fsm.state_reg[0] ));
 sg13g2_dfrbp_1 _20990_ (.CLK(net6742),
    .RESET_B(net7750),
    .D(\top1.fsm.state_next[1] ),
    .Q_N(_00067_),
    .Q(\top1.fsm.state_reg[1] ));
 sg13g2_dfrbp_1 _20991_ (.CLK(net6742),
    .RESET_B(net7741),
    .D(\top1.fsm.state_next[2] ),
    .Q_N(_00063_),
    .Q(\top1.fsm.state_reg[2] ));
 sg13g2_dfrbp_1 _20992_ (.CLK(\clknet_leaf_265_top1.acquisition_clk ),
    .RESET_B(net244),
    .D(_01164_),
    .Q_N(_08824_),
    .Q(\top1.memory1.mem1[163][0] ));
 sg13g2_dfrbp_1 _20993_ (.CLK(\clknet_leaf_279_top1.acquisition_clk ),
    .RESET_B(net243),
    .D(_01165_),
    .Q_N(_08823_),
    .Q(\top1.memory1.mem1[163][1] ));
 sg13g2_dfrbp_1 _20994_ (.CLK(\clknet_leaf_265_top1.acquisition_clk ),
    .RESET_B(net242),
    .D(_01166_),
    .Q_N(_08822_),
    .Q(\top1.memory1.mem1[163][2] ));
 sg13g2_dfrbp_1 _20995_ (.CLK(\clknet_leaf_208_top1.acquisition_clk ),
    .RESET_B(net241),
    .D(_01167_),
    .Q_N(_08821_),
    .Q(\top1.memory1.mem1[124][0] ));
 sg13g2_dfrbp_1 _20996_ (.CLK(\clknet_leaf_215_top1.acquisition_clk ),
    .RESET_B(net240),
    .D(_01168_),
    .Q_N(_08820_),
    .Q(\top1.memory1.mem1[124][1] ));
 sg13g2_dfrbp_1 _20997_ (.CLK(\clknet_leaf_204_top1.acquisition_clk ),
    .RESET_B(net239),
    .D(_01169_),
    .Q_N(_08819_),
    .Q(\top1.memory1.mem1[124][2] ));
 sg13g2_dfrbp_1 _20998_ (.CLK(\clknet_leaf_145_top1.acquisition_clk ),
    .RESET_B(net238),
    .D(_01170_),
    .Q_N(_08818_),
    .Q(\top1.memory1.mem1[32][0] ));
 sg13g2_dfrbp_1 _20999_ (.CLK(\clknet_leaf_148_top1.acquisition_clk ),
    .RESET_B(net237),
    .D(_01171_),
    .Q_N(_08817_),
    .Q(\top1.memory1.mem1[32][1] ));
 sg13g2_dfrbp_1 _21000_ (.CLK(\clknet_leaf_149_top1.acquisition_clk ),
    .RESET_B(net236),
    .D(_01172_),
    .Q_N(_08816_),
    .Q(\top1.memory1.mem1[32][2] ));
 sg13g2_dfrbp_1 _21001_ (.CLK(\clknet_leaf_214_top1.acquisition_clk ),
    .RESET_B(net235),
    .D(_01173_),
    .Q_N(_08815_),
    .Q(\top1.memory1.mem1[123][0] ));
 sg13g2_dfrbp_1 _21002_ (.CLK(\clknet_leaf_221_top1.acquisition_clk ),
    .RESET_B(net234),
    .D(_01174_),
    .Q_N(_08814_),
    .Q(\top1.memory1.mem1[123][1] ));
 sg13g2_dfrbp_1 _21003_ (.CLK(\clknet_leaf_220_top1.acquisition_clk ),
    .RESET_B(net233),
    .D(_01175_),
    .Q_N(_08813_),
    .Q(\top1.memory1.mem1[123][2] ));
 sg13g2_dfrbp_1 _21004_ (.CLK(\clknet_leaf_278_top1.acquisition_clk ),
    .RESET_B(net232),
    .D(_01176_),
    .Q_N(_08812_),
    .Q(\top1.memory1.mem1[15][0] ));
 sg13g2_dfrbp_1 _21005_ (.CLK(\clknet_leaf_272_top1.acquisition_clk ),
    .RESET_B(net231),
    .D(_01177_),
    .Q_N(_08811_),
    .Q(\top1.memory1.mem1[15][1] ));
 sg13g2_dfrbp_1 _21006_ (.CLK(\clknet_leaf_277_top1.acquisition_clk ),
    .RESET_B(net230),
    .D(_01178_),
    .Q_N(_08810_),
    .Q(\top1.memory1.mem1[15][2] ));
 sg13g2_dfrbp_1 _21007_ (.CLK(\clknet_leaf_75_top1.acquisition_clk ),
    .RESET_B(net229),
    .D(_01179_),
    .Q_N(_08809_),
    .Q(\top1.memory1.mem1[158][0] ));
 sg13g2_dfrbp_1 _21008_ (.CLK(\clknet_leaf_73_top1.acquisition_clk ),
    .RESET_B(net228),
    .D(_01180_),
    .Q_N(_08808_),
    .Q(\top1.memory1.mem1[158][1] ));
 sg13g2_dfrbp_1 _21009_ (.CLK(\clknet_leaf_59_top1.acquisition_clk ),
    .RESET_B(net227),
    .D(_01181_),
    .Q_N(_08807_),
    .Q(\top1.memory1.mem1[158][2] ));
 sg13g2_dfrbp_1 _21010_ (.CLK(\clknet_leaf_215_top1.acquisition_clk ),
    .RESET_B(net226),
    .D(_01182_),
    .Q_N(_08806_),
    .Q(\top1.memory1.mem1[118][0] ));
 sg13g2_dfrbp_1 _21011_ (.CLK(\clknet_leaf_217_top1.acquisition_clk ),
    .RESET_B(net225),
    .D(_01183_),
    .Q_N(_08805_),
    .Q(\top1.memory1.mem1[118][1] ));
 sg13g2_dfrbp_1 _21012_ (.CLK(\clknet_leaf_219_top1.acquisition_clk ),
    .RESET_B(net224),
    .D(_01184_),
    .Q_N(_08804_),
    .Q(\top1.memory1.mem1[118][2] ));
 sg13g2_dfrbp_1 _21013_ (.CLK(\clknet_leaf_214_top1.acquisition_clk ),
    .RESET_B(net223),
    .D(_01185_),
    .Q_N(_08803_),
    .Q(\top1.memory1.mem1[117][0] ));
 sg13g2_dfrbp_1 _21014_ (.CLK(\clknet_leaf_217_top1.acquisition_clk ),
    .RESET_B(net222),
    .D(_01186_),
    .Q_N(_08802_),
    .Q(\top1.memory1.mem1[117][1] ));
 sg13g2_dfrbp_1 _21015_ (.CLK(\clknet_leaf_219_top1.acquisition_clk ),
    .RESET_B(net221),
    .D(_01187_),
    .Q_N(_08801_),
    .Q(\top1.memory1.mem1[117][2] ));
 sg13g2_dfrbp_1 _21016_ (.CLK(\clknet_leaf_214_top1.acquisition_clk ),
    .RESET_B(net220),
    .D(_01188_),
    .Q_N(_08800_),
    .Q(\top1.memory1.mem1[116][0] ));
 sg13g2_dfrbp_1 _21017_ (.CLK(\clknet_leaf_217_top1.acquisition_clk ),
    .RESET_B(net219),
    .D(_01189_),
    .Q_N(_08799_),
    .Q(\top1.memory1.mem1[116][1] ));
 sg13g2_dfrbp_1 _21018_ (.CLK(\clknet_leaf_219_top1.acquisition_clk ),
    .RESET_B(net218),
    .D(_01190_),
    .Q_N(_08798_),
    .Q(\top1.memory1.mem1[116][2] ));
 sg13g2_dfrbp_1 _21019_ (.CLK(\clknet_leaf_74_top1.acquisition_clk ),
    .RESET_B(net217),
    .D(_01191_),
    .Q_N(_08797_),
    .Q(\top1.memory1.mem1[157][0] ));
 sg13g2_dfrbp_1 _21020_ (.CLK(\clknet_leaf_74_top1.acquisition_clk ),
    .RESET_B(net216),
    .D(_01192_),
    .Q_N(_08796_),
    .Q(\top1.memory1.mem1[157][1] ));
 sg13g2_dfrbp_1 _21021_ (.CLK(\clknet_leaf_59_top1.acquisition_clk ),
    .RESET_B(net215),
    .D(_01193_),
    .Q_N(_08795_),
    .Q(\top1.memory1.mem1[157][2] ));
 sg13g2_dfrbp_1 _21022_ (.CLK(\clknet_leaf_207_top1.acquisition_clk ),
    .RESET_B(net214),
    .D(_01194_),
    .Q_N(_08794_),
    .Q(\top1.memory1.mem1[115][0] ));
 sg13g2_dfrbp_1 _21023_ (.CLK(\clknet_leaf_216_top1.acquisition_clk ),
    .RESET_B(net213),
    .D(_01195_),
    .Q_N(_08793_),
    .Q(\top1.memory1.mem1[115][1] ));
 sg13g2_dfrbp_1 _21024_ (.CLK(\clknet_leaf_206_top1.acquisition_clk ),
    .RESET_B(net212),
    .D(_01196_),
    .Q_N(_08792_),
    .Q(\top1.memory1.mem1[115][2] ));
 sg13g2_dfrbp_1 _21025_ (.CLK(\clknet_leaf_69_top1.acquisition_clk ),
    .RESET_B(net211),
    .D(_01197_),
    .Q_N(_08791_),
    .Q(\top1.memory1.mem1[156][0] ));
 sg13g2_dfrbp_1 _21026_ (.CLK(\clknet_leaf_73_top1.acquisition_clk ),
    .RESET_B(net210),
    .D(_01198_),
    .Q_N(_08790_),
    .Q(\top1.memory1.mem1[156][1] ));
 sg13g2_dfrbp_1 _21027_ (.CLK(\clknet_leaf_74_top1.acquisition_clk ),
    .RESET_B(net209),
    .D(_01199_),
    .Q_N(_08789_),
    .Q(\top1.memory1.mem1[156][2] ));
 sg13g2_dfrbp_1 _21028_ (.CLK(\clknet_leaf_49_top1.acquisition_clk ),
    .RESET_B(net208),
    .D(_01200_),
    .Q_N(_08788_),
    .Q(\top1.memory1.mem1[155][0] ));
 sg13g2_dfrbp_1 _21029_ (.CLK(\clknet_leaf_45_top1.acquisition_clk ),
    .RESET_B(net207),
    .D(_01201_),
    .Q_N(_08787_),
    .Q(\top1.memory1.mem1[155][1] ));
 sg13g2_dfrbp_1 _21030_ (.CLK(\clknet_leaf_46_top1.acquisition_clk ),
    .RESET_B(net206),
    .D(_01202_),
    .Q_N(_08786_),
    .Q(\top1.memory1.mem1[155][2] ));
 sg13g2_dfrbp_1 _21031_ (.CLK(\clknet_leaf_48_top1.acquisition_clk ),
    .RESET_B(net205),
    .D(_01203_),
    .Q_N(_08785_),
    .Q(\top1.memory1.mem1[154][0] ));
 sg13g2_dfrbp_1 _21032_ (.CLK(\clknet_leaf_48_top1.acquisition_clk ),
    .RESET_B(net204),
    .D(_01204_),
    .Q_N(_08784_),
    .Q(\top1.memory1.mem1[154][1] ));
 sg13g2_dfrbp_1 _21033_ (.CLK(\clknet_leaf_48_top1.acquisition_clk ),
    .RESET_B(net203),
    .D(_01205_),
    .Q_N(_08783_),
    .Q(\top1.memory1.mem1[154][2] ));
 sg13g2_dfrbp_1 _21034_ (.CLK(\clknet_leaf_49_top1.acquisition_clk ),
    .RESET_B(net202),
    .D(_01206_),
    .Q_N(_08782_),
    .Q(\top1.memory1.mem1[153][0] ));
 sg13g2_dfrbp_1 _21035_ (.CLK(\clknet_leaf_45_top1.acquisition_clk ),
    .RESET_B(net201),
    .D(_01207_),
    .Q_N(_08781_),
    .Q(\top1.memory1.mem1[153][1] ));
 sg13g2_dfrbp_1 _21036_ (.CLK(\clknet_leaf_47_top1.acquisition_clk ),
    .RESET_B(net200),
    .D(_01208_),
    .Q_N(_08780_),
    .Q(\top1.memory1.mem1[153][2] ));
 sg13g2_dfrbp_1 _21037_ (.CLK(\clknet_leaf_48_top1.acquisition_clk ),
    .RESET_B(net199),
    .D(_01209_),
    .Q_N(_08779_),
    .Q(\top1.memory1.mem1[152][0] ));
 sg13g2_dfrbp_1 _21038_ (.CLK(\clknet_leaf_47_top1.acquisition_clk ),
    .RESET_B(net198),
    .D(_01210_),
    .Q_N(_08778_),
    .Q(\top1.memory1.mem1[152][1] ));
 sg13g2_dfrbp_1 _21039_ (.CLK(\clknet_leaf_47_top1.acquisition_clk ),
    .RESET_B(net197),
    .D(_01211_),
    .Q_N(_08777_),
    .Q(\top1.memory1.mem1[152][2] ));
 sg13g2_dfrbp_1 _21040_ (.CLK(\clknet_leaf_23_top1.acquisition_clk ),
    .RESET_B(net196),
    .D(_01212_),
    .Q_N(_08776_),
    .Q(\top1.memory1.mem1[151][0] ));
 sg13g2_dfrbp_1 _21041_ (.CLK(\clknet_leaf_23_top1.acquisition_clk ),
    .RESET_B(net195),
    .D(_01213_),
    .Q_N(_08775_),
    .Q(\top1.memory1.mem1[151][1] ));
 sg13g2_dfrbp_1 _21042_ (.CLK(\clknet_leaf_24_top1.acquisition_clk ),
    .RESET_B(net194),
    .D(_01214_),
    .Q_N(_08774_),
    .Q(\top1.memory1.mem1[151][2] ));
 sg13g2_dfrbp_1 _21043_ (.CLK(\clknet_leaf_24_top1.acquisition_clk ),
    .RESET_B(net193),
    .D(_01215_),
    .Q_N(_08773_),
    .Q(\top1.memory1.mem1[150][0] ));
 sg13g2_dfrbp_1 _21044_ (.CLK(\clknet_leaf_47_top1.acquisition_clk ),
    .RESET_B(net192),
    .D(_01216_),
    .Q_N(_08772_),
    .Q(\top1.memory1.mem1[150][1] ));
 sg13g2_dfrbp_1 _21045_ (.CLK(\clknet_leaf_24_top1.acquisition_clk ),
    .RESET_B(net191),
    .D(_01217_),
    .Q_N(_08771_),
    .Q(\top1.memory1.mem1[150][2] ));
 sg13g2_dfrbp_1 _21046_ (.CLK(\clknet_leaf_257_top1.acquisition_clk ),
    .RESET_B(net190),
    .D(_01218_),
    .Q_N(_08770_),
    .Q(\top1.memory1.mem1[30][0] ));
 sg13g2_dfrbp_1 _21047_ (.CLK(\clknet_leaf_256_top1.acquisition_clk ),
    .RESET_B(net189),
    .D(_01219_),
    .Q_N(_08769_),
    .Q(\top1.memory1.mem1[30][1] ));
 sg13g2_dfrbp_1 _21048_ (.CLK(\clknet_leaf_259_top1.acquisition_clk ),
    .RESET_B(net188),
    .D(_01220_),
    .Q_N(_08768_),
    .Q(\top1.memory1.mem1[30][2] ));
 sg13g2_dfrbp_1 _21049_ (.CLK(\clknet_leaf_275_top1.acquisition_clk ),
    .RESET_B(net187),
    .D(_01221_),
    .Q_N(_08767_),
    .Q(\top1.memory1.mem1[14][0] ));
 sg13g2_dfrbp_1 _21050_ (.CLK(\clknet_leaf_272_top1.acquisition_clk ),
    .RESET_B(net186),
    .D(_01222_),
    .Q_N(_08766_),
    .Q(\top1.memory1.mem1[14][1] ));
 sg13g2_dfrbp_1 _21051_ (.CLK(\clknet_leaf_276_top1.acquisition_clk ),
    .RESET_B(net185),
    .D(_01223_),
    .Q_N(_08765_),
    .Q(\top1.memory1.mem1[14][2] ));
 sg13g2_dfrbp_1 _21052_ (.CLK(\clknet_leaf_23_top1.acquisition_clk ),
    .RESET_B(net184),
    .D(_01224_),
    .Q_N(_08764_),
    .Q(\top1.memory1.mem1[148][0] ));
 sg13g2_dfrbp_1 _21053_ (.CLK(\clknet_leaf_23_top1.acquisition_clk ),
    .RESET_B(net183),
    .D(_01225_),
    .Q_N(_08763_),
    .Q(\top1.memory1.mem1[148][1] ));
 sg13g2_dfrbp_1 _21054_ (.CLK(\clknet_leaf_25_top1.acquisition_clk ),
    .RESET_B(net182),
    .D(_01226_),
    .Q_N(_08762_),
    .Q(\top1.memory1.mem1[148][2] ));
 sg13g2_dfrbp_1 _21055_ (.CLK(\clknet_leaf_44_top1.acquisition_clk ),
    .RESET_B(net181),
    .D(_01227_),
    .Q_N(_08761_),
    .Q(\top1.memory1.mem1[147][0] ));
 sg13g2_dfrbp_1 _21056_ (.CLK(\clknet_leaf_58_top1.acquisition_clk ),
    .RESET_B(net180),
    .D(_01228_),
    .Q_N(_08760_),
    .Q(\top1.memory1.mem1[147][1] ));
 sg13g2_dfrbp_1 _21057_ (.CLK(\clknet_leaf_46_top1.acquisition_clk ),
    .RESET_B(net179),
    .D(_01229_),
    .Q_N(_08759_),
    .Q(\top1.memory1.mem1[147][2] ));
 sg13g2_dfrbp_1 _21058_ (.CLK(\clknet_leaf_44_top1.acquisition_clk ),
    .RESET_B(net178),
    .D(_01230_),
    .Q_N(_08758_),
    .Q(\top1.memory1.mem1[146][0] ));
 sg13g2_dfrbp_1 _21059_ (.CLK(\clknet_leaf_58_top1.acquisition_clk ),
    .RESET_B(net177),
    .D(_01231_),
    .Q_N(_08757_),
    .Q(\top1.memory1.mem1[146][1] ));
 sg13g2_dfrbp_1 _21060_ (.CLK(\clknet_leaf_46_top1.acquisition_clk ),
    .RESET_B(net176),
    .D(_01232_),
    .Q_N(_08756_),
    .Q(\top1.memory1.mem1[146][2] ));
 sg13g2_dfrbp_1 _21061_ (.CLK(\clknet_leaf_44_top1.acquisition_clk ),
    .RESET_B(net175),
    .D(_01233_),
    .Q_N(_08755_),
    .Q(\top1.memory1.mem1[145][0] ));
 sg13g2_dfrbp_1 _21062_ (.CLK(\clknet_leaf_58_top1.acquisition_clk ),
    .RESET_B(net174),
    .D(_01234_),
    .Q_N(_08754_),
    .Q(\top1.memory1.mem1[145][1] ));
 sg13g2_dfrbp_1 _21063_ (.CLK(\clknet_leaf_46_top1.acquisition_clk ),
    .RESET_B(net173),
    .D(_01235_),
    .Q_N(_08753_),
    .Q(\top1.memory1.mem1[145][2] ));
 sg13g2_dfrbp_1 _21064_ (.CLK(\clknet_leaf_57_top1.acquisition_clk ),
    .RESET_B(net172),
    .D(_01236_),
    .Q_N(_08752_),
    .Q(\top1.memory1.mem1[144][0] ));
 sg13g2_dfrbp_1 _21065_ (.CLK(\clknet_leaf_58_top1.acquisition_clk ),
    .RESET_B(net171),
    .D(_01237_),
    .Q_N(_08751_),
    .Q(\top1.memory1.mem1[144][1] ));
 sg13g2_dfrbp_1 _21066_ (.CLK(\clknet_leaf_45_top1.acquisition_clk ),
    .RESET_B(net170),
    .D(_01238_),
    .Q_N(_08750_),
    .Q(\top1.memory1.mem1[144][2] ));
 sg13g2_dfrbp_1 _21067_ (.CLK(\clknet_leaf_52_top1.acquisition_clk ),
    .RESET_B(net169),
    .D(_01239_),
    .Q_N(_08749_),
    .Q(\top1.memory1.mem1[143][0] ));
 sg13g2_dfrbp_1 _21068_ (.CLK(\clknet_leaf_51_top1.acquisition_clk ),
    .RESET_B(net168),
    .D(_01240_),
    .Q_N(_08748_),
    .Q(\top1.memory1.mem1[143][1] ));
 sg13g2_dfrbp_1 _21069_ (.CLK(\clknet_leaf_51_top1.acquisition_clk ),
    .RESET_B(net167),
    .D(_01241_),
    .Q_N(_08747_),
    .Q(\top1.memory1.mem1[143][2] ));
 sg13g2_dfrbp_1 _21070_ (.CLK(\clknet_leaf_52_top1.acquisition_clk ),
    .RESET_B(net166),
    .D(_01242_),
    .Q_N(_08746_),
    .Q(\top1.memory1.mem1[142][0] ));
 sg13g2_dfrbp_1 _21071_ (.CLK(\clknet_leaf_19_top1.acquisition_clk ),
    .RESET_B(net165),
    .D(_01243_),
    .Q_N(_08745_),
    .Q(\top1.memory1.mem1[142][1] ));
 sg13g2_dfrbp_1 _21072_ (.CLK(\clknet_leaf_50_top1.acquisition_clk ),
    .RESET_B(net164),
    .D(_01244_),
    .Q_N(_08744_),
    .Q(\top1.memory1.mem1[142][2] ));
 sg13g2_dfrbp_1 _21073_ (.CLK(\clknet_leaf_182_top1.acquisition_clk ),
    .RESET_B(net163),
    .D(_01245_),
    .Q_N(_08743_),
    .Q(\top1.memory1.mem1[24][0] ));
 sg13g2_dfrbp_1 _21074_ (.CLK(\clknet_leaf_180_top1.acquisition_clk ),
    .RESET_B(net162),
    .D(_01246_),
    .Q_N(_08742_),
    .Q(\top1.memory1.mem1[24][1] ));
 sg13g2_dfrbp_1 _21075_ (.CLK(\clknet_leaf_114_top1.acquisition_clk ),
    .RESET_B(net161),
    .D(_01247_),
    .Q_N(_08741_),
    .Q(\top1.memory1.mem1[24][2] ));
 sg13g2_dfrbp_1 _21076_ (.CLK(\clknet_leaf_148_top1.acquisition_clk ),
    .RESET_B(net160),
    .D(_01248_),
    .Q_N(_08740_),
    .Q(\top1.memory1.mem1[36][0] ));
 sg13g2_dfrbp_1 _21077_ (.CLK(\clknet_leaf_148_top1.acquisition_clk ),
    .RESET_B(net159),
    .D(_01249_),
    .Q_N(_08739_),
    .Q(\top1.memory1.mem1[36][1] ));
 sg13g2_dfrbp_1 _21078_ (.CLK(\clknet_leaf_151_top1.acquisition_clk ),
    .RESET_B(net158),
    .D(_01250_),
    .Q_N(_08738_),
    .Q(\top1.memory1.mem1[36][2] ));
 sg13g2_dfrbp_1 _21079_ (.CLK(\clknet_leaf_52_top1.acquisition_clk ),
    .RESET_B(net157),
    .D(_01251_),
    .Q_N(_08737_),
    .Q(\top1.memory1.mem1[141][0] ));
 sg13g2_dfrbp_1 _21080_ (.CLK(\clknet_leaf_51_top1.acquisition_clk ),
    .RESET_B(net156),
    .D(_01252_),
    .Q_N(_08736_),
    .Q(\top1.memory1.mem1[141][1] ));
 sg13g2_dfrbp_1 _21081_ (.CLK(\clknet_leaf_53_top1.acquisition_clk ),
    .RESET_B(net155),
    .D(_01253_),
    .Q_N(_08735_),
    .Q(\top1.memory1.mem1[141][2] ));
 sg13g2_dfrbp_1 _21082_ (.CLK(\clknet_leaf_52_top1.acquisition_clk ),
    .RESET_B(net154),
    .D(_01254_),
    .Q_N(_08734_),
    .Q(\top1.memory1.mem1[140][0] ));
 sg13g2_dfrbp_1 _21083_ (.CLK(\clknet_leaf_51_top1.acquisition_clk ),
    .RESET_B(net153),
    .D(_01255_),
    .Q_N(_08733_),
    .Q(\top1.memory1.mem1[140][1] ));
 sg13g2_dfrbp_1 _21084_ (.CLK(\clknet_leaf_53_top1.acquisition_clk ),
    .RESET_B(net152),
    .D(_01256_),
    .Q_N(_08732_),
    .Q(\top1.memory1.mem1[140][2] ));
 sg13g2_dfrbp_1 _21085_ (.CLK(\clknet_leaf_274_top1.acquisition_clk ),
    .RESET_B(net151),
    .D(_01257_),
    .Q_N(_08731_),
    .Q(\top1.memory1.mem1[13][0] ));
 sg13g2_dfrbp_1 _21086_ (.CLK(\clknet_leaf_273_top1.acquisition_clk ),
    .RESET_B(net150),
    .D(_01258_),
    .Q_N(_08730_),
    .Q(\top1.memory1.mem1[13][1] ));
 sg13g2_dfrbp_1 _21087_ (.CLK(\clknet_leaf_282_top1.acquisition_clk ),
    .RESET_B(net149),
    .D(_01259_),
    .Q_N(_08729_),
    .Q(\top1.memory1.mem1[13][2] ));
 sg13g2_dfrbp_1 _21088_ (.CLK(\clknet_leaf_258_top1.acquisition_clk ),
    .RESET_B(net148),
    .D(_01260_),
    .Q_N(_08728_),
    .Q(\top1.memory1.mem1[23][0] ));
 sg13g2_dfrbp_1 _21089_ (.CLK(\clknet_leaf_258_top1.acquisition_clk ),
    .RESET_B(net147),
    .D(_01261_),
    .Q_N(_08727_),
    .Q(\top1.memory1.mem1[23][1] ));
 sg13g2_dfrbp_1 _21090_ (.CLK(\clknet_leaf_186_top1.acquisition_clk ),
    .RESET_B(net146),
    .D(_01262_),
    .Q_N(_08726_),
    .Q(\top1.memory1.mem1[23][2] ));
 sg13g2_dfrbp_1 _21091_ (.CLK(\clknet_leaf_54_top1.acquisition_clk ),
    .RESET_B(net145),
    .D(_01263_),
    .Q_N(_08725_),
    .Q(\top1.memory1.mem1[138][0] ));
 sg13g2_dfrbp_1 _21092_ (.CLK(\clknet_leaf_56_top1.acquisition_clk ),
    .RESET_B(net144),
    .D(_01264_),
    .Q_N(_08724_),
    .Q(\top1.memory1.mem1[138][1] ));
 sg13g2_dfrbp_1 _21093_ (.CLK(\clknet_leaf_50_top1.acquisition_clk ),
    .RESET_B(net143),
    .D(_01265_),
    .Q_N(_08723_),
    .Q(\top1.memory1.mem1[138][2] ));
 sg13g2_dfrbp_1 _21094_ (.CLK(\clknet_leaf_257_top1.acquisition_clk ),
    .RESET_B(net142),
    .D(_01266_),
    .Q_N(_08722_),
    .Q(\top1.memory1.mem1[22][0] ));
 sg13g2_dfrbp_1 _21095_ (.CLK(\clknet_leaf_259_top1.acquisition_clk ),
    .RESET_B(net141),
    .D(_01267_),
    .Q_N(_08721_),
    .Q(\top1.memory1.mem1[22][1] ));
 sg13g2_dfrbp_1 _21096_ (.CLK(\clknet_leaf_259_top1.acquisition_clk ),
    .RESET_B(net140),
    .D(_01268_),
    .Q_N(_08720_),
    .Q(\top1.memory1.mem1[22][2] ));
 sg13g2_dfrbp_1 _21097_ (.CLK(\clknet_leaf_54_top1.acquisition_clk ),
    .RESET_B(net139),
    .D(_01269_),
    .Q_N(_08719_),
    .Q(\top1.memory1.mem1[137][0] ));
 sg13g2_dfrbp_1 _21098_ (.CLK(\clknet_leaf_56_top1.acquisition_clk ),
    .RESET_B(net138),
    .D(_01270_),
    .Q_N(_08718_),
    .Q(\top1.memory1.mem1[137][1] ));
 sg13g2_dfrbp_1 _21099_ (.CLK(\clknet_leaf_50_top1.acquisition_clk ),
    .RESET_B(net137),
    .D(_01271_),
    .Q_N(_08717_),
    .Q(\top1.memory1.mem1[137][2] ));
 sg13g2_dfrbp_1 _21100_ (.CLK(\clknet_leaf_54_top1.acquisition_clk ),
    .RESET_B(net136),
    .D(_01272_),
    .Q_N(_08716_),
    .Q(\top1.memory1.mem1[136][0] ));
 sg13g2_dfrbp_1 _21101_ (.CLK(\clknet_leaf_54_top1.acquisition_clk ),
    .RESET_B(net135),
    .D(_01273_),
    .Q_N(_08715_),
    .Q(\top1.memory1.mem1[136][1] ));
 sg13g2_dfrbp_1 _21102_ (.CLK(\clknet_leaf_50_top1.acquisition_clk ),
    .RESET_B(net134),
    .D(_01274_),
    .Q_N(_08714_),
    .Q(\top1.memory1.mem1[136][2] ));
 sg13g2_dfrbp_1 _21103_ (.CLK(\clknet_leaf_49_top1.acquisition_clk ),
    .RESET_B(net133),
    .D(_01275_),
    .Q_N(_08713_),
    .Q(\top1.memory1.mem1[135][0] ));
 sg13g2_dfrbp_1 _21104_ (.CLK(\clknet_leaf_57_top1.acquisition_clk ),
    .RESET_B(net132),
    .D(_01276_),
    .Q_N(_08712_),
    .Q(\top1.memory1.mem1[135][1] ));
 sg13g2_dfrbp_1 _21105_ (.CLK(\clknet_leaf_49_top1.acquisition_clk ),
    .RESET_B(net131),
    .D(_01277_),
    .Q_N(_08711_),
    .Q(\top1.memory1.mem1[135][2] ));
 sg13g2_dfrbp_1 _21106_ (.CLK(\clknet_leaf_258_top1.acquisition_clk ),
    .RESET_B(net130),
    .D(_01278_),
    .Q_N(_08710_),
    .Q(\top1.memory1.mem1[21][0] ));
 sg13g2_dfrbp_1 _21107_ (.CLK(\clknet_leaf_259_top1.acquisition_clk ),
    .RESET_B(net129),
    .D(_01279_),
    .Q_N(_08709_),
    .Q(\top1.memory1.mem1[21][1] ));
 sg13g2_dfrbp_1 _21108_ (.CLK(\clknet_leaf_185_top1.acquisition_clk ),
    .RESET_B(net128),
    .D(_01280_),
    .Q_N(_08708_),
    .Q(\top1.memory1.mem1[21][2] ));
 sg13g2_dfrbp_1 _21109_ (.CLK(\clknet_leaf_45_top1.acquisition_clk ),
    .RESET_B(net127),
    .D(_01281_),
    .Q_N(_08707_),
    .Q(\top1.memory1.mem1[134][0] ));
 sg13g2_dfrbp_1 _21110_ (.CLK(\clknet_leaf_57_top1.acquisition_clk ),
    .RESET_B(net126),
    .D(_01282_),
    .Q_N(_08706_),
    .Q(\top1.memory1.mem1[134][1] ));
 sg13g2_dfrbp_1 _21111_ (.CLK(\clknet_leaf_44_top1.acquisition_clk ),
    .RESET_B(net125),
    .D(_01283_),
    .Q_N(_08705_),
    .Q(\top1.memory1.mem1[134][2] ));
 sg13g2_dfrbp_1 _21112_ (.CLK(\clknet_leaf_85_top1.acquisition_clk ),
    .RESET_B(net124),
    .D(_01284_),
    .Q_N(_08704_),
    .Q(\top1.memory2.mem2[9][0] ));
 sg13g2_dfrbp_1 _21113_ (.CLK(\clknet_leaf_86_top1.acquisition_clk ),
    .RESET_B(net123),
    .D(_01285_),
    .Q_N(_08703_),
    .Q(\top1.memory2.mem2[9][1] ));
 sg13g2_dfrbp_1 _21114_ (.CLK(\clknet_leaf_90_top1.acquisition_clk ),
    .RESET_B(net122),
    .D(_01286_),
    .Q_N(_08702_),
    .Q(\top1.memory2.mem2[9][2] ));
 sg13g2_dfrbp_1 _21115_ (.CLK(\clknet_leaf_48_top1.acquisition_clk ),
    .RESET_B(net121),
    .D(_01287_),
    .Q_N(_08701_),
    .Q(\top1.memory1.mem1[133][0] ));
 sg13g2_dfrbp_1 _21116_ (.CLK(\clknet_leaf_57_top1.acquisition_clk ),
    .RESET_B(net120),
    .D(_01288_),
    .Q_N(_08700_),
    .Q(\top1.memory1.mem1[133][1] ));
 sg13g2_dfrbp_1 _21117_ (.CLK(\clknet_leaf_22_top1.acquisition_clk ),
    .RESET_B(net119),
    .D(_01289_),
    .Q_N(_08699_),
    .Q(\top1.memory1.mem1[133][2] ));
 sg13g2_dfrbp_1 _21118_ (.CLK(\clknet_leaf_18_top1.acquisition_clk ),
    .RESET_B(net118),
    .D(_01290_),
    .Q_N(_08698_),
    .Q(\top1.memory1.mem1[131][0] ));
 sg13g2_dfrbp_1 _21119_ (.CLK(\clknet_leaf_20_top1.acquisition_clk ),
    .RESET_B(net117),
    .D(_01291_),
    .Q_N(_08697_),
    .Q(\top1.memory1.mem1[131][1] ));
 sg13g2_dfrbp_1 _21120_ (.CLK(\clknet_leaf_20_top1.acquisition_clk ),
    .RESET_B(net116),
    .D(_01292_),
    .Q_N(_08696_),
    .Q(\top1.memory1.mem1[131][2] ));
 sg13g2_dfrbp_1 _21121_ (.CLK(\clknet_leaf_18_top1.acquisition_clk ),
    .RESET_B(net115),
    .D(_01293_),
    .Q_N(_08695_),
    .Q(\top1.memory1.mem1[130][0] ));
 sg13g2_dfrbp_1 _21122_ (.CLK(\clknet_leaf_20_top1.acquisition_clk ),
    .RESET_B(net114),
    .D(_01294_),
    .Q_N(_08694_),
    .Q(\top1.memory1.mem1[130][1] ));
 sg13g2_dfrbp_1 _21123_ (.CLK(\clknet_leaf_20_top1.acquisition_clk ),
    .RESET_B(net113),
    .D(_01295_),
    .Q_N(_08693_),
    .Q(\top1.memory1.mem1[130][2] ));
 sg13g2_dfrbp_1 _21124_ (.CLK(\clknet_leaf_276_top1.acquisition_clk ),
    .RESET_B(net112),
    .D(_01296_),
    .Q_N(_08692_),
    .Q(\top1.memory1.mem1[12][0] ));
 sg13g2_dfrbp_1 _21125_ (.CLK(\clknet_leaf_273_top1.acquisition_clk ),
    .RESET_B(net111),
    .D(_01297_),
    .Q_N(_08691_),
    .Q(\top1.memory1.mem1[12][1] ));
 sg13g2_dfrbp_1 _21126_ (.CLK(\clknet_leaf_276_top1.acquisition_clk ),
    .RESET_B(net110),
    .D(_01298_),
    .Q_N(_08690_),
    .Q(\top1.memory1.mem1[12][2] ));
 sg13g2_dfrbp_1 _21127_ (.CLK(\clknet_leaf_257_top1.acquisition_clk ),
    .RESET_B(net109),
    .D(_01299_),
    .Q_N(_08689_),
    .Q(\top1.memory1.mem1[20][0] ));
 sg13g2_dfrbp_1 _21128_ (.CLK(\clknet_leaf_258_top1.acquisition_clk ),
    .RESET_B(net108),
    .D(_01300_),
    .Q_N(_08688_),
    .Q(\top1.memory1.mem1[20][1] ));
 sg13g2_dfrbp_1 _21129_ (.CLK(\clknet_leaf_185_top1.acquisition_clk ),
    .RESET_B(net107),
    .D(_01301_),
    .Q_N(_08687_),
    .Q(\top1.memory1.mem1[20][2] ));
 sg13g2_dfrbp_1 _21130_ (.CLK(\clknet_leaf_277_top1.acquisition_clk ),
    .RESET_B(net106),
    .D(_01302_),
    .Q_N(_08686_),
    .Q(\top1.memory1.mem1[1][0] ));
 sg13g2_dfrbp_1 _21131_ (.CLK(\clknet_leaf_279_top1.acquisition_clk ),
    .RESET_B(net105),
    .D(_01303_),
    .Q_N(_08685_),
    .Q(\top1.memory1.mem1[1][1] ));
 sg13g2_dfrbp_1 _21132_ (.CLK(\clknet_leaf_281_top1.acquisition_clk ),
    .RESET_B(net104),
    .D(_01304_),
    .Q_N(_08684_),
    .Q(\top1.memory1.mem1[1][2] ));
 sg13g2_dfrbp_1 _21133_ (.CLK(\clknet_leaf_39_top1.acquisition_clk ),
    .RESET_B(net103),
    .D(_01305_),
    .Q_N(_08683_),
    .Q(\top1.memory1.mem1[199][0] ));
 sg13g2_dfrbp_1 _21134_ (.CLK(\clknet_leaf_35_top1.acquisition_clk ),
    .RESET_B(net102),
    .D(_01306_),
    .Q_N(_08682_),
    .Q(\top1.memory1.mem1[199][1] ));
 sg13g2_dfrbp_1 _21135_ (.CLK(\clknet_leaf_33_top1.acquisition_clk ),
    .RESET_B(net101),
    .D(_01307_),
    .Q_N(_08681_),
    .Q(\top1.memory1.mem1[199][2] ));
 sg13g2_dfrbp_1 _21136_ (.CLK(\clknet_leaf_39_top1.acquisition_clk ),
    .RESET_B(net7742),
    .D(net4852),
    .Q_N(_00000_),
    .Q(\top1.addr_in[8] ));
 sg13g2_dfrbp_1 _21137_ (.CLK(net6745),
    .RESET_B(net7746),
    .D(_01309_),
    .Q_N(_00006_),
    .Q(\top1.addr_out[8] ));
 sg13g2_dfrbp_1 _21138_ (.CLK(\clknet_leaf_37_top1.acquisition_clk ),
    .RESET_B(net7742),
    .D(_00007_),
    .Q_N(_09933_),
    .Q(\top1.addr_in[0] ));
 sg13g2_dfrbp_1 _21139_ (.CLK(\clknet_leaf_37_top1.acquisition_clk ),
    .RESET_B(net7742),
    .D(_00008_),
    .Q_N(_09934_),
    .Q(\top1.addr_in[1] ));
 sg13g2_dfrbp_1 _21140_ (.CLK(\clknet_leaf_37_top1.acquisition_clk ),
    .RESET_B(net7742),
    .D(_00009_),
    .Q_N(_09935_),
    .Q(\top1.addr_in[2] ));
 sg13g2_dfrbp_1 _21141_ (.CLK(\clknet_leaf_37_top1.acquisition_clk ),
    .RESET_B(net7742),
    .D(_00010_),
    .Q_N(_09936_),
    .Q(\top1.addr_in[3] ));
 sg13g2_dfrbp_1 _21142_ (.CLK(\clknet_leaf_35_top1.acquisition_clk ),
    .RESET_B(net7744),
    .D(_00011_),
    .Q_N(_09937_),
    .Q(\top1.addr_in[4] ));
 sg13g2_dfrbp_1 _21143_ (.CLK(\clknet_leaf_34_top1.acquisition_clk ),
    .RESET_B(net7744),
    .D(_00012_),
    .Q_N(_09938_),
    .Q(\top1.addr_in[5] ));
 sg13g2_dfrbp_1 _21144_ (.CLK(\clknet_leaf_34_top1.acquisition_clk ),
    .RESET_B(net7744),
    .D(_00013_),
    .Q_N(_09939_),
    .Q(\top1.addr_in[6] ));
 sg13g2_dfrbp_1 _21145_ (.CLK(\clknet_leaf_35_top1.acquisition_clk ),
    .RESET_B(net7744),
    .D(_00014_),
    .Q_N(_08680_),
    .Q(\top1.addr_in[7] ));
 sg13g2_dfrbp_1 _21146_ (.CLK(\clknet_leaf_40_top1.acquisition_clk ),
    .RESET_B(net7742),
    .D(net4859),
    .Q_N(_08679_),
    .Q(\top1.bank0_full ));
 sg13g2_dfrbp_1 _21147_ (.CLK(\clknet_leaf_40_top1.acquisition_clk ),
    .RESET_B(net7743),
    .D(net4483),
    .Q_N(_08678_),
    .Q(\top1.fsm.idx_final[0] ));
 sg13g2_dfrbp_1 _21148_ (.CLK(\clknet_leaf_39_top1.acquisition_clk ),
    .RESET_B(net7746),
    .D(net4586),
    .Q_N(_08677_),
    .Q(\top1.fsm.idx_final[1] ));
 sg13g2_dfrbp_1 _21149_ (.CLK(\clknet_leaf_39_top1.acquisition_clk ),
    .RESET_B(net7745),
    .D(net4676),
    .Q_N(_08676_),
    .Q(\top1.fsm.idx_final[2] ));
 sg13g2_dfrbp_1 _21150_ (.CLK(\clknet_leaf_39_top1.acquisition_clk ),
    .RESET_B(net7746),
    .D(net4590),
    .Q_N(_08675_),
    .Q(\top1.fsm.idx_final[3] ));
 sg13g2_dfrbp_1 _21151_ (.CLK(\clknet_leaf_34_top1.acquisition_clk ),
    .RESET_B(net7744),
    .D(net4740),
    .Q_N(_08674_),
    .Q(\top1.fsm.idx_final[4] ));
 sg13g2_dfrbp_1 _21152_ (.CLK(\clknet_leaf_34_top1.acquisition_clk ),
    .RESET_B(net7744),
    .D(_01316_),
    .Q_N(_08673_),
    .Q(\top1.fsm.idx_final[5] ));
 sg13g2_dfrbp_1 _21153_ (.CLK(\clknet_leaf_34_top1.acquisition_clk ),
    .RESET_B(net7744),
    .D(net4706),
    .Q_N(_08672_),
    .Q(\top1.fsm.idx_final[6] ));
 sg13g2_dfrbp_1 _21154_ (.CLK(\clknet_leaf_39_top1.acquisition_clk ),
    .RESET_B(net7744),
    .D(net4304),
    .Q_N(_08671_),
    .Q(\top1.fsm.idx_final[7] ));
 sg13g2_dfrbp_1 _21155_ (.CLK(\clknet_leaf_40_top1.acquisition_clk ),
    .RESET_B(net7742),
    .D(net4862),
    .Q_N(_09940_),
    .Q(\top1.bank1_full ));
 sg13g2_dfrbp_1 _21156_ (.CLK(net6740),
    .RESET_B(net7740),
    .D(_00015_),
    .Q_N(_09941_),
    .Q(\top1.piso_time_reg.register[0] ));
 sg13g2_dfrbp_1 _21157_ (.CLK(net6740),
    .RESET_B(net7734),
    .D(_00026_),
    .Q_N(_09942_),
    .Q(\top1.piso_time_reg.register[1] ));
 sg13g2_dfrbp_1 _21158_ (.CLK(net6740),
    .RESET_B(net7734),
    .D(_00037_),
    .Q_N(_09943_),
    .Q(\top1.piso_time_reg.register[2] ));
 sg13g2_dfrbp_1 _21159_ (.CLK(net6740),
    .RESET_B(net7732),
    .D(_00039_),
    .Q_N(_09944_),
    .Q(\top1.piso_time_reg.register[3] ));
 sg13g2_dfrbp_1 _21160_ (.CLK(net6740),
    .RESET_B(net7737),
    .D(_00040_),
    .Q_N(_09945_),
    .Q(\top1.piso_time_reg.register[4] ));
 sg13g2_dfrbp_1 _21161_ (.CLK(net6741),
    .RESET_B(net7737),
    .D(_00041_),
    .Q_N(_09946_),
    .Q(\top1.piso_time_reg.register[5] ));
 sg13g2_dfrbp_1 _21162_ (.CLK(net6740),
    .RESET_B(net7737),
    .D(_00042_),
    .Q_N(_09947_),
    .Q(\top1.piso_time_reg.register[6] ));
 sg13g2_dfrbp_1 _21163_ (.CLK(net6740),
    .RESET_B(net7737),
    .D(_00043_),
    .Q_N(_09948_),
    .Q(\top1.piso_time_reg.register[7] ));
 sg13g2_dfrbp_1 _21164_ (.CLK(net6741),
    .RESET_B(net7737),
    .D(_00044_),
    .Q_N(_09949_),
    .Q(\top1.piso_time_reg.register[8] ));
 sg13g2_dfrbp_1 _21165_ (.CLK(net6741),
    .RESET_B(net7738),
    .D(_00045_),
    .Q_N(_09950_),
    .Q(\top1.piso_time_reg.register[9] ));
 sg13g2_dfrbp_1 _21166_ (.CLK(net6741),
    .RESET_B(net7738),
    .D(_00016_),
    .Q_N(_09951_),
    .Q(\top1.piso_time_reg.register[10] ));
 sg13g2_dfrbp_1 _21167_ (.CLK(net6741),
    .RESET_B(net7737),
    .D(_00017_),
    .Q_N(_09952_),
    .Q(\top1.piso_time_reg.register[11] ));
 sg13g2_dfrbp_1 _21168_ (.CLK(net6741),
    .RESET_B(net7735),
    .D(_00018_),
    .Q_N(_09953_),
    .Q(\top1.piso_time_reg.register[12] ));
 sg13g2_dfrbp_1 _21169_ (.CLK(net6737),
    .RESET_B(net7735),
    .D(_00019_),
    .Q_N(_09954_),
    .Q(\top1.piso_time_reg.register[13] ));
 sg13g2_dfrbp_1 _21170_ (.CLK(net6737),
    .RESET_B(net7735),
    .D(_00020_),
    .Q_N(_09955_),
    .Q(\top1.piso_time_reg.register[14] ));
 sg13g2_dfrbp_1 _21171_ (.CLK(net6737),
    .RESET_B(net7729),
    .D(_00021_),
    .Q_N(_09956_),
    .Q(\top1.piso_time_reg.register[15] ));
 sg13g2_dfrbp_1 _21172_ (.CLK(net6737),
    .RESET_B(net7730),
    .D(_00022_),
    .Q_N(_09957_),
    .Q(\top1.piso_time_reg.register[16] ));
 sg13g2_dfrbp_1 _21173_ (.CLK(net6736),
    .RESET_B(net7729),
    .D(_00023_),
    .Q_N(_09958_),
    .Q(\top1.piso_time_reg.register[17] ));
 sg13g2_dfrbp_1 _21174_ (.CLK(net6736),
    .RESET_B(net7729),
    .D(_00024_),
    .Q_N(_09959_),
    .Q(\top1.piso_time_reg.register[18] ));
 sg13g2_dfrbp_1 _21175_ (.CLK(net6736),
    .RESET_B(net7727),
    .D(_00025_),
    .Q_N(_09960_),
    .Q(\top1.piso_time_reg.register[19] ));
 sg13g2_dfrbp_1 _21176_ (.CLK(net6737),
    .RESET_B(net7726),
    .D(_00027_),
    .Q_N(_09961_),
    .Q(\top1.piso_time_reg.register[20] ));
 sg13g2_dfrbp_1 _21177_ (.CLK(net6737),
    .RESET_B(net7728),
    .D(_00028_),
    .Q_N(_09962_),
    .Q(\top1.piso_time_reg.register[21] ));
 sg13g2_dfrbp_1 _21178_ (.CLK(net6736),
    .RESET_B(net7730),
    .D(_00029_),
    .Q_N(_09963_),
    .Q(\top1.piso_time_reg.register[22] ));
 sg13g2_dfrbp_1 _21179_ (.CLK(net6736),
    .RESET_B(net7725),
    .D(_00030_),
    .Q_N(_09964_),
    .Q(\top1.piso_time_reg.register[23] ));
 sg13g2_dfrbp_1 _21180_ (.CLK(net6736),
    .RESET_B(net7725),
    .D(_00031_),
    .Q_N(_09965_),
    .Q(\top1.piso_time_reg.register[24] ));
 sg13g2_dfrbp_1 _21181_ (.CLK(net6736),
    .RESET_B(net7725),
    .D(_00032_),
    .Q_N(_09966_),
    .Q(\top1.piso_time_reg.register[25] ));
 sg13g2_dfrbp_1 _21182_ (.CLK(net6736),
    .RESET_B(net7725),
    .D(_00033_),
    .Q_N(_09967_),
    .Q(\top1.piso_time_reg.register[26] ));
 sg13g2_dfrbp_1 _21183_ (.CLK(net6738),
    .RESET_B(net7731),
    .D(_00034_),
    .Q_N(_09968_),
    .Q(\top1.piso_time_reg.register[27] ));
 sg13g2_dfrbp_1 _21184_ (.CLK(net6738),
    .RESET_B(net7725),
    .D(_00035_),
    .Q_N(_09969_),
    .Q(\top1.piso_time_reg.register[28] ));
 sg13g2_dfrbp_1 _21185_ (.CLK(net6738),
    .RESET_B(net7724),
    .D(_00036_),
    .Q_N(_09970_),
    .Q(\top1.piso_time_reg.register[29] ));
 sg13g2_dfrbp_1 _21186_ (.CLK(net6738),
    .RESET_B(net7723),
    .D(_00038_),
    .Q_N(_09971_),
    .Q(\top1.piso_time_reg.register[30] ));
 sg13g2_dfrbp_1 _21187_ (.CLK(net7571),
    .RESET_B(net7732),
    .D(\top1.event_time[0] ),
    .Q_N(_09972_),
    .Q(\top1.event_time_out[0] ));
 sg13g2_dfrbp_1 _21188_ (.CLK(net7571),
    .RESET_B(net7732),
    .D(\top1.event_time[1] ),
    .Q_N(_09973_),
    .Q(\top1.event_time_out[1] ));
 sg13g2_dfrbp_1 _21189_ (.CLK(net7571),
    .RESET_B(net7733),
    .D(\top1.event_time[2] ),
    .Q_N(_09974_),
    .Q(\top1.event_time_out[2] ));
 sg13g2_dfrbp_1 _21190_ (.CLK(net7569),
    .RESET_B(net7733),
    .D(\top1.event_time[3] ),
    .Q_N(_09975_),
    .Q(\top1.event_time_out[3] ));
 sg13g2_dfrbp_1 _21191_ (.CLK(net7569),
    .RESET_B(net7733),
    .D(\top1.event_time[4] ),
    .Q_N(_09976_),
    .Q(\top1.event_time_out[4] ));
 sg13g2_dfrbp_1 _21192_ (.CLK(net7571),
    .RESET_B(net7736),
    .D(\top1.event_time[5] ),
    .Q_N(_09977_),
    .Q(\top1.event_time_out[5] ));
 sg13g2_dfrbp_1 _21193_ (.CLK(net7571),
    .RESET_B(net7737),
    .D(\top1.event_time[6] ),
    .Q_N(_09978_),
    .Q(\top1.event_time_out[6] ));
 sg13g2_dfrbp_1 _21194_ (.CLK(net7571),
    .RESET_B(net7737),
    .D(\top1.event_time[7] ),
    .Q_N(_09979_),
    .Q(\top1.event_time_out[7] ));
 sg13g2_dfrbp_1 _21195_ (.CLK(net7571),
    .RESET_B(net7738),
    .D(\top1.event_time[8] ),
    .Q_N(_09980_),
    .Q(\top1.event_time_out[8] ));
 sg13g2_dfrbp_1 _21196_ (.CLK(net7571),
    .RESET_B(net7738),
    .D(\top1.event_time[9] ),
    .Q_N(_09981_),
    .Q(\top1.event_time_out[9] ));
 sg13g2_dfrbp_1 _21197_ (.CLK(net7572),
    .RESET_B(net7739),
    .D(\top1.event_time[10] ),
    .Q_N(_09982_),
    .Q(\top1.event_time_out[10] ));
 sg13g2_dfrbp_1 _21198_ (.CLK(net7572),
    .RESET_B(net7739),
    .D(\top1.event_time[11] ),
    .Q_N(_09983_),
    .Q(\top1.event_time_out[11] ));
 sg13g2_dfrbp_1 _21199_ (.CLK(net7572),
    .RESET_B(net7736),
    .D(\top1.event_time[12] ),
    .Q_N(_09984_),
    .Q(\top1.event_time_out[12] ));
 sg13g2_dfrbp_1 _21200_ (.CLK(net7569),
    .RESET_B(net7735),
    .D(\top1.event_time[13] ),
    .Q_N(_09985_),
    .Q(\top1.event_time_out[13] ));
 sg13g2_dfrbp_1 _21201_ (.CLK(net7569),
    .RESET_B(net7735),
    .D(\top1.event_time[14] ),
    .Q_N(_09986_),
    .Q(\top1.event_time_out[14] ));
 sg13g2_dfrbp_1 _21202_ (.CLK(net7569),
    .RESET_B(net7729),
    .D(\top1.event_time[15] ),
    .Q_N(_09987_),
    .Q(\top1.event_time_out[15] ));
 sg13g2_dfrbp_1 _21203_ (.CLK(net7568),
    .RESET_B(net7729),
    .D(\top1.event_time[16] ),
    .Q_N(_09988_),
    .Q(\top1.event_time_out[16] ));
 sg13g2_dfrbp_1 _21204_ (.CLK(net7568),
    .RESET_B(net7729),
    .D(\top1.event_time[17] ),
    .Q_N(_09989_),
    .Q(\top1.event_time_out[17] ));
 sg13g2_dfrbp_1 _21205_ (.CLK(net7568),
    .RESET_B(net7727),
    .D(\top1.event_time[18] ),
    .Q_N(_09990_),
    .Q(\top1.event_time_out[18] ));
 sg13g2_dfrbp_1 _21206_ (.CLK(net7568),
    .RESET_B(net7727),
    .D(\top1.event_time[19] ),
    .Q_N(_09991_),
    .Q(\top1.event_time_out[19] ));
 sg13g2_dfrbp_1 _21207_ (.CLK(net7567),
    .RESET_B(net7726),
    .D(\top1.event_time[20] ),
    .Q_N(_09992_),
    .Q(\top1.event_time_out[20] ));
 sg13g2_dfrbp_1 _21208_ (.CLK(net7567),
    .RESET_B(net7726),
    .D(\top1.event_time[21] ),
    .Q_N(_09993_),
    .Q(\top1.event_time_out[21] ));
 sg13g2_dfrbp_1 _21209_ (.CLK(net7567),
    .RESET_B(net7728),
    .D(\top1.event_time[22] ),
    .Q_N(_09994_),
    .Q(\top1.event_time_out[22] ));
 sg13g2_dfrbp_1 _21210_ (.CLK(net7567),
    .RESET_B(net7728),
    .D(\top1.event_time[23] ),
    .Q_N(_09995_),
    .Q(\top1.event_time_out[23] ));
 sg13g2_dfrbp_1 _21211_ (.CLK(net7567),
    .RESET_B(net7724),
    .D(\top1.event_time[24] ),
    .Q_N(_09996_),
    .Q(\top1.event_time_out[24] ));
 sg13g2_dfrbp_1 _21212_ (.CLK(net7567),
    .RESET_B(net7724),
    .D(\top1.event_time[25] ),
    .Q_N(_09997_),
    .Q(\top1.event_time_out[25] ));
 sg13g2_dfrbp_1 _21213_ (.CLK(net7567),
    .RESET_B(net7724),
    .D(\top1.event_time[26] ),
    .Q_N(_09998_),
    .Q(\top1.event_time_out[26] ));
 sg13g2_dfrbp_1 _21214_ (.CLK(net7570),
    .RESET_B(net7724),
    .D(\top1.event_time[27] ),
    .Q_N(_09999_),
    .Q(\top1.event_time_out[27] ));
 sg13g2_dfrbp_1 _21215_ (.CLK(net7570),
    .RESET_B(net7723),
    .D(\top1.event_time[28] ),
    .Q_N(_10000_),
    .Q(\top1.event_time_out[28] ));
 sg13g2_dfrbp_1 _21216_ (.CLK(net7570),
    .RESET_B(net7724),
    .D(\top1.event_time[29] ),
    .Q_N(_10001_),
    .Q(\top1.event_time_out[29] ));
 sg13g2_dfrbp_1 _21217_ (.CLK(net7570),
    .RESET_B(net7723),
    .D(\top1.event_time[30] ),
    .Q_N(_10002_),
    .Q(\top1.event_time_out[30] ));
 sg13g2_dfrbp_1 _21218_ (.CLK(net7570),
    .RESET_B(net7723),
    .D(\top1.event_time[31] ),
    .Q_N(_08670_),
    .Q(\top1.event_time_out[31] ));
 sg13g2_dfrbp_1 _21219_ (.CLK(net7718),
    .RESET_B(net7728),
    .D(_01320_),
    .Q_N(_08669_),
    .Q(\top1.event_time[22] ));
 sg13g2_dfrbp_1 _21220_ (.CLK(net7718),
    .RESET_B(net7728),
    .D(_01321_),
    .Q_N(_08668_),
    .Q(\top1.event_time[23] ));
 sg13g2_dfrbp_1 _21221_ (.CLK(net7718),
    .RESET_B(net7728),
    .D(_01322_),
    .Q_N(_08667_),
    .Q(\top1.event_time[24] ));
 sg13g2_dfrbp_1 _21222_ (.CLK(net7719),
    .RESET_B(net7725),
    .D(_01323_),
    .Q_N(_08666_),
    .Q(\top1.event_time[25] ));
 sg13g2_dfrbp_1 _21223_ (.CLK(net7719),
    .RESET_B(net7724),
    .D(_01324_),
    .Q_N(_08665_),
    .Q(\top1.event_time[26] ));
 sg13g2_dfrbp_1 _21224_ (.CLK(\clknet_leaf_252_top1.acquisition_clk ),
    .RESET_B(net100),
    .D(_01325_),
    .Q_N(_08664_),
    .Q(\top1.memory1.mem1[179][0] ));
 sg13g2_dfrbp_1 _21225_ (.CLK(\clknet_leaf_250_top1.acquisition_clk ),
    .RESET_B(net99),
    .D(_01326_),
    .Q_N(_08663_),
    .Q(\top1.memory1.mem1[179][1] ));
 sg13g2_dfrbp_1 _21226_ (.CLK(\clknet_leaf_191_top1.acquisition_clk ),
    .RESET_B(net1239),
    .D(_01327_),
    .Q_N(_10003_),
    .Q(\top1.memory1.mem1[179][2] ));
 sg13g2_dfrbp_1 _21227_ (.CLK(net6746),
    .RESET_B(net7749),
    .D(_00050_),
    .Q_N(_10004_),
    .Q(\top1.reg2.register[0] ));
 sg13g2_dfrbp_1 _21228_ (.CLK(net6746),
    .RESET_B(net7748),
    .D(_00051_),
    .Q_N(_10005_),
    .Q(\top1.reg2.register[1] ));
 sg13g2_dfrbp_1 _21229_ (.CLK(net6744),
    .RESET_B(net7748),
    .D(_00047_),
    .Q_N(_10006_),
    .Q(\top1.reg1.register[0] ));
 sg13g2_dfrbp_1 _21230_ (.CLK(net6744),
    .RESET_B(net7748),
    .D(_00048_),
    .Q_N(_08662_),
    .Q(\top1.reg1.register[1] ));
 sg13g2_dfrbp_1 _21231_ (.CLK(\clknet_leaf_86_top1.acquisition_clk ),
    .RESET_B(net98),
    .D(_01328_),
    .Q_N(_08661_),
    .Q(\top1.memory1.mem2[9][0] ));
 sg13g2_dfrbp_1 _21232_ (.CLK(\clknet_leaf_85_top1.acquisition_clk ),
    .RESET_B(net97),
    .D(_01329_),
    .Q_N(_08660_),
    .Q(\top1.memory1.mem2[9][1] ));
 sg13g2_dfrbp_1 _21233_ (.CLK(\clknet_leaf_85_top1.acquisition_clk ),
    .RESET_B(net96),
    .D(_01330_),
    .Q_N(_08659_),
    .Q(\top1.memory1.mem2[9][2] ));
 sg13g2_dfrbp_1 _21234_ (.CLK(\clknet_leaf_109_top1.acquisition_clk ),
    .RESET_B(net95),
    .D(_01331_),
    .Q_N(_08658_),
    .Q(\top1.memory2.mem1[19][0] ));
 sg13g2_dfrbp_1 _21235_ (.CLK(\clknet_leaf_113_top1.acquisition_clk ),
    .RESET_B(net94),
    .D(_01332_),
    .Q_N(_08657_),
    .Q(\top1.memory2.mem1[19][1] ));
 sg13g2_dfrbp_1 _21236_ (.CLK(\clknet_leaf_106_top1.acquisition_clk ),
    .RESET_B(net93),
    .D(_01333_),
    .Q_N(_08656_),
    .Q(\top1.memory2.mem1[19][2] ));
 sg13g2_dfrbp_1 _21237_ (.CLK(\clknet_leaf_184_top1.acquisition_clk ),
    .RESET_B(net92),
    .D(_01334_),
    .Q_N(_08655_),
    .Q(\top1.memory2.mem1[29][0] ));
 sg13g2_dfrbp_1 _21238_ (.CLK(\clknet_leaf_183_top1.acquisition_clk ),
    .RESET_B(net91),
    .D(_01335_),
    .Q_N(_08654_),
    .Q(\top1.memory2.mem1[29][1] ));
 sg13g2_dfrbp_1 _21239_ (.CLK(\clknet_leaf_256_top1.acquisition_clk ),
    .RESET_B(net90),
    .D(_01336_),
    .Q_N(_08653_),
    .Q(\top1.memory2.mem1[29][2] ));
 sg13g2_dfrbp_1 _21240_ (.CLK(\clknet_leaf_151_top1.acquisition_clk ),
    .RESET_B(net89),
    .D(_01337_),
    .Q_N(_08652_),
    .Q(\top1.memory2.mem1[39][0] ));
 sg13g2_dfrbp_1 _21241_ (.CLK(\clknet_leaf_150_top1.acquisition_clk ),
    .RESET_B(net88),
    .D(_01338_),
    .Q_N(_08651_),
    .Q(\top1.memory2.mem1[39][1] ));
 sg13g2_dfrbp_1 _21242_ (.CLK(\clknet_leaf_150_top1.acquisition_clk ),
    .RESET_B(net87),
    .D(_01339_),
    .Q_N(_08650_),
    .Q(\top1.memory2.mem1[39][2] ));
 sg13g2_dfrbp_1 _21243_ (.CLK(\clknet_leaf_164_top1.acquisition_clk ),
    .RESET_B(net86),
    .D(_01340_),
    .Q_N(_08649_),
    .Q(\top1.memory2.mem1[49][0] ));
 sg13g2_dfrbp_1 _21244_ (.CLK(\clknet_leaf_165_top1.acquisition_clk ),
    .RESET_B(net85),
    .D(_01341_),
    .Q_N(_08648_),
    .Q(\top1.memory2.mem1[49][1] ));
 sg13g2_dfrbp_1 _21245_ (.CLK(\clknet_leaf_164_top1.acquisition_clk ),
    .RESET_B(net84),
    .D(_01342_),
    .Q_N(_08647_),
    .Q(\top1.memory2.mem1[49][2] ));
 sg13g2_dfrbp_1 _21246_ (.CLK(\clknet_leaf_169_top1.acquisition_clk ),
    .RESET_B(net83),
    .D(_01343_),
    .Q_N(_08646_),
    .Q(\top1.memory2.mem1[59][0] ));
 sg13g2_dfrbp_1 _21247_ (.CLK(\clknet_leaf_168_top1.acquisition_clk ),
    .RESET_B(net82),
    .D(_01344_),
    .Q_N(_08645_),
    .Q(\top1.memory2.mem1[59][1] ));
 sg13g2_dfrbp_1 _21248_ (.CLK(\clknet_leaf_167_top1.acquisition_clk ),
    .RESET_B(net81),
    .D(_01345_),
    .Q_N(_08644_),
    .Q(\top1.memory2.mem1[59][2] ));
 sg13g2_dfrbp_1 _21249_ (.CLK(\clknet_leaf_21_top1.acquisition_clk ),
    .RESET_B(net80),
    .D(_01346_),
    .Q_N(_08643_),
    .Q(\top1.memory2.mem1[69][0] ));
 sg13g2_dfrbp_1 _21250_ (.CLK(\clknet_leaf_21_top1.acquisition_clk ),
    .RESET_B(net79),
    .D(_01347_),
    .Q_N(_08642_),
    .Q(\top1.memory2.mem1[69][1] ));
 sg13g2_dfrbp_1 _21251_ (.CLK(\clknet_leaf_16_top1.acquisition_clk ),
    .RESET_B(net78),
    .D(_01348_),
    .Q_N(_08641_),
    .Q(\top1.memory2.mem1[69][2] ));
 sg13g2_dfrbp_1 _21252_ (.CLK(\clknet_leaf_15_top1.acquisition_clk ),
    .RESET_B(net77),
    .D(_01349_),
    .Q_N(_08640_),
    .Q(\top1.memory2.mem1[79][0] ));
 sg13g2_dfrbp_1 _21253_ (.CLK(\clknet_leaf_15_top1.acquisition_clk ),
    .RESET_B(net76),
    .D(_01350_),
    .Q_N(_08639_),
    .Q(\top1.memory2.mem1[79][1] ));
 sg13g2_dfrbp_1 _21254_ (.CLK(\clknet_leaf_14_top1.acquisition_clk ),
    .RESET_B(net75),
    .D(_01351_),
    .Q_N(_08638_),
    .Q(\top1.memory2.mem1[79][2] ));
 sg13g2_dfrbp_1 _21255_ (.CLK(\clknet_leaf_268_top1.acquisition_clk ),
    .RESET_B(net74),
    .D(_01352_),
    .Q_N(_08637_),
    .Q(\top1.memory2.mem1[89][0] ));
 sg13g2_dfrbp_1 _21256_ (.CLK(\clknet_leaf_288_top1.acquisition_clk ),
    .RESET_B(net73),
    .D(_01353_),
    .Q_N(_08636_),
    .Q(\top1.memory2.mem1[89][1] ));
 sg13g2_dfrbp_1 _21257_ (.CLK(\clknet_leaf_289_top1.acquisition_clk ),
    .RESET_B(net72),
    .D(_01354_),
    .Q_N(_08635_),
    .Q(\top1.memory2.mem1[89][2] ));
 sg13g2_dfrbp_1 _21258_ (.CLK(\clknet_leaf_189_top1.acquisition_clk ),
    .RESET_B(net71),
    .D(_01355_),
    .Q_N(_08634_),
    .Q(\top1.memory2.mem1[99][0] ));
 sg13g2_dfrbp_1 _21259_ (.CLK(\clknet_leaf_189_top1.acquisition_clk ),
    .RESET_B(net70),
    .D(_01356_),
    .Q_N(_08633_),
    .Q(\top1.memory2.mem1[99][1] ));
 sg13g2_dfrbp_1 _21260_ (.CLK(\clknet_leaf_179_top1.acquisition_clk ),
    .RESET_B(net69),
    .D(_01357_),
    .Q_N(_08632_),
    .Q(\top1.memory2.mem1[99][2] ));
 sg13g2_dfrbp_1 _21261_ (.CLK(\clknet_leaf_200_top1.acquisition_clk ),
    .RESET_B(net68),
    .D(_01358_),
    .Q_N(_08631_),
    .Q(\top1.memory2.mem1[109][0] ));
 sg13g2_dfrbp_1 _21262_ (.CLK(\clknet_leaf_197_top1.acquisition_clk ),
    .RESET_B(net67),
    .D(_01359_),
    .Q_N(_08630_),
    .Q(\top1.memory2.mem1[109][1] ));
 sg13g2_dfrbp_1 _21263_ (.CLK(\clknet_leaf_198_top1.acquisition_clk ),
    .RESET_B(net66),
    .D(_01360_),
    .Q_N(_08629_),
    .Q(\top1.memory2.mem1[109][2] ));
 sg13g2_dfrbp_1 _21264_ (.CLK(\clknet_leaf_219_top1.acquisition_clk ),
    .RESET_B(net65),
    .D(_01361_),
    .Q_N(_08628_),
    .Q(\top1.memory2.mem1[119][0] ));
 sg13g2_dfrbp_1 _21265_ (.CLK(\clknet_leaf_217_top1.acquisition_clk ),
    .RESET_B(net64),
    .D(_01362_),
    .Q_N(_08627_),
    .Q(\top1.memory2.mem1[119][1] ));
 sg13g2_dfrbp_1 _21266_ (.CLK(\clknet_leaf_218_top1.acquisition_clk ),
    .RESET_B(net63),
    .D(_01363_),
    .Q_N(_08626_),
    .Q(\top1.memory2.mem1[119][2] ));
 sg13g2_dfrbp_1 _21267_ (.CLK(\clknet_leaf_17_top1.acquisition_clk ),
    .RESET_B(net62),
    .D(_01364_),
    .Q_N(_08625_),
    .Q(\top1.memory2.mem1[129][0] ));
 sg13g2_dfrbp_1 _21268_ (.CLK(\clknet_leaf_19_top1.acquisition_clk ),
    .RESET_B(net61),
    .D(_01365_),
    .Q_N(_08624_),
    .Q(\top1.memory2.mem1[129][1] ));
 sg13g2_dfrbp_1 _21269_ (.CLK(\clknet_leaf_18_top1.acquisition_clk ),
    .RESET_B(net60),
    .D(_01366_),
    .Q_N(_08623_),
    .Q(\top1.memory2.mem1[129][2] ));
 sg13g2_dfrbp_1 _21270_ (.CLK(\clknet_leaf_55_top1.acquisition_clk ),
    .RESET_B(net59),
    .D(_01367_),
    .Q_N(_08622_),
    .Q(\top1.memory2.mem1[139][0] ));
 sg13g2_dfrbp_1 _21271_ (.CLK(\clknet_leaf_50_top1.acquisition_clk ),
    .RESET_B(net58),
    .D(_01368_),
    .Q_N(_08621_),
    .Q(\top1.memory2.mem1[139][1] ));
 sg13g2_dfrbp_1 _21272_ (.CLK(\clknet_leaf_56_top1.acquisition_clk ),
    .RESET_B(net57),
    .D(_01369_),
    .Q_N(_08620_),
    .Q(\top1.memory2.mem1[139][2] ));
 sg13g2_dfrbp_1 _21273_ (.CLK(\clknet_leaf_25_top1.acquisition_clk ),
    .RESET_B(net56),
    .D(_01370_),
    .Q_N(_08619_),
    .Q(\top1.memory2.mem1[149][0] ));
 sg13g2_dfrbp_1 _21274_ (.CLK(\clknet_leaf_25_top1.acquisition_clk ),
    .RESET_B(net55),
    .D(_01371_),
    .Q_N(_08618_),
    .Q(\top1.memory2.mem1[149][1] ));
 sg13g2_dfrbp_1 _21275_ (.CLK(\clknet_leaf_23_top1.acquisition_clk ),
    .RESET_B(net54),
    .D(_01372_),
    .Q_N(_08617_),
    .Q(\top1.memory2.mem1[149][2] ));
 sg13g2_dfrbp_1 _21276_ (.CLK(\clknet_leaf_59_top1.acquisition_clk ),
    .RESET_B(net53),
    .D(_01373_),
    .Q_N(_08616_),
    .Q(\top1.memory2.mem1[159][0] ));
 sg13g2_dfrbp_1 _21277_ (.CLK(\clknet_leaf_70_top1.acquisition_clk ),
    .RESET_B(net52),
    .D(_01374_),
    .Q_N(_08615_),
    .Q(\top1.memory2.mem1[159][1] ));
 sg13g2_dfrbp_1 _21278_ (.CLK(\clknet_leaf_71_top1.acquisition_clk ),
    .RESET_B(net51),
    .D(_01375_),
    .Q_N(_08614_),
    .Q(\top1.memory2.mem1[159][2] ));
 sg13g2_dfrbp_1 _21279_ (.CLK(\clknet_leaf_245_top1.acquisition_clk ),
    .RESET_B(net50),
    .D(_01376_),
    .Q_N(_08613_),
    .Q(\top1.memory2.mem1[169][0] ));
 sg13g2_dfrbp_1 _21280_ (.CLK(\clknet_leaf_244_top1.acquisition_clk ),
    .RESET_B(net49),
    .D(_01377_),
    .Q_N(_08612_),
    .Q(\top1.memory2.mem1[169][1] ));
 sg13g2_dfrbp_1 _21281_ (.CLK(\clknet_leaf_242_top1.acquisition_clk ),
    .RESET_B(net48),
    .D(_01378_),
    .Q_N(_08611_),
    .Q(\top1.memory2.mem1[169][2] ));
 sg13g2_dfrbp_1 _21282_ (.CLK(\clknet_leaf_190_top1.acquisition_clk ),
    .RESET_B(net47),
    .D(_01379_),
    .Q_N(_08610_),
    .Q(\top1.memory2.mem1[179][0] ));
 sg13g2_dfrbp_1 _21283_ (.CLK(\clknet_leaf_250_top1.acquisition_clk ),
    .RESET_B(net46),
    .D(_01380_),
    .Q_N(_08609_),
    .Q(\top1.memory2.mem1[179][1] ));
 sg13g2_dfrbp_1 _21284_ (.CLK(\clknet_leaf_251_top1.acquisition_clk ),
    .RESET_B(net45),
    .D(_01381_),
    .Q_N(_08608_),
    .Q(\top1.memory2.mem1[179][2] ));
 sg13g2_dfrbp_1 _21285_ (.CLK(\clknet_leaf_186_top1.acquisition_clk ),
    .RESET_B(net44),
    .D(_01382_),
    .Q_N(_08607_),
    .Q(\top1.memory2.mem1[189][0] ));
 sg13g2_dfrbp_1 _21286_ (.CLK(\clknet_leaf_186_top1.acquisition_clk ),
    .RESET_B(net43),
    .D(_01383_),
    .Q_N(_08606_),
    .Q(\top1.memory2.mem1[189][1] ));
 sg13g2_dfrbp_1 _21287_ (.CLK(\clknet_leaf_254_top1.acquisition_clk ),
    .RESET_B(net42),
    .D(_01384_),
    .Q_N(_08605_),
    .Q(\top1.memory2.mem1[189][2] ));
 sg13g2_dfrbp_1 _21288_ (.CLK(\clknet_leaf_39_top1.acquisition_clk ),
    .RESET_B(net41),
    .D(_01385_),
    .Q_N(_08604_),
    .Q(\top1.memory2.mem1[199][0] ));
 sg13g2_dfrbp_1 _21289_ (.CLK(\clknet_leaf_34_top1.acquisition_clk ),
    .RESET_B(net40),
    .D(_01386_),
    .Q_N(_08603_),
    .Q(\top1.memory2.mem1[199][1] ));
 sg13g2_dfrbp_1 _21290_ (.CLK(\clknet_leaf_34_top1.acquisition_clk ),
    .RESET_B(net39),
    .D(_01387_),
    .Q_N(_08602_),
    .Q(\top1.memory2.mem1[199][2] ));
 sg13g2_dfrbp_1 _21291_ (.CLK(\clknet_leaf_281_top1.acquisition_clk ),
    .RESET_B(net38),
    .D(_01388_),
    .Q_N(_08601_),
    .Q(\top1.memory2.mem1[1][0] ));
 sg13g2_dfrbp_1 _21292_ (.CLK(\clknet_leaf_280_top1.acquisition_clk ),
    .RESET_B(net37),
    .D(_01389_),
    .Q_N(_08600_),
    .Q(\top1.memory2.mem1[1][1] ));
 sg13g2_dfrbp_1 _21293_ (.CLK(\clknet_leaf_280_top1.acquisition_clk ),
    .RESET_B(net36),
    .D(_01390_),
    .Q_N(_08599_),
    .Q(\top1.memory2.mem1[1][2] ));
 sg13g2_dfrbp_1 _21294_ (.CLK(\clknet_leaf_184_top1.acquisition_clk ),
    .RESET_B(net35),
    .D(_01391_),
    .Q_N(_08598_),
    .Q(\top1.memory2.mem1[20][0] ));
 sg13g2_dfrbp_1 _21295_ (.CLK(\clknet_leaf_183_top1.acquisition_clk ),
    .RESET_B(net34),
    .D(_01392_),
    .Q_N(_08597_),
    .Q(\top1.memory2.mem1[20][1] ));
 sg13g2_dfrbp_1 _21296_ (.CLK(\clknet_leaf_258_top1.acquisition_clk ),
    .RESET_B(net33),
    .D(_01393_),
    .Q_N(_08596_),
    .Q(\top1.memory2.mem1[20][2] ));
 sg13g2_dfrbp_1 _21297_ (.CLK(\clknet_leaf_185_top1.acquisition_clk ),
    .RESET_B(net2438),
    .D(_01394_),
    .Q_N(_08595_),
    .Q(\top1.memory2.mem1[21][0] ));
 sg13g2_dfrbp_1 _21298_ (.CLK(\clknet_leaf_184_top1.acquisition_clk ),
    .RESET_B(net2437),
    .D(_01395_),
    .Q_N(_08594_),
    .Q(\top1.memory2.mem1[21][1] ));
 sg13g2_dfrbp_1 _21299_ (.CLK(\clknet_leaf_258_top1.acquisition_clk ),
    .RESET_B(net2436),
    .D(_01396_),
    .Q_N(_08593_),
    .Q(\top1.memory2.mem1[21][2] ));
 sg13g2_dfrbp_1 _21300_ (.CLK(\clknet_leaf_184_top1.acquisition_clk ),
    .RESET_B(net2435),
    .D(_01397_),
    .Q_N(_08592_),
    .Q(\top1.memory2.mem1[22][0] ));
 sg13g2_dfrbp_1 _21301_ (.CLK(\clknet_leaf_184_top1.acquisition_clk ),
    .RESET_B(net2434),
    .D(_01398_),
    .Q_N(_08591_),
    .Q(\top1.memory2.mem1[22][1] ));
 sg13g2_dfrbp_1 _21302_ (.CLK(\clknet_leaf_184_top1.acquisition_clk ),
    .RESET_B(net2433),
    .D(_01399_),
    .Q_N(_08590_),
    .Q(\top1.memory2.mem1[22][2] ));
 sg13g2_dfrbp_1 _21303_ (.CLK(\clknet_leaf_185_top1.acquisition_clk ),
    .RESET_B(net2432),
    .D(_01400_),
    .Q_N(_08589_),
    .Q(\top1.memory2.mem1[23][0] ));
 sg13g2_dfrbp_1 _21304_ (.CLK(\clknet_leaf_185_top1.acquisition_clk ),
    .RESET_B(net2431),
    .D(_01401_),
    .Q_N(_08588_),
    .Q(\top1.memory2.mem1[23][1] ));
 sg13g2_dfrbp_1 _21305_ (.CLK(\clknet_leaf_258_top1.acquisition_clk ),
    .RESET_B(net2430),
    .D(_01402_),
    .Q_N(_08587_),
    .Q(\top1.memory2.mem1[23][2] ));
 sg13g2_dfrbp_1 _21306_ (.CLK(\clknet_leaf_185_top1.acquisition_clk ),
    .RESET_B(net2429),
    .D(_01403_),
    .Q_N(_08586_),
    .Q(\top1.memory2.mem1[24][0] ));
 sg13g2_dfrbp_1 _21307_ (.CLK(\clknet_leaf_180_top1.acquisition_clk ),
    .RESET_B(net2428),
    .D(_01404_),
    .Q_N(_08585_),
    .Q(\top1.memory2.mem1[24][1] ));
 sg13g2_dfrbp_1 _21308_ (.CLK(\clknet_leaf_187_top1.acquisition_clk ),
    .RESET_B(net2427),
    .D(_01405_),
    .Q_N(_08584_),
    .Q(\top1.memory2.mem1[24][2] ));
 sg13g2_dfrbp_1 _21309_ (.CLK(\clknet_leaf_184_top1.acquisition_clk ),
    .RESET_B(net2426),
    .D(_01406_),
    .Q_N(_08583_),
    .Q(\top1.memory2.mem1[25][0] ));
 sg13g2_dfrbp_1 _21310_ (.CLK(\clknet_leaf_180_top1.acquisition_clk ),
    .RESET_B(net2425),
    .D(_01407_),
    .Q_N(_08582_),
    .Q(\top1.memory2.mem1[25][1] ));
 sg13g2_dfrbp_1 _21311_ (.CLK(\clknet_leaf_187_top1.acquisition_clk ),
    .RESET_B(net2424),
    .D(_01408_),
    .Q_N(_08581_),
    .Q(\top1.memory2.mem1[25][2] ));
 sg13g2_dfrbp_1 _21312_ (.CLK(\clknet_leaf_182_top1.acquisition_clk ),
    .RESET_B(net2423),
    .D(_01409_),
    .Q_N(_08580_),
    .Q(\top1.memory2.mem1[26][0] ));
 sg13g2_dfrbp_1 _21313_ (.CLK(\clknet_leaf_180_top1.acquisition_clk ),
    .RESET_B(net2422),
    .D(_01410_),
    .Q_N(_08579_),
    .Q(\top1.memory2.mem1[26][1] ));
 sg13g2_dfrbp_1 _21314_ (.CLK(\clknet_leaf_187_top1.acquisition_clk ),
    .RESET_B(net2421),
    .D(_01411_),
    .Q_N(_08578_),
    .Q(\top1.memory2.mem1[26][2] ));
 sg13g2_dfrbp_1 _21315_ (.CLK(\clknet_leaf_185_top1.acquisition_clk ),
    .RESET_B(net2420),
    .D(_01412_),
    .Q_N(_08577_),
    .Q(\top1.memory2.mem1[27][0] ));
 sg13g2_dfrbp_1 _21316_ (.CLK(\clknet_leaf_180_top1.acquisition_clk ),
    .RESET_B(net2419),
    .D(_01413_),
    .Q_N(_08576_),
    .Q(\top1.memory2.mem1[27][1] ));
 sg13g2_dfrbp_1 _21317_ (.CLK(\clknet_leaf_187_top1.acquisition_clk ),
    .RESET_B(net2418),
    .D(_01414_),
    .Q_N(_08575_),
    .Q(\top1.memory2.mem1[27][2] ));
 sg13g2_dfrbp_1 _21318_ (.CLK(\clknet_leaf_260_top1.acquisition_clk ),
    .RESET_B(net2417),
    .D(_01415_),
    .Q_N(_08574_),
    .Q(\top1.memory2.mem1[28][0] ));
 sg13g2_dfrbp_1 _21319_ (.CLK(\clknet_leaf_260_top1.acquisition_clk ),
    .RESET_B(net2416),
    .D(_01416_),
    .Q_N(_08573_),
    .Q(\top1.memory2.mem1[28][1] ));
 sg13g2_dfrbp_1 _21320_ (.CLK(\clknet_leaf_257_top1.acquisition_clk ),
    .RESET_B(net2415),
    .D(_01417_),
    .Q_N(_08572_),
    .Q(\top1.memory2.mem1[28][2] ));
 sg13g2_dfrbp_1 _21321_ (.CLK(\clknet_leaf_282_top1.acquisition_clk ),
    .RESET_B(net2414),
    .D(_01418_),
    .Q_N(_08571_),
    .Q(\top1.memory2.mem1[2][0] ));
 sg13g2_dfrbp_1 _21322_ (.CLK(\clknet_leaf_281_top1.acquisition_clk ),
    .RESET_B(net2413),
    .D(_01419_),
    .Q_N(_08570_),
    .Q(\top1.memory2.mem1[2][1] ));
 sg13g2_dfrbp_1 _21323_ (.CLK(\clknet_leaf_280_top1.acquisition_clk ),
    .RESET_B(net2412),
    .D(_01420_),
    .Q_N(_08569_),
    .Q(\top1.memory2.mem1[2][2] ));
 sg13g2_dfrbp_1 _21324_ (.CLK(\clknet_leaf_183_top1.acquisition_clk ),
    .RESET_B(net2411),
    .D(_01421_),
    .Q_N(_08568_),
    .Q(\top1.memory2.mem1[30][0] ));
 sg13g2_dfrbp_1 _21325_ (.CLK(\clknet_leaf_183_top1.acquisition_clk ),
    .RESET_B(net2410),
    .D(_01422_),
    .Q_N(_08567_),
    .Q(\top1.memory2.mem1[30][1] ));
 sg13g2_dfrbp_1 _21326_ (.CLK(\clknet_leaf_256_top1.acquisition_clk ),
    .RESET_B(net2409),
    .D(_01423_),
    .Q_N(_08566_),
    .Q(\top1.memory2.mem1[30][2] ));
 sg13g2_dfrbp_1 _21327_ (.CLK(\clknet_leaf_184_top1.acquisition_clk ),
    .RESET_B(net2408),
    .D(_01424_),
    .Q_N(_08565_),
    .Q(\top1.memory2.mem1[31][0] ));
 sg13g2_dfrbp_1 _21328_ (.CLK(\clknet_leaf_183_top1.acquisition_clk ),
    .RESET_B(net2407),
    .D(_01425_),
    .Q_N(_08564_),
    .Q(\top1.memory2.mem1[31][1] ));
 sg13g2_dfrbp_1 _21329_ (.CLK(\clknet_leaf_257_top1.acquisition_clk ),
    .RESET_B(net2406),
    .D(_01426_),
    .Q_N(_08563_),
    .Q(\top1.memory2.mem1[31][2] ));
 sg13g2_dfrbp_1 _21330_ (.CLK(\clknet_leaf_146_top1.acquisition_clk ),
    .RESET_B(net2405),
    .D(_01427_),
    .Q_N(_08562_),
    .Q(\top1.memory2.mem1[32][0] ));
 sg13g2_dfrbp_1 _21331_ (.CLK(\clknet_leaf_145_top1.acquisition_clk ),
    .RESET_B(net2404),
    .D(_01428_),
    .Q_N(_08561_),
    .Q(\top1.memory2.mem1[32][1] ));
 sg13g2_dfrbp_1 _21332_ (.CLK(\clknet_leaf_149_top1.acquisition_clk ),
    .RESET_B(net2403),
    .D(_01429_),
    .Q_N(_08560_),
    .Q(\top1.memory2.mem1[32][2] ));
 sg13g2_dfrbp_1 _21333_ (.CLK(\clknet_leaf_147_top1.acquisition_clk ),
    .RESET_B(net2402),
    .D(_01430_),
    .Q_N(_08559_),
    .Q(\top1.memory2.mem1[33][0] ));
 sg13g2_dfrbp_1 _21334_ (.CLK(\clknet_leaf_145_top1.acquisition_clk ),
    .RESET_B(net2401),
    .D(_01431_),
    .Q_N(_08558_),
    .Q(\top1.memory2.mem1[33][1] ));
 sg13g2_dfrbp_1 _21335_ (.CLK(\clknet_leaf_148_top1.acquisition_clk ),
    .RESET_B(net2400),
    .D(_01432_),
    .Q_N(_08557_),
    .Q(\top1.memory2.mem1[33][2] ));
 sg13g2_dfrbp_1 _21336_ (.CLK(\clknet_leaf_147_top1.acquisition_clk ),
    .RESET_B(net2399),
    .D(_01433_),
    .Q_N(_08556_),
    .Q(\top1.memory2.mem1[34][0] ));
 sg13g2_dfrbp_1 _21337_ (.CLK(\clknet_leaf_146_top1.acquisition_clk ),
    .RESET_B(net2398),
    .D(_01434_),
    .Q_N(_08555_),
    .Q(\top1.memory2.mem1[34][1] ));
 sg13g2_dfrbp_1 _21338_ (.CLK(\clknet_leaf_149_top1.acquisition_clk ),
    .RESET_B(net2397),
    .D(_01435_),
    .Q_N(_08554_),
    .Q(\top1.memory2.mem1[34][2] ));
 sg13g2_dfrbp_1 _21339_ (.CLK(\clknet_leaf_146_top1.acquisition_clk ),
    .RESET_B(net2396),
    .D(_01436_),
    .Q_N(_08553_),
    .Q(\top1.memory2.mem1[35][0] ));
 sg13g2_dfrbp_1 _21340_ (.CLK(\clknet_leaf_146_top1.acquisition_clk ),
    .RESET_B(net2395),
    .D(_01437_),
    .Q_N(_08552_),
    .Q(\top1.memory2.mem1[35][1] ));
 sg13g2_dfrbp_1 _21341_ (.CLK(\clknet_leaf_149_top1.acquisition_clk ),
    .RESET_B(net2394),
    .D(_01438_),
    .Q_N(_08551_),
    .Q(\top1.memory2.mem1[35][2] ));
 sg13g2_dfrbp_1 _21342_ (.CLK(\clknet_leaf_152_top1.acquisition_clk ),
    .RESET_B(net2393),
    .D(_01439_),
    .Q_N(_08550_),
    .Q(\top1.memory2.mem1[36][0] ));
 sg13g2_dfrbp_1 _21343_ (.CLK(\clknet_leaf_150_top1.acquisition_clk ),
    .RESET_B(net2392),
    .D(_01440_),
    .Q_N(_08549_),
    .Q(\top1.memory2.mem1[36][1] ));
 sg13g2_dfrbp_1 _21344_ (.CLK(\clknet_leaf_150_top1.acquisition_clk ),
    .RESET_B(net2391),
    .D(_01441_),
    .Q_N(_08548_),
    .Q(\top1.memory2.mem1[36][2] ));
 sg13g2_dfrbp_1 _21345_ (.CLK(\clknet_leaf_151_top1.acquisition_clk ),
    .RESET_B(net2390),
    .D(_01442_),
    .Q_N(_08547_),
    .Q(\top1.memory2.mem1[37][0] ));
 sg13g2_dfrbp_1 _21346_ (.CLK(\clknet_leaf_150_top1.acquisition_clk ),
    .RESET_B(net2389),
    .D(_01443_),
    .Q_N(_08546_),
    .Q(\top1.memory2.mem1[37][1] ));
 sg13g2_dfrbp_1 _21347_ (.CLK(\clknet_leaf_150_top1.acquisition_clk ),
    .RESET_B(net2388),
    .D(_01444_),
    .Q_N(_08545_),
    .Q(\top1.memory2.mem1[37][2] ));
 sg13g2_dfrbp_1 _21348_ (.CLK(\clknet_leaf_151_top1.acquisition_clk ),
    .RESET_B(net2387),
    .D(_01445_),
    .Q_N(_08544_),
    .Q(\top1.memory2.mem1[38][0] ));
 sg13g2_dfrbp_1 _21349_ (.CLK(\clknet_leaf_151_top1.acquisition_clk ),
    .RESET_B(net2386),
    .D(_01446_),
    .Q_N(_08543_),
    .Q(\top1.memory2.mem1[38][1] ));
 sg13g2_dfrbp_1 _21350_ (.CLK(\clknet_leaf_150_top1.acquisition_clk ),
    .RESET_B(net2385),
    .D(_01447_),
    .Q_N(_08542_),
    .Q(\top1.memory2.mem1[38][2] ));
 sg13g2_dfrbp_1 _21351_ (.CLK(\clknet_leaf_281_top1.acquisition_clk ),
    .RESET_B(net2384),
    .D(_01448_),
    .Q_N(_08541_),
    .Q(\top1.memory2.mem1[3][0] ));
 sg13g2_dfrbp_1 _21352_ (.CLK(\clknet_leaf_281_top1.acquisition_clk ),
    .RESET_B(net2383),
    .D(_01449_),
    .Q_N(_08540_),
    .Q(\top1.memory2.mem1[3][1] ));
 sg13g2_dfrbp_1 _21353_ (.CLK(\clknet_leaf_280_top1.acquisition_clk ),
    .RESET_B(net2382),
    .D(_01450_),
    .Q_N(_08539_),
    .Q(\top1.memory2.mem1[3][2] ));
 sg13g2_dfrbp_1 _21354_ (.CLK(\clknet_leaf_159_top1.acquisition_clk ),
    .RESET_B(net2381),
    .D(_01451_),
    .Q_N(_08538_),
    .Q(\top1.memory2.mem1[40][0] ));
 sg13g2_dfrbp_1 _21355_ (.CLK(\clknet_leaf_153_top1.acquisition_clk ),
    .RESET_B(net2380),
    .D(_01452_),
    .Q_N(_08537_),
    .Q(\top1.memory2.mem1[40][1] ));
 sg13g2_dfrbp_1 _21356_ (.CLK(\clknet_leaf_158_top1.acquisition_clk ),
    .RESET_B(net2379),
    .D(_01453_),
    .Q_N(_08536_),
    .Q(\top1.memory2.mem1[40][2] ));
 sg13g2_dfrbp_1 _21357_ (.CLK(\clknet_leaf_159_top1.acquisition_clk ),
    .RESET_B(net2378),
    .D(_01454_),
    .Q_N(_08535_),
    .Q(\top1.memory2.mem1[41][0] ));
 sg13g2_dfrbp_1 _21358_ (.CLK(\clknet_leaf_152_top1.acquisition_clk ),
    .RESET_B(net2377),
    .D(_01455_),
    .Q_N(_08534_),
    .Q(\top1.memory2.mem1[41][1] ));
 sg13g2_dfrbp_1 _21359_ (.CLK(\clknet_leaf_162_top1.acquisition_clk ),
    .RESET_B(net2376),
    .D(_01456_),
    .Q_N(_08533_),
    .Q(\top1.memory2.mem1[41][2] ));
 sg13g2_dfrbp_1 _21360_ (.CLK(\clknet_leaf_159_top1.acquisition_clk ),
    .RESET_B(net2375),
    .D(_01457_),
    .Q_N(_08532_),
    .Q(\top1.memory2.mem1[42][0] ));
 sg13g2_dfrbp_1 _21361_ (.CLK(\clknet_leaf_153_top1.acquisition_clk ),
    .RESET_B(net2374),
    .D(_01458_),
    .Q_N(_08531_),
    .Q(\top1.memory2.mem1[42][1] ));
 sg13g2_dfrbp_1 _21362_ (.CLK(\clknet_leaf_158_top1.acquisition_clk ),
    .RESET_B(net2373),
    .D(_01459_),
    .Q_N(_08530_),
    .Q(\top1.memory2.mem1[42][2] ));
 sg13g2_dfrbp_1 _21363_ (.CLK(\clknet_leaf_159_top1.acquisition_clk ),
    .RESET_B(net2372),
    .D(_01460_),
    .Q_N(_08529_),
    .Q(\top1.memory2.mem1[43][0] ));
 sg13g2_dfrbp_1 _21364_ (.CLK(\clknet_leaf_152_top1.acquisition_clk ),
    .RESET_B(net2371),
    .D(_01461_),
    .Q_N(_08528_),
    .Q(\top1.memory2.mem1[43][1] ));
 sg13g2_dfrbp_1 _21365_ (.CLK(\clknet_leaf_158_top1.acquisition_clk ),
    .RESET_B(net2370),
    .D(_01462_),
    .Q_N(_08527_),
    .Q(\top1.memory2.mem1[43][2] ));
 sg13g2_dfrbp_1 _21366_ (.CLK(\clknet_leaf_159_top1.acquisition_clk ),
    .RESET_B(net2369),
    .D(_01463_),
    .Q_N(_08526_),
    .Q(\top1.memory2.mem1[44][0] ));
 sg13g2_dfrbp_1 _21367_ (.CLK(\clknet_leaf_160_top1.acquisition_clk ),
    .RESET_B(net2368),
    .D(_01464_),
    .Q_N(_08525_),
    .Q(\top1.memory2.mem1[44][1] ));
 sg13g2_dfrbp_1 _21368_ (.CLK(\clknet_leaf_161_top1.acquisition_clk ),
    .RESET_B(net2367),
    .D(_01465_),
    .Q_N(_08524_),
    .Q(\top1.memory2.mem1[44][2] ));
 sg13g2_dfrbp_1 _21369_ (.CLK(\clknet_leaf_159_top1.acquisition_clk ),
    .RESET_B(net2366),
    .D(_01466_),
    .Q_N(_08523_),
    .Q(\top1.memory2.mem1[45][0] ));
 sg13g2_dfrbp_1 _21370_ (.CLK(\clknet_leaf_160_top1.acquisition_clk ),
    .RESET_B(net2365),
    .D(_01467_),
    .Q_N(_08522_),
    .Q(\top1.memory2.mem1[45][1] ));
 sg13g2_dfrbp_1 _21371_ (.CLK(\clknet_leaf_161_top1.acquisition_clk ),
    .RESET_B(net2364),
    .D(_01468_),
    .Q_N(_08521_),
    .Q(\top1.memory2.mem1[45][2] ));
 sg13g2_dfrbp_1 _21372_ (.CLK(\clknet_leaf_160_top1.acquisition_clk ),
    .RESET_B(net2363),
    .D(_01469_),
    .Q_N(_08520_),
    .Q(\top1.memory2.mem1[46][0] ));
 sg13g2_dfrbp_1 _21373_ (.CLK(\clknet_leaf_160_top1.acquisition_clk ),
    .RESET_B(net2362),
    .D(_01470_),
    .Q_N(_08519_),
    .Q(\top1.memory2.mem1[46][1] ));
 sg13g2_dfrbp_1 _21374_ (.CLK(\clknet_leaf_161_top1.acquisition_clk ),
    .RESET_B(net2361),
    .D(_01471_),
    .Q_N(_08518_),
    .Q(\top1.memory2.mem1[46][2] ));
 sg13g2_dfrbp_1 _21375_ (.CLK(\clknet_leaf_160_top1.acquisition_clk ),
    .RESET_B(net2360),
    .D(_01472_),
    .Q_N(_08517_),
    .Q(\top1.memory2.mem1[47][0] ));
 sg13g2_dfrbp_1 _21376_ (.CLK(\clknet_leaf_160_top1.acquisition_clk ),
    .RESET_B(net2359),
    .D(_01473_),
    .Q_N(_08516_),
    .Q(\top1.memory2.mem1[47][1] ));
 sg13g2_dfrbp_1 _21377_ (.CLK(\clknet_leaf_161_top1.acquisition_clk ),
    .RESET_B(net2358),
    .D(_01474_),
    .Q_N(_08515_),
    .Q(\top1.memory2.mem1[47][2] ));
 sg13g2_dfrbp_1 _21378_ (.CLK(\clknet_leaf_164_top1.acquisition_clk ),
    .RESET_B(net2357),
    .D(_01475_),
    .Q_N(_08514_),
    .Q(\top1.memory2.mem1[48][0] ));
 sg13g2_dfrbp_1 _21379_ (.CLK(\clknet_leaf_165_top1.acquisition_clk ),
    .RESET_B(net2356),
    .D(_01476_),
    .Q_N(_08513_),
    .Q(\top1.memory2.mem1[48][1] ));
 sg13g2_dfrbp_1 _21380_ (.CLK(\clknet_leaf_164_top1.acquisition_clk ),
    .RESET_B(net2355),
    .D(_01477_),
    .Q_N(_08512_),
    .Q(\top1.memory2.mem1[48][2] ));
 sg13g2_dfrbp_1 _21381_ (.CLK(\clknet_leaf_262_top1.acquisition_clk ),
    .RESET_B(net2354),
    .D(_01478_),
    .Q_N(_08511_),
    .Q(\top1.memory2.mem1[4][0] ));
 sg13g2_dfrbp_1 _21382_ (.CLK(\clknet_leaf_36_top1.acquisition_clk ),
    .RESET_B(net2353),
    .D(_01479_),
    .Q_N(_08510_),
    .Q(\top1.memory2.mem1[4][1] ));
 sg13g2_dfrbp_1 _21383_ (.CLK(\clknet_leaf_266_top1.acquisition_clk ),
    .RESET_B(net2352),
    .D(_01480_),
    .Q_N(_08509_),
    .Q(\top1.memory2.mem1[4][2] ));
 sg13g2_dfrbp_1 _21384_ (.CLK(\clknet_leaf_163_top1.acquisition_clk ),
    .RESET_B(net2351),
    .D(_01481_),
    .Q_N(_08508_),
    .Q(\top1.memory2.mem1[50][0] ));
 sg13g2_dfrbp_1 _21385_ (.CLK(\clknet_leaf_165_top1.acquisition_clk ),
    .RESET_B(net2350),
    .D(_01482_),
    .Q_N(_08507_),
    .Q(\top1.memory2.mem1[50][1] ));
 sg13g2_dfrbp_1 _21386_ (.CLK(\clknet_leaf_164_top1.acquisition_clk ),
    .RESET_B(net2349),
    .D(_01483_),
    .Q_N(_08506_),
    .Q(\top1.memory2.mem1[50][2] ));
 sg13g2_dfrbp_1 _21387_ (.CLK(\clknet_leaf_164_top1.acquisition_clk ),
    .RESET_B(net2348),
    .D(_01484_),
    .Q_N(_08505_),
    .Q(\top1.memory2.mem1[51][0] ));
 sg13g2_dfrbp_1 _21388_ (.CLK(\clknet_leaf_165_top1.acquisition_clk ),
    .RESET_B(net2347),
    .D(_01485_),
    .Q_N(_08504_),
    .Q(\top1.memory2.mem1[51][1] ));
 sg13g2_dfrbp_1 _21389_ (.CLK(\clknet_leaf_164_top1.acquisition_clk ),
    .RESET_B(net2346),
    .D(_01486_),
    .Q_N(_08503_),
    .Q(\top1.memory2.mem1[51][2] ));
 sg13g2_dfrbp_1 _21390_ (.CLK(\clknet_leaf_199_top1.acquisition_clk ),
    .RESET_B(net2345),
    .D(_01487_),
    .Q_N(_08502_),
    .Q(\top1.memory2.mem1[52][0] ));
 sg13g2_dfrbp_1 _21391_ (.CLK(\clknet_leaf_199_top1.acquisition_clk ),
    .RESET_B(net2344),
    .D(_01488_),
    .Q_N(_08501_),
    .Q(\top1.memory2.mem1[52][1] ));
 sg13g2_dfrbp_1 _21392_ (.CLK(\clknet_leaf_166_top1.acquisition_clk ),
    .RESET_B(net2343),
    .D(_01489_),
    .Q_N(_08500_),
    .Q(\top1.memory2.mem1[52][2] ));
 sg13g2_dfrbp_1 _21393_ (.CLK(\clknet_leaf_199_top1.acquisition_clk ),
    .RESET_B(net2342),
    .D(_01490_),
    .Q_N(_08499_),
    .Q(\top1.memory2.mem1[53][0] ));
 sg13g2_dfrbp_1 _21394_ (.CLK(\clknet_leaf_199_top1.acquisition_clk ),
    .RESET_B(net2341),
    .D(_01491_),
    .Q_N(_08498_),
    .Q(\top1.memory2.mem1[53][1] ));
 sg13g2_dfrbp_1 _21395_ (.CLK(\clknet_leaf_167_top1.acquisition_clk ),
    .RESET_B(net2340),
    .D(_01492_),
    .Q_N(_08497_),
    .Q(\top1.memory2.mem1[53][2] ));
 sg13g2_dfrbp_1 _21396_ (.CLK(\clknet_leaf_200_top1.acquisition_clk ),
    .RESET_B(net2339),
    .D(_01493_),
    .Q_N(_08496_),
    .Q(\top1.memory2.mem1[54][0] ));
 sg13g2_dfrbp_1 _21397_ (.CLK(\clknet_leaf_169_top1.acquisition_clk ),
    .RESET_B(net2338),
    .D(_01494_),
    .Q_N(_08495_),
    .Q(\top1.memory2.mem1[54][1] ));
 sg13g2_dfrbp_1 _21398_ (.CLK(\clknet_leaf_166_top1.acquisition_clk ),
    .RESET_B(net2337),
    .D(_01495_),
    .Q_N(_08494_),
    .Q(\top1.memory2.mem1[54][2] ));
 sg13g2_dfrbp_1 _21399_ (.CLK(\clknet_leaf_199_top1.acquisition_clk ),
    .RESET_B(net2336),
    .D(_01496_),
    .Q_N(_08493_),
    .Q(\top1.memory2.mem1[55][0] ));
 sg13g2_dfrbp_1 _21400_ (.CLK(\clknet_leaf_199_top1.acquisition_clk ),
    .RESET_B(net2335),
    .D(_01497_),
    .Q_N(_08492_),
    .Q(\top1.memory2.mem1[55][1] ));
 sg13g2_dfrbp_1 _21401_ (.CLK(\clknet_leaf_167_top1.acquisition_clk ),
    .RESET_B(net2334),
    .D(_01498_),
    .Q_N(_08491_),
    .Q(\top1.memory2.mem1[55][2] ));
 sg13g2_dfrbp_1 _21402_ (.CLK(\clknet_leaf_168_top1.acquisition_clk ),
    .RESET_B(net2333),
    .D(_01499_),
    .Q_N(_08490_),
    .Q(\top1.memory2.mem1[56][0] ));
 sg13g2_dfrbp_1 _21403_ (.CLK(\clknet_leaf_168_top1.acquisition_clk ),
    .RESET_B(net2332),
    .D(_01500_),
    .Q_N(_08489_),
    .Q(\top1.memory2.mem1[56][1] ));
 sg13g2_dfrbp_1 _21404_ (.CLK(\clknet_leaf_168_top1.acquisition_clk ),
    .RESET_B(net2331),
    .D(_01501_),
    .Q_N(_08488_),
    .Q(\top1.memory2.mem1[56][2] ));
 sg13g2_dfrbp_1 _21405_ (.CLK(\clknet_leaf_168_top1.acquisition_clk ),
    .RESET_B(net2330),
    .D(_01502_),
    .Q_N(_08487_),
    .Q(\top1.memory2.mem1[57][0] ));
 sg13g2_dfrbp_1 _21406_ (.CLK(\clknet_leaf_168_top1.acquisition_clk ),
    .RESET_B(net2329),
    .D(_01503_),
    .Q_N(_08486_),
    .Q(\top1.memory2.mem1[57][1] ));
 sg13g2_dfrbp_1 _21407_ (.CLK(\clknet_leaf_162_top1.acquisition_clk ),
    .RESET_B(net2328),
    .D(_01504_),
    .Q_N(_08485_),
    .Q(\top1.memory2.mem1[57][2] ));
 sg13g2_dfrbp_1 _21408_ (.CLK(\clknet_leaf_169_top1.acquisition_clk ),
    .RESET_B(net2327),
    .D(_01505_),
    .Q_N(_08484_),
    .Q(\top1.memory2.mem1[58][0] ));
 sg13g2_dfrbp_1 _21409_ (.CLK(\clknet_leaf_169_top1.acquisition_clk ),
    .RESET_B(net2326),
    .D(_01506_),
    .Q_N(_08483_),
    .Q(\top1.memory2.mem1[58][1] ));
 sg13g2_dfrbp_1 _21410_ (.CLK(\clknet_leaf_167_top1.acquisition_clk ),
    .RESET_B(net2325),
    .D(_01507_),
    .Q_N(_08482_),
    .Q(\top1.memory2.mem1[58][2] ));
 sg13g2_dfrbp_1 _21411_ (.CLK(\clknet_leaf_262_top1.acquisition_clk ),
    .RESET_B(net2324),
    .D(_01508_),
    .Q_N(_08481_),
    .Q(\top1.memory2.mem1[5][0] ));
 sg13g2_dfrbp_1 _21412_ (.CLK(\clknet_leaf_36_top1.acquisition_clk ),
    .RESET_B(net2323),
    .D(_01509_),
    .Q_N(_08480_),
    .Q(\top1.memory2.mem1[5][1] ));
 sg13g2_dfrbp_1 _21413_ (.CLK(\clknet_leaf_262_top1.acquisition_clk ),
    .RESET_B(net2322),
    .D(_01510_),
    .Q_N(_08479_),
    .Q(\top1.memory2.mem1[5][2] ));
 sg13g2_dfrbp_1 _21414_ (.CLK(\clknet_leaf_203_top1.acquisition_clk ),
    .RESET_B(net2321),
    .D(_01511_),
    .Q_N(_08478_),
    .Q(\top1.memory2.mem1[60][0] ));
 sg13g2_dfrbp_1 _21415_ (.CLK(\clknet_leaf_203_top1.acquisition_clk ),
    .RESET_B(net2320),
    .D(_01512_),
    .Q_N(_08477_),
    .Q(\top1.memory2.mem1[60][1] ));
 sg13g2_dfrbp_1 _21416_ (.CLK(\clknet_leaf_202_top1.acquisition_clk ),
    .RESET_B(net2319),
    .D(_01513_),
    .Q_N(_08476_),
    .Q(\top1.memory2.mem1[60][2] ));
 sg13g2_dfrbp_1 _21417_ (.CLK(\clknet_leaf_204_top1.acquisition_clk ),
    .RESET_B(net2318),
    .D(_01514_),
    .Q_N(_08475_),
    .Q(\top1.memory2.mem1[61][0] ));
 sg13g2_dfrbp_1 _21418_ (.CLK(\clknet_leaf_202_top1.acquisition_clk ),
    .RESET_B(net2317),
    .D(_01515_),
    .Q_N(_08474_),
    .Q(\top1.memory2.mem1[61][1] ));
 sg13g2_dfrbp_1 _21419_ (.CLK(\clknet_leaf_202_top1.acquisition_clk ),
    .RESET_B(net2316),
    .D(_01516_),
    .Q_N(_08473_),
    .Q(\top1.memory2.mem1[61][2] ));
 sg13g2_dfrbp_1 _21420_ (.CLK(\clknet_leaf_203_top1.acquisition_clk ),
    .RESET_B(net2315),
    .D(_01517_),
    .Q_N(_08472_),
    .Q(\top1.memory2.mem1[62][0] ));
 sg13g2_dfrbp_1 _21421_ (.CLK(\clknet_leaf_203_top1.acquisition_clk ),
    .RESET_B(net2314),
    .D(_01518_),
    .Q_N(_08471_),
    .Q(\top1.memory2.mem1[62][1] ));
 sg13g2_dfrbp_1 _21422_ (.CLK(\clknet_leaf_202_top1.acquisition_clk ),
    .RESET_B(net2313),
    .D(_01519_),
    .Q_N(_08470_),
    .Q(\top1.memory2.mem1[62][2] ));
 sg13g2_dfrbp_1 _21423_ (.CLK(\clknet_leaf_203_top1.acquisition_clk ),
    .RESET_B(net2312),
    .D(_01520_),
    .Q_N(_08469_),
    .Q(\top1.memory2.mem1[63][0] ));
 sg13g2_dfrbp_1 _21424_ (.CLK(\clknet_leaf_203_top1.acquisition_clk ),
    .RESET_B(net2311),
    .D(_01521_),
    .Q_N(_08468_),
    .Q(\top1.memory2.mem1[63][1] ));
 sg13g2_dfrbp_1 _21425_ (.CLK(\clknet_leaf_202_top1.acquisition_clk ),
    .RESET_B(net2310),
    .D(_01522_),
    .Q_N(_08467_),
    .Q(\top1.memory2.mem1[63][2] ));
 sg13g2_dfrbp_1 _21426_ (.CLK(\clknet_leaf_4_top1.acquisition_clk ),
    .RESET_B(net2309),
    .D(_01523_),
    .Q_N(_08466_),
    .Q(\top1.memory2.mem1[64][0] ));
 sg13g2_dfrbp_1 _21427_ (.CLK(\clknet_leaf_2_top1.acquisition_clk ),
    .RESET_B(net2308),
    .D(_01524_),
    .Q_N(_08465_),
    .Q(\top1.memory2.mem1[64][1] ));
 sg13g2_dfrbp_1 _21428_ (.CLK(\clknet_leaf_4_top1.acquisition_clk ),
    .RESET_B(net2307),
    .D(_01525_),
    .Q_N(_08464_),
    .Q(\top1.memory2.mem1[64][2] ));
 sg13g2_dfrbp_1 _21429_ (.CLK(\clknet_leaf_4_top1.acquisition_clk ),
    .RESET_B(net2306),
    .D(_01526_),
    .Q_N(_08463_),
    .Q(\top1.memory2.mem1[65][0] ));
 sg13g2_dfrbp_1 _21430_ (.CLK(\clknet_leaf_2_top1.acquisition_clk ),
    .RESET_B(net2305),
    .D(_01527_),
    .Q_N(_08462_),
    .Q(\top1.memory2.mem1[65][1] ));
 sg13g2_dfrbp_1 _21431_ (.CLK(\clknet_leaf_4_top1.acquisition_clk ),
    .RESET_B(net2304),
    .D(_01528_),
    .Q_N(_08461_),
    .Q(\top1.memory2.mem1[65][2] ));
 sg13g2_dfrbp_1 _21432_ (.CLK(\clknet_leaf_13_top1.acquisition_clk ),
    .RESET_B(net2303),
    .D(_01529_),
    .Q_N(_08460_),
    .Q(\top1.memory2.mem1[66][0] ));
 sg13g2_dfrbp_1 _21433_ (.CLK(\clknet_leaf_2_top1.acquisition_clk ),
    .RESET_B(net2302),
    .D(_01530_),
    .Q_N(_08459_),
    .Q(\top1.memory2.mem1[66][1] ));
 sg13g2_dfrbp_1 _21434_ (.CLK(\clknet_leaf_13_top1.acquisition_clk ),
    .RESET_B(net2301),
    .D(_01531_),
    .Q_N(_08458_),
    .Q(\top1.memory2.mem1[66][2] ));
 sg13g2_dfrbp_1 _21435_ (.CLK(\clknet_leaf_5_top1.acquisition_clk ),
    .RESET_B(net2300),
    .D(_01532_),
    .Q_N(_08457_),
    .Q(\top1.memory2.mem1[67][0] ));
 sg13g2_dfrbp_1 _21436_ (.CLK(\clknet_leaf_2_top1.acquisition_clk ),
    .RESET_B(net2299),
    .D(_01533_),
    .Q_N(_08456_),
    .Q(\top1.memory2.mem1[67][1] ));
 sg13g2_dfrbp_1 _21437_ (.CLK(\clknet_leaf_4_top1.acquisition_clk ),
    .RESET_B(net2298),
    .D(_01534_),
    .Q_N(_08455_),
    .Q(\top1.memory2.mem1[67][2] ));
 sg13g2_dfrbp_1 _21438_ (.CLK(\clknet_leaf_21_top1.acquisition_clk ),
    .RESET_B(net2297),
    .D(_01535_),
    .Q_N(_08454_),
    .Q(\top1.memory2.mem1[68][0] ));
 sg13g2_dfrbp_1 _21439_ (.CLK(\clknet_leaf_26_top1.acquisition_clk ),
    .RESET_B(net2296),
    .D(_01536_),
    .Q_N(_08453_),
    .Q(\top1.memory2.mem1[68][1] ));
 sg13g2_dfrbp_1 _21440_ (.CLK(\clknet_leaf_11_top1.acquisition_clk ),
    .RESET_B(net2295),
    .D(_01537_),
    .Q_N(_08452_),
    .Q(\top1.memory2.mem1[68][2] ));
 sg13g2_dfrbp_1 _21441_ (.CLK(\clknet_leaf_262_top1.acquisition_clk ),
    .RESET_B(net2294),
    .D(_01538_),
    .Q_N(_08451_),
    .Q(\top1.memory2.mem1[6][0] ));
 sg13g2_dfrbp_1 _21442_ (.CLK(\clknet_leaf_262_top1.acquisition_clk ),
    .RESET_B(net2293),
    .D(_01539_),
    .Q_N(_08450_),
    .Q(\top1.memory2.mem1[6][1] ));
 sg13g2_dfrbp_1 _21443_ (.CLK(\clknet_leaf_262_top1.acquisition_clk ),
    .RESET_B(net2292),
    .D(_01540_),
    .Q_N(_08449_),
    .Q(\top1.memory2.mem1[6][2] ));
 sg13g2_dfrbp_1 _21444_ (.CLK(\clknet_leaf_20_top1.acquisition_clk ),
    .RESET_B(net2291),
    .D(_01541_),
    .Q_N(_08448_),
    .Q(\top1.memory2.mem1[70][0] ));
 sg13g2_dfrbp_1 _21445_ (.CLK(\clknet_leaf_26_top1.acquisition_clk ),
    .RESET_B(net2290),
    .D(_01542_),
    .Q_N(_08447_),
    .Q(\top1.memory2.mem1[70][1] ));
 sg13g2_dfrbp_1 _21446_ (.CLK(\clknet_leaf_16_top1.acquisition_clk ),
    .RESET_B(net2289),
    .D(_01543_),
    .Q_N(_08446_),
    .Q(\top1.memory2.mem1[70][2] ));
 sg13g2_dfrbp_1 _21447_ (.CLK(\clknet_leaf_20_top1.acquisition_clk ),
    .RESET_B(net2288),
    .D(_01544_),
    .Q_N(_08445_),
    .Q(\top1.memory2.mem1[71][0] ));
 sg13g2_dfrbp_1 _21448_ (.CLK(\clknet_leaf_25_top1.acquisition_clk ),
    .RESET_B(net2287),
    .D(_01545_),
    .Q_N(_08444_),
    .Q(\top1.memory2.mem1[71][1] ));
 sg13g2_dfrbp_1 _21449_ (.CLK(\clknet_leaf_11_top1.acquisition_clk ),
    .RESET_B(net2286),
    .D(_01546_),
    .Q_N(_08443_),
    .Q(\top1.memory2.mem1[71][2] ));
 sg13g2_dfrbp_1 _21450_ (.CLK(\clknet_leaf_16_top1.acquisition_clk ),
    .RESET_B(net2285),
    .D(_01547_),
    .Q_N(_08442_),
    .Q(\top1.memory2.mem1[72][0] ));
 sg13g2_dfrbp_1 _21451_ (.CLK(\clknet_leaf_15_top1.acquisition_clk ),
    .RESET_B(net2284),
    .D(_01548_),
    .Q_N(_08441_),
    .Q(\top1.memory2.mem1[72][1] ));
 sg13g2_dfrbp_1 _21452_ (.CLK(\clknet_leaf_11_top1.acquisition_clk ),
    .RESET_B(net2283),
    .D(_01549_),
    .Q_N(_08440_),
    .Q(\top1.memory2.mem1[72][2] ));
 sg13g2_dfrbp_1 _21453_ (.CLK(\clknet_leaf_16_top1.acquisition_clk ),
    .RESET_B(net2282),
    .D(_01550_),
    .Q_N(_08439_),
    .Q(\top1.memory2.mem1[73][0] ));
 sg13g2_dfrbp_1 _21454_ (.CLK(\clknet_leaf_16_top1.acquisition_clk ),
    .RESET_B(net2281),
    .D(_01551_),
    .Q_N(_08438_),
    .Q(\top1.memory2.mem1[73][1] ));
 sg13g2_dfrbp_1 _21455_ (.CLK(\clknet_leaf_11_top1.acquisition_clk ),
    .RESET_B(net2280),
    .D(_01552_),
    .Q_N(_08437_),
    .Q(\top1.memory2.mem1[73][2] ));
 sg13g2_dfrbp_1 _21456_ (.CLK(\clknet_leaf_16_top1.acquisition_clk ),
    .RESET_B(net2279),
    .D(_01553_),
    .Q_N(_08436_),
    .Q(\top1.memory2.mem1[74][0] ));
 sg13g2_dfrbp_1 _21457_ (.CLK(\clknet_leaf_15_top1.acquisition_clk ),
    .RESET_B(net2278),
    .D(_01554_),
    .Q_N(_08435_),
    .Q(\top1.memory2.mem1[74][1] ));
 sg13g2_dfrbp_1 _21458_ (.CLK(\clknet_leaf_15_top1.acquisition_clk ),
    .RESET_B(net2277),
    .D(_01555_),
    .Q_N(_08434_),
    .Q(\top1.memory2.mem1[74][2] ));
 sg13g2_dfrbp_1 _21459_ (.CLK(\clknet_leaf_16_top1.acquisition_clk ),
    .RESET_B(net2276),
    .D(_01556_),
    .Q_N(_08433_),
    .Q(\top1.memory2.mem1[75][0] ));
 sg13g2_dfrbp_1 _21460_ (.CLK(\clknet_leaf_16_top1.acquisition_clk ),
    .RESET_B(net2275),
    .D(_01557_),
    .Q_N(_08432_),
    .Q(\top1.memory2.mem1[75][1] ));
 sg13g2_dfrbp_1 _21461_ (.CLK(\clknet_leaf_11_top1.acquisition_clk ),
    .RESET_B(net2274),
    .D(_01558_),
    .Q_N(_08431_),
    .Q(\top1.memory2.mem1[75][2] ));
 sg13g2_dfrbp_1 _21462_ (.CLK(\clknet_leaf_17_top1.acquisition_clk ),
    .RESET_B(net2273),
    .D(_01559_),
    .Q_N(_08430_),
    .Q(\top1.memory2.mem1[76][0] ));
 sg13g2_dfrbp_1 _21463_ (.CLK(\clknet_leaf_14_top1.acquisition_clk ),
    .RESET_B(net2272),
    .D(_01560_),
    .Q_N(_08429_),
    .Q(\top1.memory2.mem1[76][1] ));
 sg13g2_dfrbp_1 _21464_ (.CLK(\clknet_leaf_12_top1.acquisition_clk ),
    .RESET_B(net2271),
    .D(_01561_),
    .Q_N(_08428_),
    .Q(\top1.memory2.mem1[76][2] ));
 sg13g2_dfrbp_1 _21465_ (.CLK(\clknet_leaf_17_top1.acquisition_clk ),
    .RESET_B(net2270),
    .D(_01562_),
    .Q_N(_08427_),
    .Q(\top1.memory2.mem1[77][0] ));
 sg13g2_dfrbp_1 _21466_ (.CLK(\clknet_leaf_14_top1.acquisition_clk ),
    .RESET_B(net2269),
    .D(_01563_),
    .Q_N(_08426_),
    .Q(\top1.memory2.mem1[77][1] ));
 sg13g2_dfrbp_1 _21467_ (.CLK(\clknet_leaf_14_top1.acquisition_clk ),
    .RESET_B(net2268),
    .D(_01564_),
    .Q_N(_08425_),
    .Q(\top1.memory2.mem1[77][2] ));
 sg13g2_dfrbp_1 _21468_ (.CLK(\clknet_leaf_17_top1.acquisition_clk ),
    .RESET_B(net2267),
    .D(_01565_),
    .Q_N(_08424_),
    .Q(\top1.memory2.mem1[78][0] ));
 sg13g2_dfrbp_1 _21469_ (.CLK(\clknet_leaf_14_top1.acquisition_clk ),
    .RESET_B(net2266),
    .D(_01566_),
    .Q_N(_08423_),
    .Q(\top1.memory2.mem1[78][1] ));
 sg13g2_dfrbp_1 _21470_ (.CLK(\clknet_leaf_14_top1.acquisition_clk ),
    .RESET_B(net2265),
    .D(_01567_),
    .Q_N(_08422_),
    .Q(\top1.memory2.mem1[78][2] ));
 sg13g2_dfrbp_1 _21471_ (.CLK(\clknet_leaf_263_top1.acquisition_clk ),
    .RESET_B(net2264),
    .D(_01568_),
    .Q_N(_08421_),
    .Q(\top1.memory2.mem1[7][0] ));
 sg13g2_dfrbp_1 _21472_ (.CLK(\clknet_leaf_36_top1.acquisition_clk ),
    .RESET_B(net2263),
    .D(_01569_),
    .Q_N(_08420_),
    .Q(\top1.memory2.mem1[7][1] ));
 sg13g2_dfrbp_1 _21473_ (.CLK(\clknet_leaf_36_top1.acquisition_clk ),
    .RESET_B(net2262),
    .D(_01570_),
    .Q_N(_08419_),
    .Q(\top1.memory2.mem1[7][2] ));
 sg13g2_dfrbp_1 _21474_ (.CLK(\clknet_leaf_287_top1.acquisition_clk ),
    .RESET_B(net2261),
    .D(_01571_),
    .Q_N(_08418_),
    .Q(\top1.memory2.mem1[80][0] ));
 sg13g2_dfrbp_1 _21475_ (.CLK(\clknet_leaf_284_top1.acquisition_clk ),
    .RESET_B(net2260),
    .D(_01572_),
    .Q_N(_08417_),
    .Q(\top1.memory2.mem1[80][1] ));
 sg13g2_dfrbp_1 _21476_ (.CLK(\clknet_leaf_284_top1.acquisition_clk ),
    .RESET_B(net2259),
    .D(_01573_),
    .Q_N(_08416_),
    .Q(\top1.memory2.mem1[80][2] ));
 sg13g2_dfrbp_1 _21477_ (.CLK(\clknet_leaf_287_top1.acquisition_clk ),
    .RESET_B(net2258),
    .D(_01574_),
    .Q_N(_08415_),
    .Q(\top1.memory2.mem1[81][0] ));
 sg13g2_dfrbp_1 _21478_ (.CLK(\clknet_leaf_284_top1.acquisition_clk ),
    .RESET_B(net2257),
    .D(_01575_),
    .Q_N(_08414_),
    .Q(\top1.memory2.mem1[81][1] ));
 sg13g2_dfrbp_1 _21479_ (.CLK(\clknet_leaf_286_top1.acquisition_clk ),
    .RESET_B(net2256),
    .D(_01576_),
    .Q_N(_08413_),
    .Q(\top1.memory2.mem1[81][2] ));
 sg13g2_dfrbp_1 _21480_ (.CLK(\clknet_leaf_290_top1.acquisition_clk ),
    .RESET_B(net2255),
    .D(_01577_),
    .Q_N(_08412_),
    .Q(\top1.memory2.mem1[82][0] ));
 sg13g2_dfrbp_1 _21481_ (.CLK(\clknet_leaf_284_top1.acquisition_clk ),
    .RESET_B(net2254),
    .D(_01578_),
    .Q_N(_08411_),
    .Q(\top1.memory2.mem1[82][1] ));
 sg13g2_dfrbp_1 _21482_ (.CLK(\clknet_leaf_285_top1.acquisition_clk ),
    .RESET_B(net2253),
    .D(_01579_),
    .Q_N(_08410_),
    .Q(\top1.memory2.mem1[82][2] ));
 sg13g2_dfrbp_1 _21483_ (.CLK(\clknet_leaf_289_top1.acquisition_clk ),
    .RESET_B(net2252),
    .D(_01580_),
    .Q_N(_08409_),
    .Q(\top1.memory2.mem1[83][0] ));
 sg13g2_dfrbp_1 _21484_ (.CLK(\clknet_leaf_284_top1.acquisition_clk ),
    .RESET_B(net2251),
    .D(_01581_),
    .Q_N(_08408_),
    .Q(\top1.memory2.mem1[83][1] ));
 sg13g2_dfrbp_1 _21485_ (.CLK(\clknet_leaf_285_top1.acquisition_clk ),
    .RESET_B(net2250),
    .D(_01582_),
    .Q_N(_08407_),
    .Q(\top1.memory2.mem1[83][2] ));
 sg13g2_dfrbp_1 _21486_ (.CLK(\clknet_leaf_30_top1.acquisition_clk ),
    .RESET_B(net2249),
    .D(_01583_),
    .Q_N(_08406_),
    .Q(\top1.memory2.mem1[84][0] ));
 sg13g2_dfrbp_1 _21487_ (.CLK(\clknet_leaf_29_top1.acquisition_clk ),
    .RESET_B(net2248),
    .D(_01584_),
    .Q_N(_08405_),
    .Q(\top1.memory2.mem1[84][1] ));
 sg13g2_dfrbp_1 _21488_ (.CLK(\clknet_leaf_269_top1.acquisition_clk ),
    .RESET_B(net2247),
    .D(_01585_),
    .Q_N(_08404_),
    .Q(\top1.memory2.mem1[84][2] ));
 sg13g2_dfrbp_1 _21489_ (.CLK(\clknet_leaf_30_top1.acquisition_clk ),
    .RESET_B(net2246),
    .D(_01586_),
    .Q_N(_08403_),
    .Q(\top1.memory2.mem1[85][0] ));
 sg13g2_dfrbp_1 _21490_ (.CLK(\clknet_leaf_29_top1.acquisition_clk ),
    .RESET_B(net2245),
    .D(_01587_),
    .Q_N(_08402_),
    .Q(\top1.memory2.mem1[85][1] ));
 sg13g2_dfrbp_1 _21491_ (.CLK(\clknet_leaf_269_top1.acquisition_clk ),
    .RESET_B(net2244),
    .D(_01588_),
    .Q_N(_08401_),
    .Q(\top1.memory2.mem1[85][2] ));
 sg13g2_dfrbp_1 _21492_ (.CLK(\clknet_leaf_30_top1.acquisition_clk ),
    .RESET_B(net2243),
    .D(_01589_),
    .Q_N(_08400_),
    .Q(\top1.memory2.mem1[86][0] ));
 sg13g2_dfrbp_1 _21493_ (.CLK(\clknet_leaf_29_top1.acquisition_clk ),
    .RESET_B(net2242),
    .D(_01590_),
    .Q_N(_08399_),
    .Q(\top1.memory2.mem1[86][1] ));
 sg13g2_dfrbp_1 _21494_ (.CLK(\clknet_leaf_269_top1.acquisition_clk ),
    .RESET_B(net2241),
    .D(_01591_),
    .Q_N(_08398_),
    .Q(\top1.memory2.mem1[86][2] ));
 sg13g2_dfrbp_1 _21495_ (.CLK(\clknet_leaf_30_top1.acquisition_clk ),
    .RESET_B(net2240),
    .D(_01592_),
    .Q_N(_08397_),
    .Q(\top1.memory2.mem1[87][0] ));
 sg13g2_dfrbp_1 _21496_ (.CLK(\clknet_leaf_29_top1.acquisition_clk ),
    .RESET_B(net2239),
    .D(_01593_),
    .Q_N(_08396_),
    .Q(\top1.memory2.mem1[87][1] ));
 sg13g2_dfrbp_1 _21497_ (.CLK(\clknet_leaf_269_top1.acquisition_clk ),
    .RESET_B(net2238),
    .D(_01594_),
    .Q_N(_08395_),
    .Q(\top1.memory2.mem1[87][2] ));
 sg13g2_dfrbp_1 _21498_ (.CLK(\clknet_leaf_270_top1.acquisition_clk ),
    .RESET_B(net2237),
    .D(_01595_),
    .Q_N(_08394_),
    .Q(\top1.memory2.mem1[88][0] ));
 sg13g2_dfrbp_1 _21499_ (.CLK(\clknet_leaf_287_top1.acquisition_clk ),
    .RESET_B(net2236),
    .D(_01596_),
    .Q_N(_08393_),
    .Q(\top1.memory2.mem1[88][1] ));
 sg13g2_dfrbp_1 _21500_ (.CLK(\clknet_leaf_288_top1.acquisition_clk ),
    .RESET_B(net2235),
    .D(_01597_),
    .Q_N(_08392_),
    .Q(\top1.memory2.mem1[88][2] ));
 sg13g2_dfrbp_1 _21501_ (.CLK(\clknet_leaf_266_top1.acquisition_clk ),
    .RESET_B(net2234),
    .D(_01598_),
    .Q_N(_08391_),
    .Q(\top1.memory2.mem1[8][0] ));
 sg13g2_dfrbp_1 _21502_ (.CLK(\clknet_leaf_272_top1.acquisition_clk ),
    .RESET_B(net2233),
    .D(_01599_),
    .Q_N(_08390_),
    .Q(\top1.memory2.mem1[8][1] ));
 sg13g2_dfrbp_1 _21503_ (.CLK(\clknet_leaf_273_top1.acquisition_clk ),
    .RESET_B(net2232),
    .D(_01600_),
    .Q_N(_08389_),
    .Q(\top1.memory2.mem1[8][2] ));
 sg13g2_dfrbp_1 _21504_ (.CLK(\clknet_leaf_270_top1.acquisition_clk ),
    .RESET_B(net2231),
    .D(_01601_),
    .Q_N(_08388_),
    .Q(\top1.memory2.mem1[90][0] ));
 sg13g2_dfrbp_1 _21505_ (.CLK(\clknet_leaf_283_top1.acquisition_clk ),
    .RESET_B(net2230),
    .D(_01602_),
    .Q_N(_08387_),
    .Q(\top1.memory2.mem1[90][1] ));
 sg13g2_dfrbp_1 _21506_ (.CLK(\clknet_leaf_288_top1.acquisition_clk ),
    .RESET_B(net2229),
    .D(_01603_),
    .Q_N(_08386_),
    .Q(\top1.memory2.mem1[90][2] ));
 sg13g2_dfrbp_1 _21507_ (.CLK(\clknet_leaf_268_top1.acquisition_clk ),
    .RESET_B(net2228),
    .D(_01604_),
    .Q_N(_08385_),
    .Q(\top1.memory2.mem1[91][0] ));
 sg13g2_dfrbp_1 _21508_ (.CLK(\clknet_leaf_287_top1.acquisition_clk ),
    .RESET_B(net2227),
    .D(_01605_),
    .Q_N(_08384_),
    .Q(\top1.memory2.mem1[91][1] ));
 sg13g2_dfrbp_1 _21509_ (.CLK(\clknet_leaf_271_top1.acquisition_clk ),
    .RESET_B(net2226),
    .D(_01606_),
    .Q_N(_08383_),
    .Q(\top1.memory2.mem1[91][2] ));
 sg13g2_dfrbp_1 _21510_ (.CLK(\clknet_leaf_270_top1.acquisition_clk ),
    .RESET_B(net2225),
    .D(_01607_),
    .Q_N(_08382_),
    .Q(\top1.memory2.mem1[92][0] ));
 sg13g2_dfrbp_1 _21511_ (.CLK(\clknet_leaf_283_top1.acquisition_clk ),
    .RESET_B(net2224),
    .D(_01608_),
    .Q_N(_08381_),
    .Q(\top1.memory2.mem1[92][1] ));
 sg13g2_dfrbp_1 _21512_ (.CLK(\clknet_leaf_288_top1.acquisition_clk ),
    .RESET_B(net2223),
    .D(_01609_),
    .Q_N(_08380_),
    .Q(\top1.memory2.mem1[92][2] ));
 sg13g2_dfrbp_1 _21513_ (.CLK(\clknet_leaf_271_top1.acquisition_clk ),
    .RESET_B(net2222),
    .D(_01610_),
    .Q_N(_08379_),
    .Q(\top1.memory2.mem1[93][0] ));
 sg13g2_dfrbp_1 _21514_ (.CLK(\clknet_leaf_282_top1.acquisition_clk ),
    .RESET_B(net2221),
    .D(_01611_),
    .Q_N(_08378_),
    .Q(\top1.memory2.mem1[93][1] ));
 sg13g2_dfrbp_1 _21515_ (.CLK(\clknet_leaf_271_top1.acquisition_clk ),
    .RESET_B(net2220),
    .D(_01612_),
    .Q_N(_08377_),
    .Q(\top1.memory2.mem1[93][2] ));
 sg13g2_dfrbp_1 _21516_ (.CLK(\clknet_leaf_268_top1.acquisition_clk ),
    .RESET_B(net2219),
    .D(_01613_),
    .Q_N(_08376_),
    .Q(\top1.memory2.mem1[94][0] ));
 sg13g2_dfrbp_1 _21517_ (.CLK(\clknet_leaf_283_top1.acquisition_clk ),
    .RESET_B(net2218),
    .D(_01614_),
    .Q_N(_08375_),
    .Q(\top1.memory2.mem1[94][1] ));
 sg13g2_dfrbp_1 _21518_ (.CLK(\clknet_leaf_271_top1.acquisition_clk ),
    .RESET_B(net2217),
    .D(_01615_),
    .Q_N(_08374_),
    .Q(\top1.memory2.mem1[94][2] ));
 sg13g2_dfrbp_1 _21519_ (.CLK(\clknet_leaf_271_top1.acquisition_clk ),
    .RESET_B(net2216),
    .D(_01616_),
    .Q_N(_08373_),
    .Q(\top1.memory2.mem1[95][0] ));
 sg13g2_dfrbp_1 _21520_ (.CLK(\clknet_leaf_282_top1.acquisition_clk ),
    .RESET_B(net2215),
    .D(_01617_),
    .Q_N(_08372_),
    .Q(\top1.memory2.mem1[95][1] ));
 sg13g2_dfrbp_1 _21521_ (.CLK(\clknet_leaf_271_top1.acquisition_clk ),
    .RESET_B(net2214),
    .D(_01618_),
    .Q_N(_08371_),
    .Q(\top1.memory2.mem1[95][2] ));
 sg13g2_dfrbp_1 _21522_ (.CLK(\clknet_leaf_188_top1.acquisition_clk ),
    .RESET_B(net2213),
    .D(_01619_),
    .Q_N(_08370_),
    .Q(\top1.memory2.mem1[96][0] ));
 sg13g2_dfrbp_1 _21523_ (.CLK(\clknet_leaf_189_top1.acquisition_clk ),
    .RESET_B(net2212),
    .D(_01620_),
    .Q_N(_08369_),
    .Q(\top1.memory2.mem1[96][1] ));
 sg13g2_dfrbp_1 _21524_ (.CLK(\clknet_leaf_179_top1.acquisition_clk ),
    .RESET_B(net2211),
    .D(_01621_),
    .Q_N(_08368_),
    .Q(\top1.memory2.mem1[96][2] ));
 sg13g2_dfrbp_1 _21525_ (.CLK(\clknet_leaf_188_top1.acquisition_clk ),
    .RESET_B(net2210),
    .D(_01622_),
    .Q_N(_08367_),
    .Q(\top1.memory2.mem1[97][0] ));
 sg13g2_dfrbp_1 _21526_ (.CLK(\clknet_leaf_189_top1.acquisition_clk ),
    .RESET_B(net2209),
    .D(_01623_),
    .Q_N(_08366_),
    .Q(\top1.memory2.mem1[97][1] ));
 sg13g2_dfrbp_1 _21527_ (.CLK(\clknet_leaf_179_top1.acquisition_clk ),
    .RESET_B(net2208),
    .D(_01624_),
    .Q_N(_08365_),
    .Q(\top1.memory2.mem1[97][2] ));
 sg13g2_dfrbp_1 _21528_ (.CLK(\clknet_leaf_189_top1.acquisition_clk ),
    .RESET_B(net2207),
    .D(_01625_),
    .Q_N(_08364_),
    .Q(\top1.memory2.mem1[98][0] ));
 sg13g2_dfrbp_1 _21529_ (.CLK(\clknet_leaf_190_top1.acquisition_clk ),
    .RESET_B(net2206),
    .D(_01626_),
    .Q_N(_08363_),
    .Q(\top1.memory2.mem1[98][1] ));
 sg13g2_dfrbp_1 _21530_ (.CLK(\clknet_leaf_180_top1.acquisition_clk ),
    .RESET_B(net2205),
    .D(_01627_),
    .Q_N(_08362_),
    .Q(\top1.memory2.mem1[98][2] ));
 sg13g2_dfrbp_1 _21531_ (.CLK(\clknet_leaf_282_top1.acquisition_clk ),
    .RESET_B(net2204),
    .D(_01628_),
    .Q_N(_08361_),
    .Q(\top1.memory2.mem1[0][0] ));
 sg13g2_dfrbp_1 _21532_ (.CLK(\clknet_leaf_280_top1.acquisition_clk ),
    .RESET_B(net2203),
    .D(_01629_),
    .Q_N(_08360_),
    .Q(\top1.memory2.mem1[0][1] ));
 sg13g2_dfrbp_1 _21533_ (.CLK(\clknet_leaf_280_top1.acquisition_clk ),
    .RESET_B(net2202),
    .D(_01630_),
    .Q_N(_08359_),
    .Q(\top1.memory2.mem1[0][2] ));
 sg13g2_dfrbp_1 _21534_ (.CLK(\clknet_leaf_193_top1.acquisition_clk ),
    .RESET_B(net2201),
    .D(_01631_),
    .Q_N(_08358_),
    .Q(\top1.memory2.mem1[100][0] ));
 sg13g2_dfrbp_1 _21535_ (.CLK(\clknet_leaf_193_top1.acquisition_clk ),
    .RESET_B(net2200),
    .D(_01632_),
    .Q_N(_08357_),
    .Q(\top1.memory2.mem1[100][1] ));
 sg13g2_dfrbp_1 _21536_ (.CLK(\clknet_leaf_189_top1.acquisition_clk ),
    .RESET_B(net2199),
    .D(_01633_),
    .Q_N(_08356_),
    .Q(\top1.memory2.mem1[100][2] ));
 sg13g2_dfrbp_1 _21537_ (.CLK(\clknet_leaf_192_top1.acquisition_clk ),
    .RESET_B(net2198),
    .D(_01634_),
    .Q_N(_08355_),
    .Q(\top1.memory2.mem1[101][0] ));
 sg13g2_dfrbp_1 _21538_ (.CLK(\clknet_leaf_193_top1.acquisition_clk ),
    .RESET_B(net2197),
    .D(_01635_),
    .Q_N(_08354_),
    .Q(\top1.memory2.mem1[101][1] ));
 sg13g2_dfrbp_1 _21539_ (.CLK(\clknet_leaf_190_top1.acquisition_clk ),
    .RESET_B(net2196),
    .D(_01636_),
    .Q_N(_08353_),
    .Q(\top1.memory2.mem1[101][2] ));
 sg13g2_dfrbp_1 _21540_ (.CLK(\clknet_leaf_192_top1.acquisition_clk ),
    .RESET_B(net2195),
    .D(_01637_),
    .Q_N(_08352_),
    .Q(\top1.memory2.mem1[102][0] ));
 sg13g2_dfrbp_1 _21541_ (.CLK(\clknet_leaf_191_top1.acquisition_clk ),
    .RESET_B(net2194),
    .D(_01638_),
    .Q_N(_08351_),
    .Q(\top1.memory2.mem1[102][1] ));
 sg13g2_dfrbp_1 _21542_ (.CLK(\clknet_leaf_197_top1.acquisition_clk ),
    .RESET_B(net2193),
    .D(_01639_),
    .Q_N(_08350_),
    .Q(\top1.memory2.mem1[102][2] ));
 sg13g2_dfrbp_1 _21543_ (.CLK(\clknet_leaf_192_top1.acquisition_clk ),
    .RESET_B(net2192),
    .D(_01640_),
    .Q_N(_08349_),
    .Q(\top1.memory2.mem1[103][0] ));
 sg13g2_dfrbp_1 _21544_ (.CLK(\clknet_leaf_193_top1.acquisition_clk ),
    .RESET_B(net2191),
    .D(_01641_),
    .Q_N(_08348_),
    .Q(\top1.memory2.mem1[103][1] ));
 sg13g2_dfrbp_1 _21545_ (.CLK(\clknet_leaf_197_top1.acquisition_clk ),
    .RESET_B(net2190),
    .D(_01642_),
    .Q_N(_08347_),
    .Q(\top1.memory2.mem1[103][2] ));
 sg13g2_dfrbp_1 _21546_ (.CLK(\clknet_leaf_170_top1.acquisition_clk ),
    .RESET_B(net2189),
    .D(_01643_),
    .Q_N(_08346_),
    .Q(\top1.memory2.mem1[104][0] ));
 sg13g2_dfrbp_1 _21547_ (.CLK(\clknet_leaf_172_top1.acquisition_clk ),
    .RESET_B(net2188),
    .D(_01644_),
    .Q_N(_08345_),
    .Q(\top1.memory2.mem1[104][1] ));
 sg13g2_dfrbp_1 _21548_ (.CLK(\clknet_leaf_170_top1.acquisition_clk ),
    .RESET_B(net2187),
    .D(_01645_),
    .Q_N(_08344_),
    .Q(\top1.memory2.mem1[104][2] ));
 sg13g2_dfrbp_1 _21549_ (.CLK(\clknet_leaf_169_top1.acquisition_clk ),
    .RESET_B(net2186),
    .D(_01646_),
    .Q_N(_08343_),
    .Q(\top1.memory2.mem1[105][0] ));
 sg13g2_dfrbp_1 _21550_ (.CLK(\clknet_leaf_172_top1.acquisition_clk ),
    .RESET_B(net2185),
    .D(_01647_),
    .Q_N(_08342_),
    .Q(\top1.memory2.mem1[105][1] ));
 sg13g2_dfrbp_1 _21551_ (.CLK(\clknet_leaf_170_top1.acquisition_clk ),
    .RESET_B(net2184),
    .D(_01648_),
    .Q_N(_08341_),
    .Q(\top1.memory2.mem1[105][2] ));
 sg13g2_dfrbp_1 _21552_ (.CLK(\clknet_leaf_169_top1.acquisition_clk ),
    .RESET_B(net2183),
    .D(_01649_),
    .Q_N(_08340_),
    .Q(\top1.memory2.mem1[106][0] ));
 sg13g2_dfrbp_1 _21553_ (.CLK(\clknet_leaf_172_top1.acquisition_clk ),
    .RESET_B(net2182),
    .D(_01650_),
    .Q_N(_08339_),
    .Q(\top1.memory2.mem1[106][1] ));
 sg13g2_dfrbp_1 _21554_ (.CLK(\clknet_leaf_170_top1.acquisition_clk ),
    .RESET_B(net2181),
    .D(_01651_),
    .Q_N(_08338_),
    .Q(\top1.memory2.mem1[106][2] ));
 sg13g2_dfrbp_1 _21555_ (.CLK(\clknet_leaf_169_top1.acquisition_clk ),
    .RESET_B(net2180),
    .D(_01652_),
    .Q_N(_08337_),
    .Q(\top1.memory2.mem1[107][0] ));
 sg13g2_dfrbp_1 _21556_ (.CLK(\clknet_leaf_171_top1.acquisition_clk ),
    .RESET_B(net2179),
    .D(_01653_),
    .Q_N(_08336_),
    .Q(\top1.memory2.mem1[107][1] ));
 sg13g2_dfrbp_1 _21557_ (.CLK(\clknet_leaf_170_top1.acquisition_clk ),
    .RESET_B(net2178),
    .D(_01654_),
    .Q_N(_08335_),
    .Q(\top1.memory2.mem1[107][2] ));
 sg13g2_dfrbp_1 _21558_ (.CLK(\clknet_leaf_196_top1.acquisition_clk ),
    .RESET_B(net2177),
    .D(_01655_),
    .Q_N(_08334_),
    .Q(\top1.memory2.mem1[108][0] ));
 sg13g2_dfrbp_1 _21559_ (.CLK(\clknet_leaf_196_top1.acquisition_clk ),
    .RESET_B(net2176),
    .D(_01656_),
    .Q_N(_08333_),
    .Q(\top1.memory2.mem1[108][1] ));
 sg13g2_dfrbp_1 _21560_ (.CLK(\clknet_leaf_198_top1.acquisition_clk ),
    .RESET_B(net2175),
    .D(_01657_),
    .Q_N(_08332_),
    .Q(\top1.memory2.mem1[108][2] ));
 sg13g2_dfrbp_1 _21561_ (.CLK(\clknet_leaf_266_top1.acquisition_clk ),
    .RESET_B(net2174),
    .D(_01658_),
    .Q_N(_08331_),
    .Q(\top1.memory2.mem1[10][0] ));
 sg13g2_dfrbp_1 _21562_ (.CLK(\clknet_leaf_272_top1.acquisition_clk ),
    .RESET_B(net2173),
    .D(_01659_),
    .Q_N(_08330_),
    .Q(\top1.memory2.mem1[10][1] ));
 sg13g2_dfrbp_1 _21563_ (.CLK(\clknet_leaf_273_top1.acquisition_clk ),
    .RESET_B(net2172),
    .D(_01660_),
    .Q_N(_08329_),
    .Q(\top1.memory2.mem1[10][2] ));
 sg13g2_dfrbp_1 _21564_ (.CLK(\clknet_leaf_198_top1.acquisition_clk ),
    .RESET_B(net2171),
    .D(_01661_),
    .Q_N(_08328_),
    .Q(\top1.memory2.mem1[110][0] ));
 sg13g2_dfrbp_1 _21565_ (.CLK(\clknet_leaf_196_top1.acquisition_clk ),
    .RESET_B(net2170),
    .D(_01662_),
    .Q_N(_08327_),
    .Q(\top1.memory2.mem1[110][1] ));
 sg13g2_dfrbp_1 _21566_ (.CLK(\clknet_leaf_198_top1.acquisition_clk ),
    .RESET_B(net2169),
    .D(_01663_),
    .Q_N(_08326_),
    .Q(\top1.memory2.mem1[110][2] ));
 sg13g2_dfrbp_1 _21567_ (.CLK(\clknet_leaf_199_top1.acquisition_clk ),
    .RESET_B(net2168),
    .D(_01664_),
    .Q_N(_08325_),
    .Q(\top1.memory2.mem1[111][0] ));
 sg13g2_dfrbp_1 _21568_ (.CLK(\clknet_leaf_197_top1.acquisition_clk ),
    .RESET_B(net2167),
    .D(_01665_),
    .Q_N(_08324_),
    .Q(\top1.memory2.mem1[111][1] ));
 sg13g2_dfrbp_1 _21569_ (.CLK(\clknet_leaf_198_top1.acquisition_clk ),
    .RESET_B(net2166),
    .D(_01666_),
    .Q_N(_08323_),
    .Q(\top1.memory2.mem1[111][2] ));
 sg13g2_dfrbp_1 _21570_ (.CLK(\clknet_leaf_216_top1.acquisition_clk ),
    .RESET_B(net2165),
    .D(_01667_),
    .Q_N(_08322_),
    .Q(\top1.memory2.mem1[112][0] ));
 sg13g2_dfrbp_1 _21571_ (.CLK(\clknet_leaf_206_top1.acquisition_clk ),
    .RESET_B(net2164),
    .D(_01668_),
    .Q_N(_08321_),
    .Q(\top1.memory2.mem1[112][1] ));
 sg13g2_dfrbp_1 _21572_ (.CLK(\clknet_leaf_216_top1.acquisition_clk ),
    .RESET_B(net2163),
    .D(_01669_),
    .Q_N(_08320_),
    .Q(\top1.memory2.mem1[112][2] ));
 sg13g2_dfrbp_1 _21573_ (.CLK(\clknet_leaf_207_top1.acquisition_clk ),
    .RESET_B(net2162),
    .D(_01670_),
    .Q_N(_08319_),
    .Q(\top1.memory2.mem1[113][0] ));
 sg13g2_dfrbp_1 _21574_ (.CLK(\clknet_leaf_206_top1.acquisition_clk ),
    .RESET_B(net2161),
    .D(_01671_),
    .Q_N(_08318_),
    .Q(\top1.memory2.mem1[113][1] ));
 sg13g2_dfrbp_1 _21575_ (.CLK(\clknet_leaf_216_top1.acquisition_clk ),
    .RESET_B(net2160),
    .D(_01672_),
    .Q_N(_08317_),
    .Q(\top1.memory2.mem1[113][2] ));
 sg13g2_dfrbp_1 _21576_ (.CLK(\clknet_leaf_216_top1.acquisition_clk ),
    .RESET_B(net2159),
    .D(_01673_),
    .Q_N(_08316_),
    .Q(\top1.memory2.mem1[114][0] ));
 sg13g2_dfrbp_1 _21577_ (.CLK(\clknet_leaf_206_top1.acquisition_clk ),
    .RESET_B(net2158),
    .D(_01674_),
    .Q_N(_08315_),
    .Q(\top1.memory2.mem1[114][1] ));
 sg13g2_dfrbp_1 _21578_ (.CLK(\clknet_leaf_216_top1.acquisition_clk ),
    .RESET_B(net2157),
    .D(_01675_),
    .Q_N(_08314_),
    .Q(\top1.memory2.mem1[114][2] ));
 sg13g2_dfrbp_1 _21579_ (.CLK(\clknet_leaf_207_top1.acquisition_clk ),
    .RESET_B(net2156),
    .D(_01676_),
    .Q_N(_08313_),
    .Q(\top1.memory2.mem1[115][0] ));
 sg13g2_dfrbp_1 _21580_ (.CLK(\clknet_leaf_206_top1.acquisition_clk ),
    .RESET_B(net2155),
    .D(_01677_),
    .Q_N(_08312_),
    .Q(\top1.memory2.mem1[115][1] ));
 sg13g2_dfrbp_1 _21581_ (.CLK(\clknet_leaf_216_top1.acquisition_clk ),
    .RESET_B(net2154),
    .D(_01678_),
    .Q_N(_08311_),
    .Q(\top1.memory2.mem1[115][2] ));
 sg13g2_dfrbp_1 _21582_ (.CLK(\clknet_leaf_221_top1.acquisition_clk ),
    .RESET_B(net2153),
    .D(_01679_),
    .Q_N(_08310_),
    .Q(\top1.memory2.mem1[116][0] ));
 sg13g2_dfrbp_1 _21583_ (.CLK(\clknet_leaf_219_top1.acquisition_clk ),
    .RESET_B(net2152),
    .D(_01680_),
    .Q_N(_08309_),
    .Q(\top1.memory2.mem1[116][1] ));
 sg13g2_dfrbp_1 _21584_ (.CLK(\clknet_leaf_218_top1.acquisition_clk ),
    .RESET_B(net2151),
    .D(_01681_),
    .Q_N(_08308_),
    .Q(\top1.memory2.mem1[116][2] ));
 sg13g2_dfrbp_1 _21585_ (.CLK(\clknet_leaf_221_top1.acquisition_clk ),
    .RESET_B(net2150),
    .D(_01682_),
    .Q_N(_08307_),
    .Q(\top1.memory2.mem1[117][0] ));
 sg13g2_dfrbp_1 _21586_ (.CLK(\clknet_leaf_217_top1.acquisition_clk ),
    .RESET_B(net2149),
    .D(_01683_),
    .Q_N(_08306_),
    .Q(\top1.memory2.mem1[117][1] ));
 sg13g2_dfrbp_1 _21587_ (.CLK(\clknet_leaf_218_top1.acquisition_clk ),
    .RESET_B(net2148),
    .D(_01684_),
    .Q_N(_08305_),
    .Q(\top1.memory2.mem1[117][2] ));
 sg13g2_dfrbp_1 _21588_ (.CLK(\clknet_leaf_219_top1.acquisition_clk ),
    .RESET_B(net2147),
    .D(_01685_),
    .Q_N(_08304_),
    .Q(\top1.memory2.mem1[118][0] ));
 sg13g2_dfrbp_1 _21589_ (.CLK(\clknet_leaf_219_top1.acquisition_clk ),
    .RESET_B(net2146),
    .D(_01686_),
    .Q_N(_08303_),
    .Q(\top1.memory2.mem1[118][1] ));
 sg13g2_dfrbp_1 _21590_ (.CLK(\clknet_leaf_218_top1.acquisition_clk ),
    .RESET_B(net2145),
    .D(_01687_),
    .Q_N(_08302_),
    .Q(\top1.memory2.mem1[118][2] ));
 sg13g2_dfrbp_1 _21591_ (.CLK(\clknet_leaf_273_top1.acquisition_clk ),
    .RESET_B(net2144),
    .D(_01688_),
    .Q_N(_08301_),
    .Q(\top1.memory2.mem1[11][0] ));
 sg13g2_dfrbp_1 _21592_ (.CLK(\clknet_leaf_272_top1.acquisition_clk ),
    .RESET_B(net2143),
    .D(_01689_),
    .Q_N(_08300_),
    .Q(\top1.memory2.mem1[11][1] ));
 sg13g2_dfrbp_1 _21593_ (.CLK(\clknet_leaf_274_top1.acquisition_clk ),
    .RESET_B(net2142),
    .D(_01690_),
    .Q_N(_08299_),
    .Q(\top1.memory2.mem1[11][2] ));
 sg13g2_dfrbp_1 _21594_ (.CLK(\clknet_leaf_220_top1.acquisition_clk ),
    .RESET_B(net2141),
    .D(_01691_),
    .Q_N(_08298_),
    .Q(\top1.memory2.mem1[120][0] ));
 sg13g2_dfrbp_1 _21595_ (.CLK(\clknet_leaf_214_top1.acquisition_clk ),
    .RESET_B(net2140),
    .D(_01692_),
    .Q_N(_08297_),
    .Q(\top1.memory2.mem1[120][1] ));
 sg13g2_dfrbp_1 _21596_ (.CLK(\clknet_leaf_221_top1.acquisition_clk ),
    .RESET_B(net2139),
    .D(_01693_),
    .Q_N(_08296_),
    .Q(\top1.memory2.mem1[120][2] ));
 sg13g2_dfrbp_1 _21597_ (.CLK(\clknet_leaf_220_top1.acquisition_clk ),
    .RESET_B(net2138),
    .D(_01694_),
    .Q_N(_08295_),
    .Q(\top1.memory2.mem1[121][0] ));
 sg13g2_dfrbp_1 _21598_ (.CLK(\clknet_leaf_214_top1.acquisition_clk ),
    .RESET_B(net2137),
    .D(_01695_),
    .Q_N(_08294_),
    .Q(\top1.memory2.mem1[121][1] ));
 sg13g2_dfrbp_1 _21599_ (.CLK(\clknet_leaf_221_top1.acquisition_clk ),
    .RESET_B(net2136),
    .D(_01696_),
    .Q_N(_08293_),
    .Q(\top1.memory2.mem1[121][2] ));
 sg13g2_dfrbp_1 _21600_ (.CLK(\clknet_leaf_220_top1.acquisition_clk ),
    .RESET_B(net2135),
    .D(_01697_),
    .Q_N(_08292_),
    .Q(\top1.memory2.mem1[122][0] ));
 sg13g2_dfrbp_1 _21601_ (.CLK(\clknet_leaf_214_top1.acquisition_clk ),
    .RESET_B(net2134),
    .D(_01698_),
    .Q_N(_08291_),
    .Q(\top1.memory2.mem1[122][1] ));
 sg13g2_dfrbp_1 _21602_ (.CLK(\clknet_leaf_218_top1.acquisition_clk ),
    .RESET_B(net2133),
    .D(_01699_),
    .Q_N(_08290_),
    .Q(\top1.memory2.mem1[122][2] ));
 sg13g2_dfrbp_1 _21603_ (.CLK(\clknet_leaf_220_top1.acquisition_clk ),
    .RESET_B(net2132),
    .D(_01700_),
    .Q_N(_08289_),
    .Q(\top1.memory2.mem1[123][0] ));
 sg13g2_dfrbp_1 _21604_ (.CLK(\clknet_leaf_214_top1.acquisition_clk ),
    .RESET_B(net2131),
    .D(_01701_),
    .Q_N(_08288_),
    .Q(\top1.memory2.mem1[123][1] ));
 sg13g2_dfrbp_1 _21605_ (.CLK(\clknet_leaf_218_top1.acquisition_clk ),
    .RESET_B(net2130),
    .D(_01702_),
    .Q_N(_08287_),
    .Q(\top1.memory2.mem1[123][2] ));
 sg13g2_dfrbp_1 _21606_ (.CLK(\clknet_leaf_215_top1.acquisition_clk ),
    .RESET_B(net2129),
    .D(_01703_),
    .Q_N(_08286_),
    .Q(\top1.memory2.mem1[124][0] ));
 sg13g2_dfrbp_1 _21607_ (.CLK(\clknet_leaf_208_top1.acquisition_clk ),
    .RESET_B(net2128),
    .D(_01704_),
    .Q_N(_08285_),
    .Q(\top1.memory2.mem1[124][1] ));
 sg13g2_dfrbp_1 _21608_ (.CLK(\clknet_leaf_204_top1.acquisition_clk ),
    .RESET_B(net2127),
    .D(_01705_),
    .Q_N(_08284_),
    .Q(\top1.memory2.mem1[124][2] ));
 sg13g2_dfrbp_1 _21609_ (.CLK(\clknet_leaf_215_top1.acquisition_clk ),
    .RESET_B(net2126),
    .D(_01706_),
    .Q_N(_08283_),
    .Q(\top1.memory2.mem1[125][0] ));
 sg13g2_dfrbp_1 _21610_ (.CLK(\clknet_leaf_208_top1.acquisition_clk ),
    .RESET_B(net2125),
    .D(_01707_),
    .Q_N(_08282_),
    .Q(\top1.memory2.mem1[125][1] ));
 sg13g2_dfrbp_1 _21611_ (.CLK(\clknet_leaf_205_top1.acquisition_clk ),
    .RESET_B(net2124),
    .D(_01708_),
    .Q_N(_08281_),
    .Q(\top1.memory2.mem1[125][2] ));
 sg13g2_dfrbp_1 _21612_ (.CLK(\clknet_leaf_207_top1.acquisition_clk ),
    .RESET_B(net2123),
    .D(_01709_),
    .Q_N(_08280_),
    .Q(\top1.memory2.mem1[126][0] ));
 sg13g2_dfrbp_1 _21613_ (.CLK(\clknet_leaf_208_top1.acquisition_clk ),
    .RESET_B(net2122),
    .D(_01710_),
    .Q_N(_08279_),
    .Q(\top1.memory2.mem1[126][1] ));
 sg13g2_dfrbp_1 _21614_ (.CLK(\clknet_leaf_200_top1.acquisition_clk ),
    .RESET_B(net2121),
    .D(_01711_),
    .Q_N(_08278_),
    .Q(\top1.memory2.mem1[126][2] ));
 sg13g2_dfrbp_1 _21615_ (.CLK(\clknet_leaf_207_top1.acquisition_clk ),
    .RESET_B(net2120),
    .D(_01712_),
    .Q_N(_08277_),
    .Q(\top1.memory2.mem1[127][0] ));
 sg13g2_dfrbp_1 _21616_ (.CLK(\clknet_leaf_208_top1.acquisition_clk ),
    .RESET_B(net2119),
    .D(_01713_),
    .Q_N(_08276_),
    .Q(\top1.memory2.mem1[127][1] ));
 sg13g2_dfrbp_1 _21617_ (.CLK(\clknet_leaf_209_top1.acquisition_clk ),
    .RESET_B(net2118),
    .D(_01714_),
    .Q_N(_08275_),
    .Q(\top1.memory2.mem1[127][2] ));
 sg13g2_dfrbp_1 _21618_ (.CLK(\clknet_leaf_17_top1.acquisition_clk ),
    .RESET_B(net2117),
    .D(_01715_),
    .Q_N(_08274_),
    .Q(\top1.memory2.mem1[128][0] ));
 sg13g2_dfrbp_1 _21619_ (.CLK(\clknet_leaf_18_top1.acquisition_clk ),
    .RESET_B(net2116),
    .D(_01716_),
    .Q_N(_08273_),
    .Q(\top1.memory2.mem1[128][1] ));
 sg13g2_dfrbp_1 _21620_ (.CLK(\clknet_leaf_18_top1.acquisition_clk ),
    .RESET_B(net2115),
    .D(_01717_),
    .Q_N(_08272_),
    .Q(\top1.memory2.mem1[128][2] ));
 sg13g2_dfrbp_1 _21621_ (.CLK(\clknet_leaf_273_top1.acquisition_clk ),
    .RESET_B(net2114),
    .D(_01718_),
    .Q_N(_08271_),
    .Q(\top1.memory2.mem1[12][0] ));
 sg13g2_dfrbp_1 _21622_ (.CLK(\clknet_leaf_276_top1.acquisition_clk ),
    .RESET_B(net2113),
    .D(_01719_),
    .Q_N(_08270_),
    .Q(\top1.memory2.mem1[12][1] ));
 sg13g2_dfrbp_1 _21623_ (.CLK(\clknet_leaf_276_top1.acquisition_clk ),
    .RESET_B(net2112),
    .D(_01720_),
    .Q_N(_08269_),
    .Q(\top1.memory2.mem1[12][2] ));
 sg13g2_dfrbp_1 _21624_ (.CLK(\clknet_leaf_17_top1.acquisition_clk ),
    .RESET_B(net2111),
    .D(_01721_),
    .Q_N(_08268_),
    .Q(\top1.memory2.mem1[130][0] ));
 sg13g2_dfrbp_1 _21625_ (.CLK(\clknet_leaf_18_top1.acquisition_clk ),
    .RESET_B(net2110),
    .D(_01722_),
    .Q_N(_08267_),
    .Q(\top1.memory2.mem1[130][1] ));
 sg13g2_dfrbp_1 _21626_ (.CLK(\clknet_leaf_18_top1.acquisition_clk ),
    .RESET_B(net2109),
    .D(_01723_),
    .Q_N(_08266_),
    .Q(\top1.memory2.mem1[130][2] ));
 sg13g2_dfrbp_1 _21627_ (.CLK(\clknet_leaf_17_top1.acquisition_clk ),
    .RESET_B(net2108),
    .D(_01724_),
    .Q_N(_08265_),
    .Q(\top1.memory2.mem1[131][0] ));
 sg13g2_dfrbp_1 _21628_ (.CLK(\clknet_leaf_19_top1.acquisition_clk ),
    .RESET_B(net2107),
    .D(_01725_),
    .Q_N(_08264_),
    .Q(\top1.memory2.mem1[131][1] ));
 sg13g2_dfrbp_1 _21629_ (.CLK(\clknet_leaf_19_top1.acquisition_clk ),
    .RESET_B(net2106),
    .D(_01726_),
    .Q_N(_08263_),
    .Q(\top1.memory2.mem1[131][2] ));
 sg13g2_dfrbp_1 _21630_ (.CLK(\clknet_leaf_22_top1.acquisition_clk ),
    .RESET_B(net2105),
    .D(_01727_),
    .Q_N(_08262_),
    .Q(\top1.memory2.mem1[132][0] ));
 sg13g2_dfrbp_1 _21631_ (.CLK(\clknet_leaf_22_top1.acquisition_clk ),
    .RESET_B(net2104),
    .D(_01728_),
    .Q_N(_08261_),
    .Q(\top1.memory2.mem1[132][1] ));
 sg13g2_dfrbp_1 _21632_ (.CLK(\clknet_leaf_56_top1.acquisition_clk ),
    .RESET_B(net2103),
    .D(_01729_),
    .Q_N(_08260_),
    .Q(\top1.memory2.mem1[132][2] ));
 sg13g2_dfrbp_1 _21633_ (.CLK(\clknet_leaf_23_top1.acquisition_clk ),
    .RESET_B(net2102),
    .D(_01730_),
    .Q_N(_08259_),
    .Q(\top1.memory2.mem1[133][0] ));
 sg13g2_dfrbp_1 _21634_ (.CLK(\clknet_leaf_48_top1.acquisition_clk ),
    .RESET_B(net2101),
    .D(_01731_),
    .Q_N(_08258_),
    .Q(\top1.memory2.mem1[133][1] ));
 sg13g2_dfrbp_1 _21635_ (.CLK(\clknet_leaf_57_top1.acquisition_clk ),
    .RESET_B(net2100),
    .D(_01732_),
    .Q_N(_08257_),
    .Q(\top1.memory2.mem1[133][2] ));
 sg13g2_dfrbp_1 _21636_ (.CLK(\clknet_leaf_48_top1.acquisition_clk ),
    .RESET_B(net2099),
    .D(_01733_),
    .Q_N(_08256_),
    .Q(\top1.memory2.mem1[134][0] ));
 sg13g2_dfrbp_1 _21637_ (.CLK(\clknet_leaf_49_top1.acquisition_clk ),
    .RESET_B(net2098),
    .D(_01734_),
    .Q_N(_08255_),
    .Q(\top1.memory2.mem1[134][1] ));
 sg13g2_dfrbp_1 _21638_ (.CLK(\clknet_leaf_44_top1.acquisition_clk ),
    .RESET_B(net2097),
    .D(_01735_),
    .Q_N(_08254_),
    .Q(\top1.memory2.mem1[134][2] ));
 sg13g2_dfrbp_1 _21639_ (.CLK(\clknet_leaf_49_top1.acquisition_clk ),
    .RESET_B(net2096),
    .D(_01736_),
    .Q_N(_08253_),
    .Q(\top1.memory2.mem1[135][0] ));
 sg13g2_dfrbp_1 _21640_ (.CLK(\clknet_leaf_49_top1.acquisition_clk ),
    .RESET_B(net2095),
    .D(_01737_),
    .Q_N(_08252_),
    .Q(\top1.memory2.mem1[135][1] ));
 sg13g2_dfrbp_1 _21641_ (.CLK(\clknet_leaf_57_top1.acquisition_clk ),
    .RESET_B(net2094),
    .D(_01738_),
    .Q_N(_08251_),
    .Q(\top1.memory2.mem1[135][2] ));
 sg13g2_dfrbp_1 _21642_ (.CLK(\clknet_leaf_53_top1.acquisition_clk ),
    .RESET_B(net2093),
    .D(_01739_),
    .Q_N(_08250_),
    .Q(\top1.memory2.mem1[136][0] ));
 sg13g2_dfrbp_1 _21643_ (.CLK(\clknet_leaf_20_top1.acquisition_clk ),
    .RESET_B(net2092),
    .D(_01740_),
    .Q_N(_08249_),
    .Q(\top1.memory2.mem1[136][1] ));
 sg13g2_dfrbp_1 _21644_ (.CLK(\clknet_leaf_53_top1.acquisition_clk ),
    .RESET_B(net2091),
    .D(_01741_),
    .Q_N(_08248_),
    .Q(\top1.memory2.mem1[136][2] ));
 sg13g2_dfrbp_1 _21645_ (.CLK(\clknet_leaf_53_top1.acquisition_clk ),
    .RESET_B(net2090),
    .D(_01742_),
    .Q_N(_08247_),
    .Q(\top1.memory2.mem1[137][0] ));
 sg13g2_dfrbp_1 _21646_ (.CLK(\clknet_leaf_20_top1.acquisition_clk ),
    .RESET_B(net2089),
    .D(_01743_),
    .Q_N(_08246_),
    .Q(\top1.memory2.mem1[137][1] ));
 sg13g2_dfrbp_1 _21647_ (.CLK(\clknet_leaf_53_top1.acquisition_clk ),
    .RESET_B(net2088),
    .D(_01744_),
    .Q_N(_08245_),
    .Q(\top1.memory2.mem1[137][2] ));
 sg13g2_dfrbp_1 _21648_ (.CLK(\clknet_leaf_56_top1.acquisition_clk ),
    .RESET_B(net2087),
    .D(_01745_),
    .Q_N(_08244_),
    .Q(\top1.memory2.mem1[138][0] ));
 sg13g2_dfrbp_1 _21649_ (.CLK(\clknet_leaf_49_top1.acquisition_clk ),
    .RESET_B(net2086),
    .D(_01746_),
    .Q_N(_08243_),
    .Q(\top1.memory2.mem1[138][1] ));
 sg13g2_dfrbp_1 _21650_ (.CLK(\clknet_leaf_56_top1.acquisition_clk ),
    .RESET_B(net2085),
    .D(_01747_),
    .Q_N(_08242_),
    .Q(\top1.memory2.mem1[138][2] ));
 sg13g2_dfrbp_1 _21651_ (.CLK(\clknet_leaf_273_top1.acquisition_clk ),
    .RESET_B(net2084),
    .D(_01748_),
    .Q_N(_08241_),
    .Q(\top1.memory2.mem1[13][0] ));
 sg13g2_dfrbp_1 _21652_ (.CLK(\clknet_leaf_277_top1.acquisition_clk ),
    .RESET_B(net2083),
    .D(_01749_),
    .Q_N(_08240_),
    .Q(\top1.memory2.mem1[13][1] ));
 sg13g2_dfrbp_1 _21653_ (.CLK(\clknet_leaf_275_top1.acquisition_clk ),
    .RESET_B(net2082),
    .D(_01750_),
    .Q_N(_08239_),
    .Q(\top1.memory2.mem1[13][2] ));
 sg13g2_dfrbp_1 _21654_ (.CLK(\clknet_leaf_53_top1.acquisition_clk ),
    .RESET_B(net2081),
    .D(_01751_),
    .Q_N(_08238_),
    .Q(\top1.memory2.mem1[140][0] ));
 sg13g2_dfrbp_1 _21655_ (.CLK(\clknet_leaf_51_top1.acquisition_clk ),
    .RESET_B(net2080),
    .D(_01752_),
    .Q_N(_08237_),
    .Q(\top1.memory2.mem1[140][1] ));
 sg13g2_dfrbp_1 _21656_ (.CLK(\clknet_leaf_52_top1.acquisition_clk ),
    .RESET_B(net2079),
    .D(_01753_),
    .Q_N(_08236_),
    .Q(\top1.memory2.mem1[140][2] ));
 sg13g2_dfrbp_1 _21657_ (.CLK(\clknet_leaf_53_top1.acquisition_clk ),
    .RESET_B(net2078),
    .D(_01754_),
    .Q_N(_08235_),
    .Q(\top1.memory2.mem1[141][0] ));
 sg13g2_dfrbp_1 _21658_ (.CLK(\clknet_leaf_51_top1.acquisition_clk ),
    .RESET_B(net2077),
    .D(_01755_),
    .Q_N(_08234_),
    .Q(\top1.memory2.mem1[141][1] ));
 sg13g2_dfrbp_1 _21659_ (.CLK(\clknet_leaf_52_top1.acquisition_clk ),
    .RESET_B(net2076),
    .D(_01756_),
    .Q_N(_08233_),
    .Q(\top1.memory2.mem1[141][2] ));
 sg13g2_dfrbp_1 _21660_ (.CLK(\clknet_leaf_50_top1.acquisition_clk ),
    .RESET_B(net2075),
    .D(_01757_),
    .Q_N(_08232_),
    .Q(\top1.memory2.mem1[142][0] ));
 sg13g2_dfrbp_1 _21661_ (.CLK(\clknet_leaf_51_top1.acquisition_clk ),
    .RESET_B(net2074),
    .D(_01758_),
    .Q_N(_08231_),
    .Q(\top1.memory2.mem1[142][1] ));
 sg13g2_dfrbp_1 _21662_ (.CLK(\clknet_leaf_52_top1.acquisition_clk ),
    .RESET_B(net2073),
    .D(_01759_),
    .Q_N(_08230_),
    .Q(\top1.memory2.mem1[142][2] ));
 sg13g2_dfrbp_1 _21663_ (.CLK(\clknet_leaf_50_top1.acquisition_clk ),
    .RESET_B(net2072),
    .D(_01760_),
    .Q_N(_08229_),
    .Q(\top1.memory2.mem1[143][0] ));
 sg13g2_dfrbp_1 _21664_ (.CLK(\clknet_leaf_19_top1.acquisition_clk ),
    .RESET_B(net2071),
    .D(_01761_),
    .Q_N(_08228_),
    .Q(\top1.memory2.mem1[143][1] ));
 sg13g2_dfrbp_1 _21665_ (.CLK(\clknet_leaf_52_top1.acquisition_clk ),
    .RESET_B(net2070),
    .D(_01762_),
    .Q_N(_08227_),
    .Q(\top1.memory2.mem1[143][2] ));
 sg13g2_dfrbp_1 _21666_ (.CLK(\clknet_leaf_43_top1.acquisition_clk ),
    .RESET_B(net2069),
    .D(_01763_),
    .Q_N(_08226_),
    .Q(\top1.memory2.mem1[144][0] ));
 sg13g2_dfrbp_1 _21667_ (.CLK(\clknet_leaf_57_top1.acquisition_clk ),
    .RESET_B(net2068),
    .D(_01764_),
    .Q_N(_08225_),
    .Q(\top1.memory2.mem1[144][1] ));
 sg13g2_dfrbp_1 _21668_ (.CLK(\clknet_leaf_43_top1.acquisition_clk ),
    .RESET_B(net2067),
    .D(_01765_),
    .Q_N(_08224_),
    .Q(\top1.memory2.mem1[144][2] ));
 sg13g2_dfrbp_1 _21669_ (.CLK(\clknet_leaf_47_top1.acquisition_clk ),
    .RESET_B(net2066),
    .D(_01766_),
    .Q_N(_08223_),
    .Q(\top1.memory2.mem1[145][0] ));
 sg13g2_dfrbp_1 _21670_ (.CLK(\clknet_leaf_58_top1.acquisition_clk ),
    .RESET_B(net2065),
    .D(_01767_),
    .Q_N(_08222_),
    .Q(\top1.memory2.mem1[145][1] ));
 sg13g2_dfrbp_1 _21671_ (.CLK(\clknet_leaf_58_top1.acquisition_clk ),
    .RESET_B(net2064),
    .D(_01768_),
    .Q_N(_08221_),
    .Q(\top1.memory2.mem1[145][2] ));
 sg13g2_dfrbp_1 _21672_ (.CLK(\clknet_leaf_43_top1.acquisition_clk ),
    .RESET_B(net2063),
    .D(_01769_),
    .Q_N(_08220_),
    .Q(\top1.memory2.mem1[146][0] ));
 sg13g2_dfrbp_1 _21673_ (.CLK(\clknet_leaf_58_top1.acquisition_clk ),
    .RESET_B(net2062),
    .D(_01770_),
    .Q_N(_08219_),
    .Q(\top1.memory2.mem1[146][1] ));
 sg13g2_dfrbp_1 _21674_ (.CLK(\clknet_leaf_44_top1.acquisition_clk ),
    .RESET_B(net2061),
    .D(_01771_),
    .Q_N(_08218_),
    .Q(\top1.memory2.mem1[146][2] ));
 sg13g2_dfrbp_1 _21675_ (.CLK(\clknet_leaf_46_top1.acquisition_clk ),
    .RESET_B(net2060),
    .D(_01772_),
    .Q_N(_08217_),
    .Q(\top1.memory2.mem1[147][0] ));
 sg13g2_dfrbp_1 _21676_ (.CLK(\clknet_leaf_57_top1.acquisition_clk ),
    .RESET_B(net2059),
    .D(_01773_),
    .Q_N(_08216_),
    .Q(\top1.memory2.mem1[147][1] ));
 sg13g2_dfrbp_1 _21677_ (.CLK(\clknet_leaf_43_top1.acquisition_clk ),
    .RESET_B(net2058),
    .D(_01774_),
    .Q_N(_08215_),
    .Q(\top1.memory2.mem1[147][2] ));
 sg13g2_dfrbp_1 _21678_ (.CLK(\clknet_leaf_24_top1.acquisition_clk ),
    .RESET_B(net2057),
    .D(_01775_),
    .Q_N(_08214_),
    .Q(\top1.memory2.mem1[148][0] ));
 sg13g2_dfrbp_1 _21679_ (.CLK(\clknet_leaf_25_top1.acquisition_clk ),
    .RESET_B(net2056),
    .D(_01776_),
    .Q_N(_08213_),
    .Q(\top1.memory2.mem1[148][1] ));
 sg13g2_dfrbp_1 _21680_ (.CLK(\clknet_leaf_25_top1.acquisition_clk ),
    .RESET_B(net2055),
    .D(_01777_),
    .Q_N(_08212_),
    .Q(\top1.memory2.mem1[148][2] ));
 sg13g2_dfrbp_1 _21681_ (.CLK(\clknet_leaf_272_top1.acquisition_clk ),
    .RESET_B(net2054),
    .D(_01778_),
    .Q_N(_08211_),
    .Q(\top1.memory2.mem1[14][0] ));
 sg13g2_dfrbp_1 _21682_ (.CLK(\clknet_leaf_277_top1.acquisition_clk ),
    .RESET_B(net2053),
    .D(_01779_),
    .Q_N(_08210_),
    .Q(\top1.memory2.mem1[14][1] ));
 sg13g2_dfrbp_1 _21683_ (.CLK(\clknet_leaf_275_top1.acquisition_clk ),
    .RESET_B(net2052),
    .D(_01780_),
    .Q_N(_08209_),
    .Q(\top1.memory2.mem1[14][2] ));
 sg13g2_dfrbp_1 _21684_ (.CLK(\clknet_leaf_24_top1.acquisition_clk ),
    .RESET_B(net2051),
    .D(_01781_),
    .Q_N(_08208_),
    .Q(\top1.memory2.mem1[150][0] ));
 sg13g2_dfrbp_1 _21685_ (.CLK(\clknet_leaf_24_top1.acquisition_clk ),
    .RESET_B(net2050),
    .D(_01782_),
    .Q_N(_08207_),
    .Q(\top1.memory2.mem1[150][1] ));
 sg13g2_dfrbp_1 _21686_ (.CLK(\clknet_leaf_23_top1.acquisition_clk ),
    .RESET_B(net2049),
    .D(_01783_),
    .Q_N(_08206_),
    .Q(\top1.memory2.mem1[150][2] ));
 sg13g2_dfrbp_1 _21687_ (.CLK(\clknet_leaf_24_top1.acquisition_clk ),
    .RESET_B(net2048),
    .D(_01784_),
    .Q_N(_08205_),
    .Q(\top1.memory2.mem1[151][0] ));
 sg13g2_dfrbp_1 _21688_ (.CLK(\clknet_leaf_25_top1.acquisition_clk ),
    .RESET_B(net2047),
    .D(_01785_),
    .Q_N(_08204_),
    .Q(\top1.memory2.mem1[151][1] ));
 sg13g2_dfrbp_1 _21689_ (.CLK(\clknet_leaf_23_top1.acquisition_clk ),
    .RESET_B(net2046),
    .D(_01786_),
    .Q_N(_08203_),
    .Q(\top1.memory2.mem1[151][2] ));
 sg13g2_dfrbp_1 _21690_ (.CLK(\clknet_leaf_47_top1.acquisition_clk ),
    .RESET_B(net2045),
    .D(_01787_),
    .Q_N(_08202_),
    .Q(\top1.memory2.mem1[152][0] ));
 sg13g2_dfrbp_1 _21691_ (.CLK(\clknet_leaf_45_top1.acquisition_clk ),
    .RESET_B(net2044),
    .D(_01788_),
    .Q_N(_08201_),
    .Q(\top1.memory2.mem1[152][1] ));
 sg13g2_dfrbp_1 _21692_ (.CLK(\clknet_leaf_44_top1.acquisition_clk ),
    .RESET_B(net2043),
    .D(_01789_),
    .Q_N(_08200_),
    .Q(\top1.memory2.mem1[152][2] ));
 sg13g2_dfrbp_1 _21693_ (.CLK(\clknet_leaf_47_top1.acquisition_clk ),
    .RESET_B(net2042),
    .D(_01790_),
    .Q_N(_08199_),
    .Q(\top1.memory2.mem1[153][0] ));
 sg13g2_dfrbp_1 _21694_ (.CLK(\clknet_leaf_45_top1.acquisition_clk ),
    .RESET_B(net2041),
    .D(_01791_),
    .Q_N(_08198_),
    .Q(\top1.memory2.mem1[153][1] ));
 sg13g2_dfrbp_1 _21695_ (.CLK(\clknet_leaf_44_top1.acquisition_clk ),
    .RESET_B(net2040),
    .D(_01792_),
    .Q_N(_08197_),
    .Q(\top1.memory2.mem1[153][2] ));
 sg13g2_dfrbp_1 _21696_ (.CLK(\clknet_leaf_47_top1.acquisition_clk ),
    .RESET_B(net2039),
    .D(_01793_),
    .Q_N(_08196_),
    .Q(\top1.memory2.mem1[154][0] ));
 sg13g2_dfrbp_1 _21697_ (.CLK(\clknet_leaf_45_top1.acquisition_clk ),
    .RESET_B(net2038),
    .D(_01794_),
    .Q_N(_08195_),
    .Q(\top1.memory2.mem1[154][1] ));
 sg13g2_dfrbp_1 _21698_ (.CLK(\clknet_leaf_46_top1.acquisition_clk ),
    .RESET_B(net2037),
    .D(_01795_),
    .Q_N(_08194_),
    .Q(\top1.memory2.mem1[154][2] ));
 sg13g2_dfrbp_1 _21699_ (.CLK(\clknet_leaf_46_top1.acquisition_clk ),
    .RESET_B(net2036),
    .D(_01796_),
    .Q_N(_08193_),
    .Q(\top1.memory2.mem1[155][0] ));
 sg13g2_dfrbp_1 _21700_ (.CLK(\clknet_leaf_45_top1.acquisition_clk ),
    .RESET_B(net2035),
    .D(_01797_),
    .Q_N(_08192_),
    .Q(\top1.memory2.mem1[155][1] ));
 sg13g2_dfrbp_1 _21701_ (.CLK(\clknet_leaf_46_top1.acquisition_clk ),
    .RESET_B(net2034),
    .D(_01798_),
    .Q_N(_08191_),
    .Q(\top1.memory2.mem1[155][2] ));
 sg13g2_dfrbp_1 _21702_ (.CLK(\clknet_leaf_75_top1.acquisition_clk ),
    .RESET_B(net2033),
    .D(_01799_),
    .Q_N(_08190_),
    .Q(\top1.memory2.mem1[156][0] ));
 sg13g2_dfrbp_1 _21703_ (.CLK(\clknet_leaf_70_top1.acquisition_clk ),
    .RESET_B(net2032),
    .D(_01800_),
    .Q_N(_08189_),
    .Q(\top1.memory2.mem1[156][1] ));
 sg13g2_dfrbp_1 _21704_ (.CLK(\clknet_leaf_70_top1.acquisition_clk ),
    .RESET_B(net2031),
    .D(_01801_),
    .Q_N(_08188_),
    .Q(\top1.memory2.mem1[156][2] ));
 sg13g2_dfrbp_1 _21705_ (.CLK(\clknet_leaf_75_top1.acquisition_clk ),
    .RESET_B(net2030),
    .D(_01802_),
    .Q_N(_08187_),
    .Q(\top1.memory2.mem1[157][0] ));
 sg13g2_dfrbp_1 _21706_ (.CLK(\clknet_leaf_70_top1.acquisition_clk ),
    .RESET_B(net2029),
    .D(_01803_),
    .Q_N(_08186_),
    .Q(\top1.memory2.mem1[157][1] ));
 sg13g2_dfrbp_1 _21707_ (.CLK(\clknet_leaf_70_top1.acquisition_clk ),
    .RESET_B(net2028),
    .D(_01804_),
    .Q_N(_08185_),
    .Q(\top1.memory2.mem1[157][2] ));
 sg13g2_dfrbp_1 _21708_ (.CLK(\clknet_leaf_59_top1.acquisition_clk ),
    .RESET_B(net2027),
    .D(_01805_),
    .Q_N(_08184_),
    .Q(\top1.memory2.mem1[158][0] ));
 sg13g2_dfrbp_1 _21709_ (.CLK(\clknet_leaf_70_top1.acquisition_clk ),
    .RESET_B(net2026),
    .D(_01806_),
    .Q_N(_08183_),
    .Q(\top1.memory2.mem1[158][1] ));
 sg13g2_dfrbp_1 _21710_ (.CLK(\clknet_leaf_70_top1.acquisition_clk ),
    .RESET_B(net2025),
    .D(_01807_),
    .Q_N(_08182_),
    .Q(\top1.memory2.mem1[158][2] ));
 sg13g2_dfrbp_1 _21711_ (.CLK(\clknet_leaf_272_top1.acquisition_clk ),
    .RESET_B(net2024),
    .D(_01808_),
    .Q_N(_08181_),
    .Q(\top1.memory2.mem1[15][0] ));
 sg13g2_dfrbp_1 _21712_ (.CLK(\clknet_leaf_277_top1.acquisition_clk ),
    .RESET_B(net2023),
    .D(_01809_),
    .Q_N(_08180_),
    .Q(\top1.memory2.mem1[15][1] ));
 sg13g2_dfrbp_1 _21713_ (.CLK(\clknet_leaf_275_top1.acquisition_clk ),
    .RESET_B(net2022),
    .D(_01810_),
    .Q_N(_08179_),
    .Q(\top1.memory2.mem1[15][2] ));
 sg13g2_dfrbp_1 _21714_ (.CLK(\clknet_leaf_279_top1.acquisition_clk ),
    .RESET_B(net2021),
    .D(_01811_),
    .Q_N(_08178_),
    .Q(\top1.memory2.mem1[160][0] ));
 sg13g2_dfrbp_1 _21715_ (.CLK(\clknet_leaf_278_top1.acquisition_clk ),
    .RESET_B(net2020),
    .D(_01812_),
    .Q_N(_08177_),
    .Q(\top1.memory2.mem1[160][1] ));
 sg13g2_dfrbp_1 _21716_ (.CLK(\clknet_leaf_278_top1.acquisition_clk ),
    .RESET_B(net2019),
    .D(_01813_),
    .Q_N(_08176_),
    .Q(\top1.memory2.mem1[160][2] ));
 sg13g2_dfrbp_1 _21717_ (.CLK(\clknet_leaf_278_top1.acquisition_clk ),
    .RESET_B(net2018),
    .D(_01814_),
    .Q_N(_08175_),
    .Q(\top1.memory2.mem1[161][0] ));
 sg13g2_dfrbp_1 _21718_ (.CLK(\clknet_leaf_275_top1.acquisition_clk ),
    .RESET_B(net2017),
    .D(_01815_),
    .Q_N(_08174_),
    .Q(\top1.memory2.mem1[161][1] ));
 sg13g2_dfrbp_1 _21719_ (.CLK(\clknet_leaf_278_top1.acquisition_clk ),
    .RESET_B(net2016),
    .D(_01816_),
    .Q_N(_08173_),
    .Q(\top1.memory2.mem1[161][2] ));
 sg13g2_dfrbp_1 _21720_ (.CLK(\clknet_leaf_279_top1.acquisition_clk ),
    .RESET_B(net2015),
    .D(_01817_),
    .Q_N(_08172_),
    .Q(\top1.memory2.mem1[162][0] ));
 sg13g2_dfrbp_1 _21721_ (.CLK(\clknet_leaf_275_top1.acquisition_clk ),
    .RESET_B(net2014),
    .D(_01818_),
    .Q_N(_08171_),
    .Q(\top1.memory2.mem1[162][1] ));
 sg13g2_dfrbp_1 _21722_ (.CLK(\clknet_leaf_278_top1.acquisition_clk ),
    .RESET_B(net2013),
    .D(_01819_),
    .Q_N(_08170_),
    .Q(\top1.memory2.mem1[162][2] ));
 sg13g2_dfrbp_1 _21723_ (.CLK(\clknet_leaf_279_top1.acquisition_clk ),
    .RESET_B(net2012),
    .D(_01820_),
    .Q_N(_08169_),
    .Q(\top1.memory2.mem1[163][0] ));
 sg13g2_dfrbp_1 _21724_ (.CLK(\clknet_leaf_275_top1.acquisition_clk ),
    .RESET_B(net2011),
    .D(_01821_),
    .Q_N(_08168_),
    .Q(\top1.memory2.mem1[163][1] ));
 sg13g2_dfrbp_1 _21725_ (.CLK(\clknet_leaf_278_top1.acquisition_clk ),
    .RESET_B(net2010),
    .D(_01822_),
    .Q_N(_08167_),
    .Q(\top1.memory2.mem1[163][2] ));
 sg13g2_dfrbp_1 _21726_ (.CLK(\clknet_leaf_247_top1.acquisition_clk ),
    .RESET_B(net2009),
    .D(_01823_),
    .Q_N(_08166_),
    .Q(\top1.memory2.mem1[164][0] ));
 sg13g2_dfrbp_1 _21727_ (.CLK(\clknet_leaf_255_top1.acquisition_clk ),
    .RESET_B(net2008),
    .D(_01824_),
    .Q_N(_08165_),
    .Q(\top1.memory2.mem1[164][1] ));
 sg13g2_dfrbp_1 _21728_ (.CLK(\clknet_leaf_243_top1.acquisition_clk ),
    .RESET_B(net2007),
    .D(_01825_),
    .Q_N(_08164_),
    .Q(\top1.memory2.mem1[164][2] ));
 sg13g2_dfrbp_1 _21729_ (.CLK(\clknet_leaf_247_top1.acquisition_clk ),
    .RESET_B(net2006),
    .D(_01826_),
    .Q_N(_08163_),
    .Q(\top1.memory2.mem1[165][0] ));
 sg13g2_dfrbp_1 _21730_ (.CLK(\clknet_leaf_247_top1.acquisition_clk ),
    .RESET_B(net2005),
    .D(_01827_),
    .Q_N(_08162_),
    .Q(\top1.memory2.mem1[165][1] ));
 sg13g2_dfrbp_1 _21731_ (.CLK(\clknet_leaf_243_top1.acquisition_clk ),
    .RESET_B(net2004),
    .D(_01828_),
    .Q_N(_08161_),
    .Q(\top1.memory2.mem1[165][2] ));
 sg13g2_dfrbp_1 _21732_ (.CLK(\clknet_leaf_247_top1.acquisition_clk ),
    .RESET_B(net2003),
    .D(_01829_),
    .Q_N(_08160_),
    .Q(\top1.memory2.mem1[166][0] ));
 sg13g2_dfrbp_1 _21733_ (.CLK(\clknet_leaf_247_top1.acquisition_clk ),
    .RESET_B(net2002),
    .D(_01830_),
    .Q_N(_08159_),
    .Q(\top1.memory2.mem1[166][1] ));
 sg13g2_dfrbp_1 _21734_ (.CLK(\clknet_leaf_238_top1.acquisition_clk ),
    .RESET_B(net2001),
    .D(_01831_),
    .Q_N(_08158_),
    .Q(\top1.memory2.mem1[166][2] ));
 sg13g2_dfrbp_1 _21735_ (.CLK(\clknet_leaf_249_top1.acquisition_clk ),
    .RESET_B(net2000),
    .D(_01832_),
    .Q_N(_08157_),
    .Q(\top1.memory2.mem1[167][0] ));
 sg13g2_dfrbp_1 _21736_ (.CLK(\clknet_leaf_247_top1.acquisition_clk ),
    .RESET_B(net1999),
    .D(_01833_),
    .Q_N(_08156_),
    .Q(\top1.memory2.mem1[167][1] ));
 sg13g2_dfrbp_1 _21737_ (.CLK(\clknet_leaf_243_top1.acquisition_clk ),
    .RESET_B(net1998),
    .D(_01834_),
    .Q_N(_08155_),
    .Q(\top1.memory2.mem1[167][2] ));
 sg13g2_dfrbp_1 _21738_ (.CLK(\clknet_leaf_246_top1.acquisition_clk ),
    .RESET_B(net1997),
    .D(_01835_),
    .Q_N(_08154_),
    .Q(\top1.memory2.mem1[168][0] ));
 sg13g2_dfrbp_1 _21739_ (.CLK(\clknet_leaf_244_top1.acquisition_clk ),
    .RESET_B(net1996),
    .D(_01836_),
    .Q_N(_08153_),
    .Q(\top1.memory2.mem1[168][1] ));
 sg13g2_dfrbp_1 _21740_ (.CLK(\clknet_leaf_243_top1.acquisition_clk ),
    .RESET_B(net1995),
    .D(_01837_),
    .Q_N(_08152_),
    .Q(\top1.memory2.mem1[168][2] ));
 sg13g2_dfrbp_1 _21741_ (.CLK(\clknet_leaf_109_top1.acquisition_clk ),
    .RESET_B(net1994),
    .D(_01838_),
    .Q_N(_08151_),
    .Q(\top1.memory2.mem1[16][0] ));
 sg13g2_dfrbp_1 _21742_ (.CLK(\clknet_leaf_109_top1.acquisition_clk ),
    .RESET_B(net1993),
    .D(_01839_),
    .Q_N(_08150_),
    .Q(\top1.memory2.mem1[16][1] ));
 sg13g2_dfrbp_1 _21743_ (.CLK(\clknet_leaf_106_top1.acquisition_clk ),
    .RESET_B(net1992),
    .D(_01840_),
    .Q_N(_08149_),
    .Q(\top1.memory2.mem1[16][2] ));
 sg13g2_dfrbp_1 _21744_ (.CLK(\clknet_leaf_245_top1.acquisition_clk ),
    .RESET_B(net1991),
    .D(_01841_),
    .Q_N(_08148_),
    .Q(\top1.memory2.mem1[170][0] ));
 sg13g2_dfrbp_1 _21745_ (.CLK(\clknet_leaf_244_top1.acquisition_clk ),
    .RESET_B(net1990),
    .D(_01842_),
    .Q_N(_08147_),
    .Q(\top1.memory2.mem1[170][1] ));
 sg13g2_dfrbp_1 _21746_ (.CLK(\clknet_leaf_243_top1.acquisition_clk ),
    .RESET_B(net1989),
    .D(_01843_),
    .Q_N(_08146_),
    .Q(\top1.memory2.mem1[170][2] ));
 sg13g2_dfrbp_1 _21747_ (.CLK(\clknet_leaf_247_top1.acquisition_clk ),
    .RESET_B(net1988),
    .D(_01844_),
    .Q_N(_08145_),
    .Q(\top1.memory2.mem1[171][0] ));
 sg13g2_dfrbp_1 _21748_ (.CLK(\clknet_leaf_244_top1.acquisition_clk ),
    .RESET_B(net1987),
    .D(_01845_),
    .Q_N(_08144_),
    .Q(\top1.memory2.mem1[171][1] ));
 sg13g2_dfrbp_1 _21749_ (.CLK(\clknet_leaf_243_top1.acquisition_clk ),
    .RESET_B(net1986),
    .D(_01846_),
    .Q_N(_08143_),
    .Q(\top1.memory2.mem1[171][2] ));
 sg13g2_dfrbp_1 _21750_ (.CLK(\clknet_leaf_242_top1.acquisition_clk ),
    .RESET_B(net1985),
    .D(_01847_),
    .Q_N(_08142_),
    .Q(\top1.memory2.mem1[172][0] ));
 sg13g2_dfrbp_1 _21751_ (.CLK(\clknet_leaf_246_top1.acquisition_clk ),
    .RESET_B(net1984),
    .D(_01848_),
    .Q_N(_08141_),
    .Q(\top1.memory2.mem1[172][1] ));
 sg13g2_dfrbp_1 _21752_ (.CLK(\clknet_leaf_241_top1.acquisition_clk ),
    .RESET_B(net1983),
    .D(_01849_),
    .Q_N(_08140_),
    .Q(\top1.memory2.mem1[172][2] ));
 sg13g2_dfrbp_1 _21753_ (.CLK(\clknet_leaf_242_top1.acquisition_clk ),
    .RESET_B(net1982),
    .D(_01850_),
    .Q_N(_08139_),
    .Q(\top1.memory2.mem1[173][0] ));
 sg13g2_dfrbp_1 _21754_ (.CLK(\clknet_leaf_246_top1.acquisition_clk ),
    .RESET_B(net1981),
    .D(_01851_),
    .Q_N(_08138_),
    .Q(\top1.memory2.mem1[173][1] ));
 sg13g2_dfrbp_1 _21755_ (.CLK(\clknet_leaf_241_top1.acquisition_clk ),
    .RESET_B(net1980),
    .D(_01852_),
    .Q_N(_08137_),
    .Q(\top1.memory2.mem1[173][2] ));
 sg13g2_dfrbp_1 _21756_ (.CLK(\clknet_leaf_242_top1.acquisition_clk ),
    .RESET_B(net1979),
    .D(_01853_),
    .Q_N(_08136_),
    .Q(\top1.memory2.mem1[174][0] ));
 sg13g2_dfrbp_1 _21757_ (.CLK(\clknet_leaf_245_top1.acquisition_clk ),
    .RESET_B(net1978),
    .D(_01854_),
    .Q_N(_08135_),
    .Q(\top1.memory2.mem1[174][1] ));
 sg13g2_dfrbp_1 _21758_ (.CLK(\clknet_leaf_241_top1.acquisition_clk ),
    .RESET_B(net1977),
    .D(_01855_),
    .Q_N(_08134_),
    .Q(\top1.memory2.mem1[174][2] ));
 sg13g2_dfrbp_1 _21759_ (.CLK(\clknet_leaf_241_top1.acquisition_clk ),
    .RESET_B(net1976),
    .D(_01856_),
    .Q_N(_08133_),
    .Q(\top1.memory2.mem1[175][0] ));
 sg13g2_dfrbp_1 _21760_ (.CLK(\clknet_leaf_246_top1.acquisition_clk ),
    .RESET_B(net1975),
    .D(_01857_),
    .Q_N(_08132_),
    .Q(\top1.memory2.mem1[175][1] ));
 sg13g2_dfrbp_1 _21761_ (.CLK(\clknet_leaf_241_top1.acquisition_clk ),
    .RESET_B(net1974),
    .D(_01858_),
    .Q_N(_08131_),
    .Q(\top1.memory2.mem1[175][2] ));
 sg13g2_dfrbp_1 _21762_ (.CLK(\clknet_leaf_191_top1.acquisition_clk ),
    .RESET_B(net1973),
    .D(_01859_),
    .Q_N(_08130_),
    .Q(\top1.memory2.mem1[176][0] ));
 sg13g2_dfrbp_1 _21763_ (.CLK(\clknet_leaf_250_top1.acquisition_clk ),
    .RESET_B(net1972),
    .D(_01860_),
    .Q_N(_08129_),
    .Q(\top1.memory2.mem1[176][1] ));
 sg13g2_dfrbp_1 _21764_ (.CLK(\clknet_leaf_250_top1.acquisition_clk ),
    .RESET_B(net1971),
    .D(_01861_),
    .Q_N(_08128_),
    .Q(\top1.memory2.mem1[176][2] ));
 sg13g2_dfrbp_1 _21765_ (.CLK(\clknet_leaf_191_top1.acquisition_clk ),
    .RESET_B(net1970),
    .D(_01862_),
    .Q_N(_08127_),
    .Q(\top1.memory2.mem1[177][0] ));
 sg13g2_dfrbp_1 _21766_ (.CLK(\clknet_leaf_253_top1.acquisition_clk ),
    .RESET_B(net1969),
    .D(_01863_),
    .Q_N(_08126_),
    .Q(\top1.memory2.mem1[177][1] ));
 sg13g2_dfrbp_1 _21767_ (.CLK(\clknet_leaf_250_top1.acquisition_clk ),
    .RESET_B(net1968),
    .D(_01864_),
    .Q_N(_08125_),
    .Q(\top1.memory2.mem1[177][2] ));
 sg13g2_dfrbp_1 _21768_ (.CLK(\clknet_leaf_190_top1.acquisition_clk ),
    .RESET_B(net1967),
    .D(_01865_),
    .Q_N(_08124_),
    .Q(\top1.memory2.mem1[178][0] ));
 sg13g2_dfrbp_1 _21769_ (.CLK(\clknet_leaf_249_top1.acquisition_clk ),
    .RESET_B(net1966),
    .D(_01866_),
    .Q_N(_08123_),
    .Q(\top1.memory2.mem1[178][1] ));
 sg13g2_dfrbp_1 _21770_ (.CLK(\clknet_leaf_250_top1.acquisition_clk ),
    .RESET_B(net1965),
    .D(_01867_),
    .Q_N(_08122_),
    .Q(\top1.memory2.mem1[178][2] ));
 sg13g2_dfrbp_1 _21771_ (.CLK(\clknet_leaf_108_top1.acquisition_clk ),
    .RESET_B(net1964),
    .D(_01868_),
    .Q_N(_08121_),
    .Q(\top1.memory2.mem1[17][0] ));
 sg13g2_dfrbp_1 _21772_ (.CLK(\clknet_leaf_109_top1.acquisition_clk ),
    .RESET_B(net1963),
    .D(_01869_),
    .Q_N(_08120_),
    .Q(\top1.memory2.mem1[17][1] ));
 sg13g2_dfrbp_1 _21773_ (.CLK(\clknet_leaf_106_top1.acquisition_clk ),
    .RESET_B(net1962),
    .D(_01870_),
    .Q_N(_08119_),
    .Q(\top1.memory2.mem1[17][2] ));
 sg13g2_dfrbp_1 _21774_ (.CLK(\clknet_leaf_238_top1.acquisition_clk ),
    .RESET_B(net1961),
    .D(_01871_),
    .Q_N(_08118_),
    .Q(\top1.memory2.mem1[180][0] ));
 sg13g2_dfrbp_1 _21775_ (.CLK(\clknet_leaf_237_top1.acquisition_clk ),
    .RESET_B(net1960),
    .D(_01872_),
    .Q_N(_08117_),
    .Q(\top1.memory2.mem1[180][1] ));
 sg13g2_dfrbp_1 _21776_ (.CLK(\clknet_leaf_237_top1.acquisition_clk ),
    .RESET_B(net1959),
    .D(_01873_),
    .Q_N(_08116_),
    .Q(\top1.memory2.mem1[180][2] ));
 sg13g2_dfrbp_1 _21777_ (.CLK(\clknet_leaf_237_top1.acquisition_clk ),
    .RESET_B(net1958),
    .D(_01874_),
    .Q_N(_08115_),
    .Q(\top1.memory2.mem1[181][0] ));
 sg13g2_dfrbp_1 _21778_ (.CLK(\clknet_leaf_237_top1.acquisition_clk ),
    .RESET_B(net1957),
    .D(_01875_),
    .Q_N(_08114_),
    .Q(\top1.memory2.mem1[181][1] ));
 sg13g2_dfrbp_1 _21779_ (.CLK(\clknet_leaf_237_top1.acquisition_clk ),
    .RESET_B(net1956),
    .D(_01876_),
    .Q_N(_08113_),
    .Q(\top1.memory2.mem1[181][2] ));
 sg13g2_dfrbp_1 _21780_ (.CLK(\clknet_leaf_232_top1.acquisition_clk ),
    .RESET_B(net1955),
    .D(_01877_),
    .Q_N(_08112_),
    .Q(\top1.memory2.mem1[182][0] ));
 sg13g2_dfrbp_1 _21781_ (.CLK(\clknet_leaf_236_top1.acquisition_clk ),
    .RESET_B(net1954),
    .D(_01878_),
    .Q_N(_08111_),
    .Q(\top1.memory2.mem1[182][1] ));
 sg13g2_dfrbp_1 _21782_ (.CLK(\clknet_leaf_239_top1.acquisition_clk ),
    .RESET_B(net1953),
    .D(_01879_),
    .Q_N(_08110_),
    .Q(\top1.memory2.mem1[182][2] ));
 sg13g2_dfrbp_1 _21783_ (.CLK(\clknet_leaf_232_top1.acquisition_clk ),
    .RESET_B(net1952),
    .D(_01880_),
    .Q_N(_08109_),
    .Q(\top1.memory2.mem1[183][0] ));
 sg13g2_dfrbp_1 _21784_ (.CLK(\clknet_leaf_236_top1.acquisition_clk ),
    .RESET_B(net1951),
    .D(_01881_),
    .Q_N(_08108_),
    .Q(\top1.memory2.mem1[183][1] ));
 sg13g2_dfrbp_1 _21785_ (.CLK(\clknet_leaf_239_top1.acquisition_clk ),
    .RESET_B(net1950),
    .D(_01882_),
    .Q_N(_08107_),
    .Q(\top1.memory2.mem1[183][2] ));
 sg13g2_dfrbp_1 _21786_ (.CLK(\clknet_leaf_254_top1.acquisition_clk ),
    .RESET_B(net1949),
    .D(_01883_),
    .Q_N(_08106_),
    .Q(\top1.memory2.mem1[184][0] ));
 sg13g2_dfrbp_1 _21787_ (.CLK(\clknet_leaf_249_top1.acquisition_clk ),
    .RESET_B(net1948),
    .D(_01884_),
    .Q_N(_08105_),
    .Q(\top1.memory2.mem1[184][1] ));
 sg13g2_dfrbp_1 _21788_ (.CLK(\clknet_leaf_248_top1.acquisition_clk ),
    .RESET_B(net1947),
    .D(_01885_),
    .Q_N(_08104_),
    .Q(\top1.memory2.mem1[184][2] ));
 sg13g2_dfrbp_1 _21789_ (.CLK(\clknet_leaf_254_top1.acquisition_clk ),
    .RESET_B(net1946),
    .D(_01886_),
    .Q_N(_08103_),
    .Q(\top1.memory2.mem1[185][0] ));
 sg13g2_dfrbp_1 _21790_ (.CLK(\clknet_leaf_244_top1.acquisition_clk ),
    .RESET_B(net1945),
    .D(_01887_),
    .Q_N(_08102_),
    .Q(\top1.memory2.mem1[185][1] ));
 sg13g2_dfrbp_1 _21791_ (.CLK(\clknet_leaf_248_top1.acquisition_clk ),
    .RESET_B(net1944),
    .D(_01888_),
    .Q_N(_08101_),
    .Q(\top1.memory2.mem1[185][2] ));
 sg13g2_dfrbp_1 _21792_ (.CLK(\clknet_leaf_247_top1.acquisition_clk ),
    .RESET_B(net1943),
    .D(_01889_),
    .Q_N(_08100_),
    .Q(\top1.memory2.mem1[186][0] ));
 sg13g2_dfrbp_1 _21793_ (.CLK(\clknet_leaf_249_top1.acquisition_clk ),
    .RESET_B(net1942),
    .D(_01890_),
    .Q_N(_08099_),
    .Q(\top1.memory2.mem1[186][1] ));
 sg13g2_dfrbp_1 _21794_ (.CLK(\clknet_leaf_249_top1.acquisition_clk ),
    .RESET_B(net1941),
    .D(_01891_),
    .Q_N(_08098_),
    .Q(\top1.memory2.mem1[186][2] ));
 sg13g2_dfrbp_1 _21795_ (.CLK(\clknet_leaf_255_top1.acquisition_clk ),
    .RESET_B(net1940),
    .D(_01892_),
    .Q_N(_08097_),
    .Q(\top1.memory2.mem1[187][0] ));
 sg13g2_dfrbp_1 _21796_ (.CLK(\clknet_leaf_249_top1.acquisition_clk ),
    .RESET_B(net1939),
    .D(_01893_),
    .Q_N(_08096_),
    .Q(\top1.memory2.mem1[187][1] ));
 sg13g2_dfrbp_1 _21797_ (.CLK(\clknet_leaf_248_top1.acquisition_clk ),
    .RESET_B(net1938),
    .D(_01894_),
    .Q_N(_08095_),
    .Q(\top1.memory2.mem1[187][2] ));
 sg13g2_dfrbp_1 _21798_ (.CLK(\clknet_leaf_185_top1.acquisition_clk ),
    .RESET_B(net1937),
    .D(_01895_),
    .Q_N(_08094_),
    .Q(\top1.memory2.mem1[188][0] ));
 sg13g2_dfrbp_1 _21799_ (.CLK(\clknet_leaf_187_top1.acquisition_clk ),
    .RESET_B(net1936),
    .D(_01896_),
    .Q_N(_08093_),
    .Q(\top1.memory2.mem1[188][1] ));
 sg13g2_dfrbp_1 _21800_ (.CLK(\clknet_leaf_254_top1.acquisition_clk ),
    .RESET_B(net1935),
    .D(_01897_),
    .Q_N(_08092_),
    .Q(\top1.memory2.mem1[188][2] ));
 sg13g2_dfrbp_1 _21801_ (.CLK(\clknet_leaf_109_top1.acquisition_clk ),
    .RESET_B(net1934),
    .D(_01898_),
    .Q_N(_08091_),
    .Q(\top1.memory2.mem1[18][0] ));
 sg13g2_dfrbp_1 _21802_ (.CLK(\clknet_leaf_113_top1.acquisition_clk ),
    .RESET_B(net1933),
    .D(_01899_),
    .Q_N(_08090_),
    .Q(\top1.memory2.mem1[18][1] ));
 sg13g2_dfrbp_1 _21803_ (.CLK(\clknet_leaf_106_top1.acquisition_clk ),
    .RESET_B(net1932),
    .D(_01900_),
    .Q_N(_08089_),
    .Q(\top1.memory2.mem1[18][2] ));
 sg13g2_dfrbp_1 _21804_ (.CLK(\clknet_leaf_187_top1.acquisition_clk ),
    .RESET_B(net1931),
    .D(_01901_),
    .Q_N(_08088_),
    .Q(\top1.memory2.mem1[190][0] ));
 sg13g2_dfrbp_1 _21805_ (.CLK(\clknet_leaf_191_top1.acquisition_clk ),
    .RESET_B(net1930),
    .D(_01902_),
    .Q_N(_08087_),
    .Q(\top1.memory2.mem1[190][1] ));
 sg13g2_dfrbp_1 _21806_ (.CLK(\clknet_leaf_254_top1.acquisition_clk ),
    .RESET_B(net1929),
    .D(_01903_),
    .Q_N(_08086_),
    .Q(\top1.memory2.mem1[190][2] ));
 sg13g2_dfrbp_1 _21807_ (.CLK(\clknet_leaf_186_top1.acquisition_clk ),
    .RESET_B(net1928),
    .D(_01904_),
    .Q_N(_08085_),
    .Q(\top1.memory2.mem1[191][0] ));
 sg13g2_dfrbp_1 _21808_ (.CLK(\clknet_leaf_191_top1.acquisition_clk ),
    .RESET_B(net1927),
    .D(_01905_),
    .Q_N(_08084_),
    .Q(\top1.memory2.mem1[191][1] ));
 sg13g2_dfrbp_1 _21809_ (.CLK(\clknet_leaf_253_top1.acquisition_clk ),
    .RESET_B(net1926),
    .D(_01906_),
    .Q_N(_08083_),
    .Q(\top1.memory2.mem1[191][2] ));
 sg13g2_dfrbp_1 _21810_ (.CLK(\clknet_leaf_267_top1.acquisition_clk ),
    .RESET_B(net1925),
    .D(_01907_),
    .Q_N(_08082_),
    .Q(\top1.memory2.mem1[192][0] ));
 sg13g2_dfrbp_1 _21811_ (.CLK(\clknet_leaf_31_top1.acquisition_clk ),
    .RESET_B(net1924),
    .D(_01908_),
    .Q_N(_08081_),
    .Q(\top1.memory2.mem1[192][1] ));
 sg13g2_dfrbp_1 _21812_ (.CLK(\clknet_leaf_267_top1.acquisition_clk ),
    .RESET_B(net1923),
    .D(_01909_),
    .Q_N(_08080_),
    .Q(\top1.memory2.mem1[192][2] ));
 sg13g2_dfrbp_1 _21813_ (.CLK(\clknet_leaf_267_top1.acquisition_clk ),
    .RESET_B(net1922),
    .D(_01910_),
    .Q_N(_08079_),
    .Q(\top1.memory2.mem1[193][0] ));
 sg13g2_dfrbp_1 _21814_ (.CLK(\clknet_leaf_31_top1.acquisition_clk ),
    .RESET_B(net1921),
    .D(_01911_),
    .Q_N(_08078_),
    .Q(\top1.memory2.mem1[193][1] ));
 sg13g2_dfrbp_1 _21815_ (.CLK(\clknet_leaf_267_top1.acquisition_clk ),
    .RESET_B(net1920),
    .D(_01912_),
    .Q_N(_08077_),
    .Q(\top1.memory2.mem1[193][2] ));
 sg13g2_dfrbp_1 _21816_ (.CLK(\clknet_leaf_30_top1.acquisition_clk ),
    .RESET_B(net1919),
    .D(_01913_),
    .Q_N(_08076_),
    .Q(\top1.memory2.mem1[194][0] ));
 sg13g2_dfrbp_1 _21817_ (.CLK(\clknet_leaf_31_top1.acquisition_clk ),
    .RESET_B(net1918),
    .D(_01914_),
    .Q_N(_08075_),
    .Q(\top1.memory2.mem1[194][1] ));
 sg13g2_dfrbp_1 _21818_ (.CLK(\clknet_leaf_31_top1.acquisition_clk ),
    .RESET_B(net1917),
    .D(_01915_),
    .Q_N(_08074_),
    .Q(\top1.memory2.mem1[194][2] ));
 sg13g2_dfrbp_1 _21819_ (.CLK(\clknet_leaf_267_top1.acquisition_clk ),
    .RESET_B(net1916),
    .D(_01916_),
    .Q_N(_08073_),
    .Q(\top1.memory2.mem1[195][0] ));
 sg13g2_dfrbp_1 _21820_ (.CLK(\clknet_leaf_35_top1.acquisition_clk ),
    .RESET_B(net1915),
    .D(_01917_),
    .Q_N(_08072_),
    .Q(\top1.memory2.mem1[195][1] ));
 sg13g2_dfrbp_1 _21821_ (.CLK(\clknet_leaf_267_top1.acquisition_clk ),
    .RESET_B(net1914),
    .D(_01918_),
    .Q_N(_08071_),
    .Q(\top1.memory2.mem1[195][2] ));
 sg13g2_dfrbp_1 _21822_ (.CLK(\clknet_leaf_33_top1.acquisition_clk ),
    .RESET_B(net1913),
    .D(_01919_),
    .Q_N(_08070_),
    .Q(\top1.memory2.mem1[196][0] ));
 sg13g2_dfrbp_1 _21823_ (.CLK(\clknet_leaf_32_top1.acquisition_clk ),
    .RESET_B(net1912),
    .D(_01920_),
    .Q_N(_08069_),
    .Q(\top1.memory2.mem1[196][1] ));
 sg13g2_dfrbp_1 _21824_ (.CLK(\clknet_leaf_32_top1.acquisition_clk ),
    .RESET_B(net1911),
    .D(_01921_),
    .Q_N(_08068_),
    .Q(\top1.memory2.mem1[196][2] ));
 sg13g2_dfrbp_1 _21825_ (.CLK(\clknet_leaf_33_top1.acquisition_clk ),
    .RESET_B(net1910),
    .D(_01922_),
    .Q_N(_08067_),
    .Q(\top1.memory2.mem1[197][0] ));
 sg13g2_dfrbp_1 _21826_ (.CLK(\clknet_leaf_32_top1.acquisition_clk ),
    .RESET_B(net1909),
    .D(_01923_),
    .Q_N(_08066_),
    .Q(\top1.memory2.mem1[197][1] ));
 sg13g2_dfrbp_1 _21827_ (.CLK(\clknet_leaf_33_top1.acquisition_clk ),
    .RESET_B(net1908),
    .D(_01924_),
    .Q_N(_08065_),
    .Q(\top1.memory2.mem1[197][2] ));
 sg13g2_dfrbp_1 _21828_ (.CLK(\clknet_leaf_33_top1.acquisition_clk ),
    .RESET_B(net1907),
    .D(_01925_),
    .Q_N(_08064_),
    .Q(\top1.memory2.mem1[198][0] ));
 sg13g2_dfrbp_1 _21829_ (.CLK(\clknet_leaf_31_top1.acquisition_clk ),
    .RESET_B(net1906),
    .D(_01926_),
    .Q_N(_08063_),
    .Q(\top1.memory2.mem1[198][1] ));
 sg13g2_dfrbp_1 _21830_ (.CLK(\clknet_leaf_32_top1.acquisition_clk ),
    .RESET_B(net1905),
    .D(_01927_),
    .Q_N(_08062_),
    .Q(\top1.memory2.mem1[198][2] ));
 sg13g2_dfrbp_1 _21831_ (.CLK(\clknet_leaf_272_top1.acquisition_clk ),
    .RESET_B(net1904),
    .D(_01928_),
    .Q_N(_08061_),
    .Q(\top1.memory2.mem1[9][0] ));
 sg13g2_dfrbp_1 _21832_ (.CLK(\clknet_leaf_276_top1.acquisition_clk ),
    .RESET_B(net1903),
    .D(_01929_),
    .Q_N(_08060_),
    .Q(\top1.memory2.mem1[9][1] ));
 sg13g2_dfrbp_1 _21833_ (.CLK(\clknet_leaf_274_top1.acquisition_clk ),
    .RESET_B(net1902),
    .D(_01930_),
    .Q_N(_08059_),
    .Q(\top1.memory2.mem1[9][2] ));
 sg13g2_dfrbp_1 _21834_ (.CLK(\clknet_leaf_113_top1.acquisition_clk ),
    .RESET_B(net1901),
    .D(_01931_),
    .Q_N(_08058_),
    .Q(\top1.memory2.mem2[19][0] ));
 sg13g2_dfrbp_1 _21835_ (.CLK(\clknet_leaf_123_top1.acquisition_clk ),
    .RESET_B(net1900),
    .D(_01932_),
    .Q_N(_08057_),
    .Q(\top1.memory2.mem2[19][1] ));
 sg13g2_dfrbp_1 _21836_ (.CLK(\clknet_leaf_112_top1.acquisition_clk ),
    .RESET_B(net1899),
    .D(_01933_),
    .Q_N(_08056_),
    .Q(\top1.memory2.mem2[19][2] ));
 sg13g2_dfrbp_1 _21837_ (.CLK(\clknet_leaf_125_top1.acquisition_clk ),
    .RESET_B(net1898),
    .D(_01934_),
    .Q_N(_08055_),
    .Q(\top1.memory2.mem2[29][0] ));
 sg13g2_dfrbp_1 _21838_ (.CLK(\clknet_leaf_87_top1.acquisition_clk ),
    .RESET_B(net1897),
    .D(_01935_),
    .Q_N(_08054_),
    .Q(\top1.memory2.mem2[29][1] ));
 sg13g2_dfrbp_1 _21839_ (.CLK(\clknet_leaf_124_top1.acquisition_clk ),
    .RESET_B(net1896),
    .D(_01936_),
    .Q_N(_08053_),
    .Q(\top1.memory2.mem2[29][2] ));
 sg13g2_dfrbp_1 _21840_ (.CLK(\clknet_leaf_136_top1.acquisition_clk ),
    .RESET_B(net1895),
    .D(_01937_),
    .Q_N(_08052_),
    .Q(\top1.memory2.mem2[39][0] ));
 sg13g2_dfrbp_1 _21841_ (.CLK(\clknet_leaf_135_top1.acquisition_clk ),
    .RESET_B(net1894),
    .D(_01938_),
    .Q_N(_08051_),
    .Q(\top1.memory2.mem2[39][1] ));
 sg13g2_dfrbp_1 _21842_ (.CLK(\clknet_leaf_116_top1.acquisition_clk ),
    .RESET_B(net1893),
    .D(_01939_),
    .Q_N(_08050_),
    .Q(\top1.memory2.mem2[39][2] ));
 sg13g2_dfrbp_1 _21843_ (.CLK(\clknet_leaf_139_top1.acquisition_clk ),
    .RESET_B(net1892),
    .D(_01940_),
    .Q_N(_08049_),
    .Q(\top1.memory2.mem2[49][0] ));
 sg13g2_dfrbp_1 _21844_ (.CLK(\clknet_leaf_143_top1.acquisition_clk ),
    .RESET_B(net1891),
    .D(_01941_),
    .Q_N(_08048_),
    .Q(\top1.memory2.mem2[49][1] ));
 sg13g2_dfrbp_1 _21845_ (.CLK(\clknet_leaf_141_top1.acquisition_clk ),
    .RESET_B(net1890),
    .D(_01942_),
    .Q_N(_08047_),
    .Q(\top1.memory2.mem2[49][2] ));
 sg13g2_dfrbp_1 _21846_ (.CLK(\clknet_leaf_157_top1.acquisition_clk ),
    .RESET_B(net1889),
    .D(_01943_),
    .Q_N(_08046_),
    .Q(\top1.memory2.mem2[59][0] ));
 sg13g2_dfrbp_1 _21847_ (.CLK(\clknet_leaf_156_top1.acquisition_clk ),
    .RESET_B(net1888),
    .D(_01944_),
    .Q_N(_08045_),
    .Q(\top1.memory2.mem2[59][1] ));
 sg13g2_dfrbp_1 _21848_ (.CLK(\clknet_leaf_156_top1.acquisition_clk ),
    .RESET_B(net1887),
    .D(_01945_),
    .Q_N(_08044_),
    .Q(\top1.memory2.mem2[59][2] ));
 sg13g2_dfrbp_1 _21849_ (.CLK(\clknet_leaf_7_top1.acquisition_clk ),
    .RESET_B(net1886),
    .D(_01946_),
    .Q_N(_08043_),
    .Q(\top1.memory2.mem2[69][0] ));
 sg13g2_dfrbp_1 _21850_ (.CLK(\clknet_leaf_10_top1.acquisition_clk ),
    .RESET_B(net1885),
    .D(_01947_),
    .Q_N(_08042_),
    .Q(\top1.memory2.mem2[69][1] ));
 sg13g2_dfrbp_1 _21851_ (.CLK(\clknet_leaf_9_top1.acquisition_clk ),
    .RESET_B(net1884),
    .D(_01948_),
    .Q_N(_08041_),
    .Q(\top1.memory2.mem2[69][2] ));
 sg13g2_dfrbp_1 _21852_ (.CLK(\clknet_leaf_302_top1.acquisition_clk ),
    .RESET_B(net1883),
    .D(_01949_),
    .Q_N(_08040_),
    .Q(\top1.memory2.mem2[79][0] ));
 sg13g2_dfrbp_1 _21853_ (.CLK(\clknet_leaf_0_top1.acquisition_clk ),
    .RESET_B(net1882),
    .D(_01950_),
    .Q_N(_08039_),
    .Q(\top1.memory2.mem2[79][1] ));
 sg13g2_dfrbp_1 _21854_ (.CLK(\clknet_leaf_301_top1.acquisition_clk ),
    .RESET_B(net1881),
    .D(_01951_),
    .Q_N(_08038_),
    .Q(\top1.memory2.mem2[79][2] ));
 sg13g2_dfrbp_1 _21855_ (.CLK(\clknet_leaf_290_top1.acquisition_clk ),
    .RESET_B(net1880),
    .D(_01952_),
    .Q_N(_08037_),
    .Q(\top1.memory2.mem2[89][0] ));
 sg13g2_dfrbp_1 _21856_ (.CLK(\clknet_leaf_291_top1.acquisition_clk ),
    .RESET_B(net1879),
    .D(_01953_),
    .Q_N(_08036_),
    .Q(\top1.memory2.mem2[89][1] ));
 sg13g2_dfrbp_1 _21857_ (.CLK(\clknet_leaf_8_top1.acquisition_clk ),
    .RESET_B(net1878),
    .D(_01954_),
    .Q_N(_08035_),
    .Q(\top1.memory2.mem2[89][2] ));
 sg13g2_dfrbp_1 _21858_ (.CLK(\clknet_leaf_231_top1.acquisition_clk ),
    .RESET_B(net1877),
    .D(_01955_),
    .Q_N(_08034_),
    .Q(\top1.memory2.mem2[99][0] ));
 sg13g2_dfrbp_1 _21859_ (.CLK(\clknet_leaf_233_top1.acquisition_clk ),
    .RESET_B(net1876),
    .D(_01956_),
    .Q_N(_08033_),
    .Q(\top1.memory2.mem2[99][1] ));
 sg13g2_dfrbp_1 _21860_ (.CLK(\clknet_leaf_251_top1.acquisition_clk ),
    .RESET_B(net1875),
    .D(_01957_),
    .Q_N(_08032_),
    .Q(\top1.memory2.mem2[99][2] ));
 sg13g2_dfrbp_1 _21861_ (.CLK(\clknet_leaf_225_top1.acquisition_clk ),
    .RESET_B(net1874),
    .D(_01958_),
    .Q_N(_08031_),
    .Q(\top1.memory2.mem2[109][0] ));
 sg13g2_dfrbp_1 _21862_ (.CLK(\clknet_leaf_226_top1.acquisition_clk ),
    .RESET_B(net1873),
    .D(_01959_),
    .Q_N(_08030_),
    .Q(\top1.memory2.mem2[109][1] ));
 sg13g2_dfrbp_1 _21863_ (.CLK(\clknet_leaf_235_top1.acquisition_clk ),
    .RESET_B(net1872),
    .D(_01960_),
    .Q_N(_08029_),
    .Q(\top1.memory2.mem2[109][2] ));
 sg13g2_dfrbp_1 _21864_ (.CLK(\clknet_leaf_223_top1.acquisition_clk ),
    .RESET_B(net1871),
    .D(_01961_),
    .Q_N(_08028_),
    .Q(\top1.memory2.mem2[119][0] ));
 sg13g2_dfrbp_1 _21865_ (.CLK(\clknet_leaf_213_top1.acquisition_clk ),
    .RESET_B(net1870),
    .D(_01962_),
    .Q_N(_08027_),
    .Q(\top1.memory2.mem2[119][1] ));
 sg13g2_dfrbp_1 _21866_ (.CLK(\clknet_leaf_223_top1.acquisition_clk ),
    .RESET_B(net1869),
    .D(_01963_),
    .Q_N(_08026_),
    .Q(\top1.memory2.mem2[119][2] ));
 sg13g2_dfrbp_1 _21867_ (.CLK(\clknet_leaf_66_top1.acquisition_clk ),
    .RESET_B(net1868),
    .D(_01964_),
    .Q_N(_08025_),
    .Q(\top1.memory2.mem2[129][0] ));
 sg13g2_dfrbp_1 _21868_ (.CLK(\clknet_leaf_65_top1.acquisition_clk ),
    .RESET_B(net1867),
    .D(_01965_),
    .Q_N(_08024_),
    .Q(\top1.memory2.mem2[129][1] ));
 sg13g2_dfrbp_1 _21869_ (.CLK(\clknet_leaf_66_top1.acquisition_clk ),
    .RESET_B(net1866),
    .D(_01966_),
    .Q_N(_08023_),
    .Q(\top1.memory2.mem2[129][2] ));
 sg13g2_dfrbp_1 _21870_ (.CLK(\clknet_leaf_67_top1.acquisition_clk ),
    .RESET_B(net1865),
    .D(_01967_),
    .Q_N(_08022_),
    .Q(\top1.memory2.mem2[139][0] ));
 sg13g2_dfrbp_1 _21871_ (.CLK(\clknet_leaf_68_top1.acquisition_clk ),
    .RESET_B(net1864),
    .D(_01968_),
    .Q_N(_08021_),
    .Q(\top1.memory2.mem2[139][1] ));
 sg13g2_dfrbp_1 _21872_ (.CLK(\clknet_leaf_70_top1.acquisition_clk ),
    .RESET_B(net1863),
    .D(_01969_),
    .Q_N(_08020_),
    .Q(\top1.memory2.mem2[139][2] ));
 sg13g2_dfrbp_1 _21873_ (.CLK(\clknet_leaf_76_top1.acquisition_clk ),
    .RESET_B(net1862),
    .D(_01970_),
    .Q_N(_08019_),
    .Q(\top1.memory2.mem2[149][0] ));
 sg13g2_dfrbp_1 _21874_ (.CLK(\clknet_leaf_42_top1.acquisition_clk ),
    .RESET_B(net1861),
    .D(_01971_),
    .Q_N(_08018_),
    .Q(\top1.memory2.mem2[149][1] ));
 sg13g2_dfrbp_1 _21875_ (.CLK(\clknet_leaf_42_top1.acquisition_clk ),
    .RESET_B(net1860),
    .D(_01972_),
    .Q_N(_08017_),
    .Q(\top1.memory2.mem2[149][2] ));
 sg13g2_dfrbp_1 _21876_ (.CLK(\clknet_leaf_71_top1.acquisition_clk ),
    .RESET_B(net1859),
    .D(_01973_),
    .Q_N(_08016_),
    .Q(\top1.memory2.mem2[159][0] ));
 sg13g2_dfrbp_1 _21877_ (.CLK(\clknet_leaf_81_top1.acquisition_clk ),
    .RESET_B(net1858),
    .D(_01974_),
    .Q_N(_08015_),
    .Q(\top1.memory2.mem2[159][1] ));
 sg13g2_dfrbp_1 _21878_ (.CLK(\clknet_leaf_71_top1.acquisition_clk ),
    .RESET_B(net1857),
    .D(_01975_),
    .Q_N(_08014_),
    .Q(\top1.memory2.mem2[159][2] ));
 sg13g2_dfrbp_1 _21879_ (.CLK(\clknet_leaf_107_top1.acquisition_clk ),
    .RESET_B(net1856),
    .D(_01976_),
    .Q_N(_08013_),
    .Q(\top1.memory2.mem2[169][0] ));
 sg13g2_dfrbp_1 _21880_ (.CLK(\clknet_leaf_110_top1.acquisition_clk ),
    .RESET_B(net1855),
    .D(_01977_),
    .Q_N(_08012_),
    .Q(\top1.memory2.mem2[169][1] ));
 sg13g2_dfrbp_1 _21881_ (.CLK(\clknet_leaf_105_top1.acquisition_clk ),
    .RESET_B(net1854),
    .D(_01978_),
    .Q_N(_08011_),
    .Q(\top1.memory2.mem2[169][2] ));
 sg13g2_dfrbp_1 _21882_ (.CLK(\clknet_leaf_134_top1.acquisition_clk ),
    .RESET_B(net1853),
    .D(_01979_),
    .Q_N(_08010_),
    .Q(\top1.memory2.mem2[179][0] ));
 sg13g2_dfrbp_1 _21883_ (.CLK(\clknet_leaf_131_top1.acquisition_clk ),
    .RESET_B(net1852),
    .D(_01980_),
    .Q_N(_08009_),
    .Q(\top1.memory2.mem2[179][1] ));
 sg13g2_dfrbp_1 _21884_ (.CLK(\clknet_leaf_130_top1.acquisition_clk ),
    .RESET_B(net1851),
    .D(_01981_),
    .Q_N(_08008_),
    .Q(\top1.memory2.mem2[179][2] ));
 sg13g2_dfrbp_1 _21885_ (.CLK(\clknet_leaf_117_top1.acquisition_clk ),
    .RESET_B(net1850),
    .D(_01982_),
    .Q_N(_08007_),
    .Q(\top1.memory2.mem2[189][0] ));
 sg13g2_dfrbp_1 _21886_ (.CLK(\clknet_leaf_115_top1.acquisition_clk ),
    .RESET_B(net1849),
    .D(_01983_),
    .Q_N(_08006_),
    .Q(\top1.memory2.mem2[189][1] ));
 sg13g2_dfrbp_1 _21887_ (.CLK(\clknet_leaf_118_top1.acquisition_clk ),
    .RESET_B(net1848),
    .D(_01984_),
    .Q_N(_08005_),
    .Q(\top1.memory2.mem2[189][2] ));
 sg13g2_dfrbp_1 _21888_ (.CLK(\clknet_leaf_41_top1.acquisition_clk ),
    .RESET_B(net1847),
    .D(_01985_),
    .Q_N(_08004_),
    .Q(\top1.memory2.mem2[199][0] ));
 sg13g2_dfrbp_1 _21889_ (.CLK(\clknet_leaf_38_top1.acquisition_clk ),
    .RESET_B(net1846),
    .D(_01986_),
    .Q_N(_08003_),
    .Q(\top1.memory2.mem2[199][1] ));
 sg13g2_dfrbp_1 _21890_ (.CLK(\clknet_leaf_99_top1.acquisition_clk ),
    .RESET_B(net1845),
    .D(_01987_),
    .Q_N(_08002_),
    .Q(\top1.memory2.mem2[199][2] ));
 sg13g2_dfrbp_1 _21891_ (.CLK(\clknet_leaf_88_top1.acquisition_clk ),
    .RESET_B(net1844),
    .D(_01988_),
    .Q_N(_08001_),
    .Q(\top1.memory2.mem2[1][0] ));
 sg13g2_dfrbp_1 _21892_ (.CLK(\clknet_leaf_86_top1.acquisition_clk ),
    .RESET_B(net1843),
    .D(_01989_),
    .Q_N(_08000_),
    .Q(\top1.memory2.mem2[1][1] ));
 sg13g2_dfrbp_1 _21893_ (.CLK(\clknet_leaf_90_top1.acquisition_clk ),
    .RESET_B(net1842),
    .D(_01990_),
    .Q_N(_07999_),
    .Q(\top1.memory2.mem2[1][2] ));
 sg13g2_dfrbp_1 _21894_ (.CLK(\clknet_leaf_111_top1.acquisition_clk ),
    .RESET_B(net1841),
    .D(_01991_),
    .Q_N(_07998_),
    .Q(\top1.memory2.mem2[20][0] ));
 sg13g2_dfrbp_1 _21895_ (.CLK(\clknet_leaf_111_top1.acquisition_clk ),
    .RESET_B(net1840),
    .D(_01992_),
    .Q_N(_07997_),
    .Q(\top1.memory2.mem2[20][1] ));
 sg13g2_dfrbp_1 _21896_ (.CLK(\clknet_leaf_112_top1.acquisition_clk ),
    .RESET_B(net1839),
    .D(_01993_),
    .Q_N(_07996_),
    .Q(\top1.memory2.mem2[20][2] ));
 sg13g2_dfrbp_1 _21897_ (.CLK(\clknet_leaf_111_top1.acquisition_clk ),
    .RESET_B(net1838),
    .D(_01994_),
    .Q_N(_07995_),
    .Q(\top1.memory2.mem2[21][0] ));
 sg13g2_dfrbp_1 _21898_ (.CLK(\clknet_leaf_121_top1.acquisition_clk ),
    .RESET_B(net1837),
    .D(_01995_),
    .Q_N(_07994_),
    .Q(\top1.memory2.mem2[21][1] ));
 sg13g2_dfrbp_1 _21899_ (.CLK(\clknet_leaf_111_top1.acquisition_clk ),
    .RESET_B(net1836),
    .D(_01996_),
    .Q_N(_07993_),
    .Q(\top1.memory2.mem2[21][2] ));
 sg13g2_dfrbp_1 _21900_ (.CLK(\clknet_leaf_110_top1.acquisition_clk ),
    .RESET_B(net1835),
    .D(_01997_),
    .Q_N(_07992_),
    .Q(\top1.memory2.mem2[22][0] ));
 sg13g2_dfrbp_1 _21901_ (.CLK(\clknet_leaf_110_top1.acquisition_clk ),
    .RESET_B(net1834),
    .D(_01998_),
    .Q_N(_07991_),
    .Q(\top1.memory2.mem2[22][1] ));
 sg13g2_dfrbp_1 _21902_ (.CLK(\clknet_leaf_110_top1.acquisition_clk ),
    .RESET_B(net1833),
    .D(_01999_),
    .Q_N(_07990_),
    .Q(\top1.memory2.mem2[22][2] ));
 sg13g2_dfrbp_1 _21903_ (.CLK(\clknet_leaf_112_top1.acquisition_clk ),
    .RESET_B(net1832),
    .D(_02000_),
    .Q_N(_07989_),
    .Q(\top1.memory2.mem2[23][0] ));
 sg13g2_dfrbp_1 _21904_ (.CLK(\clknet_leaf_111_top1.acquisition_clk ),
    .RESET_B(net1831),
    .D(_02001_),
    .Q_N(_07988_),
    .Q(\top1.memory2.mem2[23][1] ));
 sg13g2_dfrbp_1 _21905_ (.CLK(\clknet_leaf_110_top1.acquisition_clk ),
    .RESET_B(net1830),
    .D(_02002_),
    .Q_N(_07987_),
    .Q(\top1.memory2.mem2[23][2] ));
 sg13g2_dfrbp_1 _21906_ (.CLK(\clknet_leaf_124_top1.acquisition_clk ),
    .RESET_B(net1829),
    .D(_02003_),
    .Q_N(_07986_),
    .Q(\top1.memory2.mem2[24][0] ));
 sg13g2_dfrbp_1 _21907_ (.CLK(\clknet_leaf_127_top1.acquisition_clk ),
    .RESET_B(net1828),
    .D(_02004_),
    .Q_N(_07985_),
    .Q(\top1.memory2.mem2[24][1] ));
 sg13g2_dfrbp_1 _21908_ (.CLK(\clknet_leaf_127_top1.acquisition_clk ),
    .RESET_B(net1827),
    .D(_02005_),
    .Q_N(_07984_),
    .Q(\top1.memory2.mem2[24][2] ));
 sg13g2_dfrbp_1 _21909_ (.CLK(\clknet_leaf_124_top1.acquisition_clk ),
    .RESET_B(net1826),
    .D(_02006_),
    .Q_N(_07983_),
    .Q(\top1.memory2.mem2[25][0] ));
 sg13g2_dfrbp_1 _21910_ (.CLK(\clknet_leaf_126_top1.acquisition_clk ),
    .RESET_B(net1825),
    .D(_02007_),
    .Q_N(_07982_),
    .Q(\top1.memory2.mem2[25][1] ));
 sg13g2_dfrbp_1 _21911_ (.CLK(\clknet_leaf_123_top1.acquisition_clk ),
    .RESET_B(net1824),
    .D(_02008_),
    .Q_N(_07981_),
    .Q(\top1.memory2.mem2[25][2] ));
 sg13g2_dfrbp_1 _21912_ (.CLK(\clknet_leaf_125_top1.acquisition_clk ),
    .RESET_B(net1823),
    .D(_02009_),
    .Q_N(_07980_),
    .Q(\top1.memory2.mem2[26][0] ));
 sg13g2_dfrbp_1 _21913_ (.CLK(\clknet_leaf_127_top1.acquisition_clk ),
    .RESET_B(net1822),
    .D(_02010_),
    .Q_N(_07979_),
    .Q(\top1.memory2.mem2[26][1] ));
 sg13g2_dfrbp_1 _21914_ (.CLK(\clknet_leaf_127_top1.acquisition_clk ),
    .RESET_B(net1821),
    .D(_02011_),
    .Q_N(_07978_),
    .Q(\top1.memory2.mem2[26][2] ));
 sg13g2_dfrbp_1 _21915_ (.CLK(\clknet_leaf_124_top1.acquisition_clk ),
    .RESET_B(net1820),
    .D(_02012_),
    .Q_N(_07977_),
    .Q(\top1.memory2.mem2[27][0] ));
 sg13g2_dfrbp_1 _21916_ (.CLK(\clknet_leaf_127_top1.acquisition_clk ),
    .RESET_B(net1819),
    .D(_02013_),
    .Q_N(_07976_),
    .Q(\top1.memory2.mem2[27][1] ));
 sg13g2_dfrbp_1 _21917_ (.CLK(\clknet_leaf_126_top1.acquisition_clk ),
    .RESET_B(net1818),
    .D(_02014_),
    .Q_N(_07975_),
    .Q(\top1.memory2.mem2[27][2] ));
 sg13g2_dfrbp_1 _21918_ (.CLK(\clknet_leaf_124_top1.acquisition_clk ),
    .RESET_B(net1817),
    .D(_02015_),
    .Q_N(_07974_),
    .Q(\top1.memory2.mem2[28][0] ));
 sg13g2_dfrbp_1 _21919_ (.CLK(\clknet_leaf_125_top1.acquisition_clk ),
    .RESET_B(net1816),
    .D(_02016_),
    .Q_N(_07973_),
    .Q(\top1.memory2.mem2[28][1] ));
 sg13g2_dfrbp_1 _21920_ (.CLK(\clknet_leaf_89_top1.acquisition_clk ),
    .RESET_B(net1815),
    .D(_02017_),
    .Q_N(_07972_),
    .Q(\top1.memory2.mem2[28][2] ));
 sg13g2_dfrbp_1 _21921_ (.CLK(\clknet_leaf_89_top1.acquisition_clk ),
    .RESET_B(net1814),
    .D(_02018_),
    .Q_N(_07971_),
    .Q(\top1.memory2.mem2[2][0] ));
 sg13g2_dfrbp_1 _21922_ (.CLK(\clknet_leaf_87_top1.acquisition_clk ),
    .RESET_B(net1813),
    .D(_02019_),
    .Q_N(_07970_),
    .Q(\top1.memory2.mem2[2][1] ));
 sg13g2_dfrbp_1 _21923_ (.CLK(\clknet_leaf_91_top1.acquisition_clk ),
    .RESET_B(net1812),
    .D(_02020_),
    .Q_N(_07969_),
    .Q(\top1.memory2.mem2[2][2] ));
 sg13g2_dfrbp_1 _21924_ (.CLK(\clknet_leaf_121_top1.acquisition_clk ),
    .RESET_B(net1811),
    .D(_02021_),
    .Q_N(_07968_),
    .Q(\top1.memory2.mem2[30][0] ));
 sg13g2_dfrbp_1 _21925_ (.CLK(\clknet_leaf_88_top1.acquisition_clk ),
    .RESET_B(net1810),
    .D(_02022_),
    .Q_N(_07967_),
    .Q(\top1.memory2.mem2[30][1] ));
 sg13g2_dfrbp_1 _21926_ (.CLK(\clknet_leaf_91_top1.acquisition_clk ),
    .RESET_B(net1809),
    .D(_02023_),
    .Q_N(_07966_),
    .Q(\top1.memory2.mem2[30][2] ));
 sg13g2_dfrbp_1 _21927_ (.CLK(\clknet_leaf_122_top1.acquisition_clk ),
    .RESET_B(net1808),
    .D(_02024_),
    .Q_N(_07965_),
    .Q(\top1.memory2.mem2[31][0] ));
 sg13g2_dfrbp_1 _21928_ (.CLK(\clknet_leaf_125_top1.acquisition_clk ),
    .RESET_B(net1807),
    .D(_02025_),
    .Q_N(_07964_),
    .Q(\top1.memory2.mem2[31][1] ));
 sg13g2_dfrbp_1 _21929_ (.CLK(\clknet_leaf_92_top1.acquisition_clk ),
    .RESET_B(net1806),
    .D(_02026_),
    .Q_N(_07963_),
    .Q(\top1.memory2.mem2[31][2] ));
 sg13g2_dfrbp_1 _21930_ (.CLK(\clknet_leaf_176_top1.acquisition_clk ),
    .RESET_B(net1805),
    .D(_02027_),
    .Q_N(_07962_),
    .Q(\top1.memory2.mem2[32][0] ));
 sg13g2_dfrbp_1 _21931_ (.CLK(\clknet_leaf_178_top1.acquisition_clk ),
    .RESET_B(net1804),
    .D(_02028_),
    .Q_N(_07961_),
    .Q(\top1.memory2.mem2[32][1] ));
 sg13g2_dfrbp_1 _21932_ (.CLK(\clknet_leaf_176_top1.acquisition_clk ),
    .RESET_B(net1803),
    .D(_02029_),
    .Q_N(_07960_),
    .Q(\top1.memory2.mem2[32][2] ));
 sg13g2_dfrbp_1 _21933_ (.CLK(\clknet_leaf_176_top1.acquisition_clk ),
    .RESET_B(net1802),
    .D(_02030_),
    .Q_N(_07959_),
    .Q(\top1.memory2.mem2[33][0] ));
 sg13g2_dfrbp_1 _21934_ (.CLK(\clknet_leaf_178_top1.acquisition_clk ),
    .RESET_B(net1801),
    .D(_02031_),
    .Q_N(_07958_),
    .Q(\top1.memory2.mem2[33][1] ));
 sg13g2_dfrbp_1 _21935_ (.CLK(\clknet_leaf_176_top1.acquisition_clk ),
    .RESET_B(net1800),
    .D(_02032_),
    .Q_N(_07957_),
    .Q(\top1.memory2.mem2[33][2] ));
 sg13g2_dfrbp_1 _21936_ (.CLK(\clknet_leaf_116_top1.acquisition_clk ),
    .RESET_B(net1799),
    .D(_02033_),
    .Q_N(_07956_),
    .Q(\top1.memory2.mem2[34][0] ));
 sg13g2_dfrbp_1 _21937_ (.CLK(\clknet_leaf_178_top1.acquisition_clk ),
    .RESET_B(net1798),
    .D(_02034_),
    .Q_N(_07955_),
    .Q(\top1.memory2.mem2[34][1] ));
 sg13g2_dfrbp_1 _21938_ (.CLK(\clknet_leaf_175_top1.acquisition_clk ),
    .RESET_B(net1797),
    .D(_02035_),
    .Q_N(_07954_),
    .Q(\top1.memory2.mem2[34][2] ));
 sg13g2_dfrbp_1 _21939_ (.CLK(\clknet_leaf_116_top1.acquisition_clk ),
    .RESET_B(net1796),
    .D(_02036_),
    .Q_N(_07953_),
    .Q(\top1.memory2.mem2[35][0] ));
 sg13g2_dfrbp_1 _21940_ (.CLK(\clknet_leaf_178_top1.acquisition_clk ),
    .RESET_B(net1795),
    .D(_02037_),
    .Q_N(_07952_),
    .Q(\top1.memory2.mem2[35][1] ));
 sg13g2_dfrbp_1 _21941_ (.CLK(\clknet_leaf_175_top1.acquisition_clk ),
    .RESET_B(net1794),
    .D(_02038_),
    .Q_N(_07951_),
    .Q(\top1.memory2.mem2[35][2] ));
 sg13g2_dfrbp_1 _21942_ (.CLK(\clknet_leaf_133_top1.acquisition_clk ),
    .RESET_B(net1793),
    .D(_02039_),
    .Q_N(_07950_),
    .Q(\top1.memory2.mem2[36][0] ));
 sg13g2_dfrbp_1 _21943_ (.CLK(\clknet_leaf_136_top1.acquisition_clk ),
    .RESET_B(net1792),
    .D(_02040_),
    .Q_N(_07949_),
    .Q(\top1.memory2.mem2[36][1] ));
 sg13g2_dfrbp_1 _21944_ (.CLK(\clknet_leaf_117_top1.acquisition_clk ),
    .RESET_B(net1791),
    .D(_02041_),
    .Q_N(_07948_),
    .Q(\top1.memory2.mem2[36][2] ));
 sg13g2_dfrbp_1 _21945_ (.CLK(\clknet_leaf_133_top1.acquisition_clk ),
    .RESET_B(net1790),
    .D(_02042_),
    .Q_N(_07947_),
    .Q(\top1.memory2.mem2[37][0] ));
 sg13g2_dfrbp_1 _21946_ (.CLK(\clknet_leaf_136_top1.acquisition_clk ),
    .RESET_B(net1789),
    .D(_02043_),
    .Q_N(_07946_),
    .Q(\top1.memory2.mem2[37][1] ));
 sg13g2_dfrbp_1 _21947_ (.CLK(\clknet_leaf_117_top1.acquisition_clk ),
    .RESET_B(net1788),
    .D(_02044_),
    .Q_N(_07945_),
    .Q(\top1.memory2.mem2[37][2] ));
 sg13g2_dfrbp_1 _21948_ (.CLK(\clknet_leaf_135_top1.acquisition_clk ),
    .RESET_B(net1787),
    .D(_02045_),
    .Q_N(_07944_),
    .Q(\top1.memory2.mem2[38][0] ));
 sg13g2_dfrbp_1 _21949_ (.CLK(\clknet_leaf_136_top1.acquisition_clk ),
    .RESET_B(net1786),
    .D(_02046_),
    .Q_N(_07943_),
    .Q(\top1.memory2.mem2[38][1] ));
 sg13g2_dfrbp_1 _21950_ (.CLK(\clknet_leaf_116_top1.acquisition_clk ),
    .RESET_B(net1785),
    .D(_02047_),
    .Q_N(_07942_),
    .Q(\top1.memory2.mem2[38][2] ));
 sg13g2_dfrbp_1 _21951_ (.CLK(\clknet_leaf_89_top1.acquisition_clk ),
    .RESET_B(net1784),
    .D(_02048_),
    .Q_N(_07941_),
    .Q(\top1.memory2.mem2[3][0] ));
 sg13g2_dfrbp_1 _21952_ (.CLK(\clknet_leaf_87_top1.acquisition_clk ),
    .RESET_B(net1783),
    .D(_02049_),
    .Q_N(_07940_),
    .Q(\top1.memory2.mem2[3][1] ));
 sg13g2_dfrbp_1 _21953_ (.CLK(\clknet_leaf_91_top1.acquisition_clk ),
    .RESET_B(net1782),
    .D(_02050_),
    .Q_N(_07939_),
    .Q(\top1.memory2.mem2[3][2] ));
 sg13g2_dfrbp_1 _21954_ (.CLK(\clknet_leaf_136_top1.acquisition_clk ),
    .RESET_B(net1781),
    .D(_02051_),
    .Q_N(_07938_),
    .Q(\top1.memory2.mem2[40][0] ));
 sg13g2_dfrbp_1 _21955_ (.CLK(\clknet_leaf_175_top1.acquisition_clk ),
    .RESET_B(net1780),
    .D(_02052_),
    .Q_N(_07937_),
    .Q(\top1.memory2.mem2[40][1] ));
 sg13g2_dfrbp_1 _21956_ (.CLK(\clknet_leaf_174_top1.acquisition_clk ),
    .RESET_B(net1779),
    .D(_02053_),
    .Q_N(_07936_),
    .Q(\top1.memory2.mem2[40][2] ));
 sg13g2_dfrbp_1 _21957_ (.CLK(\clknet_leaf_136_top1.acquisition_clk ),
    .RESET_B(net1778),
    .D(_02054_),
    .Q_N(_07935_),
    .Q(\top1.memory2.mem2[41][0] ));
 sg13g2_dfrbp_1 _21958_ (.CLK(\clknet_leaf_175_top1.acquisition_clk ),
    .RESET_B(net1777),
    .D(_02055_),
    .Q_N(_07934_),
    .Q(\top1.memory2.mem2[41][1] ));
 sg13g2_dfrbp_1 _21959_ (.CLK(\clknet_leaf_174_top1.acquisition_clk ),
    .RESET_B(net1776),
    .D(_02056_),
    .Q_N(_07933_),
    .Q(\top1.memory2.mem2[41][2] ));
 sg13g2_dfrbp_1 _21960_ (.CLK(\clknet_leaf_137_top1.acquisition_clk ),
    .RESET_B(net1775),
    .D(_02057_),
    .Q_N(_07932_),
    .Q(\top1.memory2.mem2[42][0] ));
 sg13g2_dfrbp_1 _21961_ (.CLK(\clknet_leaf_155_top1.acquisition_clk ),
    .RESET_B(net1774),
    .D(_02058_),
    .Q_N(_07931_),
    .Q(\top1.memory2.mem2[42][1] ));
 sg13g2_dfrbp_1 _21962_ (.CLK(\clknet_leaf_174_top1.acquisition_clk ),
    .RESET_B(net1773),
    .D(_02059_),
    .Q_N(_07930_),
    .Q(\top1.memory2.mem2[42][2] ));
 sg13g2_dfrbp_1 _21963_ (.CLK(\clknet_leaf_136_top1.acquisition_clk ),
    .RESET_B(net1772),
    .D(_02060_),
    .Q_N(_07929_),
    .Q(\top1.memory2.mem2[43][0] ));
 sg13g2_dfrbp_1 _21964_ (.CLK(\clknet_leaf_155_top1.acquisition_clk ),
    .RESET_B(net1771),
    .D(_02061_),
    .Q_N(_07928_),
    .Q(\top1.memory2.mem2[43][1] ));
 sg13g2_dfrbp_1 _21965_ (.CLK(\clknet_leaf_174_top1.acquisition_clk ),
    .RESET_B(net1770),
    .D(_02062_),
    .Q_N(_07927_),
    .Q(\top1.memory2.mem2[43][2] ));
 sg13g2_dfrbp_1 _21966_ (.CLK(\clknet_leaf_133_top1.acquisition_clk ),
    .RESET_B(net1769),
    .D(_02063_),
    .Q_N(_07926_),
    .Q(\top1.memory2.mem2[44][0] ));
 sg13g2_dfrbp_1 _21967_ (.CLK(\clknet_leaf_142_top1.acquisition_clk ),
    .RESET_B(net1768),
    .D(_02064_),
    .Q_N(_07925_),
    .Q(\top1.memory2.mem2[44][1] ));
 sg13g2_dfrbp_1 _21968_ (.CLK(\clknet_leaf_132_top1.acquisition_clk ),
    .RESET_B(net1767),
    .D(_02065_),
    .Q_N(_07924_),
    .Q(\top1.memory2.mem2[44][2] ));
 sg13g2_dfrbp_1 _21969_ (.CLK(\clknet_leaf_135_top1.acquisition_clk ),
    .RESET_B(net1766),
    .D(_02066_),
    .Q_N(_07923_),
    .Q(\top1.memory2.mem2[45][0] ));
 sg13g2_dfrbp_1 _21970_ (.CLK(\clknet_leaf_142_top1.acquisition_clk ),
    .RESET_B(net1765),
    .D(_02067_),
    .Q_N(_07922_),
    .Q(\top1.memory2.mem2[45][1] ));
 sg13g2_dfrbp_1 _21971_ (.CLK(\clknet_leaf_132_top1.acquisition_clk ),
    .RESET_B(net1764),
    .D(_02068_),
    .Q_N(_07921_),
    .Q(\top1.memory2.mem2[45][2] ));
 sg13g2_dfrbp_1 _21972_ (.CLK(\clknet_leaf_133_top1.acquisition_clk ),
    .RESET_B(net1763),
    .D(_02069_),
    .Q_N(_07920_),
    .Q(\top1.memory2.mem2[46][0] ));
 sg13g2_dfrbp_1 _21973_ (.CLK(\clknet_leaf_142_top1.acquisition_clk ),
    .RESET_B(net1762),
    .D(_02070_),
    .Q_N(_07919_),
    .Q(\top1.memory2.mem2[46][1] ));
 sg13g2_dfrbp_1 _21974_ (.CLK(\clknet_leaf_133_top1.acquisition_clk ),
    .RESET_B(net1761),
    .D(_02071_),
    .Q_N(_07918_),
    .Q(\top1.memory2.mem2[46][2] ));
 sg13g2_dfrbp_1 _21975_ (.CLK(\clknet_leaf_133_top1.acquisition_clk ),
    .RESET_B(net1760),
    .D(_02072_),
    .Q_N(_07917_),
    .Q(\top1.memory2.mem2[47][0] ));
 sg13g2_dfrbp_1 _21976_ (.CLK(\clknet_leaf_142_top1.acquisition_clk ),
    .RESET_B(net1759),
    .D(_02073_),
    .Q_N(_07916_),
    .Q(\top1.memory2.mem2[47][1] ));
 sg13g2_dfrbp_1 _21977_ (.CLK(\clknet_leaf_132_top1.acquisition_clk ),
    .RESET_B(net1758),
    .D(_02074_),
    .Q_N(_07915_),
    .Q(\top1.memory2.mem2[47][2] ));
 sg13g2_dfrbp_1 _21978_ (.CLK(\clknet_leaf_139_top1.acquisition_clk ),
    .RESET_B(net1757),
    .D(_02075_),
    .Q_N(_07914_),
    .Q(\top1.memory2.mem2[48][0] ));
 sg13g2_dfrbp_1 _21979_ (.CLK(\clknet_leaf_143_top1.acquisition_clk ),
    .RESET_B(net1756),
    .D(_02076_),
    .Q_N(_07913_),
    .Q(\top1.memory2.mem2[48][1] ));
 sg13g2_dfrbp_1 _21980_ (.CLK(\clknet_leaf_141_top1.acquisition_clk ),
    .RESET_B(net1755),
    .D(_02077_),
    .Q_N(_07912_),
    .Q(\top1.memory2.mem2[48][2] ));
 sg13g2_dfrbp_1 _21981_ (.CLK(\clknet_leaf_100_top1.acquisition_clk ),
    .RESET_B(net1754),
    .D(_02078_),
    .Q_N(_07911_),
    .Q(\top1.memory2.mem2[4][0] ));
 sg13g2_dfrbp_1 _21982_ (.CLK(\clknet_leaf_90_top1.acquisition_clk ),
    .RESET_B(net1753),
    .D(_02079_),
    .Q_N(_07910_),
    .Q(\top1.memory2.mem2[4][1] ));
 sg13g2_dfrbp_1 _21983_ (.CLK(\clknet_leaf_93_top1.acquisition_clk ),
    .RESET_B(net1752),
    .D(_02080_),
    .Q_N(_07909_),
    .Q(\top1.memory2.mem2[4][2] ));
 sg13g2_dfrbp_1 _21984_ (.CLK(\clknet_leaf_139_top1.acquisition_clk ),
    .RESET_B(net1751),
    .D(_02081_),
    .Q_N(_07908_),
    .Q(\top1.memory2.mem2[50][0] ));
 sg13g2_dfrbp_1 _21985_ (.CLK(\clknet_leaf_143_top1.acquisition_clk ),
    .RESET_B(net1750),
    .D(_02082_),
    .Q_N(_07907_),
    .Q(\top1.memory2.mem2[50][1] ));
 sg13g2_dfrbp_1 _21986_ (.CLK(\clknet_leaf_140_top1.acquisition_clk ),
    .RESET_B(net1749),
    .D(_02083_),
    .Q_N(_07906_),
    .Q(\top1.memory2.mem2[50][2] ));
 sg13g2_dfrbp_1 _21987_ (.CLK(\clknet_leaf_140_top1.acquisition_clk ),
    .RESET_B(net1748),
    .D(_02084_),
    .Q_N(_07905_),
    .Q(\top1.memory2.mem2[51][0] ));
 sg13g2_dfrbp_1 _21988_ (.CLK(\clknet_leaf_143_top1.acquisition_clk ),
    .RESET_B(net1747),
    .D(_02085_),
    .Q_N(_07904_),
    .Q(\top1.memory2.mem2[51][1] ));
 sg13g2_dfrbp_1 _21989_ (.CLK(\clknet_leaf_140_top1.acquisition_clk ),
    .RESET_B(net1746),
    .D(_02086_),
    .Q_N(_07903_),
    .Q(\top1.memory2.mem2[51][2] ));
 sg13g2_dfrbp_1 _21990_ (.CLK(\clknet_leaf_138_top1.acquisition_clk ),
    .RESET_B(net1745),
    .D(_02087_),
    .Q_N(_07902_),
    .Q(\top1.memory2.mem2[52][0] ));
 sg13g2_dfrbp_1 _21991_ (.CLK(\clknet_leaf_173_top1.acquisition_clk ),
    .RESET_B(net1744),
    .D(_02088_),
    .Q_N(_07901_),
    .Q(\top1.memory2.mem2[52][1] ));
 sg13g2_dfrbp_1 _21992_ (.CLK(\clknet_leaf_155_top1.acquisition_clk ),
    .RESET_B(net1743),
    .D(_02089_),
    .Q_N(_07900_),
    .Q(\top1.memory2.mem2[52][2] ));
 sg13g2_dfrbp_1 _21993_ (.CLK(\clknet_leaf_137_top1.acquisition_clk ),
    .RESET_B(net1742),
    .D(_02090_),
    .Q_N(_07899_),
    .Q(\top1.memory2.mem2[53][0] ));
 sg13g2_dfrbp_1 _21994_ (.CLK(\clknet_leaf_174_top1.acquisition_clk ),
    .RESET_B(net1741),
    .D(_02091_),
    .Q_N(_07898_),
    .Q(\top1.memory2.mem2[53][1] ));
 sg13g2_dfrbp_1 _21995_ (.CLK(\clknet_leaf_155_top1.acquisition_clk ),
    .RESET_B(net1740),
    .D(_02092_),
    .Q_N(_07897_),
    .Q(\top1.memory2.mem2[53][2] ));
 sg13g2_dfrbp_1 _21996_ (.CLK(\clknet_leaf_138_top1.acquisition_clk ),
    .RESET_B(net1739),
    .D(_02093_),
    .Q_N(_07896_),
    .Q(\top1.memory2.mem2[54][0] ));
 sg13g2_dfrbp_1 _21997_ (.CLK(\clknet_leaf_173_top1.acquisition_clk ),
    .RESET_B(net1738),
    .D(_02094_),
    .Q_N(_07895_),
    .Q(\top1.memory2.mem2[54][1] ));
 sg13g2_dfrbp_1 _21998_ (.CLK(\clknet_leaf_155_top1.acquisition_clk ),
    .RESET_B(net1737),
    .D(_02095_),
    .Q_N(_07894_),
    .Q(\top1.memory2.mem2[54][2] ));
 sg13g2_dfrbp_1 _21999_ (.CLK(\clknet_leaf_138_top1.acquisition_clk ),
    .RESET_B(net1736),
    .D(_02096_),
    .Q_N(_07893_),
    .Q(\top1.memory2.mem2[55][0] ));
 sg13g2_dfrbp_1 _22000_ (.CLK(\clknet_leaf_155_top1.acquisition_clk ),
    .RESET_B(net1735),
    .D(_02097_),
    .Q_N(_07892_),
    .Q(\top1.memory2.mem2[55][1] ));
 sg13g2_dfrbp_1 _22001_ (.CLK(\clknet_leaf_155_top1.acquisition_clk ),
    .RESET_B(net1734),
    .D(_02098_),
    .Q_N(_07891_),
    .Q(\top1.memory2.mem2[55][2] ));
 sg13g2_dfrbp_1 _22002_ (.CLK(\clknet_leaf_157_top1.acquisition_clk ),
    .RESET_B(net1733),
    .D(_02099_),
    .Q_N(_07890_),
    .Q(\top1.memory2.mem2[56][0] ));
 sg13g2_dfrbp_1 _22003_ (.CLK(\clknet_leaf_156_top1.acquisition_clk ),
    .RESET_B(net1732),
    .D(_02100_),
    .Q_N(_07889_),
    .Q(\top1.memory2.mem2[56][1] ));
 sg13g2_dfrbp_1 _22004_ (.CLK(\clknet_leaf_156_top1.acquisition_clk ),
    .RESET_B(net1731),
    .D(_02101_),
    .Q_N(_07888_),
    .Q(\top1.memory2.mem2[56][2] ));
 sg13g2_dfrbp_1 _22005_ (.CLK(\clknet_leaf_157_top1.acquisition_clk ),
    .RESET_B(net1730),
    .D(_02102_),
    .Q_N(_07887_),
    .Q(\top1.memory2.mem2[57][0] ));
 sg13g2_dfrbp_1 _22006_ (.CLK(\clknet_leaf_156_top1.acquisition_clk ),
    .RESET_B(net1729),
    .D(_02103_),
    .Q_N(_07886_),
    .Q(\top1.memory2.mem2[57][1] ));
 sg13g2_dfrbp_1 _22007_ (.CLK(\clknet_leaf_156_top1.acquisition_clk ),
    .RESET_B(net1728),
    .D(_02104_),
    .Q_N(_07885_),
    .Q(\top1.memory2.mem2[57][2] ));
 sg13g2_dfrbp_1 _22008_ (.CLK(\clknet_leaf_157_top1.acquisition_clk ),
    .RESET_B(net1727),
    .D(_02105_),
    .Q_N(_07884_),
    .Q(\top1.memory2.mem2[58][0] ));
 sg13g2_dfrbp_1 _22009_ (.CLK(\clknet_leaf_156_top1.acquisition_clk ),
    .RESET_B(net1726),
    .D(_02106_),
    .Q_N(_07883_),
    .Q(\top1.memory2.mem2[58][1] ));
 sg13g2_dfrbp_1 _22010_ (.CLK(\clknet_leaf_156_top1.acquisition_clk ),
    .RESET_B(net1725),
    .D(_02107_),
    .Q_N(_07882_),
    .Q(\top1.memory2.mem2[58][2] ));
 sg13g2_dfrbp_1 _22011_ (.CLK(\clknet_leaf_100_top1.acquisition_clk ),
    .RESET_B(net1724),
    .D(_02108_),
    .Q_N(_07881_),
    .Q(\top1.memory2.mem2[5][0] ));
 sg13g2_dfrbp_1 _22012_ (.CLK(\clknet_leaf_90_top1.acquisition_clk ),
    .RESET_B(net1723),
    .D(_02109_),
    .Q_N(_07880_),
    .Q(\top1.memory2.mem2[5][1] ));
 sg13g2_dfrbp_1 _22013_ (.CLK(\clknet_leaf_100_top1.acquisition_clk ),
    .RESET_B(net1722),
    .D(_02110_),
    .Q_N(_07879_),
    .Q(\top1.memory2.mem2[5][2] ));
 sg13g2_dfrbp_1 _22014_ (.CLK(\clknet_leaf_144_top1.acquisition_clk ),
    .RESET_B(net1721),
    .D(_02111_),
    .Q_N(_07878_),
    .Q(\top1.memory2.mem2[60][0] ));
 sg13g2_dfrbp_1 _22015_ (.CLK(\clknet_leaf_153_top1.acquisition_clk ),
    .RESET_B(net1720),
    .D(_02112_),
    .Q_N(_07877_),
    .Q(\top1.memory2.mem2[60][1] ));
 sg13g2_dfrbp_1 _22016_ (.CLK(\clknet_leaf_153_top1.acquisition_clk ),
    .RESET_B(net1719),
    .D(_02113_),
    .Q_N(_07876_),
    .Q(\top1.memory2.mem2[60][2] ));
 sg13g2_dfrbp_1 _22017_ (.CLK(\clknet_leaf_144_top1.acquisition_clk ),
    .RESET_B(net1718),
    .D(_02114_),
    .Q_N(_07875_),
    .Q(\top1.memory2.mem2[61][0] ));
 sg13g2_dfrbp_1 _22018_ (.CLK(\clknet_leaf_153_top1.acquisition_clk ),
    .RESET_B(net1717),
    .D(_02115_),
    .Q_N(_07874_),
    .Q(\top1.memory2.mem2[61][1] ));
 sg13g2_dfrbp_1 _22019_ (.CLK(\clknet_leaf_154_top1.acquisition_clk ),
    .RESET_B(net1716),
    .D(_02116_),
    .Q_N(_07873_),
    .Q(\top1.memory2.mem2[61][2] ));
 sg13g2_dfrbp_1 _22020_ (.CLK(\clknet_leaf_144_top1.acquisition_clk ),
    .RESET_B(net1715),
    .D(_02117_),
    .Q_N(_07872_),
    .Q(\top1.memory2.mem2[62][0] ));
 sg13g2_dfrbp_1 _22021_ (.CLK(\clknet_leaf_153_top1.acquisition_clk ),
    .RESET_B(net1714),
    .D(_02118_),
    .Q_N(_07871_),
    .Q(\top1.memory2.mem2[62][1] ));
 sg13g2_dfrbp_1 _22022_ (.CLK(\clknet_leaf_153_top1.acquisition_clk ),
    .RESET_B(net1713),
    .D(_02119_),
    .Q_N(_07870_),
    .Q(\top1.memory2.mem2[62][2] ));
 sg13g2_dfrbp_1 _22023_ (.CLK(\clknet_leaf_144_top1.acquisition_clk ),
    .RESET_B(net1712),
    .D(_02120_),
    .Q_N(_07869_),
    .Q(\top1.memory2.mem2[63][0] ));
 sg13g2_dfrbp_1 _22024_ (.CLK(\clknet_leaf_139_top1.acquisition_clk ),
    .RESET_B(net1711),
    .D(_02121_),
    .Q_N(_07868_),
    .Q(\top1.memory2.mem2[63][1] ));
 sg13g2_dfrbp_1 _22025_ (.CLK(\clknet_leaf_153_top1.acquisition_clk ),
    .RESET_B(net1710),
    .D(_02122_),
    .Q_N(_07867_),
    .Q(\top1.memory2.mem2[63][2] ));
 sg13g2_dfrbp_1 _22026_ (.CLK(\clknet_leaf_300_top1.acquisition_clk ),
    .RESET_B(net1709),
    .D(_02123_),
    .Q_N(_07866_),
    .Q(\top1.memory2.mem2[64][0] ));
 sg13g2_dfrbp_1 _22027_ (.CLK(\clknet_leaf_0_top1.acquisition_clk ),
    .RESET_B(net1708),
    .D(_02124_),
    .Q_N(_07865_),
    .Q(\top1.memory2.mem2[64][1] ));
 sg13g2_dfrbp_1 _22028_ (.CLK(\clknet_leaf_301_top1.acquisition_clk ),
    .RESET_B(net1707),
    .D(_02125_),
    .Q_N(_07864_),
    .Q(\top1.memory2.mem2[64][2] ));
 sg13g2_dfrbp_1 _22029_ (.CLK(\clknet_leaf_301_top1.acquisition_clk ),
    .RESET_B(net1706),
    .D(_02126_),
    .Q_N(_07863_),
    .Q(\top1.memory2.mem2[65][0] ));
 sg13g2_dfrbp_1 _22030_ (.CLK(\clknet_leaf_299_top1.acquisition_clk ),
    .RESET_B(net1705),
    .D(_02127_),
    .Q_N(_07862_),
    .Q(\top1.memory2.mem2[65][1] ));
 sg13g2_dfrbp_1 _22031_ (.CLK(\clknet_leaf_301_top1.acquisition_clk ),
    .RESET_B(net1704),
    .D(_02128_),
    .Q_N(_07861_),
    .Q(\top1.memory2.mem2[65][2] ));
 sg13g2_dfrbp_1 _22032_ (.CLK(\clknet_leaf_301_top1.acquisition_clk ),
    .RESET_B(net1703),
    .D(_02129_),
    .Q_N(_07860_),
    .Q(\top1.memory2.mem2[66][0] ));
 sg13g2_dfrbp_1 _22033_ (.CLK(\clknet_leaf_0_top1.acquisition_clk ),
    .RESET_B(net1702),
    .D(_02130_),
    .Q_N(_07859_),
    .Q(\top1.memory2.mem2[66][1] ));
 sg13g2_dfrbp_1 _22034_ (.CLK(\clknet_leaf_301_top1.acquisition_clk ),
    .RESET_B(net1701),
    .D(_02131_),
    .Q_N(_07858_),
    .Q(\top1.memory2.mem2[66][2] ));
 sg13g2_dfrbp_1 _22035_ (.CLK(\clknet_leaf_300_top1.acquisition_clk ),
    .RESET_B(net1700),
    .D(_02132_),
    .Q_N(_07857_),
    .Q(\top1.memory2.mem2[67][0] ));
 sg13g2_dfrbp_1 _22036_ (.CLK(\clknet_leaf_1_top1.acquisition_clk ),
    .RESET_B(net1699),
    .D(_02133_),
    .Q_N(_07856_),
    .Q(\top1.memory2.mem2[67][1] ));
 sg13g2_dfrbp_1 _22037_ (.CLK(\clknet_leaf_301_top1.acquisition_clk ),
    .RESET_B(net1698),
    .D(_02134_),
    .Q_N(_07855_),
    .Q(\top1.memory2.mem2[67][2] ));
 sg13g2_dfrbp_1 _22038_ (.CLK(\clknet_leaf_292_top1.acquisition_clk ),
    .RESET_B(net1697),
    .D(_02135_),
    .Q_N(_07854_),
    .Q(\top1.memory2.mem2[68][0] ));
 sg13g2_dfrbp_1 _22039_ (.CLK(\clknet_leaf_10_top1.acquisition_clk ),
    .RESET_B(net1696),
    .D(_02136_),
    .Q_N(_07853_),
    .Q(\top1.memory2.mem2[68][1] ));
 sg13g2_dfrbp_1 _22040_ (.CLK(\clknet_leaf_10_top1.acquisition_clk ),
    .RESET_B(net1695),
    .D(_02137_),
    .Q_N(_07852_),
    .Q(\top1.memory2.mem2[68][2] ));
 sg13g2_dfrbp_1 _22041_ (.CLK(\clknet_leaf_93_top1.acquisition_clk ),
    .RESET_B(net1694),
    .D(_02138_),
    .Q_N(_07851_),
    .Q(\top1.memory2.mem2[6][0] ));
 sg13g2_dfrbp_1 _22042_ (.CLK(\clknet_leaf_94_top1.acquisition_clk ),
    .RESET_B(net1693),
    .D(_02139_),
    .Q_N(_07850_),
    .Q(\top1.memory2.mem2[6][1] ));
 sg13g2_dfrbp_1 _22043_ (.CLK(\clknet_leaf_100_top1.acquisition_clk ),
    .RESET_B(net1692),
    .D(_02140_),
    .Q_N(_07849_),
    .Q(\top1.memory2.mem2[6][2] ));
 sg13g2_dfrbp_1 _22044_ (.CLK(\clknet_leaf_292_top1.acquisition_clk ),
    .RESET_B(net1691),
    .D(_02141_),
    .Q_N(_07848_),
    .Q(\top1.memory2.mem2[70][0] ));
 sg13g2_dfrbp_1 _22045_ (.CLK(\clknet_leaf_10_top1.acquisition_clk ),
    .RESET_B(net1690),
    .D(_02142_),
    .Q_N(_07847_),
    .Q(\top1.memory2.mem2[70][1] ));
 sg13g2_dfrbp_1 _22046_ (.CLK(\clknet_leaf_10_top1.acquisition_clk ),
    .RESET_B(net1689),
    .D(_02143_),
    .Q_N(_07846_),
    .Q(\top1.memory2.mem2[70][2] ));
 sg13g2_dfrbp_1 _22047_ (.CLK(\clknet_leaf_292_top1.acquisition_clk ),
    .RESET_B(net1688),
    .D(_02144_),
    .Q_N(_07845_),
    .Q(\top1.memory2.mem2[71][0] ));
 sg13g2_dfrbp_1 _22048_ (.CLK(\clknet_leaf_26_top1.acquisition_clk ),
    .RESET_B(net1687),
    .D(_02145_),
    .Q_N(_07844_),
    .Q(\top1.memory2.mem2[71][1] ));
 sg13g2_dfrbp_1 _22049_ (.CLK(\clknet_leaf_26_top1.acquisition_clk ),
    .RESET_B(net1686),
    .D(_02146_),
    .Q_N(_07843_),
    .Q(\top1.memory2.mem2[71][2] ));
 sg13g2_dfrbp_1 _22050_ (.CLK(\clknet_leaf_297_top1.acquisition_clk ),
    .RESET_B(net1685),
    .D(_02147_),
    .Q_N(_07842_),
    .Q(\top1.memory2.mem2[72][0] ));
 sg13g2_dfrbp_1 _22051_ (.CLK(\clknet_leaf_299_top1.acquisition_clk ),
    .RESET_B(net1684),
    .D(_02148_),
    .Q_N(_07841_),
    .Q(\top1.memory2.mem2[72][1] ));
 sg13g2_dfrbp_1 _22052_ (.CLK(\clknet_leaf_300_top1.acquisition_clk ),
    .RESET_B(net1683),
    .D(_02149_),
    .Q_N(_07840_),
    .Q(\top1.memory2.mem2[72][2] ));
 sg13g2_dfrbp_1 _22053_ (.CLK(\clknet_leaf_297_top1.acquisition_clk ),
    .RESET_B(net1682),
    .D(_02150_),
    .Q_N(_07839_),
    .Q(\top1.memory2.mem2[73][0] ));
 sg13g2_dfrbp_1 _22054_ (.CLK(\clknet_leaf_299_top1.acquisition_clk ),
    .RESET_B(net1681),
    .D(_02151_),
    .Q_N(_07838_),
    .Q(\top1.memory2.mem2[73][1] ));
 sg13g2_dfrbp_1 _22055_ (.CLK(\clknet_leaf_297_top1.acquisition_clk ),
    .RESET_B(net1680),
    .D(_02152_),
    .Q_N(_07837_),
    .Q(\top1.memory2.mem2[73][2] ));
 sg13g2_dfrbp_1 _22056_ (.CLK(\clknet_leaf_297_top1.acquisition_clk ),
    .RESET_B(net1679),
    .D(_02153_),
    .Q_N(_07836_),
    .Q(\top1.memory2.mem2[74][0] ));
 sg13g2_dfrbp_1 _22057_ (.CLK(\clknet_leaf_299_top1.acquisition_clk ),
    .RESET_B(net1678),
    .D(_02154_),
    .Q_N(_07835_),
    .Q(\top1.memory2.mem2[74][1] ));
 sg13g2_dfrbp_1 _22058_ (.CLK(\clknet_leaf_300_top1.acquisition_clk ),
    .RESET_B(net1677),
    .D(_02155_),
    .Q_N(_07834_),
    .Q(\top1.memory2.mem2[74][2] ));
 sg13g2_dfrbp_1 _22059_ (.CLK(\clknet_leaf_296_top1.acquisition_clk ),
    .RESET_B(net1676),
    .D(_02156_),
    .Q_N(_07833_),
    .Q(\top1.memory2.mem2[75][0] ));
 sg13g2_dfrbp_1 _22060_ (.CLK(\clknet_leaf_298_top1.acquisition_clk ),
    .RESET_B(net1675),
    .D(_02157_),
    .Q_N(_07832_),
    .Q(\top1.memory2.mem2[75][1] ));
 sg13g2_dfrbp_1 _22061_ (.CLK(\clknet_leaf_300_top1.acquisition_clk ),
    .RESET_B(net1674),
    .D(_02158_),
    .Q_N(_07831_),
    .Q(\top1.memory2.mem2[75][2] ));
 sg13g2_dfrbp_1 _22062_ (.CLK(\clknet_leaf_302_top1.acquisition_clk ),
    .RESET_B(net1673),
    .D(_02159_),
    .Q_N(_07830_),
    .Q(\top1.memory2.mem2[76][0] ));
 sg13g2_dfrbp_1 _22063_ (.CLK(\clknet_leaf_2_top1.acquisition_clk ),
    .RESET_B(net1672),
    .D(_02160_),
    .Q_N(_07829_),
    .Q(\top1.memory2.mem2[76][1] ));
 sg13g2_dfrbp_1 _22064_ (.CLK(\clknet_leaf_302_top1.acquisition_clk ),
    .RESET_B(net1671),
    .D(_02161_),
    .Q_N(_07828_),
    .Q(\top1.memory2.mem2[76][2] ));
 sg13g2_dfrbp_1 _22065_ (.CLK(\clknet_leaf_0_top1.acquisition_clk ),
    .RESET_B(net1670),
    .D(_02162_),
    .Q_N(_07827_),
    .Q(\top1.memory2.mem2[77][0] ));
 sg13g2_dfrbp_1 _22066_ (.CLK(\clknet_leaf_2_top1.acquisition_clk ),
    .RESET_B(net1669),
    .D(_02163_),
    .Q_N(_07826_),
    .Q(\top1.memory2.mem2[77][1] ));
 sg13g2_dfrbp_1 _22067_ (.CLK(\clknet_leaf_301_top1.acquisition_clk ),
    .RESET_B(net1668),
    .D(_02164_),
    .Q_N(_07825_),
    .Q(\top1.memory2.mem2[77][2] ));
 sg13g2_dfrbp_1 _22068_ (.CLK(\clknet_leaf_302_top1.acquisition_clk ),
    .RESET_B(net1667),
    .D(_02165_),
    .Q_N(_07824_),
    .Q(\top1.memory2.mem2[78][0] ));
 sg13g2_dfrbp_1 _22069_ (.CLK(\clknet_leaf_3_top1.acquisition_clk ),
    .RESET_B(net1666),
    .D(_02166_),
    .Q_N(_07823_),
    .Q(\top1.memory2.mem2[78][1] ));
 sg13g2_dfrbp_1 _22070_ (.CLK(\clknet_leaf_302_top1.acquisition_clk ),
    .RESET_B(net1665),
    .D(_02167_),
    .Q_N(_07822_),
    .Q(\top1.memory2.mem2[78][2] ));
 sg13g2_dfrbp_1 _22071_ (.CLK(\clknet_leaf_100_top1.acquisition_clk ),
    .RESET_B(net1664),
    .D(_02168_),
    .Q_N(_07821_),
    .Q(\top1.memory2.mem2[7][0] ));
 sg13g2_dfrbp_1 _22072_ (.CLK(\clknet_leaf_92_top1.acquisition_clk ),
    .RESET_B(net1663),
    .D(_02169_),
    .Q_N(_07820_),
    .Q(\top1.memory2.mem2[7][1] ));
 sg13g2_dfrbp_1 _22073_ (.CLK(\clknet_leaf_93_top1.acquisition_clk ),
    .RESET_B(net1662),
    .D(_02170_),
    .Q_N(_07819_),
    .Q(\top1.memory2.mem2[7][2] ));
 sg13g2_dfrbp_1 _22074_ (.CLK(\clknet_leaf_295_top1.acquisition_clk ),
    .RESET_B(net1661),
    .D(_02171_),
    .Q_N(_07818_),
    .Q(\top1.memory2.mem2[80][0] ));
 sg13g2_dfrbp_1 _22075_ (.CLK(\clknet_leaf_297_top1.acquisition_clk ),
    .RESET_B(net1660),
    .D(_02172_),
    .Q_N(_07817_),
    .Q(\top1.memory2.mem2[80][1] ));
 sg13g2_dfrbp_1 _22076_ (.CLK(\clknet_leaf_296_top1.acquisition_clk ),
    .RESET_B(net1659),
    .D(_02173_),
    .Q_N(_07816_),
    .Q(\top1.memory2.mem2[80][2] ));
 sg13g2_dfrbp_1 _22077_ (.CLK(\clknet_leaf_295_top1.acquisition_clk ),
    .RESET_B(net1658),
    .D(_02174_),
    .Q_N(_07815_),
    .Q(\top1.memory2.mem2[81][0] ));
 sg13g2_dfrbp_1 _22078_ (.CLK(\clknet_leaf_297_top1.acquisition_clk ),
    .RESET_B(net1657),
    .D(_02175_),
    .Q_N(_07814_),
    .Q(\top1.memory2.mem2[81][1] ));
 sg13g2_dfrbp_1 _22079_ (.CLK(\clknet_leaf_296_top1.acquisition_clk ),
    .RESET_B(net1656),
    .D(_02176_),
    .Q_N(_07813_),
    .Q(\top1.memory2.mem2[81][2] ));
 sg13g2_dfrbp_1 _22080_ (.CLK(\clknet_leaf_294_top1.acquisition_clk ),
    .RESET_B(net1655),
    .D(_02177_),
    .Q_N(_07812_),
    .Q(\top1.memory2.mem2[82][0] ));
 sg13g2_dfrbp_1 _22081_ (.CLK(\clknet_leaf_297_top1.acquisition_clk ),
    .RESET_B(net1654),
    .D(_02178_),
    .Q_N(_07811_),
    .Q(\top1.memory2.mem2[82][1] ));
 sg13g2_dfrbp_1 _22082_ (.CLK(\clknet_leaf_296_top1.acquisition_clk ),
    .RESET_B(net1653),
    .D(_02179_),
    .Q_N(_07810_),
    .Q(\top1.memory2.mem2[82][2] ));
 sg13g2_dfrbp_1 _22083_ (.CLK(\clknet_leaf_295_top1.acquisition_clk ),
    .RESET_B(net1652),
    .D(_02180_),
    .Q_N(_07809_),
    .Q(\top1.memory2.mem2[83][0] ));
 sg13g2_dfrbp_1 _22084_ (.CLK(\clknet_leaf_293_top1.acquisition_clk ),
    .RESET_B(net1651),
    .D(_02181_),
    .Q_N(_07808_),
    .Q(\top1.memory2.mem2[83][1] ));
 sg13g2_dfrbp_1 _22085_ (.CLK(\clknet_leaf_296_top1.acquisition_clk ),
    .RESET_B(net1650),
    .D(_02182_),
    .Q_N(_07807_),
    .Q(\top1.memory2.mem2[83][2] ));
 sg13g2_dfrbp_1 _22086_ (.CLK(\clknet_leaf_28_top1.acquisition_clk ),
    .RESET_B(net1649),
    .D(_02183_),
    .Q_N(_07806_),
    .Q(\top1.memory2.mem2[84][0] ));
 sg13g2_dfrbp_1 _22087_ (.CLK(\clknet_leaf_9_top1.acquisition_clk ),
    .RESET_B(net1648),
    .D(_02184_),
    .Q_N(_07805_),
    .Q(\top1.memory2.mem2[84][1] ));
 sg13g2_dfrbp_1 _22088_ (.CLK(\clknet_leaf_9_top1.acquisition_clk ),
    .RESET_B(net1647),
    .D(_02185_),
    .Q_N(_07804_),
    .Q(\top1.memory2.mem2[84][2] ));
 sg13g2_dfrbp_1 _22089_ (.CLK(\clknet_leaf_28_top1.acquisition_clk ),
    .RESET_B(net1646),
    .D(_02186_),
    .Q_N(_07803_),
    .Q(\top1.memory2.mem2[85][0] ));
 sg13g2_dfrbp_1 _22090_ (.CLK(\clknet_leaf_26_top1.acquisition_clk ),
    .RESET_B(net1645),
    .D(_02187_),
    .Q_N(_07802_),
    .Q(\top1.memory2.mem2[85][1] ));
 sg13g2_dfrbp_1 _22091_ (.CLK(\clknet_leaf_26_top1.acquisition_clk ),
    .RESET_B(net1644),
    .D(_02188_),
    .Q_N(_07801_),
    .Q(\top1.memory2.mem2[85][2] ));
 sg13g2_dfrbp_1 _22092_ (.CLK(\clknet_leaf_25_top1.acquisition_clk ),
    .RESET_B(net1643),
    .D(_02189_),
    .Q_N(_07800_),
    .Q(\top1.memory2.mem2[86][0] ));
 sg13g2_dfrbp_1 _22093_ (.CLK(\clknet_leaf_27_top1.acquisition_clk ),
    .RESET_B(net1642),
    .D(_02190_),
    .Q_N(_07799_),
    .Q(\top1.memory2.mem2[86][1] ));
 sg13g2_dfrbp_1 _22094_ (.CLK(\clknet_leaf_28_top1.acquisition_clk ),
    .RESET_B(net1641),
    .D(_02191_),
    .Q_N(_07798_),
    .Q(\top1.memory2.mem2[86][2] ));
 sg13g2_dfrbp_1 _22095_ (.CLK(\clknet_leaf_27_top1.acquisition_clk ),
    .RESET_B(net1640),
    .D(_02192_),
    .Q_N(_07797_),
    .Q(\top1.memory2.mem2[87][0] ));
 sg13g2_dfrbp_1 _22096_ (.CLK(\clknet_leaf_27_top1.acquisition_clk ),
    .RESET_B(net1639),
    .D(_02193_),
    .Q_N(_07796_),
    .Q(\top1.memory2.mem2[87][1] ));
 sg13g2_dfrbp_1 _22097_ (.CLK(\clknet_leaf_26_top1.acquisition_clk ),
    .RESET_B(net1638),
    .D(_02194_),
    .Q_N(_07795_),
    .Q(\top1.memory2.mem2[87][2] ));
 sg13g2_dfrbp_1 _22098_ (.CLK(\clknet_leaf_9_top1.acquisition_clk ),
    .RESET_B(net1637),
    .D(_02195_),
    .Q_N(_07794_),
    .Q(\top1.memory2.mem2[88][0] ));
 sg13g2_dfrbp_1 _22099_ (.CLK(\clknet_leaf_7_top1.acquisition_clk ),
    .RESET_B(net1636),
    .D(_02196_),
    .Q_N(_07793_),
    .Q(\top1.memory2.mem2[88][1] ));
 sg13g2_dfrbp_1 _22100_ (.CLK(\clknet_leaf_8_top1.acquisition_clk ),
    .RESET_B(net1635),
    .D(_02197_),
    .Q_N(_07792_),
    .Q(\top1.memory2.mem2[88][2] ));
 sg13g2_dfrbp_1 _22101_ (.CLK(\clknet_leaf_94_top1.acquisition_clk ),
    .RESET_B(net1634),
    .D(_02198_),
    .Q_N(_07791_),
    .Q(\top1.memory2.mem2[8][0] ));
 sg13g2_dfrbp_1 _22102_ (.CLK(\clknet_leaf_86_top1.acquisition_clk ),
    .RESET_B(net1633),
    .D(_02199_),
    .Q_N(_07790_),
    .Q(\top1.memory2.mem2[8][1] ));
 sg13g2_dfrbp_1 _22103_ (.CLK(\clknet_leaf_84_top1.acquisition_clk ),
    .RESET_B(net1632),
    .D(_02200_),
    .Q_N(_07789_),
    .Q(\top1.memory2.mem2[8][2] ));
 sg13g2_dfrbp_1 _22104_ (.CLK(\clknet_leaf_290_top1.acquisition_clk ),
    .RESET_B(net1631),
    .D(_02201_),
    .Q_N(_07788_),
    .Q(\top1.memory2.mem2[90][0] ));
 sg13g2_dfrbp_1 _22105_ (.CLK(\clknet_leaf_292_top1.acquisition_clk ),
    .RESET_B(net1630),
    .D(_02202_),
    .Q_N(_07787_),
    .Q(\top1.memory2.mem2[90][1] ));
 sg13g2_dfrbp_1 _22106_ (.CLK(\clknet_leaf_8_top1.acquisition_clk ),
    .RESET_B(net1629),
    .D(_02203_),
    .Q_N(_07786_),
    .Q(\top1.memory2.mem2[90][2] ));
 sg13g2_dfrbp_1 _22107_ (.CLK(\clknet_leaf_269_top1.acquisition_clk ),
    .RESET_B(net1628),
    .D(_02204_),
    .Q_N(_07785_),
    .Q(\top1.memory2.mem2[91][0] ));
 sg13g2_dfrbp_1 _22108_ (.CLK(\clknet_leaf_291_top1.acquisition_clk ),
    .RESET_B(net1627),
    .D(_02205_),
    .Q_N(_07784_),
    .Q(\top1.memory2.mem2[91][1] ));
 sg13g2_dfrbp_1 _22109_ (.CLK(\clknet_leaf_8_top1.acquisition_clk ),
    .RESET_B(net1626),
    .D(_02206_),
    .Q_N(_07783_),
    .Q(\top1.memory2.mem2[91][2] ));
 sg13g2_dfrbp_1 _22110_ (.CLK(\clknet_leaf_294_top1.acquisition_clk ),
    .RESET_B(net1625),
    .D(_02207_),
    .Q_N(_07782_),
    .Q(\top1.memory2.mem2[92][0] ));
 sg13g2_dfrbp_1 _22111_ (.CLK(\clknet_leaf_291_top1.acquisition_clk ),
    .RESET_B(net1624),
    .D(_02208_),
    .Q_N(_07781_),
    .Q(\top1.memory2.mem2[92][1] ));
 sg13g2_dfrbp_1 _22112_ (.CLK(\clknet_leaf_291_top1.acquisition_clk ),
    .RESET_B(net1623),
    .D(_02209_),
    .Q_N(_07780_),
    .Q(\top1.memory2.mem2[92][2] ));
 sg13g2_dfrbp_1 _22113_ (.CLK(\clknet_leaf_294_top1.acquisition_clk ),
    .RESET_B(net1622),
    .D(_02210_),
    .Q_N(_07779_),
    .Q(\top1.memory2.mem2[93][0] ));
 sg13g2_dfrbp_1 _22114_ (.CLK(\clknet_leaf_291_top1.acquisition_clk ),
    .RESET_B(net1621),
    .D(_02211_),
    .Q_N(_07778_),
    .Q(\top1.memory2.mem2[93][1] ));
 sg13g2_dfrbp_1 _22115_ (.CLK(\clknet_leaf_291_top1.acquisition_clk ),
    .RESET_B(net1620),
    .D(_02212_),
    .Q_N(_07777_),
    .Q(\top1.memory2.mem2[93][2] ));
 sg13g2_dfrbp_1 _22116_ (.CLK(\clknet_leaf_294_top1.acquisition_clk ),
    .RESET_B(net1619),
    .D(_02213_),
    .Q_N(_07776_),
    .Q(\top1.memory2.mem2[94][0] ));
 sg13g2_dfrbp_1 _22117_ (.CLK(\clknet_leaf_293_top1.acquisition_clk ),
    .RESET_B(net1618),
    .D(_02214_),
    .Q_N(_07775_),
    .Q(\top1.memory2.mem2[94][1] ));
 sg13g2_dfrbp_1 _22118_ (.CLK(\clknet_leaf_293_top1.acquisition_clk ),
    .RESET_B(net1617),
    .D(_02215_),
    .Q_N(_07774_),
    .Q(\top1.memory2.mem2[94][2] ));
 sg13g2_dfrbp_1 _22119_ (.CLK(\clknet_leaf_294_top1.acquisition_clk ),
    .RESET_B(net1616),
    .D(_02216_),
    .Q_N(_07773_),
    .Q(\top1.memory2.mem2[95][0] ));
 sg13g2_dfrbp_1 _22120_ (.CLK(\clknet_leaf_293_top1.acquisition_clk ),
    .RESET_B(net1615),
    .D(_02217_),
    .Q_N(_07772_),
    .Q(\top1.memory2.mem2[95][1] ));
 sg13g2_dfrbp_1 _22121_ (.CLK(\clknet_leaf_291_top1.acquisition_clk ),
    .RESET_B(net1614),
    .D(_02218_),
    .Q_N(_07771_),
    .Q(\top1.memory2.mem2[95][2] ));
 sg13g2_dfrbp_1 _22122_ (.CLK(\clknet_leaf_231_top1.acquisition_clk ),
    .RESET_B(net1613),
    .D(_02219_),
    .Q_N(_07770_),
    .Q(\top1.memory2.mem2[96][0] ));
 sg13g2_dfrbp_1 _22123_ (.CLK(\clknet_leaf_232_top1.acquisition_clk ),
    .RESET_B(net1612),
    .D(_02220_),
    .Q_N(_07769_),
    .Q(\top1.memory2.mem2[96][1] ));
 sg13g2_dfrbp_1 _22124_ (.CLK(\clknet_leaf_231_top1.acquisition_clk ),
    .RESET_B(net1611),
    .D(_02221_),
    .Q_N(_07768_),
    .Q(\top1.memory2.mem2[96][2] ));
 sg13g2_dfrbp_1 _22125_ (.CLK(\clknet_leaf_231_top1.acquisition_clk ),
    .RESET_B(net1610),
    .D(_02222_),
    .Q_N(_07767_),
    .Q(\top1.memory2.mem2[97][0] ));
 sg13g2_dfrbp_1 _22126_ (.CLK(\clknet_leaf_233_top1.acquisition_clk ),
    .RESET_B(net1609),
    .D(_02223_),
    .Q_N(_07766_),
    .Q(\top1.memory2.mem2[97][1] ));
 sg13g2_dfrbp_1 _22127_ (.CLK(\clknet_leaf_230_top1.acquisition_clk ),
    .RESET_B(net1608),
    .D(_02224_),
    .Q_N(_07765_),
    .Q(\top1.memory2.mem2[97][2] ));
 sg13g2_dfrbp_1 _22128_ (.CLK(\clknet_leaf_231_top1.acquisition_clk ),
    .RESET_B(net1607),
    .D(_02225_),
    .Q_N(_07764_),
    .Q(\top1.memory2.mem2[98][0] ));
 sg13g2_dfrbp_1 _22129_ (.CLK(\clknet_leaf_233_top1.acquisition_clk ),
    .RESET_B(net1606),
    .D(_02226_),
    .Q_N(_07763_),
    .Q(\top1.memory2.mem2[98][1] ));
 sg13g2_dfrbp_1 _22130_ (.CLK(\clknet_leaf_230_top1.acquisition_clk ),
    .RESET_B(net1605),
    .D(_02227_),
    .Q_N(_07762_),
    .Q(\top1.memory2.mem2[98][2] ));
 sg13g2_dfrbp_1 _22131_ (.CLK(\clknet_leaf_89_top1.acquisition_clk ),
    .RESET_B(net1604),
    .D(_02228_),
    .Q_N(_07761_),
    .Q(\top1.memory2.mem2[0][0] ));
 sg13g2_dfrbp_1 _22132_ (.CLK(\clknet_leaf_87_top1.acquisition_clk ),
    .RESET_B(net1603),
    .D(_02229_),
    .Q_N(_07760_),
    .Q(\top1.memory2.mem2[0][1] ));
 sg13g2_dfrbp_1 _22133_ (.CLK(\clknet_leaf_91_top1.acquisition_clk ),
    .RESET_B(net1602),
    .D(_02230_),
    .Q_N(_07759_),
    .Q(\top1.memory2.mem2[0][2] ));
 sg13g2_dfrbp_1 _22134_ (.CLK(\clknet_leaf_234_top1.acquisition_clk ),
    .RESET_B(net1601),
    .D(_02231_),
    .Q_N(_07758_),
    .Q(\top1.memory2.mem2[100][0] ));
 sg13g2_dfrbp_1 _22135_ (.CLK(\clknet_leaf_233_top1.acquisition_clk ),
    .RESET_B(net1600),
    .D(_02232_),
    .Q_N(_07757_),
    .Q(\top1.memory2.mem2[100][1] ));
 sg13g2_dfrbp_1 _22136_ (.CLK(\clknet_leaf_235_top1.acquisition_clk ),
    .RESET_B(net1599),
    .D(_02233_),
    .Q_N(_07756_),
    .Q(\top1.memory2.mem2[100][2] ));
 sg13g2_dfrbp_1 _22137_ (.CLK(\clknet_leaf_234_top1.acquisition_clk ),
    .RESET_B(net1598),
    .D(_02234_),
    .Q_N(_07755_),
    .Q(\top1.memory2.mem2[101][0] ));
 sg13g2_dfrbp_1 _22138_ (.CLK(\clknet_leaf_233_top1.acquisition_clk ),
    .RESET_B(net1597),
    .D(_02235_),
    .Q_N(_07754_),
    .Q(\top1.memory2.mem2[101][1] ));
 sg13g2_dfrbp_1 _22139_ (.CLK(\clknet_leaf_235_top1.acquisition_clk ),
    .RESET_B(net1596),
    .D(_02236_),
    .Q_N(_07753_),
    .Q(\top1.memory2.mem2[101][2] ));
 sg13g2_dfrbp_1 _22140_ (.CLK(\clknet_leaf_234_top1.acquisition_clk ),
    .RESET_B(net1595),
    .D(_02237_),
    .Q_N(_07752_),
    .Q(\top1.memory2.mem2[102][0] ));
 sg13g2_dfrbp_1 _22141_ (.CLK(\clknet_leaf_233_top1.acquisition_clk ),
    .RESET_B(net1594),
    .D(_02238_),
    .Q_N(_07751_),
    .Q(\top1.memory2.mem2[102][1] ));
 sg13g2_dfrbp_1 _22142_ (.CLK(\clknet_leaf_235_top1.acquisition_clk ),
    .RESET_B(net1593),
    .D(_02239_),
    .Q_N(_07750_),
    .Q(\top1.memory2.mem2[102][2] ));
 sg13g2_dfrbp_1 _22143_ (.CLK(\clknet_leaf_234_top1.acquisition_clk ),
    .RESET_B(net1592),
    .D(_02240_),
    .Q_N(_07749_),
    .Q(\top1.memory2.mem2[103][0] ));
 sg13g2_dfrbp_1 _22144_ (.CLK(\clknet_leaf_231_top1.acquisition_clk ),
    .RESET_B(net1591),
    .D(_02241_),
    .Q_N(_07748_),
    .Q(\top1.memory2.mem2[103][1] ));
 sg13g2_dfrbp_1 _22145_ (.CLK(\clknet_leaf_235_top1.acquisition_clk ),
    .RESET_B(net1590),
    .D(_02242_),
    .Q_N(_07747_),
    .Q(\top1.memory2.mem2[103][2] ));
 sg13g2_dfrbp_1 _22146_ (.CLK(\clknet_leaf_230_top1.acquisition_clk ),
    .RESET_B(net1589),
    .D(_02243_),
    .Q_N(_07746_),
    .Q(\top1.memory2.mem2[104][0] ));
 sg13g2_dfrbp_1 _22147_ (.CLK(\clknet_leaf_192_top1.acquisition_clk ),
    .RESET_B(net1588),
    .D(_02244_),
    .Q_N(_07745_),
    .Q(\top1.memory2.mem2[104][1] ));
 sg13g2_dfrbp_1 _22148_ (.CLK(\clknet_leaf_252_top1.acquisition_clk ),
    .RESET_B(net1587),
    .D(_02245_),
    .Q_N(_07744_),
    .Q(\top1.memory2.mem2[104][2] ));
 sg13g2_dfrbp_1 _22149_ (.CLK(\clknet_leaf_230_top1.acquisition_clk ),
    .RESET_B(net1586),
    .D(_02246_),
    .Q_N(_07743_),
    .Q(\top1.memory2.mem2[105][0] ));
 sg13g2_dfrbp_1 _22150_ (.CLK(\clknet_leaf_193_top1.acquisition_clk ),
    .RESET_B(net1585),
    .D(_02247_),
    .Q_N(_07742_),
    .Q(\top1.memory2.mem2[105][1] ));
 sg13g2_dfrbp_1 _22151_ (.CLK(\clknet_leaf_230_top1.acquisition_clk ),
    .RESET_B(net1584),
    .D(_02248_),
    .Q_N(_07741_),
    .Q(\top1.memory2.mem2[105][2] ));
 sg13g2_dfrbp_1 _22152_ (.CLK(\clknet_leaf_231_top1.acquisition_clk ),
    .RESET_B(net1583),
    .D(_02249_),
    .Q_N(_07740_),
    .Q(\top1.memory2.mem2[106][0] ));
 sg13g2_dfrbp_1 _22153_ (.CLK(\clknet_leaf_194_top1.acquisition_clk ),
    .RESET_B(net1582),
    .D(_02250_),
    .Q_N(_07739_),
    .Q(\top1.memory2.mem2[106][1] ));
 sg13g2_dfrbp_1 _22154_ (.CLK(\clknet_leaf_230_top1.acquisition_clk ),
    .RESET_B(net1581),
    .D(_02251_),
    .Q_N(_07738_),
    .Q(\top1.memory2.mem2[106][2] ));
 sg13g2_dfrbp_1 _22155_ (.CLK(\clknet_leaf_231_top1.acquisition_clk ),
    .RESET_B(net1580),
    .D(_02252_),
    .Q_N(_07737_),
    .Q(\top1.memory2.mem2[107][0] ));
 sg13g2_dfrbp_1 _22156_ (.CLK(\clknet_leaf_194_top1.acquisition_clk ),
    .RESET_B(net1579),
    .D(_02253_),
    .Q_N(_07736_),
    .Q(\top1.memory2.mem2[107][1] ));
 sg13g2_dfrbp_1 _22157_ (.CLK(\clknet_leaf_230_top1.acquisition_clk ),
    .RESET_B(net1578),
    .D(_02254_),
    .Q_N(_07735_),
    .Q(\top1.memory2.mem2[107][2] ));
 sg13g2_dfrbp_1 _22158_ (.CLK(\clknet_leaf_225_top1.acquisition_clk ),
    .RESET_B(net1577),
    .D(_02255_),
    .Q_N(_07734_),
    .Q(\top1.memory2.mem2[108][0] ));
 sg13g2_dfrbp_1 _22159_ (.CLK(\clknet_leaf_226_top1.acquisition_clk ),
    .RESET_B(net1576),
    .D(_02256_),
    .Q_N(_07733_),
    .Q(\top1.memory2.mem2[108][1] ));
 sg13g2_dfrbp_1 _22160_ (.CLK(\clknet_leaf_235_top1.acquisition_clk ),
    .RESET_B(net1575),
    .D(_02257_),
    .Q_N(_07732_),
    .Q(\top1.memory2.mem2[108][2] ));
 sg13g2_dfrbp_1 _22161_ (.CLK(\clknet_leaf_89_top1.acquisition_clk ),
    .RESET_B(net1574),
    .D(_02258_),
    .Q_N(_07731_),
    .Q(\top1.memory2.mem2[10][0] ));
 sg13g2_dfrbp_1 _22162_ (.CLK(\clknet_leaf_85_top1.acquisition_clk ),
    .RESET_B(net1573),
    .D(_02259_),
    .Q_N(_07730_),
    .Q(\top1.memory2.mem2[10][1] ));
 sg13g2_dfrbp_1 _22163_ (.CLK(\clknet_leaf_94_top1.acquisition_clk ),
    .RESET_B(net1572),
    .D(_02260_),
    .Q_N(_07729_),
    .Q(\top1.memory2.mem2[10][2] ));
 sg13g2_dfrbp_1 _22164_ (.CLK(\clknet_leaf_225_top1.acquisition_clk ),
    .RESET_B(net1571),
    .D(_02261_),
    .Q_N(_07728_),
    .Q(\top1.memory2.mem2[110][0] ));
 sg13g2_dfrbp_1 _22165_ (.CLK(\clknet_leaf_226_top1.acquisition_clk ),
    .RESET_B(net1570),
    .D(_02262_),
    .Q_N(_07727_),
    .Q(\top1.memory2.mem2[110][1] ));
 sg13g2_dfrbp_1 _22166_ (.CLK(\clknet_leaf_234_top1.acquisition_clk ),
    .RESET_B(net1569),
    .D(_02263_),
    .Q_N(_07726_),
    .Q(\top1.memory2.mem2[110][2] ));
 sg13g2_dfrbp_1 _22167_ (.CLK(\clknet_leaf_224_top1.acquisition_clk ),
    .RESET_B(net1568),
    .D(_02264_),
    .Q_N(_07725_),
    .Q(\top1.memory2.mem2[111][0] ));
 sg13g2_dfrbp_1 _22168_ (.CLK(\clknet_leaf_226_top1.acquisition_clk ),
    .RESET_B(net1567),
    .D(_02265_),
    .Q_N(_07724_),
    .Q(\top1.memory2.mem2[111][1] ));
 sg13g2_dfrbp_1 _22169_ (.CLK(\clknet_leaf_225_top1.acquisition_clk ),
    .RESET_B(net1566),
    .D(_02266_),
    .Q_N(_07723_),
    .Q(\top1.memory2.mem2[111][2] ));
 sg13g2_dfrbp_1 _22170_ (.CLK(\clknet_leaf_213_top1.acquisition_clk ),
    .RESET_B(net1565),
    .D(_02267_),
    .Q_N(_07722_),
    .Q(\top1.memory2.mem2[112][0] ));
 sg13g2_dfrbp_1 _22171_ (.CLK(\clknet_leaf_196_top1.acquisition_clk ),
    .RESET_B(net1564),
    .D(_02268_),
    .Q_N(_07721_),
    .Q(\top1.memory2.mem2[112][1] ));
 sg13g2_dfrbp_1 _22172_ (.CLK(\clknet_leaf_209_top1.acquisition_clk ),
    .RESET_B(net1563),
    .D(_02269_),
    .Q_N(_07720_),
    .Q(\top1.memory2.mem2[112][2] ));
 sg13g2_dfrbp_1 _22173_ (.CLK(\clknet_leaf_215_top1.acquisition_clk ),
    .RESET_B(net1562),
    .D(_02270_),
    .Q_N(_07719_),
    .Q(\top1.memory2.mem2[113][0] ));
 sg13g2_dfrbp_1 _22174_ (.CLK(\clknet_leaf_200_top1.acquisition_clk ),
    .RESET_B(net1561),
    .D(_02271_),
    .Q_N(_07718_),
    .Q(\top1.memory2.mem2[113][1] ));
 sg13g2_dfrbp_1 _22175_ (.CLK(\clknet_leaf_209_top1.acquisition_clk ),
    .RESET_B(net1560),
    .D(_02272_),
    .Q_N(_07717_),
    .Q(\top1.memory2.mem2[113][2] ));
 sg13g2_dfrbp_1 _22176_ (.CLK(\clknet_leaf_212_top1.acquisition_clk ),
    .RESET_B(net1559),
    .D(_02273_),
    .Q_N(_07716_),
    .Q(\top1.memory2.mem2[114][0] ));
 sg13g2_dfrbp_1 _22177_ (.CLK(\clknet_leaf_196_top1.acquisition_clk ),
    .RESET_B(net1558),
    .D(_02274_),
    .Q_N(_07715_),
    .Q(\top1.memory2.mem2[114][1] ));
 sg13g2_dfrbp_1 _22178_ (.CLK(\clknet_leaf_209_top1.acquisition_clk ),
    .RESET_B(net1557),
    .D(_02275_),
    .Q_N(_07714_),
    .Q(\top1.memory2.mem2[114][2] ));
 sg13g2_dfrbp_1 _22179_ (.CLK(\clknet_leaf_215_top1.acquisition_clk ),
    .RESET_B(net1556),
    .D(_02276_),
    .Q_N(_07713_),
    .Q(\top1.memory2.mem2[115][0] ));
 sg13g2_dfrbp_1 _22180_ (.CLK(\clknet_leaf_200_top1.acquisition_clk ),
    .RESET_B(net1555),
    .D(_02277_),
    .Q_N(_07712_),
    .Q(\top1.memory2.mem2[115][1] ));
 sg13g2_dfrbp_1 _22181_ (.CLK(\clknet_leaf_209_top1.acquisition_clk ),
    .RESET_B(net1554),
    .D(_02278_),
    .Q_N(_07711_),
    .Q(\top1.memory2.mem2[115][2] ));
 sg13g2_dfrbp_1 _22182_ (.CLK(\clknet_leaf_223_top1.acquisition_clk ),
    .RESET_B(net1553),
    .D(_02279_),
    .Q_N(_07710_),
    .Q(\top1.memory2.mem2[116][0] ));
 sg13g2_dfrbp_1 _22183_ (.CLK(\clknet_leaf_228_top1.acquisition_clk ),
    .RESET_B(net1552),
    .D(_02280_),
    .Q_N(_07709_),
    .Q(\top1.memory2.mem2[116][1] ));
 sg13g2_dfrbp_1 _22184_ (.CLK(\clknet_leaf_223_top1.acquisition_clk ),
    .RESET_B(net1551),
    .D(_02281_),
    .Q_N(_07708_),
    .Q(\top1.memory2.mem2[116][2] ));
 sg13g2_dfrbp_1 _22185_ (.CLK(\clknet_leaf_222_top1.acquisition_clk ),
    .RESET_B(net1550),
    .D(_02282_),
    .Q_N(_07707_),
    .Q(\top1.memory2.mem2[117][0] ));
 sg13g2_dfrbp_1 _22186_ (.CLK(\clknet_leaf_213_top1.acquisition_clk ),
    .RESET_B(net1549),
    .D(_02283_),
    .Q_N(_07706_),
    .Q(\top1.memory2.mem2[117][1] ));
 sg13g2_dfrbp_1 _22187_ (.CLK(\clknet_leaf_222_top1.acquisition_clk ),
    .RESET_B(net1548),
    .D(_02284_),
    .Q_N(_07705_),
    .Q(\top1.memory2.mem2[117][2] ));
 sg13g2_dfrbp_1 _22188_ (.CLK(\clknet_leaf_223_top1.acquisition_clk ),
    .RESET_B(net1547),
    .D(_02285_),
    .Q_N(_07704_),
    .Q(\top1.memory2.mem2[118][0] ));
 sg13g2_dfrbp_1 _22189_ (.CLK(\clknet_leaf_228_top1.acquisition_clk ),
    .RESET_B(net1546),
    .D(_02286_),
    .Q_N(_07703_),
    .Q(\top1.memory2.mem2[118][1] ));
 sg13g2_dfrbp_1 _22190_ (.CLK(\clknet_leaf_222_top1.acquisition_clk ),
    .RESET_B(net1545),
    .D(_02287_),
    .Q_N(_07702_),
    .Q(\top1.memory2.mem2[118][2] ));
 sg13g2_dfrbp_1 _22191_ (.CLK(\clknet_leaf_90_top1.acquisition_clk ),
    .RESET_B(net1544),
    .D(_02288_),
    .Q_N(_07701_),
    .Q(\top1.memory2.mem2[11][0] ));
 sg13g2_dfrbp_1 _22192_ (.CLK(\clknet_leaf_86_top1.acquisition_clk ),
    .RESET_B(net1543),
    .D(_02289_),
    .Q_N(_07700_),
    .Q(\top1.memory2.mem2[11][1] ));
 sg13g2_dfrbp_1 _22193_ (.CLK(\clknet_leaf_90_top1.acquisition_clk ),
    .RESET_B(net1542),
    .D(_02290_),
    .Q_N(_07699_),
    .Q(\top1.memory2.mem2[11][2] ));
 sg13g2_dfrbp_1 _22194_ (.CLK(\clknet_leaf_212_top1.acquisition_clk ),
    .RESET_B(net1541),
    .D(_02291_),
    .Q_N(_07698_),
    .Q(\top1.memory2.mem2[120][0] ));
 sg13g2_dfrbp_1 _22195_ (.CLK(\clknet_leaf_210_top1.acquisition_clk ),
    .RESET_B(net1540),
    .D(_02292_),
    .Q_N(_07697_),
    .Q(\top1.memory2.mem2[120][1] ));
 sg13g2_dfrbp_1 _22196_ (.CLK(\clknet_leaf_210_top1.acquisition_clk ),
    .RESET_B(net1539),
    .D(_02293_),
    .Q_N(_07696_),
    .Q(\top1.memory2.mem2[120][2] ));
 sg13g2_dfrbp_1 _22197_ (.CLK(\clknet_leaf_212_top1.acquisition_clk ),
    .RESET_B(net1538),
    .D(_02294_),
    .Q_N(_07695_),
    .Q(\top1.memory2.mem2[121][0] ));
 sg13g2_dfrbp_1 _22198_ (.CLK(\clknet_leaf_210_top1.acquisition_clk ),
    .RESET_B(net1537),
    .D(_02295_),
    .Q_N(_07694_),
    .Q(\top1.memory2.mem2[121][1] ));
 sg13g2_dfrbp_1 _22199_ (.CLK(\clknet_leaf_209_top1.acquisition_clk ),
    .RESET_B(net1536),
    .D(_02296_),
    .Q_N(_07693_),
    .Q(\top1.memory2.mem2[121][2] ));
 sg13g2_dfrbp_1 _22200_ (.CLK(\clknet_leaf_212_top1.acquisition_clk ),
    .RESET_B(net1535),
    .D(_02297_),
    .Q_N(_07692_),
    .Q(\top1.memory2.mem2[122][0] ));
 sg13g2_dfrbp_1 _22201_ (.CLK(\clknet_leaf_212_top1.acquisition_clk ),
    .RESET_B(net1534),
    .D(_02298_),
    .Q_N(_07691_),
    .Q(\top1.memory2.mem2[122][1] ));
 sg13g2_dfrbp_1 _22202_ (.CLK(\clknet_leaf_210_top1.acquisition_clk ),
    .RESET_B(net1533),
    .D(_02299_),
    .Q_N(_07690_),
    .Q(\top1.memory2.mem2[122][2] ));
 sg13g2_dfrbp_1 _22203_ (.CLK(\clknet_leaf_212_top1.acquisition_clk ),
    .RESET_B(net1532),
    .D(_02300_),
    .Q_N(_07689_),
    .Q(\top1.memory2.mem2[123][0] ));
 sg13g2_dfrbp_1 _22204_ (.CLK(\clknet_leaf_194_top1.acquisition_clk ),
    .RESET_B(net1531),
    .D(_02301_),
    .Q_N(_07688_),
    .Q(\top1.memory2.mem2[123][1] ));
 sg13g2_dfrbp_1 _22205_ (.CLK(\clknet_leaf_210_top1.acquisition_clk ),
    .RESET_B(net1530),
    .D(_02302_),
    .Q_N(_07687_),
    .Q(\top1.memory2.mem2[123][2] ));
 sg13g2_dfrbp_1 _22206_ (.CLK(\clknet_leaf_228_top1.acquisition_clk ),
    .RESET_B(net1529),
    .D(_02303_),
    .Q_N(_07686_),
    .Q(\top1.memory2.mem2[124][0] ));
 sg13g2_dfrbp_1 _22207_ (.CLK(\clknet_leaf_227_top1.acquisition_clk ),
    .RESET_B(net1528),
    .D(_02304_),
    .Q_N(_07685_),
    .Q(\top1.memory2.mem2[124][1] ));
 sg13g2_dfrbp_1 _22208_ (.CLK(\clknet_leaf_224_top1.acquisition_clk ),
    .RESET_B(net1527),
    .D(_02305_),
    .Q_N(_07684_),
    .Q(\top1.memory2.mem2[124][2] ));
 sg13g2_dfrbp_1 _22209_ (.CLK(\clknet_leaf_228_top1.acquisition_clk ),
    .RESET_B(net1526),
    .D(_02306_),
    .Q_N(_07683_),
    .Q(\top1.memory2.mem2[125][0] ));
 sg13g2_dfrbp_1 _22210_ (.CLK(\clknet_leaf_227_top1.acquisition_clk ),
    .RESET_B(net1525),
    .D(_02307_),
    .Q_N(_07682_),
    .Q(\top1.memory2.mem2[125][1] ));
 sg13g2_dfrbp_1 _22211_ (.CLK(\clknet_leaf_224_top1.acquisition_clk ),
    .RESET_B(net1524),
    .D(_02308_),
    .Q_N(_07681_),
    .Q(\top1.memory2.mem2[125][2] ));
 sg13g2_dfrbp_1 _22212_ (.CLK(\clknet_leaf_213_top1.acquisition_clk ),
    .RESET_B(net1523),
    .D(_02309_),
    .Q_N(_07680_),
    .Q(\top1.memory2.mem2[126][0] ));
 sg13g2_dfrbp_1 _22213_ (.CLK(\clknet_leaf_227_top1.acquisition_clk ),
    .RESET_B(net1522),
    .D(_02310_),
    .Q_N(_07679_),
    .Q(\top1.memory2.mem2[126][1] ));
 sg13g2_dfrbp_1 _22214_ (.CLK(\clknet_leaf_224_top1.acquisition_clk ),
    .RESET_B(net1521),
    .D(_02311_),
    .Q_N(_07678_),
    .Q(\top1.memory2.mem2[126][2] ));
 sg13g2_dfrbp_1 _22215_ (.CLK(\clknet_leaf_213_top1.acquisition_clk ),
    .RESET_B(net1520),
    .D(_02312_),
    .Q_N(_07677_),
    .Q(\top1.memory2.mem2[127][0] ));
 sg13g2_dfrbp_1 _22216_ (.CLK(\clknet_leaf_227_top1.acquisition_clk ),
    .RESET_B(net1519),
    .D(_02313_),
    .Q_N(_07676_),
    .Q(\top1.memory2.mem2[127][1] ));
 sg13g2_dfrbp_1 _22217_ (.CLK(\clknet_leaf_224_top1.acquisition_clk ),
    .RESET_B(net1518),
    .D(_02314_),
    .Q_N(_07675_),
    .Q(\top1.memory2.mem2[127][2] ));
 sg13g2_dfrbp_1 _22218_ (.CLK(\clknet_leaf_66_top1.acquisition_clk ),
    .RESET_B(net1517),
    .D(_02315_),
    .Q_N(_07674_),
    .Q(\top1.memory2.mem2[128][0] ));
 sg13g2_dfrbp_1 _22219_ (.CLK(\clknet_leaf_65_top1.acquisition_clk ),
    .RESET_B(net1516),
    .D(_02316_),
    .Q_N(_07673_),
    .Q(\top1.memory2.mem2[128][1] ));
 sg13g2_dfrbp_1 _22220_ (.CLK(\clknet_leaf_66_top1.acquisition_clk ),
    .RESET_B(net1515),
    .D(_02317_),
    .Q_N(_07672_),
    .Q(\top1.memory2.mem2[128][2] ));
 sg13g2_dfrbp_1 _22221_ (.CLK(\clknet_leaf_79_top1.acquisition_clk ),
    .RESET_B(net1514),
    .D(_02318_),
    .Q_N(_07671_),
    .Q(\top1.memory2.mem2[12][0] ));
 sg13g2_dfrbp_1 _22222_ (.CLK(\clknet_leaf_79_top1.acquisition_clk ),
    .RESET_B(net1513),
    .D(_02319_),
    .Q_N(_07670_),
    .Q(\top1.memory2.mem2[12][1] ));
 sg13g2_dfrbp_1 _22223_ (.CLK(\clknet_leaf_95_top1.acquisition_clk ),
    .RESET_B(net1512),
    .D(_02320_),
    .Q_N(_07669_),
    .Q(\top1.memory2.mem2[12][2] ));
 sg13g2_dfrbp_1 _22224_ (.CLK(\clknet_leaf_66_top1.acquisition_clk ),
    .RESET_B(net1511),
    .D(_02321_),
    .Q_N(_07668_),
    .Q(\top1.memory2.mem2[130][0] ));
 sg13g2_dfrbp_1 _22225_ (.CLK(\clknet_leaf_68_top1.acquisition_clk ),
    .RESET_B(net1510),
    .D(_02322_),
    .Q_N(_07667_),
    .Q(\top1.memory2.mem2[130][1] ));
 sg13g2_dfrbp_1 _22226_ (.CLK(\clknet_leaf_66_top1.acquisition_clk ),
    .RESET_B(net1509),
    .D(_02323_),
    .Q_N(_07666_),
    .Q(\top1.memory2.mem2[130][2] ));
 sg13g2_dfrbp_1 _22227_ (.CLK(\clknet_leaf_67_top1.acquisition_clk ),
    .RESET_B(net1508),
    .D(_02324_),
    .Q_N(_07665_),
    .Q(\top1.memory2.mem2[131][0] ));
 sg13g2_dfrbp_1 _22228_ (.CLK(\clknet_leaf_68_top1.acquisition_clk ),
    .RESET_B(net1507),
    .D(_02325_),
    .Q_N(_07664_),
    .Q(\top1.memory2.mem2[131][1] ));
 sg13g2_dfrbp_1 _22229_ (.CLK(\clknet_leaf_66_top1.acquisition_clk ),
    .RESET_B(net1506),
    .D(_02326_),
    .Q_N(_07663_),
    .Q(\top1.memory2.mem2[131][2] ));
 sg13g2_dfrbp_1 _22230_ (.CLK(\clknet_leaf_61_top1.acquisition_clk ),
    .RESET_B(net1505),
    .D(_02327_),
    .Q_N(_07662_),
    .Q(\top1.memory2.mem2[132][0] ));
 sg13g2_dfrbp_1 _22231_ (.CLK(\clknet_leaf_61_top1.acquisition_clk ),
    .RESET_B(net1504),
    .D(_02328_),
    .Q_N(_07661_),
    .Q(\top1.memory2.mem2[132][1] ));
 sg13g2_dfrbp_1 _22232_ (.CLK(\clknet_leaf_68_top1.acquisition_clk ),
    .RESET_B(net1503),
    .D(_02329_),
    .Q_N(_07660_),
    .Q(\top1.memory2.mem2[132][2] ));
 sg13g2_dfrbp_1 _22233_ (.CLK(\clknet_leaf_59_top1.acquisition_clk ),
    .RESET_B(net1502),
    .D(_02330_),
    .Q_N(_07659_),
    .Q(\top1.memory2.mem2[133][0] ));
 sg13g2_dfrbp_1 _22234_ (.CLK(\clknet_leaf_61_top1.acquisition_clk ),
    .RESET_B(net1501),
    .D(_02331_),
    .Q_N(_07658_),
    .Q(\top1.memory2.mem2[133][1] ));
 sg13g2_dfrbp_1 _22235_ (.CLK(\clknet_leaf_60_top1.acquisition_clk ),
    .RESET_B(net1500),
    .D(_02332_),
    .Q_N(_07657_),
    .Q(\top1.memory2.mem2[133][2] ));
 sg13g2_dfrbp_1 _22236_ (.CLK(\clknet_leaf_60_top1.acquisition_clk ),
    .RESET_B(net1499),
    .D(_02333_),
    .Q_N(_07656_),
    .Q(\top1.memory2.mem2[134][0] ));
 sg13g2_dfrbp_1 _22237_ (.CLK(\clknet_leaf_62_top1.acquisition_clk ),
    .RESET_B(net1498),
    .D(_02334_),
    .Q_N(_07655_),
    .Q(\top1.memory2.mem2[134][1] ));
 sg13g2_dfrbp_1 _22238_ (.CLK(\clknet_leaf_74_top1.acquisition_clk ),
    .RESET_B(net1497),
    .D(_02335_),
    .Q_N(_07654_),
    .Q(\top1.memory2.mem2[134][2] ));
 sg13g2_dfrbp_1 _22239_ (.CLK(\clknet_leaf_60_top1.acquisition_clk ),
    .RESET_B(net1496),
    .D(_02336_),
    .Q_N(_07653_),
    .Q(\top1.memory2.mem2[135][0] ));
 sg13g2_dfrbp_1 _22240_ (.CLK(\clknet_leaf_61_top1.acquisition_clk ),
    .RESET_B(net1495),
    .D(_02337_),
    .Q_N(_07652_),
    .Q(\top1.memory2.mem2[135][1] ));
 sg13g2_dfrbp_1 _22241_ (.CLK(\clknet_leaf_60_top1.acquisition_clk ),
    .RESET_B(net1494),
    .D(_02338_),
    .Q_N(_07651_),
    .Q(\top1.memory2.mem2[135][2] ));
 sg13g2_dfrbp_1 _22242_ (.CLK(\clknet_leaf_67_top1.acquisition_clk ),
    .RESET_B(net1493),
    .D(_02339_),
    .Q_N(_07650_),
    .Q(\top1.memory2.mem2[136][0] ));
 sg13g2_dfrbp_1 _22243_ (.CLK(\clknet_leaf_64_top1.acquisition_clk ),
    .RESET_B(net1492),
    .D(_02340_),
    .Q_N(_07649_),
    .Q(\top1.memory2.mem2[136][1] ));
 sg13g2_dfrbp_1 _22244_ (.CLK(\clknet_leaf_69_top1.acquisition_clk ),
    .RESET_B(net1491),
    .D(_02341_),
    .Q_N(_07648_),
    .Q(\top1.memory2.mem2[136][2] ));
 sg13g2_dfrbp_1 _22245_ (.CLK(\clknet_leaf_67_top1.acquisition_clk ),
    .RESET_B(net1490),
    .D(_02342_),
    .Q_N(_07647_),
    .Q(\top1.memory2.mem2[137][0] ));
 sg13g2_dfrbp_1 _22246_ (.CLK(\clknet_leaf_68_top1.acquisition_clk ),
    .RESET_B(net1489),
    .D(_02343_),
    .Q_N(_07646_),
    .Q(\top1.memory2.mem2[137][1] ));
 sg13g2_dfrbp_1 _22247_ (.CLK(\clknet_leaf_69_top1.acquisition_clk ),
    .RESET_B(net1488),
    .D(_02344_),
    .Q_N(_07645_),
    .Q(\top1.memory2.mem2[137][2] ));
 sg13g2_dfrbp_1 _22248_ (.CLK(\clknet_leaf_67_top1.acquisition_clk ),
    .RESET_B(net1487),
    .D(_02345_),
    .Q_N(_07644_),
    .Q(\top1.memory2.mem2[138][0] ));
 sg13g2_dfrbp_1 _22249_ (.CLK(\clknet_leaf_64_top1.acquisition_clk ),
    .RESET_B(net1486),
    .D(_02346_),
    .Q_N(_07643_),
    .Q(\top1.memory2.mem2[138][1] ));
 sg13g2_dfrbp_1 _22250_ (.CLK(\clknet_leaf_69_top1.acquisition_clk ),
    .RESET_B(net1485),
    .D(_02347_),
    .Q_N(_07642_),
    .Q(\top1.memory2.mem2[138][2] ));
 sg13g2_dfrbp_1 _22251_ (.CLK(\clknet_leaf_79_top1.acquisition_clk ),
    .RESET_B(net1484),
    .D(_02348_),
    .Q_N(_07641_),
    .Q(\top1.memory2.mem2[13][0] ));
 sg13g2_dfrbp_1 _22252_ (.CLK(\clknet_leaf_79_top1.acquisition_clk ),
    .RESET_B(net1483),
    .D(_02349_),
    .Q_N(_07640_),
    .Q(\top1.memory2.mem2[13][1] ));
 sg13g2_dfrbp_1 _22253_ (.CLK(\clknet_leaf_94_top1.acquisition_clk ),
    .RESET_B(net1482),
    .D(_02350_),
    .Q_N(_07639_),
    .Q(\top1.memory2.mem2[13][2] ));
 sg13g2_dfrbp_1 _22254_ (.CLK(\clknet_leaf_63_top1.acquisition_clk ),
    .RESET_B(net1481),
    .D(_02351_),
    .Q_N(_07638_),
    .Q(\top1.memory2.mem2[140][0] ));
 sg13g2_dfrbp_1 _22255_ (.CLK(\clknet_leaf_64_top1.acquisition_clk ),
    .RESET_B(net1480),
    .D(_02352_),
    .Q_N(_07637_),
    .Q(\top1.memory2.mem2[140][1] ));
 sg13g2_dfrbp_1 _22256_ (.CLK(\clknet_leaf_55_top1.acquisition_clk ),
    .RESET_B(net1479),
    .D(_02353_),
    .Q_N(_07636_),
    .Q(\top1.memory2.mem2[140][2] ));
 sg13g2_dfrbp_1 _22257_ (.CLK(\clknet_leaf_63_top1.acquisition_clk ),
    .RESET_B(net1478),
    .D(_02354_),
    .Q_N(_07635_),
    .Q(\top1.memory2.mem2[141][0] ));
 sg13g2_dfrbp_1 _22258_ (.CLK(\clknet_leaf_63_top1.acquisition_clk ),
    .RESET_B(net1477),
    .D(_02355_),
    .Q_N(_07634_),
    .Q(\top1.memory2.mem2[141][1] ));
 sg13g2_dfrbp_1 _22259_ (.CLK(\clknet_leaf_54_top1.acquisition_clk ),
    .RESET_B(net1476),
    .D(_02356_),
    .Q_N(_07633_),
    .Q(\top1.memory2.mem2[141][2] ));
 sg13g2_dfrbp_1 _22260_ (.CLK(\clknet_leaf_62_top1.acquisition_clk ),
    .RESET_B(net1475),
    .D(_02357_),
    .Q_N(_07632_),
    .Q(\top1.memory2.mem2[142][0] ));
 sg13g2_dfrbp_1 _22261_ (.CLK(\clknet_leaf_63_top1.acquisition_clk ),
    .RESET_B(net1474),
    .D(_02358_),
    .Q_N(_07631_),
    .Q(\top1.memory2.mem2[142][1] ));
 sg13g2_dfrbp_1 _22262_ (.CLK(\clknet_leaf_54_top1.acquisition_clk ),
    .RESET_B(net1473),
    .D(_02359_),
    .Q_N(_07630_),
    .Q(\top1.memory2.mem2[142][2] ));
 sg13g2_dfrbp_1 _22263_ (.CLK(\clknet_leaf_63_top1.acquisition_clk ),
    .RESET_B(net1472),
    .D(_02360_),
    .Q_N(_07629_),
    .Q(\top1.memory2.mem2[143][0] ));
 sg13g2_dfrbp_1 _22264_ (.CLK(\clknet_leaf_64_top1.acquisition_clk ),
    .RESET_B(net1471),
    .D(_02361_),
    .Q_N(_07628_),
    .Q(\top1.memory2.mem2[143][1] ));
 sg13g2_dfrbp_1 _22265_ (.CLK(\clknet_leaf_54_top1.acquisition_clk ),
    .RESET_B(net1470),
    .D(_02362_),
    .Q_N(_07627_),
    .Q(\top1.memory2.mem2[143][2] ));
 sg13g2_dfrbp_1 _22266_ (.CLK(\clknet_leaf_75_top1.acquisition_clk ),
    .RESET_B(net1469),
    .D(_02363_),
    .Q_N(_07626_),
    .Q(\top1.memory2.mem2[144][0] ));
 sg13g2_dfrbp_1 _22267_ (.CLK(\clknet_leaf_80_top1.acquisition_clk ),
    .RESET_B(net1468),
    .D(_02364_),
    .Q_N(_07625_),
    .Q(\top1.memory2.mem2[144][1] ));
 sg13g2_dfrbp_1 _22268_ (.CLK(\clknet_leaf_76_top1.acquisition_clk ),
    .RESET_B(net1467),
    .D(_02365_),
    .Q_N(_07624_),
    .Q(\top1.memory2.mem2[144][2] ));
 sg13g2_dfrbp_1 _22269_ (.CLK(\clknet_leaf_75_top1.acquisition_clk ),
    .RESET_B(net1466),
    .D(_02366_),
    .Q_N(_07623_),
    .Q(\top1.memory2.mem2[145][0] ));
 sg13g2_dfrbp_1 _22270_ (.CLK(\clknet_leaf_80_top1.acquisition_clk ),
    .RESET_B(net1465),
    .D(_02367_),
    .Q_N(_07622_),
    .Q(\top1.memory2.mem2[145][1] ));
 sg13g2_dfrbp_1 _22271_ (.CLK(\clknet_leaf_78_top1.acquisition_clk ),
    .RESET_B(net1464),
    .D(_02368_),
    .Q_N(_07621_),
    .Q(\top1.memory2.mem2[145][2] ));
 sg13g2_dfrbp_1 _22272_ (.CLK(\clknet_leaf_76_top1.acquisition_clk ),
    .RESET_B(net1463),
    .D(_02369_),
    .Q_N(_07620_),
    .Q(\top1.memory2.mem2[146][0] ));
 sg13g2_dfrbp_1 _22273_ (.CLK(\clknet_leaf_78_top1.acquisition_clk ),
    .RESET_B(net1462),
    .D(_02370_),
    .Q_N(_07619_),
    .Q(\top1.memory2.mem2[146][1] ));
 sg13g2_dfrbp_1 _22274_ (.CLK(\clknet_leaf_76_top1.acquisition_clk ),
    .RESET_B(net1461),
    .D(_02371_),
    .Q_N(_07618_),
    .Q(\top1.memory2.mem2[146][2] ));
 sg13g2_dfrbp_1 _22275_ (.CLK(\clknet_leaf_76_top1.acquisition_clk ),
    .RESET_B(net1460),
    .D(_02372_),
    .Q_N(_07617_),
    .Q(\top1.memory2.mem2[147][0] ));
 sg13g2_dfrbp_1 _22276_ (.CLK(\clknet_leaf_78_top1.acquisition_clk ),
    .RESET_B(net1459),
    .D(_02373_),
    .Q_N(_07616_),
    .Q(\top1.memory2.mem2[147][1] ));
 sg13g2_dfrbp_1 _22277_ (.CLK(\clknet_leaf_76_top1.acquisition_clk ),
    .RESET_B(net1458),
    .D(_02374_),
    .Q_N(_07615_),
    .Q(\top1.memory2.mem2[147][2] ));
 sg13g2_dfrbp_1 _22278_ (.CLK(\clknet_leaf_77_top1.acquisition_clk ),
    .RESET_B(net1457),
    .D(_02375_),
    .Q_N(_07614_),
    .Q(\top1.memory2.mem2[148][0] ));
 sg13g2_dfrbp_1 _22279_ (.CLK(\clknet_leaf_41_top1.acquisition_clk ),
    .RESET_B(net1456),
    .D(_02376_),
    .Q_N(_07613_),
    .Q(\top1.memory2.mem2[148][1] ));
 sg13g2_dfrbp_1 _22280_ (.CLK(\clknet_leaf_97_top1.acquisition_clk ),
    .RESET_B(net1455),
    .D(_02377_),
    .Q_N(_07612_),
    .Q(\top1.memory2.mem2[148][2] ));
 sg13g2_dfrbp_1 _22281_ (.CLK(\clknet_leaf_84_top1.acquisition_clk ),
    .RESET_B(net1454),
    .D(_02378_),
    .Q_N(_07611_),
    .Q(\top1.memory2.mem2[14][0] ));
 sg13g2_dfrbp_1 _22282_ (.CLK(\clknet_leaf_84_top1.acquisition_clk ),
    .RESET_B(net1453),
    .D(_02379_),
    .Q_N(_07610_),
    .Q(\top1.memory2.mem2[14][1] ));
 sg13g2_dfrbp_1 _22283_ (.CLK(\clknet_leaf_84_top1.acquisition_clk ),
    .RESET_B(net1452),
    .D(_02380_),
    .Q_N(_07609_),
    .Q(\top1.memory2.mem2[14][2] ));
 sg13g2_dfrbp_1 _22284_ (.CLK(\clknet_leaf_97_top1.acquisition_clk ),
    .RESET_B(net1451),
    .D(_02381_),
    .Q_N(_07608_),
    .Q(\top1.memory2.mem2[150][0] ));
 sg13g2_dfrbp_1 _22285_ (.CLK(\clknet_leaf_41_top1.acquisition_clk ),
    .RESET_B(net1450),
    .D(_02382_),
    .Q_N(_07607_),
    .Q(\top1.memory2.mem2[150][1] ));
 sg13g2_dfrbp_1 _22286_ (.CLK(\clknet_leaf_43_top1.acquisition_clk ),
    .RESET_B(net1449),
    .D(_02383_),
    .Q_N(_07606_),
    .Q(\top1.memory2.mem2[150][2] ));
 sg13g2_dfrbp_1 _22287_ (.CLK(\clknet_leaf_77_top1.acquisition_clk ),
    .RESET_B(net1448),
    .D(_02384_),
    .Q_N(_07605_),
    .Q(\top1.memory2.mem2[151][0] ));
 sg13g2_dfrbp_1 _22288_ (.CLK(\clknet_leaf_42_top1.acquisition_clk ),
    .RESET_B(net1447),
    .D(_02385_),
    .Q_N(_07604_),
    .Q(\top1.memory2.mem2[151][1] ));
 sg13g2_dfrbp_1 _22289_ (.CLK(\clknet_leaf_42_top1.acquisition_clk ),
    .RESET_B(net1446),
    .D(_02386_),
    .Q_N(_07603_),
    .Q(\top1.memory2.mem2[151][2] ));
 sg13g2_dfrbp_1 _22290_ (.CLK(\clknet_leaf_78_top1.acquisition_clk ),
    .RESET_B(net1445),
    .D(_02387_),
    .Q_N(_07602_),
    .Q(\top1.memory2.mem2[152][0] ));
 sg13g2_dfrbp_1 _22291_ (.CLK(\clknet_leaf_82_top1.acquisition_clk ),
    .RESET_B(net1444),
    .D(_02388_),
    .Q_N(_07601_),
    .Q(\top1.memory2.mem2[152][1] ));
 sg13g2_dfrbp_1 _22292_ (.CLK(\clknet_leaf_80_top1.acquisition_clk ),
    .RESET_B(net1443),
    .D(_02389_),
    .Q_N(_07600_),
    .Q(\top1.memory2.mem2[152][2] ));
 sg13g2_dfrbp_1 _22293_ (.CLK(\clknet_leaf_78_top1.acquisition_clk ),
    .RESET_B(net1442),
    .D(_02390_),
    .Q_N(_07599_),
    .Q(\top1.memory2.mem2[153][0] ));
 sg13g2_dfrbp_1 _22294_ (.CLK(\clknet_leaf_82_top1.acquisition_clk ),
    .RESET_B(net1441),
    .D(_02391_),
    .Q_N(_07598_),
    .Q(\top1.memory2.mem2[153][1] ));
 sg13g2_dfrbp_1 _22295_ (.CLK(\clknet_leaf_80_top1.acquisition_clk ),
    .RESET_B(net1440),
    .D(_02392_),
    .Q_N(_07597_),
    .Q(\top1.memory2.mem2[153][2] ));
 sg13g2_dfrbp_1 _22296_ (.CLK(\clknet_leaf_79_top1.acquisition_clk ),
    .RESET_B(net1439),
    .D(_02393_),
    .Q_N(_07596_),
    .Q(\top1.memory2.mem2[154][0] ));
 sg13g2_dfrbp_1 _22297_ (.CLK(\clknet_leaf_81_top1.acquisition_clk ),
    .RESET_B(net1438),
    .D(_02394_),
    .Q_N(_07595_),
    .Q(\top1.memory2.mem2[154][1] ));
 sg13g2_dfrbp_1 _22298_ (.CLK(\clknet_leaf_84_top1.acquisition_clk ),
    .RESET_B(net1437),
    .D(_02395_),
    .Q_N(_07594_),
    .Q(\top1.memory2.mem2[154][2] ));
 sg13g2_dfrbp_1 _22299_ (.CLK(\clknet_leaf_79_top1.acquisition_clk ),
    .RESET_B(net1436),
    .D(_02396_),
    .Q_N(_07593_),
    .Q(\top1.memory2.mem2[155][0] ));
 sg13g2_dfrbp_1 _22300_ (.CLK(\clknet_leaf_81_top1.acquisition_clk ),
    .RESET_B(net1435),
    .D(_02397_),
    .Q_N(_07592_),
    .Q(\top1.memory2.mem2[155][1] ));
 sg13g2_dfrbp_1 _22301_ (.CLK(\clknet_leaf_80_top1.acquisition_clk ),
    .RESET_B(net1434),
    .D(_02398_),
    .Q_N(_07591_),
    .Q(\top1.memory2.mem2[155][2] ));
 sg13g2_dfrbp_1 _22302_ (.CLK(\clknet_leaf_71_top1.acquisition_clk ),
    .RESET_B(net1433),
    .D(_02399_),
    .Q_N(_07590_),
    .Q(\top1.memory2.mem2[156][0] ));
 sg13g2_dfrbp_1 _22303_ (.CLK(\clknet_leaf_81_top1.acquisition_clk ),
    .RESET_B(net1432),
    .D(_02400_),
    .Q_N(_07589_),
    .Q(\top1.memory2.mem2[156][1] ));
 sg13g2_dfrbp_1 _22304_ (.CLK(\clknet_leaf_72_top1.acquisition_clk ),
    .RESET_B(net1431),
    .D(_02401_),
    .Q_N(_07588_),
    .Q(\top1.memory2.mem2[156][2] ));
 sg13g2_dfrbp_1 _22305_ (.CLK(\clknet_leaf_71_top1.acquisition_clk ),
    .RESET_B(net1430),
    .D(_02402_),
    .Q_N(_07587_),
    .Q(\top1.memory2.mem2[157][0] ));
 sg13g2_dfrbp_1 _22306_ (.CLK(\clknet_leaf_81_top1.acquisition_clk ),
    .RESET_B(net1429),
    .D(_02403_),
    .Q_N(_07586_),
    .Q(\top1.memory2.mem2[157][1] ));
 sg13g2_dfrbp_1 _22307_ (.CLK(\clknet_leaf_72_top1.acquisition_clk ),
    .RESET_B(net1428),
    .D(_02404_),
    .Q_N(_07585_),
    .Q(\top1.memory2.mem2[157][2] ));
 sg13g2_dfrbp_1 _22308_ (.CLK(\clknet_leaf_71_top1.acquisition_clk ),
    .RESET_B(net1427),
    .D(_02405_),
    .Q_N(_07584_),
    .Q(\top1.memory2.mem2[158][0] ));
 sg13g2_dfrbp_1 _22309_ (.CLK(\clknet_leaf_80_top1.acquisition_clk ),
    .RESET_B(net1426),
    .D(_02406_),
    .Q_N(_07583_),
    .Q(\top1.memory2.mem2[158][1] ));
 sg13g2_dfrbp_1 _22310_ (.CLK(\clknet_leaf_72_top1.acquisition_clk ),
    .RESET_B(net1425),
    .D(_02407_),
    .Q_N(_07582_),
    .Q(\top1.memory2.mem2[158][2] ));
 sg13g2_dfrbp_1 _22311_ (.CLK(\clknet_leaf_84_top1.acquisition_clk ),
    .RESET_B(net1424),
    .D(_02408_),
    .Q_N(_07581_),
    .Q(\top1.memory2.mem2[15][0] ));
 sg13g2_dfrbp_1 _22312_ (.CLK(\clknet_leaf_79_top1.acquisition_clk ),
    .RESET_B(net1423),
    .D(_02409_),
    .Q_N(_07580_),
    .Q(\top1.memory2.mem2[15][1] ));
 sg13g2_dfrbp_1 _22313_ (.CLK(\clknet_leaf_84_top1.acquisition_clk ),
    .RESET_B(net1422),
    .D(_02410_),
    .Q_N(_07579_),
    .Q(\top1.memory2.mem2[15][2] ));
 sg13g2_dfrbp_1 _22314_ (.CLK(\clknet_leaf_104_top1.acquisition_clk ),
    .RESET_B(net1421),
    .D(_02411_),
    .Q_N(_07578_),
    .Q(\top1.memory2.mem2[160][0] ));
 sg13g2_dfrbp_1 _22315_ (.CLK(\clknet_leaf_103_top1.acquisition_clk ),
    .RESET_B(net1420),
    .D(_02412_),
    .Q_N(_07577_),
    .Q(\top1.memory2.mem2[160][1] ));
 sg13g2_dfrbp_1 _22316_ (.CLK(\clknet_leaf_105_top1.acquisition_clk ),
    .RESET_B(net1419),
    .D(_02413_),
    .Q_N(_07576_),
    .Q(\top1.memory2.mem2[160][2] ));
 sg13g2_dfrbp_1 _22317_ (.CLK(\clknet_leaf_104_top1.acquisition_clk ),
    .RESET_B(net1418),
    .D(_02414_),
    .Q_N(_07575_),
    .Q(\top1.memory2.mem2[161][0] ));
 sg13g2_dfrbp_1 _22318_ (.CLK(\clknet_leaf_103_top1.acquisition_clk ),
    .RESET_B(net1417),
    .D(_02415_),
    .Q_N(_07574_),
    .Q(\top1.memory2.mem2[161][1] ));
 sg13g2_dfrbp_1 _22319_ (.CLK(\clknet_leaf_37_top1.acquisition_clk ),
    .RESET_B(net1416),
    .D(_02416_),
    .Q_N(_07573_),
    .Q(\top1.memory2.mem2[161][2] ));
 sg13g2_dfrbp_1 _22320_ (.CLK(\clknet_leaf_104_top1.acquisition_clk ),
    .RESET_B(net1415),
    .D(_02417_),
    .Q_N(_07572_),
    .Q(\top1.memory2.mem2[162][0] ));
 sg13g2_dfrbp_1 _22321_ (.CLK(\clknet_leaf_104_top1.acquisition_clk ),
    .RESET_B(net1414),
    .D(_02418_),
    .Q_N(_07571_),
    .Q(\top1.memory2.mem2[162][1] ));
 sg13g2_dfrbp_1 _22322_ (.CLK(\clknet_leaf_37_top1.acquisition_clk ),
    .RESET_B(net1413),
    .D(_02419_),
    .Q_N(_07570_),
    .Q(\top1.memory2.mem2[162][2] ));
 sg13g2_dfrbp_1 _22323_ (.CLK(\clknet_leaf_102_top1.acquisition_clk ),
    .RESET_B(net1412),
    .D(_02420_),
    .Q_N(_07569_),
    .Q(\top1.memory2.mem2[163][0] ));
 sg13g2_dfrbp_1 _22324_ (.CLK(\clknet_leaf_105_top1.acquisition_clk ),
    .RESET_B(net1411),
    .D(_02421_),
    .Q_N(_07568_),
    .Q(\top1.memory2.mem2[163][1] ));
 sg13g2_dfrbp_1 _22325_ (.CLK(\clknet_leaf_105_top1.acquisition_clk ),
    .RESET_B(net1410),
    .D(_02422_),
    .Q_N(_07567_),
    .Q(\top1.memory2.mem2[163][2] ));
 sg13g2_dfrbp_1 _22326_ (.CLK(\clknet_leaf_103_top1.acquisition_clk ),
    .RESET_B(net1409),
    .D(_02423_),
    .Q_N(_07566_),
    .Q(\top1.memory2.mem2[164][0] ));
 sg13g2_dfrbp_1 _22327_ (.CLK(\clknet_leaf_101_top1.acquisition_clk ),
    .RESET_B(net1408),
    .D(_02424_),
    .Q_N(_07565_),
    .Q(\top1.memory2.mem2[164][1] ));
 sg13g2_dfrbp_1 _22328_ (.CLK(\clknet_leaf_92_top1.acquisition_clk ),
    .RESET_B(net1407),
    .D(_02425_),
    .Q_N(_07564_),
    .Q(\top1.memory2.mem2[164][2] ));
 sg13g2_dfrbp_1 _22329_ (.CLK(\clknet_leaf_103_top1.acquisition_clk ),
    .RESET_B(net1406),
    .D(_02426_),
    .Q_N(_07563_),
    .Q(\top1.memory2.mem2[165][0] ));
 sg13g2_dfrbp_1 _22330_ (.CLK(\clknet_leaf_102_top1.acquisition_clk ),
    .RESET_B(net1405),
    .D(_02427_),
    .Q_N(_07562_),
    .Q(\top1.memory2.mem2[165][1] ));
 sg13g2_dfrbp_1 _22331_ (.CLK(\clknet_leaf_92_top1.acquisition_clk ),
    .RESET_B(net1404),
    .D(_02428_),
    .Q_N(_07561_),
    .Q(\top1.memory2.mem2[165][2] ));
 sg13g2_dfrbp_1 _22332_ (.CLK(\clknet_leaf_103_top1.acquisition_clk ),
    .RESET_B(net1403),
    .D(_02429_),
    .Q_N(_07560_),
    .Q(\top1.memory2.mem2[166][0] ));
 sg13g2_dfrbp_1 _22333_ (.CLK(\clknet_leaf_100_top1.acquisition_clk ),
    .RESET_B(net1402),
    .D(_02430_),
    .Q_N(_07559_),
    .Q(\top1.memory2.mem2[166][1] ));
 sg13g2_dfrbp_1 _22334_ (.CLK(\clknet_leaf_92_top1.acquisition_clk ),
    .RESET_B(net1401),
    .D(_02431_),
    .Q_N(_07558_),
    .Q(\top1.memory2.mem2[166][2] ));
 sg13g2_dfrbp_1 _22335_ (.CLK(\clknet_leaf_102_top1.acquisition_clk ),
    .RESET_B(net1400),
    .D(_02432_),
    .Q_N(_07557_),
    .Q(\top1.memory2.mem2[167][0] ));
 sg13g2_dfrbp_1 _22336_ (.CLK(\clknet_leaf_102_top1.acquisition_clk ),
    .RESET_B(net1399),
    .D(_02433_),
    .Q_N(_07556_),
    .Q(\top1.memory2.mem2[167][1] ));
 sg13g2_dfrbp_1 _22337_ (.CLK(\clknet_leaf_92_top1.acquisition_clk ),
    .RESET_B(net1398),
    .D(_02434_),
    .Q_N(_07555_),
    .Q(\top1.memory2.mem2[167][2] ));
 sg13g2_dfrbp_1 _22338_ (.CLK(\clknet_leaf_107_top1.acquisition_clk ),
    .RESET_B(net1397),
    .D(_02435_),
    .Q_N(_07554_),
    .Q(\top1.memory2.mem2[168][0] ));
 sg13g2_dfrbp_1 _22339_ (.CLK(\clknet_leaf_110_top1.acquisition_clk ),
    .RESET_B(net1396),
    .D(_02436_),
    .Q_N(_07553_),
    .Q(\top1.memory2.mem2[168][1] ));
 sg13g2_dfrbp_1 _22340_ (.CLK(\clknet_leaf_105_top1.acquisition_clk ),
    .RESET_B(net1395),
    .D(_02437_),
    .Q_N(_07552_),
    .Q(\top1.memory2.mem2[168][2] ));
 sg13g2_dfrbp_1 _22341_ (.CLK(\clknet_leaf_112_top1.acquisition_clk ),
    .RESET_B(net1394),
    .D(_02438_),
    .Q_N(_07551_),
    .Q(\top1.memory2.mem2[16][0] ));
 sg13g2_dfrbp_1 _22342_ (.CLK(\clknet_leaf_119_top1.acquisition_clk ),
    .RESET_B(net1393),
    .D(_02439_),
    .Q_N(_07550_),
    .Q(\top1.memory2.mem2[16][1] ));
 sg13g2_dfrbp_1 _22343_ (.CLK(\clknet_leaf_112_top1.acquisition_clk ),
    .RESET_B(net1392),
    .D(_02440_),
    .Q_N(_07549_),
    .Q(\top1.memory2.mem2[16][2] ));
 sg13g2_dfrbp_1 _22344_ (.CLK(\clknet_leaf_106_top1.acquisition_clk ),
    .RESET_B(net1391),
    .D(_02441_),
    .Q_N(_07548_),
    .Q(\top1.memory2.mem2[170][0] ));
 sg13g2_dfrbp_1 _22345_ (.CLK(\clknet_leaf_111_top1.acquisition_clk ),
    .RESET_B(net1390),
    .D(_02442_),
    .Q_N(_07547_),
    .Q(\top1.memory2.mem2[170][1] ));
 sg13g2_dfrbp_1 _22346_ (.CLK(\clknet_leaf_107_top1.acquisition_clk ),
    .RESET_B(net1389),
    .D(_02443_),
    .Q_N(_07546_),
    .Q(\top1.memory2.mem2[170][2] ));
 sg13g2_dfrbp_1 _22347_ (.CLK(\clknet_leaf_106_top1.acquisition_clk ),
    .RESET_B(net1388),
    .D(_02444_),
    .Q_N(_07545_),
    .Q(\top1.memory2.mem2[171][0] ));
 sg13g2_dfrbp_1 _22348_ (.CLK(\clknet_leaf_110_top1.acquisition_clk ),
    .RESET_B(net1387),
    .D(_02445_),
    .Q_N(_07544_),
    .Q(\top1.memory2.mem2[171][1] ));
 sg13g2_dfrbp_1 _22349_ (.CLK(\clknet_leaf_107_top1.acquisition_clk ),
    .RESET_B(net1386),
    .D(_02446_),
    .Q_N(_07543_),
    .Q(\top1.memory2.mem2[171][2] ));
 sg13g2_dfrbp_1 _22350_ (.CLK(\clknet_leaf_260_top1.acquisition_clk ),
    .RESET_B(net1385),
    .D(_02447_),
    .Q_N(_07542_),
    .Q(\top1.memory2.mem2[172][0] ));
 sg13g2_dfrbp_1 _22351_ (.CLK(\clknet_leaf_264_top1.acquisition_clk ),
    .RESET_B(net1384),
    .D(_02448_),
    .Q_N(_07541_),
    .Q(\top1.memory2.mem2[172][1] ));
 sg13g2_dfrbp_1 _22352_ (.CLK(\clknet_leaf_261_top1.acquisition_clk ),
    .RESET_B(net1383),
    .D(_02449_),
    .Q_N(_07540_),
    .Q(\top1.memory2.mem2[172][2] ));
 sg13g2_dfrbp_1 _22353_ (.CLK(\clknet_leaf_259_top1.acquisition_clk ),
    .RESET_B(net1382),
    .D(_02450_),
    .Q_N(_07539_),
    .Q(\top1.memory2.mem2[173][0] ));
 sg13g2_dfrbp_1 _22354_ (.CLK(\clknet_leaf_264_top1.acquisition_clk ),
    .RESET_B(net1381),
    .D(_02451_),
    .Q_N(_07538_),
    .Q(\top1.memory2.mem2[173][1] ));
 sg13g2_dfrbp_1 _22355_ (.CLK(\clknet_leaf_260_top1.acquisition_clk ),
    .RESET_B(net1380),
    .D(_02452_),
    .Q_N(_07537_),
    .Q(\top1.memory2.mem2[173][2] ));
 sg13g2_dfrbp_1 _22356_ (.CLK(\clknet_leaf_260_top1.acquisition_clk ),
    .RESET_B(net1379),
    .D(_02453_),
    .Q_N(_07536_),
    .Q(\top1.memory2.mem2[174][0] ));
 sg13g2_dfrbp_1 _22357_ (.CLK(\clknet_leaf_263_top1.acquisition_clk ),
    .RESET_B(net1378),
    .D(_02454_),
    .Q_N(_07535_),
    .Q(\top1.memory2.mem2[174][1] ));
 sg13g2_dfrbp_1 _22358_ (.CLK(\clknet_leaf_261_top1.acquisition_clk ),
    .RESET_B(net1377),
    .D(_02455_),
    .Q_N(_07534_),
    .Q(\top1.memory2.mem2[174][2] ));
 sg13g2_dfrbp_1 _22359_ (.CLK(\clknet_leaf_261_top1.acquisition_clk ),
    .RESET_B(net1376),
    .D(_02456_),
    .Q_N(_07533_),
    .Q(\top1.memory2.mem2[175][0] ));
 sg13g2_dfrbp_1 _22360_ (.CLK(\clknet_leaf_263_top1.acquisition_clk ),
    .RESET_B(net1375),
    .D(_02457_),
    .Q_N(_07532_),
    .Q(\top1.memory2.mem2[175][1] ));
 sg13g2_dfrbp_1 _22361_ (.CLK(\clknet_leaf_261_top1.acquisition_clk ),
    .RESET_B(net1374),
    .D(_02458_),
    .Q_N(_07531_),
    .Q(\top1.memory2.mem2[175][2] ));
 sg13g2_dfrbp_1 _22362_ (.CLK(\clknet_leaf_134_top1.acquisition_clk ),
    .RESET_B(net1373),
    .D(_02459_),
    .Q_N(_07530_),
    .Q(\top1.memory2.mem2[176][0] ));
 sg13g2_dfrbp_1 _22363_ (.CLK(\clknet_leaf_130_top1.acquisition_clk ),
    .RESET_B(net1372),
    .D(_02460_),
    .Q_N(_07529_),
    .Q(\top1.memory2.mem2[176][1] ));
 sg13g2_dfrbp_1 _22364_ (.CLK(\clknet_leaf_130_top1.acquisition_clk ),
    .RESET_B(net1371),
    .D(_02461_),
    .Q_N(_07528_),
    .Q(\top1.memory2.mem2[176][2] ));
 sg13g2_dfrbp_1 _22365_ (.CLK(\clknet_leaf_133_top1.acquisition_clk ),
    .RESET_B(net1370),
    .D(_02462_),
    .Q_N(_07527_),
    .Q(\top1.memory2.mem2[177][0] ));
 sg13g2_dfrbp_1 _22366_ (.CLK(\clknet_leaf_131_top1.acquisition_clk ),
    .RESET_B(net1369),
    .D(_02463_),
    .Q_N(_07526_),
    .Q(\top1.memory2.mem2[177][1] ));
 sg13g2_dfrbp_1 _22367_ (.CLK(\clknet_leaf_129_top1.acquisition_clk ),
    .RESET_B(net1368),
    .D(_02464_),
    .Q_N(_07525_),
    .Q(\top1.memory2.mem2[177][2] ));
 sg13g2_dfrbp_1 _22368_ (.CLK(\clknet_leaf_134_top1.acquisition_clk ),
    .RESET_B(net1367),
    .D(_02465_),
    .Q_N(_07524_),
    .Q(\top1.memory2.mem2[178][0] ));
 sg13g2_dfrbp_1 _22369_ (.CLK(\clknet_leaf_131_top1.acquisition_clk ),
    .RESET_B(net1366),
    .D(_02466_),
    .Q_N(_07523_),
    .Q(\top1.memory2.mem2[178][1] ));
 sg13g2_dfrbp_1 _22370_ (.CLK(\clknet_leaf_130_top1.acquisition_clk ),
    .RESET_B(net1365),
    .D(_02467_),
    .Q_N(_07522_),
    .Q(\top1.memory2.mem2[178][2] ));
 sg13g2_dfrbp_1 _22371_ (.CLK(\clknet_leaf_112_top1.acquisition_clk ),
    .RESET_B(net1364),
    .D(_02468_),
    .Q_N(_07521_),
    .Q(\top1.memory2.mem2[17][0] ));
 sg13g2_dfrbp_1 _22372_ (.CLK(\clknet_leaf_119_top1.acquisition_clk ),
    .RESET_B(net1363),
    .D(_02469_),
    .Q_N(_07520_),
    .Q(\top1.memory2.mem2[17][1] ));
 sg13g2_dfrbp_1 _22373_ (.CLK(\clknet_leaf_120_top1.acquisition_clk ),
    .RESET_B(net1362),
    .D(_02470_),
    .Q_N(_07519_),
    .Q(\top1.memory2.mem2[17][2] ));
 sg13g2_dfrbp_1 _22374_ (.CLK(\clknet_leaf_114_top1.acquisition_clk ),
    .RESET_B(net1361),
    .D(_02471_),
    .Q_N(_07518_),
    .Q(\top1.memory2.mem2[180][0] ));
 sg13g2_dfrbp_1 _22375_ (.CLK(\clknet_leaf_181_top1.acquisition_clk ),
    .RESET_B(net1360),
    .D(_02472_),
    .Q_N(_07517_),
    .Q(\top1.memory2.mem2[180][1] ));
 sg13g2_dfrbp_1 _22376_ (.CLK(\clknet_leaf_176_top1.acquisition_clk ),
    .RESET_B(net1359),
    .D(_02473_),
    .Q_N(_07516_),
    .Q(\top1.memory2.mem2[180][2] ));
 sg13g2_dfrbp_1 _22377_ (.CLK(\clknet_leaf_114_top1.acquisition_clk ),
    .RESET_B(net1358),
    .D(_02474_),
    .Q_N(_07515_),
    .Q(\top1.memory2.mem2[181][0] ));
 sg13g2_dfrbp_1 _22378_ (.CLK(\clknet_leaf_181_top1.acquisition_clk ),
    .RESET_B(net1357),
    .D(_02475_),
    .Q_N(_07514_),
    .Q(\top1.memory2.mem2[181][1] ));
 sg13g2_dfrbp_1 _22379_ (.CLK(\clknet_leaf_181_top1.acquisition_clk ),
    .RESET_B(net1356),
    .D(_02476_),
    .Q_N(_07513_),
    .Q(\top1.memory2.mem2[181][2] ));
 sg13g2_dfrbp_1 _22380_ (.CLK(\clknet_leaf_176_top1.acquisition_clk ),
    .RESET_B(net1355),
    .D(_02477_),
    .Q_N(_07512_),
    .Q(\top1.memory2.mem2[182][0] ));
 sg13g2_dfrbp_1 _22381_ (.CLK(\clknet_leaf_177_top1.acquisition_clk ),
    .RESET_B(net1354),
    .D(_02478_),
    .Q_N(_07511_),
    .Q(\top1.memory2.mem2[182][1] ));
 sg13g2_dfrbp_1 _22382_ (.CLK(\clknet_leaf_177_top1.acquisition_clk ),
    .RESET_B(net1353),
    .D(_02479_),
    .Q_N(_07510_),
    .Q(\top1.memory2.mem2[182][2] ));
 sg13g2_dfrbp_1 _22383_ (.CLK(\clknet_leaf_176_top1.acquisition_clk ),
    .RESET_B(net1352),
    .D(_02480_),
    .Q_N(_07509_),
    .Q(\top1.memory2.mem2[183][0] ));
 sg13g2_dfrbp_1 _22384_ (.CLK(\clknet_leaf_177_top1.acquisition_clk ),
    .RESET_B(net1351),
    .D(_02481_),
    .Q_N(_07508_),
    .Q(\top1.memory2.mem2[183][1] ));
 sg13g2_dfrbp_1 _22385_ (.CLK(\clknet_leaf_177_top1.acquisition_clk ),
    .RESET_B(net1350),
    .D(_02482_),
    .Q_N(_07507_),
    .Q(\top1.memory2.mem2[183][2] ));
 sg13g2_dfrbp_1 _22386_ (.CLK(\clknet_leaf_112_top1.acquisition_clk ),
    .RESET_B(net1349),
    .D(_02483_),
    .Q_N(_07506_),
    .Q(\top1.memory2.mem2[184][0] ));
 sg13g2_dfrbp_1 _22387_ (.CLK(\clknet_leaf_128_top1.acquisition_clk ),
    .RESET_B(net1348),
    .D(_02484_),
    .Q_N(_07505_),
    .Q(\top1.memory2.mem2[184][1] ));
 sg13g2_dfrbp_1 _22388_ (.CLK(\clknet_leaf_127_top1.acquisition_clk ),
    .RESET_B(net1347),
    .D(_02485_),
    .Q_N(_07504_),
    .Q(\top1.memory2.mem2[184][2] ));
 sg13g2_dfrbp_1 _22389_ (.CLK(\clknet_leaf_112_top1.acquisition_clk ),
    .RESET_B(net1346),
    .D(_02486_),
    .Q_N(_07503_),
    .Q(\top1.memory2.mem2[185][0] ));
 sg13g2_dfrbp_1 _22390_ (.CLK(\clknet_leaf_128_top1.acquisition_clk ),
    .RESET_B(net1345),
    .D(_02487_),
    .Q_N(_07502_),
    .Q(\top1.memory2.mem2[185][1] ));
 sg13g2_dfrbp_1 _22391_ (.CLK(\clknet_leaf_127_top1.acquisition_clk ),
    .RESET_B(net1344),
    .D(_02488_),
    .Q_N(_07501_),
    .Q(\top1.memory2.mem2[185][2] ));
 sg13g2_dfrbp_1 _22392_ (.CLK(\clknet_leaf_115_top1.acquisition_clk ),
    .RESET_B(net1343),
    .D(_02489_),
    .Q_N(_07500_),
    .Q(\top1.memory2.mem2[186][0] ));
 sg13g2_dfrbp_1 _22393_ (.CLK(\clknet_leaf_129_top1.acquisition_clk ),
    .RESET_B(net1342),
    .D(_02490_),
    .Q_N(_07499_),
    .Q(\top1.memory2.mem2[186][1] ));
 sg13g2_dfrbp_1 _22394_ (.CLK(\clknet_leaf_129_top1.acquisition_clk ),
    .RESET_B(net1341),
    .D(_02491_),
    .Q_N(_07498_),
    .Q(\top1.memory2.mem2[186][2] ));
 sg13g2_dfrbp_1 _22395_ (.CLK(\clknet_leaf_115_top1.acquisition_clk ),
    .RESET_B(net1340),
    .D(_02492_),
    .Q_N(_07497_),
    .Q(\top1.memory2.mem2[187][0] ));
 sg13g2_dfrbp_1 _22396_ (.CLK(\clknet_leaf_129_top1.acquisition_clk ),
    .RESET_B(net1339),
    .D(_02493_),
    .Q_N(_07496_),
    .Q(\top1.memory2.mem2[187][1] ));
 sg13g2_dfrbp_1 _22397_ (.CLK(\clknet_leaf_130_top1.acquisition_clk ),
    .RESET_B(net1338),
    .D(_02494_),
    .Q_N(_07495_),
    .Q(\top1.memory2.mem2[187][2] ));
 sg13g2_dfrbp_1 _22398_ (.CLK(\clknet_leaf_118_top1.acquisition_clk ),
    .RESET_B(net1337),
    .D(_02495_),
    .Q_N(_07494_),
    .Q(\top1.memory2.mem2[188][0] ));
 sg13g2_dfrbp_1 _22399_ (.CLK(\clknet_leaf_116_top1.acquisition_clk ),
    .RESET_B(net1336),
    .D(_02496_),
    .Q_N(_07493_),
    .Q(\top1.memory2.mem2[188][1] ));
 sg13g2_dfrbp_1 _22400_ (.CLK(\clknet_leaf_118_top1.acquisition_clk ),
    .RESET_B(net1335),
    .D(_02497_),
    .Q_N(_07492_),
    .Q(\top1.memory2.mem2[188][2] ));
 sg13g2_dfrbp_1 _22401_ (.CLK(\clknet_leaf_113_top1.acquisition_clk ),
    .RESET_B(net1334),
    .D(_02498_),
    .Q_N(_07491_),
    .Q(\top1.memory2.mem2[18][0] ));
 sg13g2_dfrbp_1 _22402_ (.CLK(\clknet_leaf_119_top1.acquisition_clk ),
    .RESET_B(net1333),
    .D(_02499_),
    .Q_N(_07490_),
    .Q(\top1.memory2.mem2[18][1] ));
 sg13g2_dfrbp_1 _22403_ (.CLK(\clknet_leaf_113_top1.acquisition_clk ),
    .RESET_B(net1332),
    .D(_02500_),
    .Q_N(_07489_),
    .Q(\top1.memory2.mem2[18][2] ));
 sg13g2_dfrbp_1 _22404_ (.CLK(\clknet_leaf_135_top1.acquisition_clk ),
    .RESET_B(net1331),
    .D(_02501_),
    .Q_N(_07488_),
    .Q(\top1.memory2.mem2[190][0] ));
 sg13g2_dfrbp_1 _22405_ (.CLK(\clknet_leaf_116_top1.acquisition_clk ),
    .RESET_B(net1330),
    .D(_02502_),
    .Q_N(_07487_),
    .Q(\top1.memory2.mem2[190][1] ));
 sg13g2_dfrbp_1 _22406_ (.CLK(\clknet_leaf_118_top1.acquisition_clk ),
    .RESET_B(net1329),
    .D(_02503_),
    .Q_N(_07486_),
    .Q(\top1.memory2.mem2[190][2] ));
 sg13g2_dfrbp_1 _22407_ (.CLK(\clknet_leaf_135_top1.acquisition_clk ),
    .RESET_B(net1328),
    .D(_02504_),
    .Q_N(_07485_),
    .Q(\top1.memory2.mem2[191][0] ));
 sg13g2_dfrbp_1 _22408_ (.CLK(\clknet_leaf_116_top1.acquisition_clk ),
    .RESET_B(net1327),
    .D(_02505_),
    .Q_N(_07484_),
    .Q(\top1.memory2.mem2[191][1] ));
 sg13g2_dfrbp_1 _22409_ (.CLK(\clknet_leaf_118_top1.acquisition_clk ),
    .RESET_B(net1326),
    .D(_02506_),
    .Q_N(_07483_),
    .Q(\top1.memory2.mem2[191][2] ));
 sg13g2_dfrbp_1 _22410_ (.CLK(\clknet_leaf_98_top1.acquisition_clk ),
    .RESET_B(net1325),
    .D(_02507_),
    .Q_N(_07482_),
    .Q(\top1.memory2.mem2[192][0] ));
 sg13g2_dfrbp_1 _22411_ (.CLK(\clknet_leaf_98_top1.acquisition_clk ),
    .RESET_B(net1324),
    .D(_02508_),
    .Q_N(_07481_),
    .Q(\top1.memory2.mem2[192][1] ));
 sg13g2_dfrbp_1 _22412_ (.CLK(\clknet_leaf_95_top1.acquisition_clk ),
    .RESET_B(net1323),
    .D(_02509_),
    .Q_N(_07480_),
    .Q(\top1.memory2.mem2[192][2] ));
 sg13g2_dfrbp_1 _22413_ (.CLK(\clknet_leaf_96_top1.acquisition_clk ),
    .RESET_B(net1322),
    .D(_02510_),
    .Q_N(_07479_),
    .Q(\top1.memory2.mem2[193][0] ));
 sg13g2_dfrbp_1 _22414_ (.CLK(\clknet_leaf_99_top1.acquisition_clk ),
    .RESET_B(net1321),
    .D(_02511_),
    .Q_N(_07478_),
    .Q(\top1.memory2.mem2[193][1] ));
 sg13g2_dfrbp_1 _22415_ (.CLK(\clknet_leaf_95_top1.acquisition_clk ),
    .RESET_B(net1320),
    .D(_02512_),
    .Q_N(_07477_),
    .Q(\top1.memory2.mem2[193][2] ));
 sg13g2_dfrbp_1 _22416_ (.CLK(\clknet_leaf_97_top1.acquisition_clk ),
    .RESET_B(net1319),
    .D(_02513_),
    .Q_N(_07476_),
    .Q(\top1.memory2.mem2[194][0] ));
 sg13g2_dfrbp_1 _22417_ (.CLK(\clknet_leaf_98_top1.acquisition_clk ),
    .RESET_B(net1318),
    .D(_02514_),
    .Q_N(_07475_),
    .Q(\top1.memory2.mem2[194][1] ));
 sg13g2_dfrbp_1 _22418_ (.CLK(\clknet_leaf_95_top1.acquisition_clk ),
    .RESET_B(net1317),
    .D(_02515_),
    .Q_N(_07474_),
    .Q(\top1.memory2.mem2[194][2] ));
 sg13g2_dfrbp_1 _22419_ (.CLK(\clknet_leaf_97_top1.acquisition_clk ),
    .RESET_B(net1316),
    .D(_02516_),
    .Q_N(_07473_),
    .Q(\top1.memory2.mem2[195][0] ));
 sg13g2_dfrbp_1 _22420_ (.CLK(\clknet_leaf_98_top1.acquisition_clk ),
    .RESET_B(net1315),
    .D(_02517_),
    .Q_N(_07472_),
    .Q(\top1.memory2.mem2[195][1] ));
 sg13g2_dfrbp_1 _22421_ (.CLK(\clknet_leaf_98_top1.acquisition_clk ),
    .RESET_B(net1314),
    .D(_02518_),
    .Q_N(_07471_),
    .Q(\top1.memory2.mem2[195][2] ));
 sg13g2_dfrbp_1 _22422_ (.CLK(\clknet_leaf_99_top1.acquisition_clk ),
    .RESET_B(net1313),
    .D(_02519_),
    .Q_N(_07470_),
    .Q(\top1.memory2.mem2[196][0] ));
 sg13g2_dfrbp_1 _22423_ (.CLK(\clknet_leaf_38_top1.acquisition_clk ),
    .RESET_B(net1312),
    .D(_02520_),
    .Q_N(_07469_),
    .Q(\top1.memory2.mem2[196][1] ));
 sg13g2_dfrbp_1 _22424_ (.CLK(\clknet_leaf_98_top1.acquisition_clk ),
    .RESET_B(net1311),
    .D(_02521_),
    .Q_N(_07468_),
    .Q(\top1.memory2.mem2[196][2] ));
 sg13g2_dfrbp_1 _22425_ (.CLK(\clknet_leaf_99_top1.acquisition_clk ),
    .RESET_B(net1310),
    .D(_02522_),
    .Q_N(_07467_),
    .Q(\top1.memory2.mem2[197][0] ));
 sg13g2_dfrbp_1 _22426_ (.CLK(\clknet_leaf_38_top1.acquisition_clk ),
    .RESET_B(net1309),
    .D(_02523_),
    .Q_N(_07466_),
    .Q(\top1.memory2.mem2[197][1] ));
 sg13g2_dfrbp_1 _22427_ (.CLK(\clknet_leaf_99_top1.acquisition_clk ),
    .RESET_B(net1308),
    .D(_02524_),
    .Q_N(_07465_),
    .Q(\top1.memory2.mem2[197][2] ));
 sg13g2_dfrbp_1 _22428_ (.CLK(\clknet_leaf_41_top1.acquisition_clk ),
    .RESET_B(net1307),
    .D(_02525_),
    .Q_N(_07464_),
    .Q(\top1.memory2.mem2[198][0] ));
 sg13g2_dfrbp_1 _22429_ (.CLK(\clknet_leaf_39_top1.acquisition_clk ),
    .RESET_B(net1306),
    .D(_02526_),
    .Q_N(_07463_),
    .Q(\top1.memory2.mem2[198][1] ));
 sg13g2_dfrbp_1 _22430_ (.CLK(\clknet_leaf_98_top1.acquisition_clk ),
    .RESET_B(net1305),
    .D(_02527_),
    .Q_N(_07462_),
    .Q(\top1.memory2.mem2[198][2] ));
 sg13g2_tiehi _21295__34 (.L_HI(net34));
 sg13g2_tiehi _21294__35 (.L_HI(net35));
 sg13g2_tiehi _21293__36 (.L_HI(net36));
 sg13g2_tiehi _21292__37 (.L_HI(net37));
 sg13g2_tiehi _21291__38 (.L_HI(net38));
 sg13g2_tiehi _21290__39 (.L_HI(net39));
 sg13g2_tiehi _21289__40 (.L_HI(net40));
 sg13g2_tiehi _21288__41 (.L_HI(net41));
 sg13g2_tiehi _21287__42 (.L_HI(net42));
 sg13g2_tiehi _21286__43 (.L_HI(net43));
 sg13g2_tiehi _21285__44 (.L_HI(net44));
 sg13g2_tiehi _21284__45 (.L_HI(net45));
 sg13g2_tiehi _21283__46 (.L_HI(net46));
 sg13g2_tiehi _21282__47 (.L_HI(net47));
 sg13g2_tiehi _21281__48 (.L_HI(net48));
 sg13g2_tiehi _21280__49 (.L_HI(net49));
 sg13g2_tiehi _21279__50 (.L_HI(net50));
 sg13g2_tiehi _21278__51 (.L_HI(net51));
 sg13g2_tiehi _21277__52 (.L_HI(net52));
 sg13g2_tiehi _21276__53 (.L_HI(net53));
 sg13g2_tiehi _21275__54 (.L_HI(net54));
 sg13g2_tiehi _21274__55 (.L_HI(net55));
 sg13g2_tiehi _21273__56 (.L_HI(net56));
 sg13g2_tiehi _21272__57 (.L_HI(net57));
 sg13g2_tiehi _21271__58 (.L_HI(net58));
 sg13g2_tiehi _21270__59 (.L_HI(net59));
 sg13g2_tiehi _21269__60 (.L_HI(net60));
 sg13g2_tiehi _21268__61 (.L_HI(net61));
 sg13g2_tiehi _21267__62 (.L_HI(net62));
 sg13g2_tiehi _21266__63 (.L_HI(net63));
 sg13g2_tiehi _21265__64 (.L_HI(net64));
 sg13g2_tiehi _21264__65 (.L_HI(net65));
 sg13g2_tiehi _21263__66 (.L_HI(net66));
 sg13g2_tiehi _21262__67 (.L_HI(net67));
 sg13g2_tiehi _21261__68 (.L_HI(net68));
 sg13g2_tiehi _21260__69 (.L_HI(net69));
 sg13g2_tiehi _21259__70 (.L_HI(net70));
 sg13g2_tiehi _21258__71 (.L_HI(net71));
 sg13g2_tiehi _21257__72 (.L_HI(net72));
 sg13g2_tiehi _21256__73 (.L_HI(net73));
 sg13g2_tiehi _21255__74 (.L_HI(net74));
 sg13g2_tiehi _21254__75 (.L_HI(net75));
 sg13g2_tiehi _21253__76 (.L_HI(net76));
 sg13g2_tiehi _21252__77 (.L_HI(net77));
 sg13g2_tiehi _21251__78 (.L_HI(net78));
 sg13g2_tiehi _21250__79 (.L_HI(net79));
 sg13g2_tiehi _21249__80 (.L_HI(net80));
 sg13g2_tiehi _21248__81 (.L_HI(net81));
 sg13g2_tiehi _21247__82 (.L_HI(net82));
 sg13g2_tiehi _21246__83 (.L_HI(net83));
 sg13g2_tiehi _21245__84 (.L_HI(net84));
 sg13g2_tiehi _21244__85 (.L_HI(net85));
 sg13g2_tiehi _21243__86 (.L_HI(net86));
 sg13g2_tiehi _21242__87 (.L_HI(net87));
 sg13g2_tiehi _21241__88 (.L_HI(net88));
 sg13g2_tiehi _21240__89 (.L_HI(net89));
 sg13g2_tiehi _21239__90 (.L_HI(net90));
 sg13g2_tiehi _21238__91 (.L_HI(net91));
 sg13g2_tiehi _21237__92 (.L_HI(net92));
 sg13g2_tiehi _21236__93 (.L_HI(net93));
 sg13g2_tiehi _21235__94 (.L_HI(net94));
 sg13g2_tiehi _21234__95 (.L_HI(net95));
 sg13g2_tiehi _21233__96 (.L_HI(net96));
 sg13g2_tiehi _21232__97 (.L_HI(net97));
 sg13g2_tiehi _21231__98 (.L_HI(net98));
 sg13g2_tiehi _21225__99 (.L_HI(net99));
 sg13g2_tiehi _21224__100 (.L_HI(net100));
 sg13g2_tiehi _21135__101 (.L_HI(net101));
 sg13g2_tiehi _21134__102 (.L_HI(net102));
 sg13g2_tiehi _21133__103 (.L_HI(net103));
 sg13g2_tiehi _21132__104 (.L_HI(net104));
 sg13g2_tiehi _21131__105 (.L_HI(net105));
 sg13g2_tiehi _21130__106 (.L_HI(net106));
 sg13g2_tiehi _21129__107 (.L_HI(net107));
 sg13g2_tiehi _21128__108 (.L_HI(net108));
 sg13g2_tiehi _21127__109 (.L_HI(net109));
 sg13g2_tiehi _21126__110 (.L_HI(net110));
 sg13g2_tiehi _21125__111 (.L_HI(net111));
 sg13g2_tiehi _21124__112 (.L_HI(net112));
 sg13g2_tiehi _21123__113 (.L_HI(net113));
 sg13g2_tiehi _21122__114 (.L_HI(net114));
 sg13g2_tiehi _21121__115 (.L_HI(net115));
 sg13g2_tiehi _21120__116 (.L_HI(net116));
 sg13g2_tiehi _21119__117 (.L_HI(net117));
 sg13g2_tiehi _21118__118 (.L_HI(net118));
 sg13g2_tiehi _21117__119 (.L_HI(net119));
 sg13g2_tiehi _21116__120 (.L_HI(net120));
 sg13g2_tiehi _21115__121 (.L_HI(net121));
 sg13g2_tiehi _21114__122 (.L_HI(net122));
 sg13g2_tiehi _21113__123 (.L_HI(net123));
 sg13g2_tiehi _21112__124 (.L_HI(net124));
 sg13g2_tiehi _21111__125 (.L_HI(net125));
 sg13g2_tiehi _21110__126 (.L_HI(net126));
 sg13g2_tiehi _21109__127 (.L_HI(net127));
 sg13g2_tiehi _21108__128 (.L_HI(net128));
 sg13g2_tiehi _21107__129 (.L_HI(net129));
 sg13g2_tiehi _21106__130 (.L_HI(net130));
 sg13g2_tiehi _21105__131 (.L_HI(net131));
 sg13g2_tiehi _21104__132 (.L_HI(net132));
 sg13g2_tiehi _21103__133 (.L_HI(net133));
 sg13g2_tiehi _21102__134 (.L_HI(net134));
 sg13g2_tiehi _21101__135 (.L_HI(net135));
 sg13g2_tiehi _21100__136 (.L_HI(net136));
 sg13g2_tiehi _21099__137 (.L_HI(net137));
 sg13g2_tiehi _21098__138 (.L_HI(net138));
 sg13g2_tiehi _21097__139 (.L_HI(net139));
 sg13g2_tiehi _21096__140 (.L_HI(net140));
 sg13g2_tiehi _21095__141 (.L_HI(net141));
 sg13g2_tiehi _21094__142 (.L_HI(net142));
 sg13g2_tiehi _21093__143 (.L_HI(net143));
 sg13g2_tiehi _21092__144 (.L_HI(net144));
 sg13g2_tiehi _21091__145 (.L_HI(net145));
 sg13g2_tiehi _21090__146 (.L_HI(net146));
 sg13g2_tiehi _21089__147 (.L_HI(net147));
 sg13g2_tiehi _21088__148 (.L_HI(net148));
 sg13g2_tiehi _21087__149 (.L_HI(net149));
 sg13g2_tiehi _21086__150 (.L_HI(net150));
 sg13g2_tiehi _21085__151 (.L_HI(net151));
 sg13g2_tiehi _21084__152 (.L_HI(net152));
 sg13g2_tiehi _21083__153 (.L_HI(net153));
 sg13g2_tiehi _21082__154 (.L_HI(net154));
 sg13g2_tiehi _21081__155 (.L_HI(net155));
 sg13g2_tiehi _21080__156 (.L_HI(net156));
 sg13g2_tiehi _21079__157 (.L_HI(net157));
 sg13g2_tiehi _21078__158 (.L_HI(net158));
 sg13g2_tiehi _21077__159 (.L_HI(net159));
 sg13g2_tiehi _21076__160 (.L_HI(net160));
 sg13g2_tiehi _21075__161 (.L_HI(net161));
 sg13g2_tiehi _21074__162 (.L_HI(net162));
 sg13g2_tiehi _21073__163 (.L_HI(net163));
 sg13g2_tiehi _21072__164 (.L_HI(net164));
 sg13g2_tiehi _21071__165 (.L_HI(net165));
 sg13g2_tiehi _21070__166 (.L_HI(net166));
 sg13g2_tiehi _21069__167 (.L_HI(net167));
 sg13g2_tiehi _21068__168 (.L_HI(net168));
 sg13g2_tiehi _21067__169 (.L_HI(net169));
 sg13g2_tiehi _21066__170 (.L_HI(net170));
 sg13g2_tiehi _21065__171 (.L_HI(net171));
 sg13g2_tiehi _21064__172 (.L_HI(net172));
 sg13g2_tiehi _21063__173 (.L_HI(net173));
 sg13g2_tiehi _21062__174 (.L_HI(net174));
 sg13g2_tiehi _21061__175 (.L_HI(net175));
 sg13g2_tiehi _21060__176 (.L_HI(net176));
 sg13g2_tiehi _21059__177 (.L_HI(net177));
 sg13g2_tiehi _21058__178 (.L_HI(net178));
 sg13g2_tiehi _21057__179 (.L_HI(net179));
 sg13g2_tiehi _21056__180 (.L_HI(net180));
 sg13g2_tiehi _21055__181 (.L_HI(net181));
 sg13g2_tiehi _21054__182 (.L_HI(net182));
 sg13g2_tiehi _21053__183 (.L_HI(net183));
 sg13g2_tiehi _21052__184 (.L_HI(net184));
 sg13g2_tiehi _21051__185 (.L_HI(net185));
 sg13g2_tiehi _21050__186 (.L_HI(net186));
 sg13g2_tiehi _21049__187 (.L_HI(net187));
 sg13g2_tiehi _21048__188 (.L_HI(net188));
 sg13g2_tiehi _21047__189 (.L_HI(net189));
 sg13g2_tiehi _21046__190 (.L_HI(net190));
 sg13g2_tiehi _21045__191 (.L_HI(net191));
 sg13g2_tiehi _21044__192 (.L_HI(net192));
 sg13g2_tiehi _21043__193 (.L_HI(net193));
 sg13g2_tiehi _21042__194 (.L_HI(net194));
 sg13g2_tiehi _21041__195 (.L_HI(net195));
 sg13g2_tiehi _21040__196 (.L_HI(net196));
 sg13g2_tiehi _21039__197 (.L_HI(net197));
 sg13g2_tiehi _21038__198 (.L_HI(net198));
 sg13g2_tiehi _21037__199 (.L_HI(net199));
 sg13g2_tiehi _21036__200 (.L_HI(net200));
 sg13g2_tiehi _21035__201 (.L_HI(net201));
 sg13g2_tiehi _21034__202 (.L_HI(net202));
 sg13g2_tiehi _21033__203 (.L_HI(net203));
 sg13g2_tiehi _21032__204 (.L_HI(net204));
 sg13g2_tiehi _21031__205 (.L_HI(net205));
 sg13g2_tiehi _21030__206 (.L_HI(net206));
 sg13g2_tiehi _21029__207 (.L_HI(net207));
 sg13g2_tiehi _21028__208 (.L_HI(net208));
 sg13g2_tiehi _21027__209 (.L_HI(net209));
 sg13g2_tiehi _21026__210 (.L_HI(net210));
 sg13g2_tiehi _21025__211 (.L_HI(net211));
 sg13g2_tiehi _21024__212 (.L_HI(net212));
 sg13g2_tiehi _21023__213 (.L_HI(net213));
 sg13g2_tiehi _21022__214 (.L_HI(net214));
 sg13g2_tiehi _21021__215 (.L_HI(net215));
 sg13g2_tiehi _21020__216 (.L_HI(net216));
 sg13g2_tiehi _21019__217 (.L_HI(net217));
 sg13g2_tiehi _21018__218 (.L_HI(net218));
 sg13g2_tiehi _21017__219 (.L_HI(net219));
 sg13g2_tiehi _21016__220 (.L_HI(net220));
 sg13g2_tiehi _21015__221 (.L_HI(net221));
 sg13g2_tiehi _21014__222 (.L_HI(net222));
 sg13g2_tiehi _21013__223 (.L_HI(net223));
 sg13g2_tiehi _21012__224 (.L_HI(net224));
 sg13g2_tiehi _21011__225 (.L_HI(net225));
 sg13g2_tiehi _21010__226 (.L_HI(net226));
 sg13g2_tiehi _21009__227 (.L_HI(net227));
 sg13g2_tiehi _21008__228 (.L_HI(net228));
 sg13g2_tiehi _21007__229 (.L_HI(net229));
 sg13g2_tiehi _21006__230 (.L_HI(net230));
 sg13g2_tiehi _21005__231 (.L_HI(net231));
 sg13g2_tiehi _21004__232 (.L_HI(net232));
 sg13g2_tiehi _21003__233 (.L_HI(net233));
 sg13g2_tiehi _21002__234 (.L_HI(net234));
 sg13g2_tiehi _21001__235 (.L_HI(net235));
 sg13g2_tiehi _21000__236 (.L_HI(net236));
 sg13g2_tiehi _20999__237 (.L_HI(net237));
 sg13g2_tiehi _20998__238 (.L_HI(net238));
 sg13g2_tiehi _20997__239 (.L_HI(net239));
 sg13g2_tiehi _20996__240 (.L_HI(net240));
 sg13g2_tiehi _20995__241 (.L_HI(net241));
 sg13g2_tiehi _20994__242 (.L_HI(net242));
 sg13g2_tiehi _20993__243 (.L_HI(net243));
 sg13g2_tiehi _20992__244 (.L_HI(net244));
 sg13g2_tiehi _20980__245 (.L_HI(net245));
 sg13g2_tiehi _20979__246 (.L_HI(net246));
 sg13g2_tiehi _20978__247 (.L_HI(net247));
 sg13g2_tiehi _20971__248 (.L_HI(net248));
 sg13g2_tiehi _20970__249 (.L_HI(net249));
 sg13g2_tiehi _20969__250 (.L_HI(net250));
 sg13g2_tiehi _20968__251 (.L_HI(net251));
 sg13g2_tiehi _20967__252 (.L_HI(net252));
 sg13g2_tiehi _20964__253 (.L_HI(net253));
 sg13g2_tiehi _20963__254 (.L_HI(net254));
 sg13g2_tiehi _20962__255 (.L_HI(net255));
 sg13g2_tiehi _20951__256 (.L_HI(net256));
 sg13g2_tiehi _20950__257 (.L_HI(net257));
 sg13g2_tiehi _20949__258 (.L_HI(net258));
 sg13g2_tiehi _20948__259 (.L_HI(net259));
 sg13g2_tiehi _20947__260 (.L_HI(net260));
 sg13g2_tiehi _20946__261 (.L_HI(net261));
 sg13g2_tiehi _20945__262 (.L_HI(net262));
 sg13g2_tiehi _20944__263 (.L_HI(net263));
 sg13g2_tiehi _20943__264 (.L_HI(net264));
 sg13g2_tiehi _20942__265 (.L_HI(net265));
 sg13g2_tiehi _20941__266 (.L_HI(net266));
 sg13g2_tiehi _20940__267 (.L_HI(net267));
 sg13g2_tiehi _20939__268 (.L_HI(net268));
 sg13g2_tiehi _20938__269 (.L_HI(net269));
 sg13g2_tiehi _20937__270 (.L_HI(net270));
 sg13g2_tiehi _20936__271 (.L_HI(net271));
 sg13g2_tiehi _20935__272 (.L_HI(net272));
 sg13g2_tiehi _20934__273 (.L_HI(net273));
 sg13g2_tiehi _20933__274 (.L_HI(net274));
 sg13g2_tiehi _20932__275 (.L_HI(net275));
 sg13g2_tiehi _20931__276 (.L_HI(net276));
 sg13g2_tiehi _20930__277 (.L_HI(net277));
 sg13g2_tiehi _20929__278 (.L_HI(net278));
 sg13g2_tiehi _20928__279 (.L_HI(net279));
 sg13g2_tiehi _20927__280 (.L_HI(net280));
 sg13g2_tiehi _20926__281 (.L_HI(net281));
 sg13g2_tiehi _20925__282 (.L_HI(net282));
 sg13g2_tiehi _20924__283 (.L_HI(net283));
 sg13g2_tiehi _20923__284 (.L_HI(net284));
 sg13g2_tiehi _20922__285 (.L_HI(net285));
 sg13g2_tiehi _20921__286 (.L_HI(net286));
 sg13g2_tiehi _20920__287 (.L_HI(net287));
 sg13g2_tiehi _20919__288 (.L_HI(net288));
 sg13g2_tiehi _20918__289 (.L_HI(net289));
 sg13g2_tiehi _20917__290 (.L_HI(net290));
 sg13g2_tiehi _20916__291 (.L_HI(net291));
 sg13g2_tiehi _20915__292 (.L_HI(net292));
 sg13g2_tiehi _20914__293 (.L_HI(net293));
 sg13g2_tiehi _20913__294 (.L_HI(net294));
 sg13g2_tiehi _20912__295 (.L_HI(net295));
 sg13g2_tiehi _20911__296 (.L_HI(net296));
 sg13g2_tiehi _20910__297 (.L_HI(net297));
 sg13g2_tiehi _20909__298 (.L_HI(net298));
 sg13g2_tiehi _20908__299 (.L_HI(net299));
 sg13g2_tiehi _20907__300 (.L_HI(net300));
 sg13g2_tiehi _20906__301 (.L_HI(net301));
 sg13g2_tiehi _20905__302 (.L_HI(net302));
 sg13g2_tiehi _20904__303 (.L_HI(net303));
 sg13g2_tiehi _20903__304 (.L_HI(net304));
 sg13g2_tiehi _20902__305 (.L_HI(net305));
 sg13g2_tiehi _20901__306 (.L_HI(net306));
 sg13g2_tiehi _20900__307 (.L_HI(net307));
 sg13g2_tiehi _20899__308 (.L_HI(net308));
 sg13g2_tiehi _20898__309 (.L_HI(net309));
 sg13g2_tiehi _20897__310 (.L_HI(net310));
 sg13g2_tiehi _20896__311 (.L_HI(net311));
 sg13g2_tiehi _20895__312 (.L_HI(net312));
 sg13g2_tiehi _20892__313 (.L_HI(net313));
 sg13g2_tiehi _20891__314 (.L_HI(net314));
 sg13g2_tiehi _20890__315 (.L_HI(net315));
 sg13g2_tiehi _20889__316 (.L_HI(net316));
 sg13g2_tiehi _20888__317 (.L_HI(net317));
 sg13g2_tiehi _20887__318 (.L_HI(net318));
 sg13g2_tiehi _20886__319 (.L_HI(net319));
 sg13g2_tiehi _20885__320 (.L_HI(net320));
 sg13g2_tiehi _20884__321 (.L_HI(net321));
 sg13g2_tiehi _20883__322 (.L_HI(net322));
 sg13g2_tiehi _20882__323 (.L_HI(net323));
 sg13g2_tiehi _20881__324 (.L_HI(net324));
 sg13g2_tiehi _20880__325 (.L_HI(net325));
 sg13g2_tiehi _20879__326 (.L_HI(net326));
 sg13g2_tiehi _20878__327 (.L_HI(net327));
 sg13g2_tiehi _20877__328 (.L_HI(net328));
 sg13g2_tiehi _20876__329 (.L_HI(net329));
 sg13g2_tiehi _20875__330 (.L_HI(net330));
 sg13g2_tiehi _20874__331 (.L_HI(net331));
 sg13g2_tiehi _20873__332 (.L_HI(net332));
 sg13g2_tiehi _20872__333 (.L_HI(net333));
 sg13g2_tiehi _20871__334 (.L_HI(net334));
 sg13g2_tiehi _20870__335 (.L_HI(net335));
 sg13g2_tiehi _20869__336 (.L_HI(net336));
 sg13g2_tiehi _20868__337 (.L_HI(net337));
 sg13g2_tiehi _20867__338 (.L_HI(net338));
 sg13g2_tiehi _20866__339 (.L_HI(net339));
 sg13g2_tiehi _20865__340 (.L_HI(net340));
 sg13g2_tiehi _20864__341 (.L_HI(net341));
 sg13g2_tiehi _20863__342 (.L_HI(net342));
 sg13g2_tiehi _20862__343 (.L_HI(net343));
 sg13g2_tiehi _20861__344 (.L_HI(net344));
 sg13g2_tiehi _20860__345 (.L_HI(net345));
 sg13g2_tiehi _20859__346 (.L_HI(net346));
 sg13g2_tiehi _20858__347 (.L_HI(net347));
 sg13g2_tiehi _20857__348 (.L_HI(net348));
 sg13g2_tiehi _20856__349 (.L_HI(net349));
 sg13g2_tiehi _20855__350 (.L_HI(net350));
 sg13g2_tiehi _20854__351 (.L_HI(net351));
 sg13g2_tiehi _20853__352 (.L_HI(net352));
 sg13g2_tiehi _20852__353 (.L_HI(net353));
 sg13g2_tiehi _20851__354 (.L_HI(net354));
 sg13g2_tiehi _20850__355 (.L_HI(net355));
 sg13g2_tiehi _20849__356 (.L_HI(net356));
 sg13g2_tiehi _20848__357 (.L_HI(net357));
 sg13g2_tiehi _20847__358 (.L_HI(net358));
 sg13g2_tiehi _20846__359 (.L_HI(net359));
 sg13g2_tiehi _20845__360 (.L_HI(net360));
 sg13g2_tiehi _20844__361 (.L_HI(net361));
 sg13g2_tiehi _20843__362 (.L_HI(net362));
 sg13g2_tiehi _20842__363 (.L_HI(net363));
 sg13g2_tiehi _20839__364 (.L_HI(net364));
 sg13g2_tiehi _20838__365 (.L_HI(net365));
 sg13g2_tiehi _20820__366 (.L_HI(net366));
 sg13g2_tiehi _20819__367 (.L_HI(net367));
 sg13g2_tiehi _20818__368 (.L_HI(net368));
 sg13g2_tiehi _20811__369 (.L_HI(net369));
 sg13g2_tiehi _20810__370 (.L_HI(net370));
 sg13g2_tiehi _20809__371 (.L_HI(net371));
 sg13g2_tiehi _20808__372 (.L_HI(net372));
 sg13g2_tiehi _20807__373 (.L_HI(net373));
 sg13g2_tiehi _20806__374 (.L_HI(net374));
 sg13g2_tiehi _20805__375 (.L_HI(net375));
 sg13g2_tiehi _20804__376 (.L_HI(net376));
 sg13g2_tiehi _20803__377 (.L_HI(net377));
 sg13g2_tiehi _20802__378 (.L_HI(net378));
 sg13g2_tiehi _20801__379 (.L_HI(net379));
 sg13g2_tiehi _20800__380 (.L_HI(net380));
 sg13g2_tiehi _20799__381 (.L_HI(net381));
 sg13g2_tiehi _20798__382 (.L_HI(net382));
 sg13g2_tiehi _20797__383 (.L_HI(net383));
 sg13g2_tiehi _20794__384 (.L_HI(net384));
 sg13g2_tiehi _20793__385 (.L_HI(net385));
 sg13g2_tiehi _20792__386 (.L_HI(net386));
 sg13g2_tiehi _20791__387 (.L_HI(net387));
 sg13g2_tiehi _20790__388 (.L_HI(net388));
 sg13g2_tiehi _20789__389 (.L_HI(net389));
 sg13g2_tiehi _20788__390 (.L_HI(net390));
 sg13g2_tiehi _20787__391 (.L_HI(net391));
 sg13g2_tiehi _20786__392 (.L_HI(net392));
 sg13g2_tiehi _20785__393 (.L_HI(net393));
 sg13g2_tiehi _20784__394 (.L_HI(net394));
 sg13g2_tiehi _20783__395 (.L_HI(net395));
 sg13g2_tiehi _20782__396 (.L_HI(net396));
 sg13g2_tiehi _20781__397 (.L_HI(net397));
 sg13g2_tiehi _20780__398 (.L_HI(net398));
 sg13g2_tiehi _20779__399 (.L_HI(net399));
 sg13g2_tiehi _20778__400 (.L_HI(net400));
 sg13g2_tiehi _20777__401 (.L_HI(net401));
 sg13g2_tiehi _20776__402 (.L_HI(net402));
 sg13g2_tiehi _20775__403 (.L_HI(net403));
 sg13g2_tiehi _20774__404 (.L_HI(net404));
 sg13g2_tiehi _20773__405 (.L_HI(net405));
 sg13g2_tiehi _20772__406 (.L_HI(net406));
 sg13g2_tiehi _20771__407 (.L_HI(net407));
 sg13g2_tiehi _20770__408 (.L_HI(net408));
 sg13g2_tiehi _20769__409 (.L_HI(net409));
 sg13g2_tiehi _20768__410 (.L_HI(net410));
 sg13g2_tiehi _20767__411 (.L_HI(net411));
 sg13g2_tiehi _20766__412 (.L_HI(net412));
 sg13g2_tiehi _20765__413 (.L_HI(net413));
 sg13g2_tiehi _20764__414 (.L_HI(net414));
 sg13g2_tiehi _20763__415 (.L_HI(net415));
 sg13g2_tiehi _20762__416 (.L_HI(net416));
 sg13g2_tiehi _20761__417 (.L_HI(net417));
 sg13g2_tiehi _20760__418 (.L_HI(net418));
 sg13g2_tiehi _20759__419 (.L_HI(net419));
 sg13g2_tiehi _20758__420 (.L_HI(net420));
 sg13g2_tiehi _20757__421 (.L_HI(net421));
 sg13g2_tiehi _20756__422 (.L_HI(net422));
 sg13g2_tiehi _20755__423 (.L_HI(net423));
 sg13g2_tiehi _20754__424 (.L_HI(net424));
 sg13g2_tiehi _20753__425 (.L_HI(net425));
 sg13g2_tiehi _20752__426 (.L_HI(net426));
 sg13g2_tiehi _20751__427 (.L_HI(net427));
 sg13g2_tiehi _20750__428 (.L_HI(net428));
 sg13g2_tiehi _20749__429 (.L_HI(net429));
 sg13g2_tiehi _20748__430 (.L_HI(net430));
 sg13g2_tiehi _20747__431 (.L_HI(net431));
 sg13g2_tiehi _20746__432 (.L_HI(net432));
 sg13g2_tiehi _20745__433 (.L_HI(net433));
 sg13g2_tiehi _20744__434 (.L_HI(net434));
 sg13g2_tiehi _20743__435 (.L_HI(net435));
 sg13g2_tiehi _20742__436 (.L_HI(net436));
 sg13g2_tiehi _20741__437 (.L_HI(net437));
 sg13g2_tiehi _20740__438 (.L_HI(net438));
 sg13g2_tiehi _20739__439 (.L_HI(net439));
 sg13g2_tiehi _20738__440 (.L_HI(net440));
 sg13g2_tiehi _20737__441 (.L_HI(net441));
 sg13g2_tiehi _20736__442 (.L_HI(net442));
 sg13g2_tiehi _20735__443 (.L_HI(net443));
 sg13g2_tiehi _20734__444 (.L_HI(net444));
 sg13g2_tiehi _20733__445 (.L_HI(net445));
 sg13g2_tiehi _20732__446 (.L_HI(net446));
 sg13g2_tiehi _20731__447 (.L_HI(net447));
 sg13g2_tiehi _20730__448 (.L_HI(net448));
 sg13g2_tiehi _20729__449 (.L_HI(net449));
 sg13g2_tiehi _20728__450 (.L_HI(net450));
 sg13g2_tiehi _20727__451 (.L_HI(net451));
 sg13g2_tiehi _20726__452 (.L_HI(net452));
 sg13g2_tiehi _20725__453 (.L_HI(net453));
 sg13g2_tiehi _20724__454 (.L_HI(net454));
 sg13g2_tiehi _20723__455 (.L_HI(net455));
 sg13g2_tiehi _20722__456 (.L_HI(net456));
 sg13g2_tiehi _20721__457 (.L_HI(net457));
 sg13g2_tiehi _20720__458 (.L_HI(net458));
 sg13g2_tiehi _20719__459 (.L_HI(net459));
 sg13g2_tiehi _20718__460 (.L_HI(net460));
 sg13g2_tiehi _20717__461 (.L_HI(net461));
 sg13g2_tiehi _20716__462 (.L_HI(net462));
 sg13g2_tiehi _20715__463 (.L_HI(net463));
 sg13g2_tiehi _20714__464 (.L_HI(net464));
 sg13g2_tiehi _20713__465 (.L_HI(net465));
 sg13g2_tiehi _20712__466 (.L_HI(net466));
 sg13g2_tiehi _20711__467 (.L_HI(net467));
 sg13g2_tiehi _20710__468 (.L_HI(net468));
 sg13g2_tiehi _20709__469 (.L_HI(net469));
 sg13g2_tiehi _20708__470 (.L_HI(net470));
 sg13g2_tiehi _20707__471 (.L_HI(net471));
 sg13g2_tiehi _20706__472 (.L_HI(net472));
 sg13g2_tiehi _20705__473 (.L_HI(net473));
 sg13g2_tiehi _20704__474 (.L_HI(net474));
 sg13g2_tiehi _20703__475 (.L_HI(net475));
 sg13g2_tiehi _20702__476 (.L_HI(net476));
 sg13g2_tiehi _20701__477 (.L_HI(net477));
 sg13g2_tiehi _20700__478 (.L_HI(net478));
 sg13g2_tiehi _20699__479 (.L_HI(net479));
 sg13g2_tiehi _20698__480 (.L_HI(net480));
 sg13g2_tiehi _20697__481 (.L_HI(net481));
 sg13g2_tiehi _20696__482 (.L_HI(net482));
 sg13g2_tiehi _20695__483 (.L_HI(net483));
 sg13g2_tiehi _20694__484 (.L_HI(net484));
 sg13g2_tiehi _20693__485 (.L_HI(net485));
 sg13g2_tiehi _20692__486 (.L_HI(net486));
 sg13g2_tiehi _20691__487 (.L_HI(net487));
 sg13g2_tiehi _20690__488 (.L_HI(net488));
 sg13g2_tiehi _20689__489 (.L_HI(net489));
 sg13g2_tiehi _20688__490 (.L_HI(net490));
 sg13g2_tiehi _20687__491 (.L_HI(net491));
 sg13g2_tiehi _20686__492 (.L_HI(net492));
 sg13g2_tiehi _20685__493 (.L_HI(net493));
 sg13g2_tiehi _20684__494 (.L_HI(net494));
 sg13g2_tiehi _20683__495 (.L_HI(net495));
 sg13g2_tiehi _20682__496 (.L_HI(net496));
 sg13g2_tiehi _20681__497 (.L_HI(net497));
 sg13g2_tiehi _20680__498 (.L_HI(net498));
 sg13g2_tiehi _20679__499 (.L_HI(net499));
 sg13g2_tiehi _20678__500 (.L_HI(net500));
 sg13g2_tiehi _20677__501 (.L_HI(net501));
 sg13g2_tiehi _20676__502 (.L_HI(net502));
 sg13g2_tiehi _20675__503 (.L_HI(net503));
 sg13g2_tiehi _20674__504 (.L_HI(net504));
 sg13g2_tiehi _20673__505 (.L_HI(net505));
 sg13g2_tiehi _20672__506 (.L_HI(net506));
 sg13g2_tiehi _20671__507 (.L_HI(net507));
 sg13g2_tiehi _20670__508 (.L_HI(net508));
 sg13g2_tiehi _20669__509 (.L_HI(net509));
 sg13g2_tiehi _20668__510 (.L_HI(net510));
 sg13g2_tiehi _20667__511 (.L_HI(net511));
 sg13g2_tiehi _20666__512 (.L_HI(net512));
 sg13g2_tiehi _20665__513 (.L_HI(net513));
 sg13g2_tiehi _20664__514 (.L_HI(net514));
 sg13g2_tiehi _20663__515 (.L_HI(net515));
 sg13g2_tiehi _20662__516 (.L_HI(net516));
 sg13g2_tiehi _20661__517 (.L_HI(net517));
 sg13g2_tiehi _20660__518 (.L_HI(net518));
 sg13g2_tiehi _20659__519 (.L_HI(net519));
 sg13g2_tiehi _20658__520 (.L_HI(net520));
 sg13g2_tiehi _20657__521 (.L_HI(net521));
 sg13g2_tiehi _20656__522 (.L_HI(net522));
 sg13g2_tiehi _20655__523 (.L_HI(net523));
 sg13g2_tiehi _20654__524 (.L_HI(net524));
 sg13g2_tiehi _20653__525 (.L_HI(net525));
 sg13g2_tiehi _20652__526 (.L_HI(net526));
 sg13g2_tiehi _20651__527 (.L_HI(net527));
 sg13g2_tiehi _20650__528 (.L_HI(net528));
 sg13g2_tiehi _20649__529 (.L_HI(net529));
 sg13g2_tiehi _20648__530 (.L_HI(net530));
 sg13g2_tiehi _20647__531 (.L_HI(net531));
 sg13g2_tiehi _20646__532 (.L_HI(net532));
 sg13g2_tiehi _20645__533 (.L_HI(net533));
 sg13g2_tiehi _20644__534 (.L_HI(net534));
 sg13g2_tiehi _20643__535 (.L_HI(net535));
 sg13g2_tiehi _20642__536 (.L_HI(net536));
 sg13g2_tiehi _20641__537 (.L_HI(net537));
 sg13g2_tiehi _20640__538 (.L_HI(net538));
 sg13g2_tiehi _20639__539 (.L_HI(net539));
 sg13g2_tiehi _20638__540 (.L_HI(net540));
 sg13g2_tiehi _20637__541 (.L_HI(net541));
 sg13g2_tiehi _20636__542 (.L_HI(net542));
 sg13g2_tiehi _20635__543 (.L_HI(net543));
 sg13g2_tiehi _20634__544 (.L_HI(net544));
 sg13g2_tiehi _20633__545 (.L_HI(net545));
 sg13g2_tiehi _20632__546 (.L_HI(net546));
 sg13g2_tiehi _20631__547 (.L_HI(net547));
 sg13g2_tiehi _20630__548 (.L_HI(net548));
 sg13g2_tiehi _20629__549 (.L_HI(net549));
 sg13g2_tiehi _20628__550 (.L_HI(net550));
 sg13g2_tiehi _20627__551 (.L_HI(net551));
 sg13g2_tiehi _20626__552 (.L_HI(net552));
 sg13g2_tiehi _20625__553 (.L_HI(net553));
 sg13g2_tiehi _20624__554 (.L_HI(net554));
 sg13g2_tiehi _20623__555 (.L_HI(net555));
 sg13g2_tiehi _20622__556 (.L_HI(net556));
 sg13g2_tiehi _20621__557 (.L_HI(net557));
 sg13g2_tiehi _20620__558 (.L_HI(net558));
 sg13g2_tiehi _20619__559 (.L_HI(net559));
 sg13g2_tiehi _20618__560 (.L_HI(net560));
 sg13g2_tiehi _20617__561 (.L_HI(net561));
 sg13g2_tiehi _20616__562 (.L_HI(net562));
 sg13g2_tiehi _20615__563 (.L_HI(net563));
 sg13g2_tiehi _20614__564 (.L_HI(net564));
 sg13g2_tiehi _20613__565 (.L_HI(net565));
 sg13g2_tiehi _20612__566 (.L_HI(net566));
 sg13g2_tiehi _20611__567 (.L_HI(net567));
 sg13g2_tiehi _20610__568 (.L_HI(net568));
 sg13g2_tiehi _20609__569 (.L_HI(net569));
 sg13g2_tiehi _20608__570 (.L_HI(net570));
 sg13g2_tiehi _20607__571 (.L_HI(net571));
 sg13g2_tiehi _20606__572 (.L_HI(net572));
 sg13g2_tiehi _20605__573 (.L_HI(net573));
 sg13g2_tiehi _20604__574 (.L_HI(net574));
 sg13g2_tiehi _20603__575 (.L_HI(net575));
 sg13g2_tiehi _20602__576 (.L_HI(net576));
 sg13g2_tiehi _20601__577 (.L_HI(net577));
 sg13g2_tiehi _20600__578 (.L_HI(net578));
 sg13g2_tiehi _20599__579 (.L_HI(net579));
 sg13g2_tiehi _20598__580 (.L_HI(net580));
 sg13g2_tiehi _20597__581 (.L_HI(net581));
 sg13g2_tiehi _20596__582 (.L_HI(net582));
 sg13g2_tiehi _20595__583 (.L_HI(net583));
 sg13g2_tiehi _20594__584 (.L_HI(net584));
 sg13g2_tiehi _20593__585 (.L_HI(net585));
 sg13g2_tiehi _20592__586 (.L_HI(net586));
 sg13g2_tiehi _20591__587 (.L_HI(net587));
 sg13g2_tiehi _20590__588 (.L_HI(net588));
 sg13g2_tiehi _20589__589 (.L_HI(net589));
 sg13g2_tiehi _20588__590 (.L_HI(net590));
 sg13g2_tiehi _20587__591 (.L_HI(net591));
 sg13g2_tiehi _20586__592 (.L_HI(net592));
 sg13g2_tiehi _20585__593 (.L_HI(net593));
 sg13g2_tiehi _20584__594 (.L_HI(net594));
 sg13g2_tiehi _20583__595 (.L_HI(net595));
 sg13g2_tiehi _20582__596 (.L_HI(net596));
 sg13g2_tiehi _20581__597 (.L_HI(net597));
 sg13g2_tiehi _20580__598 (.L_HI(net598));
 sg13g2_tiehi _20579__599 (.L_HI(net599));
 sg13g2_tiehi _20578__600 (.L_HI(net600));
 sg13g2_tiehi _20577__601 (.L_HI(net601));
 sg13g2_tiehi _20576__602 (.L_HI(net602));
 sg13g2_tiehi _20575__603 (.L_HI(net603));
 sg13g2_tiehi _20574__604 (.L_HI(net604));
 sg13g2_tiehi _20573__605 (.L_HI(net605));
 sg13g2_tiehi _20572__606 (.L_HI(net606));
 sg13g2_tiehi _20571__607 (.L_HI(net607));
 sg13g2_tiehi _20570__608 (.L_HI(net608));
 sg13g2_tiehi _20569__609 (.L_HI(net609));
 sg13g2_tiehi _20568__610 (.L_HI(net610));
 sg13g2_tiehi _20567__611 (.L_HI(net611));
 sg13g2_tiehi _20566__612 (.L_HI(net612));
 sg13g2_tiehi _20565__613 (.L_HI(net613));
 sg13g2_tiehi _20564__614 (.L_HI(net614));
 sg13g2_tiehi _20563__615 (.L_HI(net615));
 sg13g2_tiehi _20562__616 (.L_HI(net616));
 sg13g2_tiehi _20561__617 (.L_HI(net617));
 sg13g2_tiehi _20560__618 (.L_HI(net618));
 sg13g2_tiehi _20559__619 (.L_HI(net619));
 sg13g2_tiehi _20553__620 (.L_HI(net620));
 sg13g2_tiehi _20552__621 (.L_HI(net621));
 sg13g2_tiehi _20551__622 (.L_HI(net622));
 sg13g2_tiehi _20550__623 (.L_HI(net623));
 sg13g2_tiehi _20549__624 (.L_HI(net624));
 sg13g2_tiehi _20548__625 (.L_HI(net625));
 sg13g2_tiehi _20547__626 (.L_HI(net626));
 sg13g2_tiehi _20546__627 (.L_HI(net627));
 sg13g2_tiehi _20545__628 (.L_HI(net628));
 sg13g2_tiehi _20544__629 (.L_HI(net629));
 sg13g2_tiehi _20543__630 (.L_HI(net630));
 sg13g2_tiehi _20542__631 (.L_HI(net631));
 sg13g2_tiehi _20541__632 (.L_HI(net632));
 sg13g2_tiehi _20540__633 (.L_HI(net633));
 sg13g2_tiehi _20539__634 (.L_HI(net634));
 sg13g2_tiehi _20538__635 (.L_HI(net635));
 sg13g2_tiehi _20537__636 (.L_HI(net636));
 sg13g2_tiehi _20536__637 (.L_HI(net637));
 sg13g2_tiehi _20535__638 (.L_HI(net638));
 sg13g2_tiehi _20534__639 (.L_HI(net639));
 sg13g2_tiehi _20533__640 (.L_HI(net640));
 sg13g2_tiehi _20532__641 (.L_HI(net641));
 sg13g2_tiehi _20531__642 (.L_HI(net642));
 sg13g2_tiehi _20530__643 (.L_HI(net643));
 sg13g2_tiehi _20529__644 (.L_HI(net644));
 sg13g2_tiehi _20528__645 (.L_HI(net645));
 sg13g2_tiehi _20527__646 (.L_HI(net646));
 sg13g2_tiehi _20526__647 (.L_HI(net647));
 sg13g2_tiehi _20525__648 (.L_HI(net648));
 sg13g2_tiehi _20524__649 (.L_HI(net649));
 sg13g2_tiehi _20523__650 (.L_HI(net650));
 sg13g2_tiehi _20522__651 (.L_HI(net651));
 sg13g2_tiehi _20521__652 (.L_HI(net652));
 sg13g2_tiehi _20520__653 (.L_HI(net653));
 sg13g2_tiehi _20519__654 (.L_HI(net654));
 sg13g2_tiehi _20518__655 (.L_HI(net655));
 sg13g2_tiehi _20517__656 (.L_HI(net656));
 sg13g2_tiehi _20516__657 (.L_HI(net657));
 sg13g2_tiehi _20515__658 (.L_HI(net658));
 sg13g2_tiehi _20514__659 (.L_HI(net659));
 sg13g2_tiehi _20513__660 (.L_HI(net660));
 sg13g2_tiehi _20512__661 (.L_HI(net661));
 sg13g2_tiehi _20511__662 (.L_HI(net662));
 sg13g2_tiehi _20510__663 (.L_HI(net663));
 sg13g2_tiehi _20509__664 (.L_HI(net664));
 sg13g2_tiehi _20508__665 (.L_HI(net665));
 sg13g2_tiehi _20507__666 (.L_HI(net666));
 sg13g2_tiehi _20506__667 (.L_HI(net667));
 sg13g2_tiehi _20505__668 (.L_HI(net668));
 sg13g2_tiehi _20504__669 (.L_HI(net669));
 sg13g2_tiehi _20503__670 (.L_HI(net670));
 sg13g2_tiehi _20502__671 (.L_HI(net671));
 sg13g2_tiehi _20501__672 (.L_HI(net672));
 sg13g2_tiehi _20500__673 (.L_HI(net673));
 sg13g2_tiehi _20499__674 (.L_HI(net674));
 sg13g2_tiehi _20498__675 (.L_HI(net675));
 sg13g2_tiehi _20497__676 (.L_HI(net676));
 sg13g2_tiehi _20496__677 (.L_HI(net677));
 sg13g2_tiehi _20495__678 (.L_HI(net678));
 sg13g2_tiehi _20494__679 (.L_HI(net679));
 sg13g2_tiehi _20493__680 (.L_HI(net680));
 sg13g2_tiehi _20492__681 (.L_HI(net681));
 sg13g2_tiehi _20491__682 (.L_HI(net682));
 sg13g2_tiehi _20490__683 (.L_HI(net683));
 sg13g2_tiehi _20489__684 (.L_HI(net684));
 sg13g2_tiehi _20488__685 (.L_HI(net685));
 sg13g2_tiehi _20487__686 (.L_HI(net686));
 sg13g2_tiehi _20486__687 (.L_HI(net687));
 sg13g2_tiehi _20485__688 (.L_HI(net688));
 sg13g2_tiehi _20484__689 (.L_HI(net689));
 sg13g2_tiehi _20483__690 (.L_HI(net690));
 sg13g2_tiehi _20482__691 (.L_HI(net691));
 sg13g2_tiehi _20481__692 (.L_HI(net692));
 sg13g2_tiehi _20480__693 (.L_HI(net693));
 sg13g2_tiehi _20479__694 (.L_HI(net694));
 sg13g2_tiehi _20478__695 (.L_HI(net695));
 sg13g2_tiehi _20477__696 (.L_HI(net696));
 sg13g2_tiehi _20476__697 (.L_HI(net697));
 sg13g2_tiehi _20475__698 (.L_HI(net698));
 sg13g2_tiehi _20474__699 (.L_HI(net699));
 sg13g2_tiehi _20473__700 (.L_HI(net700));
 sg13g2_tiehi _20472__701 (.L_HI(net701));
 sg13g2_tiehi _20471__702 (.L_HI(net702));
 sg13g2_tiehi _20470__703 (.L_HI(net703));
 sg13g2_tiehi _20469__704 (.L_HI(net704));
 sg13g2_tiehi _20468__705 (.L_HI(net705));
 sg13g2_tiehi _20467__706 (.L_HI(net706));
 sg13g2_tiehi _20466__707 (.L_HI(net707));
 sg13g2_tiehi _20465__708 (.L_HI(net708));
 sg13g2_tiehi _20464__709 (.L_HI(net709));
 sg13g2_tiehi _20463__710 (.L_HI(net710));
 sg13g2_tiehi _20462__711 (.L_HI(net711));
 sg13g2_tiehi _20461__712 (.L_HI(net712));
 sg13g2_tiehi _20460__713 (.L_HI(net713));
 sg13g2_tiehi _20459__714 (.L_HI(net714));
 sg13g2_tiehi _20458__715 (.L_HI(net715));
 sg13g2_tiehi _20457__716 (.L_HI(net716));
 sg13g2_tiehi _20456__717 (.L_HI(net717));
 sg13g2_tiehi _20455__718 (.L_HI(net718));
 sg13g2_tiehi _20454__719 (.L_HI(net719));
 sg13g2_tiehi _20453__720 (.L_HI(net720));
 sg13g2_tiehi _20452__721 (.L_HI(net721));
 sg13g2_tiehi _20451__722 (.L_HI(net722));
 sg13g2_tiehi _20450__723 (.L_HI(net723));
 sg13g2_tiehi _20449__724 (.L_HI(net724));
 sg13g2_tiehi _20448__725 (.L_HI(net725));
 sg13g2_tiehi _20447__726 (.L_HI(net726));
 sg13g2_tiehi _20446__727 (.L_HI(net727));
 sg13g2_tiehi _20445__728 (.L_HI(net728));
 sg13g2_tiehi _20444__729 (.L_HI(net729));
 sg13g2_tiehi _20443__730 (.L_HI(net730));
 sg13g2_tiehi _20442__731 (.L_HI(net731));
 sg13g2_tiehi _20441__732 (.L_HI(net732));
 sg13g2_tiehi _20440__733 (.L_HI(net733));
 sg13g2_tiehi _20439__734 (.L_HI(net734));
 sg13g2_tiehi _20438__735 (.L_HI(net735));
 sg13g2_tiehi _20437__736 (.L_HI(net736));
 sg13g2_tiehi _20436__737 (.L_HI(net737));
 sg13g2_tiehi _20435__738 (.L_HI(net738));
 sg13g2_tiehi _20434__739 (.L_HI(net739));
 sg13g2_tiehi _20433__740 (.L_HI(net740));
 sg13g2_tiehi _20432__741 (.L_HI(net741));
 sg13g2_tiehi _20431__742 (.L_HI(net742));
 sg13g2_tiehi _20430__743 (.L_HI(net743));
 sg13g2_tiehi _20429__744 (.L_HI(net744));
 sg13g2_tiehi _20428__745 (.L_HI(net745));
 sg13g2_tiehi _20427__746 (.L_HI(net746));
 sg13g2_tiehi _20426__747 (.L_HI(net747));
 sg13g2_tiehi _20425__748 (.L_HI(net748));
 sg13g2_tiehi _20424__749 (.L_HI(net749));
 sg13g2_tiehi _20423__750 (.L_HI(net750));
 sg13g2_tiehi _20422__751 (.L_HI(net751));
 sg13g2_tiehi _20421__752 (.L_HI(net752));
 sg13g2_tiehi _20420__753 (.L_HI(net753));
 sg13g2_tiehi _20419__754 (.L_HI(net754));
 sg13g2_tiehi _20418__755 (.L_HI(net755));
 sg13g2_tiehi _20417__756 (.L_HI(net756));
 sg13g2_tiehi _20416__757 (.L_HI(net757));
 sg13g2_tiehi _20415__758 (.L_HI(net758));
 sg13g2_tiehi _20414__759 (.L_HI(net759));
 sg13g2_tiehi _20413__760 (.L_HI(net760));
 sg13g2_tiehi _20412__761 (.L_HI(net761));
 sg13g2_tiehi _20411__762 (.L_HI(net762));
 sg13g2_tiehi _20410__763 (.L_HI(net763));
 sg13g2_tiehi _20409__764 (.L_HI(net764));
 sg13g2_tiehi _20408__765 (.L_HI(net765));
 sg13g2_tiehi _20407__766 (.L_HI(net766));
 sg13g2_tiehi _20406__767 (.L_HI(net767));
 sg13g2_tiehi _20405__768 (.L_HI(net768));
 sg13g2_tiehi _20404__769 (.L_HI(net769));
 sg13g2_tiehi _20403__770 (.L_HI(net770));
 sg13g2_tiehi _20402__771 (.L_HI(net771));
 sg13g2_tiehi _20401__772 (.L_HI(net772));
 sg13g2_tiehi _20400__773 (.L_HI(net773));
 sg13g2_tiehi _20399__774 (.L_HI(net774));
 sg13g2_tiehi _20398__775 (.L_HI(net775));
 sg13g2_tiehi _20397__776 (.L_HI(net776));
 sg13g2_tiehi _20396__777 (.L_HI(net777));
 sg13g2_tiehi _20395__778 (.L_HI(net778));
 sg13g2_tiehi _20394__779 (.L_HI(net779));
 sg13g2_tiehi _20393__780 (.L_HI(net780));
 sg13g2_tiehi _20392__781 (.L_HI(net781));
 sg13g2_tiehi _20391__782 (.L_HI(net782));
 sg13g2_tiehi _20390__783 (.L_HI(net783));
 sg13g2_tiehi _20389__784 (.L_HI(net784));
 sg13g2_tiehi _20388__785 (.L_HI(net785));
 sg13g2_tiehi _20387__786 (.L_HI(net786));
 sg13g2_tiehi _20386__787 (.L_HI(net787));
 sg13g2_tiehi _20385__788 (.L_HI(net788));
 sg13g2_tiehi _20384__789 (.L_HI(net789));
 sg13g2_tiehi _20383__790 (.L_HI(net790));
 sg13g2_tiehi _20382__791 (.L_HI(net791));
 sg13g2_tiehi _20381__792 (.L_HI(net792));
 sg13g2_tiehi _20380__793 (.L_HI(net793));
 sg13g2_tiehi _20379__794 (.L_HI(net794));
 sg13g2_tiehi _20378__795 (.L_HI(net795));
 sg13g2_tiehi _20377__796 (.L_HI(net796));
 sg13g2_tiehi _20376__797 (.L_HI(net797));
 sg13g2_tiehi _20375__798 (.L_HI(net798));
 sg13g2_tiehi _20374__799 (.L_HI(net799));
 sg13g2_tiehi _20373__800 (.L_HI(net800));
 sg13g2_tiehi _20372__801 (.L_HI(net801));
 sg13g2_tiehi _20371__802 (.L_HI(net802));
 sg13g2_tiehi _20370__803 (.L_HI(net803));
 sg13g2_tiehi _20369__804 (.L_HI(net804));
 sg13g2_tiehi _20368__805 (.L_HI(net805));
 sg13g2_tiehi _20367__806 (.L_HI(net806));
 sg13g2_tiehi _20366__807 (.L_HI(net807));
 sg13g2_tiehi _20365__808 (.L_HI(net808));
 sg13g2_tiehi _20364__809 (.L_HI(net809));
 sg13g2_tiehi _20363__810 (.L_HI(net810));
 sg13g2_tiehi _20362__811 (.L_HI(net811));
 sg13g2_tiehi _20361__812 (.L_HI(net812));
 sg13g2_tiehi _20360__813 (.L_HI(net813));
 sg13g2_tiehi _20359__814 (.L_HI(net814));
 sg13g2_tiehi _20358__815 (.L_HI(net815));
 sg13g2_tiehi _20357__816 (.L_HI(net816));
 sg13g2_tiehi _20356__817 (.L_HI(net817));
 sg13g2_tiehi _20355__818 (.L_HI(net818));
 sg13g2_tiehi _20354__819 (.L_HI(net819));
 sg13g2_tiehi _20353__820 (.L_HI(net820));
 sg13g2_tiehi _20352__821 (.L_HI(net821));
 sg13g2_tiehi _20351__822 (.L_HI(net822));
 sg13g2_tiehi _20350__823 (.L_HI(net823));
 sg13g2_tiehi _20349__824 (.L_HI(net824));
 sg13g2_tiehi _20348__825 (.L_HI(net825));
 sg13g2_tiehi _20347__826 (.L_HI(net826));
 sg13g2_tiehi _20346__827 (.L_HI(net827));
 sg13g2_tiehi _20345__828 (.L_HI(net828));
 sg13g2_tiehi _20344__829 (.L_HI(net829));
 sg13g2_tiehi _20343__830 (.L_HI(net830));
 sg13g2_tiehi _20342__831 (.L_HI(net831));
 sg13g2_tiehi _20341__832 (.L_HI(net832));
 sg13g2_tiehi _20340__833 (.L_HI(net833));
 sg13g2_tiehi _20339__834 (.L_HI(net834));
 sg13g2_tiehi _20338__835 (.L_HI(net835));
 sg13g2_tiehi _20337__836 (.L_HI(net836));
 sg13g2_tiehi _20336__837 (.L_HI(net837));
 sg13g2_tiehi _20335__838 (.L_HI(net838));
 sg13g2_tiehi _20334__839 (.L_HI(net839));
 sg13g2_tiehi _20333__840 (.L_HI(net840));
 sg13g2_tiehi _20332__841 (.L_HI(net841));
 sg13g2_tiehi _20331__842 (.L_HI(net842));
 sg13g2_tiehi _20330__843 (.L_HI(net843));
 sg13g2_tiehi _20329__844 (.L_HI(net844));
 sg13g2_tiehi _20328__845 (.L_HI(net845));
 sg13g2_tiehi _20327__846 (.L_HI(net846));
 sg13g2_tiehi _20326__847 (.L_HI(net847));
 sg13g2_tiehi _20325__848 (.L_HI(net848));
 sg13g2_tiehi _20324__849 (.L_HI(net849));
 sg13g2_tiehi _20323__850 (.L_HI(net850));
 sg13g2_tiehi _20322__851 (.L_HI(net851));
 sg13g2_tiehi _20321__852 (.L_HI(net852));
 sg13g2_tiehi _20320__853 (.L_HI(net853));
 sg13g2_tiehi _20319__854 (.L_HI(net854));
 sg13g2_tiehi _20318__855 (.L_HI(net855));
 sg13g2_tiehi _20317__856 (.L_HI(net856));
 sg13g2_tiehi _20316__857 (.L_HI(net857));
 sg13g2_tiehi _20315__858 (.L_HI(net858));
 sg13g2_tiehi _20314__859 (.L_HI(net859));
 sg13g2_tiehi _20313__860 (.L_HI(net860));
 sg13g2_tiehi _20312__861 (.L_HI(net861));
 sg13g2_tiehi _20311__862 (.L_HI(net862));
 sg13g2_tiehi _20310__863 (.L_HI(net863));
 sg13g2_tiehi _20309__864 (.L_HI(net864));
 sg13g2_tiehi _20308__865 (.L_HI(net865));
 sg13g2_tiehi _20307__866 (.L_HI(net866));
 sg13g2_tiehi _20306__867 (.L_HI(net867));
 sg13g2_tiehi _20305__868 (.L_HI(net868));
 sg13g2_tiehi _20304__869 (.L_HI(net869));
 sg13g2_tiehi _20303__870 (.L_HI(net870));
 sg13g2_tiehi _20302__871 (.L_HI(net871));
 sg13g2_tiehi _20301__872 (.L_HI(net872));
 sg13g2_tiehi _20300__873 (.L_HI(net873));
 sg13g2_tiehi _20299__874 (.L_HI(net874));
 sg13g2_tiehi _20298__875 (.L_HI(net875));
 sg13g2_tiehi _20297__876 (.L_HI(net876));
 sg13g2_tiehi _20296__877 (.L_HI(net877));
 sg13g2_tiehi _20295__878 (.L_HI(net878));
 sg13g2_tiehi _20294__879 (.L_HI(net879));
 sg13g2_tiehi _20293__880 (.L_HI(net880));
 sg13g2_tiehi _20292__881 (.L_HI(net881));
 sg13g2_tiehi _20291__882 (.L_HI(net882));
 sg13g2_tiehi _20290__883 (.L_HI(net883));
 sg13g2_tiehi _20289__884 (.L_HI(net884));
 sg13g2_tiehi _20288__885 (.L_HI(net885));
 sg13g2_tiehi _20287__886 (.L_HI(net886));
 sg13g2_tiehi _20286__887 (.L_HI(net887));
 sg13g2_tiehi _20285__888 (.L_HI(net888));
 sg13g2_tiehi _20284__889 (.L_HI(net889));
 sg13g2_tiehi _20283__890 (.L_HI(net890));
 sg13g2_tiehi _20282__891 (.L_HI(net891));
 sg13g2_tiehi _20281__892 (.L_HI(net892));
 sg13g2_tiehi _20280__893 (.L_HI(net893));
 sg13g2_tiehi _20279__894 (.L_HI(net894));
 sg13g2_tiehi _20278__895 (.L_HI(net895));
 sg13g2_tiehi _20277__896 (.L_HI(net896));
 sg13g2_tiehi _20276__897 (.L_HI(net897));
 sg13g2_tiehi _20275__898 (.L_HI(net898));
 sg13g2_tiehi _20274__899 (.L_HI(net899));
 sg13g2_tiehi _20273__900 (.L_HI(net900));
 sg13g2_tiehi _20272__901 (.L_HI(net901));
 sg13g2_tiehi _20271__902 (.L_HI(net902));
 sg13g2_tiehi _20270__903 (.L_HI(net903));
 sg13g2_tiehi _19873__904 (.L_HI(net904));
 sg13g2_tiehi _20269__905 (.L_HI(net905));
 sg13g2_tiehi _20268__906 (.L_HI(net906));
 sg13g2_tiehi _20267__907 (.L_HI(net907));
 sg13g2_tiehi _20266__908 (.L_HI(net908));
 sg13g2_tiehi _20265__909 (.L_HI(net909));
 sg13g2_tiehi _20264__910 (.L_HI(net910));
 sg13g2_tiehi _20263__911 (.L_HI(net911));
 sg13g2_tiehi _20262__912 (.L_HI(net912));
 sg13g2_tiehi _20261__913 (.L_HI(net913));
 sg13g2_tiehi _20260__914 (.L_HI(net914));
 sg13g2_tiehi _20259__915 (.L_HI(net915));
 sg13g2_tiehi _20258__916 (.L_HI(net916));
 sg13g2_tiehi _20257__917 (.L_HI(net917));
 sg13g2_tiehi _20256__918 (.L_HI(net918));
 sg13g2_tiehi _20255__919 (.L_HI(net919));
 sg13g2_tiehi _20254__920 (.L_HI(net920));
 sg13g2_tiehi _20253__921 (.L_HI(net921));
 sg13g2_tiehi _20252__922 (.L_HI(net922));
 sg13g2_tiehi _20251__923 (.L_HI(net923));
 sg13g2_tiehi _20250__924 (.L_HI(net924));
 sg13g2_tiehi _20249__925 (.L_HI(net925));
 sg13g2_tiehi _20248__926 (.L_HI(net926));
 sg13g2_tiehi _20247__927 (.L_HI(net927));
 sg13g2_tiehi _20246__928 (.L_HI(net928));
 sg13g2_tiehi _20245__929 (.L_HI(net929));
 sg13g2_tiehi _20244__930 (.L_HI(net930));
 sg13g2_tiehi _20243__931 (.L_HI(net931));
 sg13g2_tiehi _20242__932 (.L_HI(net932));
 sg13g2_tiehi _20241__933 (.L_HI(net933));
 sg13g2_tiehi _20240__934 (.L_HI(net934));
 sg13g2_tiehi _20795__935 (.L_HI(net935));
 sg13g2_tiehi _20239__936 (.L_HI(net936));
 sg13g2_tiehi _20238__937 (.L_HI(net937));
 sg13g2_tiehi _20237__938 (.L_HI(net938));
 sg13g2_tiehi _20236__939 (.L_HI(net939));
 sg13g2_tiehi _20235__940 (.L_HI(net940));
 sg13g2_tiehi _20234__941 (.L_HI(net941));
 sg13g2_tiehi _20233__942 (.L_HI(net942));
 sg13g2_tiehi _20232__943 (.L_HI(net943));
 sg13g2_tiehi _20231__944 (.L_HI(net944));
 sg13g2_tiehi _20230__945 (.L_HI(net945));
 sg13g2_tiehi _20229__946 (.L_HI(net946));
 sg13g2_tiehi _20228__947 (.L_HI(net947));
 sg13g2_tiehi _20227__948 (.L_HI(net948));
 sg13g2_tiehi _20226__949 (.L_HI(net949));
 sg13g2_tiehi _20225__950 (.L_HI(net950));
 sg13g2_tiehi _20224__951 (.L_HI(net951));
 sg13g2_tiehi _20223__952 (.L_HI(net952));
 sg13g2_tiehi _20222__953 (.L_HI(net953));
 sg13g2_tiehi _20221__954 (.L_HI(net954));
 sg13g2_tiehi _20220__955 (.L_HI(net955));
 sg13g2_tiehi _20219__956 (.L_HI(net956));
 sg13g2_tiehi _20218__957 (.L_HI(net957));
 sg13g2_tiehi _20217__958 (.L_HI(net958));
 sg13g2_tiehi _20216__959 (.L_HI(net959));
 sg13g2_tiehi _20215__960 (.L_HI(net960));
 sg13g2_tiehi _20214__961 (.L_HI(net961));
 sg13g2_tiehi _20213__962 (.L_HI(net962));
 sg13g2_tiehi _20212__963 (.L_HI(net963));
 sg13g2_tiehi _20211__964 (.L_HI(net964));
 sg13g2_tiehi _20210__965 (.L_HI(net965));
 sg13g2_tiehi _20209__966 (.L_HI(net966));
 sg13g2_tiehi _20208__967 (.L_HI(net967));
 sg13g2_tiehi _20207__968 (.L_HI(net968));
 sg13g2_tiehi _20206__969 (.L_HI(net969));
 sg13g2_tiehi _20205__970 (.L_HI(net970));
 sg13g2_tiehi _20204__971 (.L_HI(net971));
 sg13g2_tiehi _20203__972 (.L_HI(net972));
 sg13g2_tiehi _20202__973 (.L_HI(net973));
 sg13g2_tiehi _20201__974 (.L_HI(net974));
 sg13g2_tiehi _20200__975 (.L_HI(net975));
 sg13g2_tiehi _20199__976 (.L_HI(net976));
 sg13g2_tiehi _20198__977 (.L_HI(net977));
 sg13g2_tiehi _20197__978 (.L_HI(net978));
 sg13g2_tiehi _20196__979 (.L_HI(net979));
 sg13g2_tiehi _20195__980 (.L_HI(net980));
 sg13g2_tiehi _20194__981 (.L_HI(net981));
 sg13g2_tiehi _20193__982 (.L_HI(net982));
 sg13g2_tiehi _20192__983 (.L_HI(net983));
 sg13g2_tiehi _20191__984 (.L_HI(net984));
 sg13g2_tiehi _20190__985 (.L_HI(net985));
 sg13g2_tiehi _20189__986 (.L_HI(net986));
 sg13g2_tiehi _20188__987 (.L_HI(net987));
 sg13g2_tiehi _20187__988 (.L_HI(net988));
 sg13g2_tiehi _20186__989 (.L_HI(net989));
 sg13g2_tiehi _20185__990 (.L_HI(net990));
 sg13g2_tiehi _20184__991 (.L_HI(net991));
 sg13g2_tiehi _20183__992 (.L_HI(net992));
 sg13g2_tiehi _20182__993 (.L_HI(net993));
 sg13g2_tiehi _20181__994 (.L_HI(net994));
 sg13g2_tiehi _20180__995 (.L_HI(net995));
 sg13g2_tiehi _20179__996 (.L_HI(net996));
 sg13g2_tiehi _20178__997 (.L_HI(net997));
 sg13g2_tiehi _20177__998 (.L_HI(net998));
 sg13g2_tiehi _20176__999 (.L_HI(net999));
 sg13g2_tiehi _20175__1000 (.L_HI(net1000));
 sg13g2_tiehi _20174__1001 (.L_HI(net1001));
 sg13g2_tiehi _20173__1002 (.L_HI(net1002));
 sg13g2_tiehi _20172__1003 (.L_HI(net1003));
 sg13g2_tiehi _20171__1004 (.L_HI(net1004));
 sg13g2_tiehi _20170__1005 (.L_HI(net1005));
 sg13g2_tiehi _20169__1006 (.L_HI(net1006));
 sg13g2_tiehi _20168__1007 (.L_HI(net1007));
 sg13g2_tiehi _20167__1008 (.L_HI(net1008));
 sg13g2_tiehi _20166__1009 (.L_HI(net1009));
 sg13g2_tiehi _20165__1010 (.L_HI(net1010));
 sg13g2_tiehi _20164__1011 (.L_HI(net1011));
 sg13g2_tiehi _20163__1012 (.L_HI(net1012));
 sg13g2_tiehi _20162__1013 (.L_HI(net1013));
 sg13g2_tiehi _20161__1014 (.L_HI(net1014));
 sg13g2_tiehi _20160__1015 (.L_HI(net1015));
 sg13g2_tiehi _20159__1016 (.L_HI(net1016));
 sg13g2_tiehi _20158__1017 (.L_HI(net1017));
 sg13g2_tiehi _20157__1018 (.L_HI(net1018));
 sg13g2_tiehi _20156__1019 (.L_HI(net1019));
 sg13g2_tiehi _20155__1020 (.L_HI(net1020));
 sg13g2_tiehi _20154__1021 (.L_HI(net1021));
 sg13g2_tiehi _20153__1022 (.L_HI(net1022));
 sg13g2_tiehi _20152__1023 (.L_HI(net1023));
 sg13g2_tiehi _20151__1024 (.L_HI(net1024));
 sg13g2_tiehi _20150__1025 (.L_HI(net1025));
 sg13g2_tiehi _20149__1026 (.L_HI(net1026));
 sg13g2_tiehi _20148__1027 (.L_HI(net1027));
 sg13g2_tiehi _20147__1028 (.L_HI(net1028));
 sg13g2_tiehi _20146__1029 (.L_HI(net1029));
 sg13g2_tiehi _20145__1030 (.L_HI(net1030));
 sg13g2_tiehi _20144__1031 (.L_HI(net1031));
 sg13g2_tiehi _20143__1032 (.L_HI(net1032));
 sg13g2_tiehi _20142__1033 (.L_HI(net1033));
 sg13g2_tiehi _20141__1034 (.L_HI(net1034));
 sg13g2_tiehi _20140__1035 (.L_HI(net1035));
 sg13g2_tiehi _20139__1036 (.L_HI(net1036));
 sg13g2_tiehi _20138__1037 (.L_HI(net1037));
 sg13g2_tiehi _20137__1038 (.L_HI(net1038));
 sg13g2_tiehi _20136__1039 (.L_HI(net1039));
 sg13g2_tiehi _20135__1040 (.L_HI(net1040));
 sg13g2_tiehi _20134__1041 (.L_HI(net1041));
 sg13g2_tiehi _20133__1042 (.L_HI(net1042));
 sg13g2_tiehi _20132__1043 (.L_HI(net1043));
 sg13g2_tiehi _20131__1044 (.L_HI(net1044));
 sg13g2_tiehi _20130__1045 (.L_HI(net1045));
 sg13g2_tiehi _20129__1046 (.L_HI(net1046));
 sg13g2_tiehi _20128__1047 (.L_HI(net1047));
 sg13g2_tiehi _20127__1048 (.L_HI(net1048));
 sg13g2_tiehi _20126__1049 (.L_HI(net1049));
 sg13g2_tiehi _20840__1050 (.L_HI(net1050));
 sg13g2_tiehi _20125__1051 (.L_HI(net1051));
 sg13g2_tiehi _20124__1052 (.L_HI(net1052));
 sg13g2_tiehi _20123__1053 (.L_HI(net1053));
 sg13g2_tiehi _20122__1054 (.L_HI(net1054));
 sg13g2_tiehi _20121__1055 (.L_HI(net1055));
 sg13g2_tiehi _20120__1056 (.L_HI(net1056));
 sg13g2_tiehi _20119__1057 (.L_HI(net1057));
 sg13g2_tiehi _20118__1058 (.L_HI(net1058));
 sg13g2_tiehi _20117__1059 (.L_HI(net1059));
 sg13g2_tiehi _20116__1060 (.L_HI(net1060));
 sg13g2_tiehi _20115__1061 (.L_HI(net1061));
 sg13g2_tiehi _20114__1062 (.L_HI(net1062));
 sg13g2_tiehi _20972__1063 (.L_HI(net1063));
 sg13g2_tiehi _20113__1064 (.L_HI(net1064));
 sg13g2_tiehi _20112__1065 (.L_HI(net1065));
 sg13g2_tiehi _20111__1066 (.L_HI(net1066));
 sg13g2_tiehi _20110__1067 (.L_HI(net1067));
 sg13g2_tiehi _20109__1068 (.L_HI(net1068));
 sg13g2_tiehi _20108__1069 (.L_HI(net1069));
 sg13g2_tiehi _20107__1070 (.L_HI(net1070));
 sg13g2_tiehi _20106__1071 (.L_HI(net1071));
 sg13g2_tiehi _20105__1072 (.L_HI(net1072));
 sg13g2_tiehi _20104__1073 (.L_HI(net1073));
 sg13g2_tiehi _20103__1074 (.L_HI(net1074));
 sg13g2_tiehi _20102__1075 (.L_HI(net1075));
 sg13g2_tiehi _20101__1076 (.L_HI(net1076));
 sg13g2_tiehi _20100__1077 (.L_HI(net1077));
 sg13g2_tiehi _20099__1078 (.L_HI(net1078));
 sg13g2_tiehi _20098__1079 (.L_HI(net1079));
 sg13g2_tiehi _20097__1080 (.L_HI(net1080));
 sg13g2_tiehi _20096__1081 (.L_HI(net1081));
 sg13g2_tiehi _20095__1082 (.L_HI(net1082));
 sg13g2_tiehi _20094__1083 (.L_HI(net1083));
 sg13g2_tiehi _20093__1084 (.L_HI(net1084));
 sg13g2_tiehi _20092__1085 (.L_HI(net1085));
 sg13g2_tiehi _20091__1086 (.L_HI(net1086));
 sg13g2_tiehi _20090__1087 (.L_HI(net1087));
 sg13g2_tiehi _20089__1088 (.L_HI(net1088));
 sg13g2_tiehi _20088__1089 (.L_HI(net1089));
 sg13g2_tiehi _20087__1090 (.L_HI(net1090));
 sg13g2_tiehi _20086__1091 (.L_HI(net1091));
 sg13g2_tiehi _20085__1092 (.L_HI(net1092));
 sg13g2_tiehi _20084__1093 (.L_HI(net1093));
 sg13g2_tiehi _20083__1094 (.L_HI(net1094));
 sg13g2_tiehi _20082__1095 (.L_HI(net1095));
 sg13g2_tiehi _20081__1096 (.L_HI(net1096));
 sg13g2_tiehi _20080__1097 (.L_HI(net1097));
 sg13g2_tiehi _20079__1098 (.L_HI(net1098));
 sg13g2_tiehi _20078__1099 (.L_HI(net1099));
 sg13g2_tiehi _20077__1100 (.L_HI(net1100));
 sg13g2_tiehi _20076__1101 (.L_HI(net1101));
 sg13g2_tiehi _20075__1102 (.L_HI(net1102));
 sg13g2_tiehi _20074__1103 (.L_HI(net1103));
 sg13g2_tiehi _20073__1104 (.L_HI(net1104));
 sg13g2_tiehi _20072__1105 (.L_HI(net1105));
 sg13g2_tiehi _20071__1106 (.L_HI(net1106));
 sg13g2_tiehi _20070__1107 (.L_HI(net1107));
 sg13g2_tiehi _20069__1108 (.L_HI(net1108));
 sg13g2_tiehi _20068__1109 (.L_HI(net1109));
 sg13g2_tiehi _20067__1110 (.L_HI(net1110));
 sg13g2_tiehi _20066__1111 (.L_HI(net1111));
 sg13g2_tiehi _20065__1112 (.L_HI(net1112));
 sg13g2_tiehi _20064__1113 (.L_HI(net1113));
 sg13g2_tiehi _20063__1114 (.L_HI(net1114));
 sg13g2_tiehi _20062__1115 (.L_HI(net1115));
 sg13g2_tiehi _20061__1116 (.L_HI(net1116));
 sg13g2_tiehi _20060__1117 (.L_HI(net1117));
 sg13g2_tiehi _20059__1118 (.L_HI(net1118));
 sg13g2_tiehi _20058__1119 (.L_HI(net1119));
 sg13g2_tiehi _20057__1120 (.L_HI(net1120));
 sg13g2_tiehi _20056__1121 (.L_HI(net1121));
 sg13g2_tiehi _20055__1122 (.L_HI(net1122));
 sg13g2_tiehi _20054__1123 (.L_HI(net1123));
 sg13g2_tiehi _20053__1124 (.L_HI(net1124));
 sg13g2_tiehi _20052__1125 (.L_HI(net1125));
 sg13g2_tiehi _20051__1126 (.L_HI(net1126));
 sg13g2_tiehi _20050__1127 (.L_HI(net1127));
 sg13g2_tiehi _20049__1128 (.L_HI(net1128));
 sg13g2_tiehi _20048__1129 (.L_HI(net1129));
 sg13g2_tiehi _20047__1130 (.L_HI(net1130));
 sg13g2_tiehi _20046__1131 (.L_HI(net1131));
 sg13g2_tiehi _20045__1132 (.L_HI(net1132));
 sg13g2_tiehi _20044__1133 (.L_HI(net1133));
 sg13g2_tiehi _20043__1134 (.L_HI(net1134));
 sg13g2_tiehi _20042__1135 (.L_HI(net1135));
 sg13g2_tiehi _20041__1136 (.L_HI(net1136));
 sg13g2_tiehi _20040__1137 (.L_HI(net1137));
 sg13g2_tiehi _20039__1138 (.L_HI(net1138));
 sg13g2_tiehi _20038__1139 (.L_HI(net1139));
 sg13g2_tiehi _20037__1140 (.L_HI(net1140));
 sg13g2_tiehi _20036__1141 (.L_HI(net1141));
 sg13g2_tiehi _20035__1142 (.L_HI(net1142));
 sg13g2_tiehi _20034__1143 (.L_HI(net1143));
 sg13g2_tiehi _20033__1144 (.L_HI(net1144));
 sg13g2_tiehi _20032__1145 (.L_HI(net1145));
 sg13g2_tiehi _20031__1146 (.L_HI(net1146));
 sg13g2_tiehi _20030__1147 (.L_HI(net1147));
 sg13g2_tiehi _20029__1148 (.L_HI(net1148));
 sg13g2_tiehi _20028__1149 (.L_HI(net1149));
 sg13g2_tiehi _20027__1150 (.L_HI(net1150));
 sg13g2_tiehi _20026__1151 (.L_HI(net1151));
 sg13g2_tiehi _20025__1152 (.L_HI(net1152));
 sg13g2_tiehi _20024__1153 (.L_HI(net1153));
 sg13g2_tiehi _20023__1154 (.L_HI(net1154));
 sg13g2_tiehi _20022__1155 (.L_HI(net1155));
 sg13g2_tiehi _20021__1156 (.L_HI(net1156));
 sg13g2_tiehi _20020__1157 (.L_HI(net1157));
 sg13g2_tiehi _20019__1158 (.L_HI(net1158));
 sg13g2_tiehi _20018__1159 (.L_HI(net1159));
 sg13g2_tiehi _20017__1160 (.L_HI(net1160));
 sg13g2_tiehi _20016__1161 (.L_HI(net1161));
 sg13g2_tiehi _20015__1162 (.L_HI(net1162));
 sg13g2_tiehi _20014__1163 (.L_HI(net1163));
 sg13g2_tiehi _20013__1164 (.L_HI(net1164));
 sg13g2_tiehi _20012__1165 (.L_HI(net1165));
 sg13g2_tiehi _20011__1166 (.L_HI(net1166));
 sg13g2_tiehi _20010__1167 (.L_HI(net1167));
 sg13g2_tiehi _20009__1168 (.L_HI(net1168));
 sg13g2_tiehi _20008__1169 (.L_HI(net1169));
 sg13g2_tiehi _20007__1170 (.L_HI(net1170));
 sg13g2_tiehi _20006__1171 (.L_HI(net1171));
 sg13g2_tiehi _20005__1172 (.L_HI(net1172));
 sg13g2_tiehi _20004__1173 (.L_HI(net1173));
 sg13g2_tiehi _20003__1174 (.L_HI(net1174));
 sg13g2_tiehi _20002__1175 (.L_HI(net1175));
 sg13g2_tiehi _20001__1176 (.L_HI(net1176));
 sg13g2_tiehi _20000__1177 (.L_HI(net1177));
 sg13g2_tiehi _19999__1178 (.L_HI(net1178));
 sg13g2_tiehi _19998__1179 (.L_HI(net1179));
 sg13g2_tiehi _19997__1180 (.L_HI(net1180));
 sg13g2_tiehi _19996__1181 (.L_HI(net1181));
 sg13g2_tiehi _19995__1182 (.L_HI(net1182));
 sg13g2_tiehi _19994__1183 (.L_HI(net1183));
 sg13g2_tiehi _19993__1184 (.L_HI(net1184));
 sg13g2_tiehi _19992__1185 (.L_HI(net1185));
 sg13g2_tiehi _19991__1186 (.L_HI(net1186));
 sg13g2_tiehi _19990__1187 (.L_HI(net1187));
 sg13g2_tiehi _19989__1188 (.L_HI(net1188));
 sg13g2_tiehi _19988__1189 (.L_HI(net1189));
 sg13g2_tiehi _19987__1190 (.L_HI(net1190));
 sg13g2_tiehi _19986__1191 (.L_HI(net1191));
 sg13g2_tiehi _19985__1192 (.L_HI(net1192));
 sg13g2_tiehi _19984__1193 (.L_HI(net1193));
 sg13g2_tiehi _19983__1194 (.L_HI(net1194));
 sg13g2_tiehi _19982__1195 (.L_HI(net1195));
 sg13g2_tiehi _19981__1196 (.L_HI(net1196));
 sg13g2_tiehi _19980__1197 (.L_HI(net1197));
 sg13g2_tiehi _19979__1198 (.L_HI(net1198));
 sg13g2_tiehi _19978__1199 (.L_HI(net1199));
 sg13g2_tiehi _19977__1200 (.L_HI(net1200));
 sg13g2_tiehi _19976__1201 (.L_HI(net1201));
 sg13g2_tiehi _19975__1202 (.L_HI(net1202));
 sg13g2_tiehi _19974__1203 (.L_HI(net1203));
 sg13g2_tiehi _19973__1204 (.L_HI(net1204));
 sg13g2_tiehi _19972__1205 (.L_HI(net1205));
 sg13g2_tiehi _19971__1206 (.L_HI(net1206));
 sg13g2_tiehi _19970__1207 (.L_HI(net1207));
 sg13g2_tiehi _19969__1208 (.L_HI(net1208));
 sg13g2_tiehi _19968__1209 (.L_HI(net1209));
 sg13g2_tiehi _19967__1210 (.L_HI(net1210));
 sg13g2_tiehi _19966__1211 (.L_HI(net1211));
 sg13g2_tiehi _19965__1212 (.L_HI(net1212));
 sg13g2_tiehi _19964__1213 (.L_HI(net1213));
 sg13g2_tiehi _19963__1214 (.L_HI(net1214));
 sg13g2_tiehi _19962__1215 (.L_HI(net1215));
 sg13g2_tiehi _19961__1216 (.L_HI(net1216));
 sg13g2_tiehi _19960__1217 (.L_HI(net1217));
 sg13g2_tiehi _19959__1218 (.L_HI(net1218));
 sg13g2_tiehi _19958__1219 (.L_HI(net1219));
 sg13g2_tiehi _19957__1220 (.L_HI(net1220));
 sg13g2_tiehi _19956__1221 (.L_HI(net1221));
 sg13g2_tiehi _19955__1222 (.L_HI(net1222));
 sg13g2_tiehi _19954__1223 (.L_HI(net1223));
 sg13g2_tiehi _19953__1224 (.L_HI(net1224));
 sg13g2_tiehi _19952__1225 (.L_HI(net1225));
 sg13g2_tiehi _19951__1226 (.L_HI(net1226));
 sg13g2_tiehi _19950__1227 (.L_HI(net1227));
 sg13g2_tiehi _19949__1228 (.L_HI(net1228));
 sg13g2_tiehi _19948__1229 (.L_HI(net1229));
 sg13g2_tiehi _19947__1230 (.L_HI(net1230));
 sg13g2_tiehi _19946__1231 (.L_HI(net1231));
 sg13g2_tiehi _19945__1232 (.L_HI(net1232));
 sg13g2_tiehi _19944__1233 (.L_HI(net1233));
 sg13g2_tiehi _19943__1234 (.L_HI(net1234));
 sg13g2_tiehi _19942__1235 (.L_HI(net1235));
 sg13g2_tiehi _19941__1236 (.L_HI(net1236));
 sg13g2_tiehi _19940__1237 (.L_HI(net1237));
 sg13g2_tiehi _19939__1238 (.L_HI(net1238));
 sg13g2_tiehi _21226__1239 (.L_HI(net1239));
 sg13g2_tiehi _19938__1240 (.L_HI(net1240));
 sg13g2_tiehi _19937__1241 (.L_HI(net1241));
 sg13g2_tiehi _19936__1242 (.L_HI(net1242));
 sg13g2_tiehi _19935__1243 (.L_HI(net1243));
 sg13g2_tiehi _19934__1244 (.L_HI(net1244));
 sg13g2_tiehi _19933__1245 (.L_HI(net1245));
 sg13g2_tiehi _19932__1246 (.L_HI(net1246));
 sg13g2_tiehi _19931__1247 (.L_HI(net1247));
 sg13g2_tiehi _19930__1248 (.L_HI(net1248));
 sg13g2_tiehi _19929__1249 (.L_HI(net1249));
 sg13g2_tiehi _19928__1250 (.L_HI(net1250));
 sg13g2_tiehi _19927__1251 (.L_HI(net1251));
 sg13g2_tiehi _19926__1252 (.L_HI(net1252));
 sg13g2_tiehi _19925__1253 (.L_HI(net1253));
 sg13g2_tiehi _19924__1254 (.L_HI(net1254));
 sg13g2_tiehi _19923__1255 (.L_HI(net1255));
 sg13g2_tiehi _19922__1256 (.L_HI(net1256));
 sg13g2_tiehi _19921__1257 (.L_HI(net1257));
 sg13g2_tiehi _19920__1258 (.L_HI(net1258));
 sg13g2_tiehi _19919__1259 (.L_HI(net1259));
 sg13g2_tiehi _19918__1260 (.L_HI(net1260));
 sg13g2_tiehi _19917__1261 (.L_HI(net1261));
 sg13g2_tiehi _19916__1262 (.L_HI(net1262));
 sg13g2_tiehi _19915__1263 (.L_HI(net1263));
 sg13g2_tiehi _19914__1264 (.L_HI(net1264));
 sg13g2_tiehi _19913__1265 (.L_HI(net1265));
 sg13g2_tiehi _19912__1266 (.L_HI(net1266));
 sg13g2_tiehi _19911__1267 (.L_HI(net1267));
 sg13g2_tiehi _19910__1268 (.L_HI(net1268));
 sg13g2_tiehi _19909__1269 (.L_HI(net1269));
 sg13g2_tiehi _19908__1270 (.L_HI(net1270));
 sg13g2_tiehi _19907__1271 (.L_HI(net1271));
 sg13g2_tiehi _19906__1272 (.L_HI(net1272));
 sg13g2_tiehi _19905__1273 (.L_HI(net1273));
 sg13g2_tiehi _19904__1274 (.L_HI(net1274));
 sg13g2_tiehi _19903__1275 (.L_HI(net1275));
 sg13g2_tiehi _19902__1276 (.L_HI(net1276));
 sg13g2_tiehi _19901__1277 (.L_HI(net1277));
 sg13g2_tiehi _19900__1278 (.L_HI(net1278));
 sg13g2_tiehi _19899__1279 (.L_HI(net1279));
 sg13g2_tiehi _19898__1280 (.L_HI(net1280));
 sg13g2_tiehi _19897__1281 (.L_HI(net1281));
 sg13g2_tiehi _19896__1282 (.L_HI(net1282));
 sg13g2_tiehi _19895__1283 (.L_HI(net1283));
 sg13g2_tiehi _19894__1284 (.L_HI(net1284));
 sg13g2_tiehi _19893__1285 (.L_HI(net1285));
 sg13g2_tiehi _19892__1286 (.L_HI(net1286));
 sg13g2_tiehi _19891__1287 (.L_HI(net1287));
 sg13g2_tiehi _19890__1288 (.L_HI(net1288));
 sg13g2_tiehi _19889__1289 (.L_HI(net1289));
 sg13g2_tiehi _19888__1290 (.L_HI(net1290));
 sg13g2_tiehi _19887__1291 (.L_HI(net1291));
 sg13g2_tiehi _19886__1292 (.L_HI(net1292));
 sg13g2_tiehi _19885__1293 (.L_HI(net1293));
 sg13g2_tiehi _19884__1294 (.L_HI(net1294));
 sg13g2_tiehi _19883__1295 (.L_HI(net1295));
 sg13g2_tiehi _19882__1296 (.L_HI(net1296));
 sg13g2_tiehi _19881__1297 (.L_HI(net1297));
 sg13g2_tiehi _19880__1298 (.L_HI(net1298));
 sg13g2_tiehi _19879__1299 (.L_HI(net1299));
 sg13g2_tiehi _19878__1300 (.L_HI(net1300));
 sg13g2_tiehi _19877__1301 (.L_HI(net1301));
 sg13g2_tiehi _19876__1302 (.L_HI(net1302));
 sg13g2_tiehi _19875__1303 (.L_HI(net1303));
 sg13g2_tiehi _19874__1304 (.L_HI(net1304));
 sg13g2_tiehi _22430__1305 (.L_HI(net1305));
 sg13g2_tiehi _22429__1306 (.L_HI(net1306));
 sg13g2_tiehi _22428__1307 (.L_HI(net1307));
 sg13g2_tiehi _22427__1308 (.L_HI(net1308));
 sg13g2_tiehi _22426__1309 (.L_HI(net1309));
 sg13g2_tiehi _22425__1310 (.L_HI(net1310));
 sg13g2_tiehi _22424__1311 (.L_HI(net1311));
 sg13g2_tiehi _22423__1312 (.L_HI(net1312));
 sg13g2_tiehi _22422__1313 (.L_HI(net1313));
 sg13g2_tiehi _22421__1314 (.L_HI(net1314));
 sg13g2_tiehi _22420__1315 (.L_HI(net1315));
 sg13g2_tiehi _22419__1316 (.L_HI(net1316));
 sg13g2_tiehi _22418__1317 (.L_HI(net1317));
 sg13g2_tiehi _22417__1318 (.L_HI(net1318));
 sg13g2_tiehi _22416__1319 (.L_HI(net1319));
 sg13g2_tiehi _22415__1320 (.L_HI(net1320));
 sg13g2_tiehi _22414__1321 (.L_HI(net1321));
 sg13g2_tiehi _22413__1322 (.L_HI(net1322));
 sg13g2_tiehi _22412__1323 (.L_HI(net1323));
 sg13g2_tiehi _22411__1324 (.L_HI(net1324));
 sg13g2_tiehi _22410__1325 (.L_HI(net1325));
 sg13g2_tiehi _22409__1326 (.L_HI(net1326));
 sg13g2_tiehi _22408__1327 (.L_HI(net1327));
 sg13g2_tiehi _22407__1328 (.L_HI(net1328));
 sg13g2_tiehi _22406__1329 (.L_HI(net1329));
 sg13g2_tiehi _22405__1330 (.L_HI(net1330));
 sg13g2_tiehi _22404__1331 (.L_HI(net1331));
 sg13g2_tiehi _22403__1332 (.L_HI(net1332));
 sg13g2_tiehi _22402__1333 (.L_HI(net1333));
 sg13g2_tiehi _22401__1334 (.L_HI(net1334));
 sg13g2_tiehi _22400__1335 (.L_HI(net1335));
 sg13g2_tiehi _22399__1336 (.L_HI(net1336));
 sg13g2_tiehi _22398__1337 (.L_HI(net1337));
 sg13g2_tiehi _22397__1338 (.L_HI(net1338));
 sg13g2_tiehi _22396__1339 (.L_HI(net1339));
 sg13g2_tiehi _22395__1340 (.L_HI(net1340));
 sg13g2_tiehi _22394__1341 (.L_HI(net1341));
 sg13g2_tiehi _22393__1342 (.L_HI(net1342));
 sg13g2_tiehi _22392__1343 (.L_HI(net1343));
 sg13g2_tiehi _22391__1344 (.L_HI(net1344));
 sg13g2_tiehi _22390__1345 (.L_HI(net1345));
 sg13g2_tiehi _22389__1346 (.L_HI(net1346));
 sg13g2_tiehi _22388__1347 (.L_HI(net1347));
 sg13g2_tiehi _22387__1348 (.L_HI(net1348));
 sg13g2_tiehi _22386__1349 (.L_HI(net1349));
 sg13g2_tiehi _22385__1350 (.L_HI(net1350));
 sg13g2_tiehi _22384__1351 (.L_HI(net1351));
 sg13g2_tiehi _22383__1352 (.L_HI(net1352));
 sg13g2_tiehi _22382__1353 (.L_HI(net1353));
 sg13g2_tiehi _22381__1354 (.L_HI(net1354));
 sg13g2_tiehi _22380__1355 (.L_HI(net1355));
 sg13g2_tiehi _22379__1356 (.L_HI(net1356));
 sg13g2_tiehi _22378__1357 (.L_HI(net1357));
 sg13g2_tiehi _22377__1358 (.L_HI(net1358));
 sg13g2_tiehi _22376__1359 (.L_HI(net1359));
 sg13g2_tiehi _22375__1360 (.L_HI(net1360));
 sg13g2_tiehi _22374__1361 (.L_HI(net1361));
 sg13g2_tiehi _22373__1362 (.L_HI(net1362));
 sg13g2_tiehi _22372__1363 (.L_HI(net1363));
 sg13g2_tiehi _22371__1364 (.L_HI(net1364));
 sg13g2_tiehi _22370__1365 (.L_HI(net1365));
 sg13g2_tiehi _22369__1366 (.L_HI(net1366));
 sg13g2_tiehi _22368__1367 (.L_HI(net1367));
 sg13g2_tiehi _22367__1368 (.L_HI(net1368));
 sg13g2_tiehi _22366__1369 (.L_HI(net1369));
 sg13g2_tiehi _22365__1370 (.L_HI(net1370));
 sg13g2_tiehi _22364__1371 (.L_HI(net1371));
 sg13g2_tiehi _22363__1372 (.L_HI(net1372));
 sg13g2_tiehi _22362__1373 (.L_HI(net1373));
 sg13g2_tiehi _22361__1374 (.L_HI(net1374));
 sg13g2_tiehi _22360__1375 (.L_HI(net1375));
 sg13g2_tiehi _22359__1376 (.L_HI(net1376));
 sg13g2_tiehi _22358__1377 (.L_HI(net1377));
 sg13g2_tiehi _22357__1378 (.L_HI(net1378));
 sg13g2_tiehi _22356__1379 (.L_HI(net1379));
 sg13g2_tiehi _22355__1380 (.L_HI(net1380));
 sg13g2_tiehi _22354__1381 (.L_HI(net1381));
 sg13g2_tiehi _22353__1382 (.L_HI(net1382));
 sg13g2_tiehi _22352__1383 (.L_HI(net1383));
 sg13g2_tiehi _22351__1384 (.L_HI(net1384));
 sg13g2_tiehi _22350__1385 (.L_HI(net1385));
 sg13g2_tiehi _22349__1386 (.L_HI(net1386));
 sg13g2_tiehi _22348__1387 (.L_HI(net1387));
 sg13g2_tiehi _22347__1388 (.L_HI(net1388));
 sg13g2_tiehi _22346__1389 (.L_HI(net1389));
 sg13g2_tiehi _22345__1390 (.L_HI(net1390));
 sg13g2_tiehi _22344__1391 (.L_HI(net1391));
 sg13g2_tiehi _22343__1392 (.L_HI(net1392));
 sg13g2_tiehi _22342__1393 (.L_HI(net1393));
 sg13g2_tiehi _22341__1394 (.L_HI(net1394));
 sg13g2_tiehi _22340__1395 (.L_HI(net1395));
 sg13g2_tiehi _22339__1396 (.L_HI(net1396));
 sg13g2_tiehi _22338__1397 (.L_HI(net1397));
 sg13g2_tiehi _22337__1398 (.L_HI(net1398));
 sg13g2_tiehi _22336__1399 (.L_HI(net1399));
 sg13g2_tiehi _22335__1400 (.L_HI(net1400));
 sg13g2_tiehi _22334__1401 (.L_HI(net1401));
 sg13g2_tiehi _22333__1402 (.L_HI(net1402));
 sg13g2_tiehi _22332__1403 (.L_HI(net1403));
 sg13g2_tiehi _22331__1404 (.L_HI(net1404));
 sg13g2_tiehi _22330__1405 (.L_HI(net1405));
 sg13g2_tiehi _22329__1406 (.L_HI(net1406));
 sg13g2_tiehi _22328__1407 (.L_HI(net1407));
 sg13g2_tiehi _22327__1408 (.L_HI(net1408));
 sg13g2_tiehi _22326__1409 (.L_HI(net1409));
 sg13g2_tiehi _22325__1410 (.L_HI(net1410));
 sg13g2_tiehi _22324__1411 (.L_HI(net1411));
 sg13g2_tiehi _22323__1412 (.L_HI(net1412));
 sg13g2_tiehi _22322__1413 (.L_HI(net1413));
 sg13g2_tiehi _22321__1414 (.L_HI(net1414));
 sg13g2_tiehi _22320__1415 (.L_HI(net1415));
 sg13g2_tiehi _22319__1416 (.L_HI(net1416));
 sg13g2_tiehi _22318__1417 (.L_HI(net1417));
 sg13g2_tiehi _22317__1418 (.L_HI(net1418));
 sg13g2_tiehi _22316__1419 (.L_HI(net1419));
 sg13g2_tiehi _22315__1420 (.L_HI(net1420));
 sg13g2_tiehi _22314__1421 (.L_HI(net1421));
 sg13g2_tiehi _22313__1422 (.L_HI(net1422));
 sg13g2_tiehi _22312__1423 (.L_HI(net1423));
 sg13g2_tiehi _22311__1424 (.L_HI(net1424));
 sg13g2_tiehi _22310__1425 (.L_HI(net1425));
 sg13g2_tiehi _22309__1426 (.L_HI(net1426));
 sg13g2_tiehi _22308__1427 (.L_HI(net1427));
 sg13g2_tiehi _22307__1428 (.L_HI(net1428));
 sg13g2_tiehi _22306__1429 (.L_HI(net1429));
 sg13g2_tiehi _22305__1430 (.L_HI(net1430));
 sg13g2_tiehi _22304__1431 (.L_HI(net1431));
 sg13g2_tiehi _22303__1432 (.L_HI(net1432));
 sg13g2_tiehi _22302__1433 (.L_HI(net1433));
 sg13g2_tiehi _22301__1434 (.L_HI(net1434));
 sg13g2_tiehi _22300__1435 (.L_HI(net1435));
 sg13g2_tiehi _22299__1436 (.L_HI(net1436));
 sg13g2_tiehi _22298__1437 (.L_HI(net1437));
 sg13g2_tiehi _22297__1438 (.L_HI(net1438));
 sg13g2_tiehi _22296__1439 (.L_HI(net1439));
 sg13g2_tiehi _22295__1440 (.L_HI(net1440));
 sg13g2_tiehi _22294__1441 (.L_HI(net1441));
 sg13g2_tiehi _22293__1442 (.L_HI(net1442));
 sg13g2_tiehi _22292__1443 (.L_HI(net1443));
 sg13g2_tiehi _22291__1444 (.L_HI(net1444));
 sg13g2_tiehi _22290__1445 (.L_HI(net1445));
 sg13g2_tiehi _22289__1446 (.L_HI(net1446));
 sg13g2_tiehi _22288__1447 (.L_HI(net1447));
 sg13g2_tiehi _22287__1448 (.L_HI(net1448));
 sg13g2_tiehi _22286__1449 (.L_HI(net1449));
 sg13g2_tiehi _22285__1450 (.L_HI(net1450));
 sg13g2_tiehi _22284__1451 (.L_HI(net1451));
 sg13g2_tiehi _22283__1452 (.L_HI(net1452));
 sg13g2_tiehi _22282__1453 (.L_HI(net1453));
 sg13g2_tiehi _22281__1454 (.L_HI(net1454));
 sg13g2_tiehi _22280__1455 (.L_HI(net1455));
 sg13g2_tiehi _22279__1456 (.L_HI(net1456));
 sg13g2_tiehi _22278__1457 (.L_HI(net1457));
 sg13g2_tiehi _22277__1458 (.L_HI(net1458));
 sg13g2_tiehi _22276__1459 (.L_HI(net1459));
 sg13g2_tiehi _22275__1460 (.L_HI(net1460));
 sg13g2_tiehi _22274__1461 (.L_HI(net1461));
 sg13g2_tiehi _22273__1462 (.L_HI(net1462));
 sg13g2_tiehi _22272__1463 (.L_HI(net1463));
 sg13g2_tiehi _22271__1464 (.L_HI(net1464));
 sg13g2_tiehi _22270__1465 (.L_HI(net1465));
 sg13g2_tiehi _22269__1466 (.L_HI(net1466));
 sg13g2_tiehi _22268__1467 (.L_HI(net1467));
 sg13g2_tiehi _22267__1468 (.L_HI(net1468));
 sg13g2_tiehi _22266__1469 (.L_HI(net1469));
 sg13g2_tiehi _22265__1470 (.L_HI(net1470));
 sg13g2_tiehi _22264__1471 (.L_HI(net1471));
 sg13g2_tiehi _22263__1472 (.L_HI(net1472));
 sg13g2_tiehi _22262__1473 (.L_HI(net1473));
 sg13g2_tiehi _22261__1474 (.L_HI(net1474));
 sg13g2_tiehi _22260__1475 (.L_HI(net1475));
 sg13g2_tiehi _22259__1476 (.L_HI(net1476));
 sg13g2_tiehi _22258__1477 (.L_HI(net1477));
 sg13g2_tiehi _22257__1478 (.L_HI(net1478));
 sg13g2_tiehi _22256__1479 (.L_HI(net1479));
 sg13g2_tiehi _22255__1480 (.L_HI(net1480));
 sg13g2_tiehi _22254__1481 (.L_HI(net1481));
 sg13g2_tiehi _22253__1482 (.L_HI(net1482));
 sg13g2_tiehi _22252__1483 (.L_HI(net1483));
 sg13g2_tiehi _22251__1484 (.L_HI(net1484));
 sg13g2_tiehi _22250__1485 (.L_HI(net1485));
 sg13g2_tiehi _22249__1486 (.L_HI(net1486));
 sg13g2_tiehi _22248__1487 (.L_HI(net1487));
 sg13g2_tiehi _22247__1488 (.L_HI(net1488));
 sg13g2_tiehi _22246__1489 (.L_HI(net1489));
 sg13g2_tiehi _22245__1490 (.L_HI(net1490));
 sg13g2_tiehi _22244__1491 (.L_HI(net1491));
 sg13g2_tiehi _22243__1492 (.L_HI(net1492));
 sg13g2_tiehi _22242__1493 (.L_HI(net1493));
 sg13g2_tiehi _22241__1494 (.L_HI(net1494));
 sg13g2_tiehi _22240__1495 (.L_HI(net1495));
 sg13g2_tiehi _22239__1496 (.L_HI(net1496));
 sg13g2_tiehi _22238__1497 (.L_HI(net1497));
 sg13g2_tiehi _22237__1498 (.L_HI(net1498));
 sg13g2_tiehi _22236__1499 (.L_HI(net1499));
 sg13g2_tiehi _22235__1500 (.L_HI(net1500));
 sg13g2_tiehi _22234__1501 (.L_HI(net1501));
 sg13g2_tiehi _22233__1502 (.L_HI(net1502));
 sg13g2_tiehi _22232__1503 (.L_HI(net1503));
 sg13g2_tiehi _22231__1504 (.L_HI(net1504));
 sg13g2_tiehi _22230__1505 (.L_HI(net1505));
 sg13g2_tiehi _22229__1506 (.L_HI(net1506));
 sg13g2_tiehi _22228__1507 (.L_HI(net1507));
 sg13g2_tiehi _22227__1508 (.L_HI(net1508));
 sg13g2_tiehi _22226__1509 (.L_HI(net1509));
 sg13g2_tiehi _22225__1510 (.L_HI(net1510));
 sg13g2_tiehi _22224__1511 (.L_HI(net1511));
 sg13g2_tiehi _22223__1512 (.L_HI(net1512));
 sg13g2_tiehi _22222__1513 (.L_HI(net1513));
 sg13g2_tiehi _22221__1514 (.L_HI(net1514));
 sg13g2_tiehi _22220__1515 (.L_HI(net1515));
 sg13g2_tiehi _22219__1516 (.L_HI(net1516));
 sg13g2_tiehi _22218__1517 (.L_HI(net1517));
 sg13g2_tiehi _22217__1518 (.L_HI(net1518));
 sg13g2_tiehi _22216__1519 (.L_HI(net1519));
 sg13g2_tiehi _22215__1520 (.L_HI(net1520));
 sg13g2_tiehi _22214__1521 (.L_HI(net1521));
 sg13g2_tiehi _22213__1522 (.L_HI(net1522));
 sg13g2_tiehi _22212__1523 (.L_HI(net1523));
 sg13g2_tiehi _22211__1524 (.L_HI(net1524));
 sg13g2_tiehi _22210__1525 (.L_HI(net1525));
 sg13g2_tiehi _22209__1526 (.L_HI(net1526));
 sg13g2_tiehi _22208__1527 (.L_HI(net1527));
 sg13g2_tiehi _22207__1528 (.L_HI(net1528));
 sg13g2_tiehi _22206__1529 (.L_HI(net1529));
 sg13g2_tiehi _22205__1530 (.L_HI(net1530));
 sg13g2_tiehi _22204__1531 (.L_HI(net1531));
 sg13g2_tiehi _22203__1532 (.L_HI(net1532));
 sg13g2_tiehi _22202__1533 (.L_HI(net1533));
 sg13g2_tiehi _22201__1534 (.L_HI(net1534));
 sg13g2_tiehi _22200__1535 (.L_HI(net1535));
 sg13g2_tiehi _22199__1536 (.L_HI(net1536));
 sg13g2_tiehi _22198__1537 (.L_HI(net1537));
 sg13g2_tiehi _22197__1538 (.L_HI(net1538));
 sg13g2_tiehi _22196__1539 (.L_HI(net1539));
 sg13g2_tiehi _22195__1540 (.L_HI(net1540));
 sg13g2_tiehi _22194__1541 (.L_HI(net1541));
 sg13g2_tiehi _22193__1542 (.L_HI(net1542));
 sg13g2_tiehi _22192__1543 (.L_HI(net1543));
 sg13g2_tiehi _22191__1544 (.L_HI(net1544));
 sg13g2_tiehi _22190__1545 (.L_HI(net1545));
 sg13g2_tiehi _22189__1546 (.L_HI(net1546));
 sg13g2_tiehi _22188__1547 (.L_HI(net1547));
 sg13g2_tiehi _22187__1548 (.L_HI(net1548));
 sg13g2_tiehi _22186__1549 (.L_HI(net1549));
 sg13g2_tiehi _22185__1550 (.L_HI(net1550));
 sg13g2_tiehi _22184__1551 (.L_HI(net1551));
 sg13g2_tiehi _22183__1552 (.L_HI(net1552));
 sg13g2_tiehi _22182__1553 (.L_HI(net1553));
 sg13g2_tiehi _22181__1554 (.L_HI(net1554));
 sg13g2_tiehi _22180__1555 (.L_HI(net1555));
 sg13g2_tiehi _22179__1556 (.L_HI(net1556));
 sg13g2_tiehi _22178__1557 (.L_HI(net1557));
 sg13g2_tiehi _22177__1558 (.L_HI(net1558));
 sg13g2_tiehi _22176__1559 (.L_HI(net1559));
 sg13g2_tiehi _22175__1560 (.L_HI(net1560));
 sg13g2_tiehi _22174__1561 (.L_HI(net1561));
 sg13g2_tiehi _22173__1562 (.L_HI(net1562));
 sg13g2_tiehi _22172__1563 (.L_HI(net1563));
 sg13g2_tiehi _22171__1564 (.L_HI(net1564));
 sg13g2_tiehi _22170__1565 (.L_HI(net1565));
 sg13g2_tiehi _22169__1566 (.L_HI(net1566));
 sg13g2_tiehi _22168__1567 (.L_HI(net1567));
 sg13g2_tiehi _22167__1568 (.L_HI(net1568));
 sg13g2_tiehi _22166__1569 (.L_HI(net1569));
 sg13g2_tiehi _22165__1570 (.L_HI(net1570));
 sg13g2_tiehi _22164__1571 (.L_HI(net1571));
 sg13g2_tiehi _22163__1572 (.L_HI(net1572));
 sg13g2_tiehi _22162__1573 (.L_HI(net1573));
 sg13g2_tiehi _22161__1574 (.L_HI(net1574));
 sg13g2_tiehi _22160__1575 (.L_HI(net1575));
 sg13g2_tiehi _22159__1576 (.L_HI(net1576));
 sg13g2_tiehi _22158__1577 (.L_HI(net1577));
 sg13g2_tiehi _22157__1578 (.L_HI(net1578));
 sg13g2_tiehi _22156__1579 (.L_HI(net1579));
 sg13g2_tiehi _22155__1580 (.L_HI(net1580));
 sg13g2_tiehi _22154__1581 (.L_HI(net1581));
 sg13g2_tiehi _22153__1582 (.L_HI(net1582));
 sg13g2_tiehi _22152__1583 (.L_HI(net1583));
 sg13g2_tiehi _22151__1584 (.L_HI(net1584));
 sg13g2_tiehi _22150__1585 (.L_HI(net1585));
 sg13g2_tiehi _22149__1586 (.L_HI(net1586));
 sg13g2_tiehi _22148__1587 (.L_HI(net1587));
 sg13g2_tiehi _22147__1588 (.L_HI(net1588));
 sg13g2_tiehi _22146__1589 (.L_HI(net1589));
 sg13g2_tiehi _22145__1590 (.L_HI(net1590));
 sg13g2_tiehi _22144__1591 (.L_HI(net1591));
 sg13g2_tiehi _22143__1592 (.L_HI(net1592));
 sg13g2_tiehi _22142__1593 (.L_HI(net1593));
 sg13g2_tiehi _22141__1594 (.L_HI(net1594));
 sg13g2_tiehi _22140__1595 (.L_HI(net1595));
 sg13g2_tiehi _22139__1596 (.L_HI(net1596));
 sg13g2_tiehi _22138__1597 (.L_HI(net1597));
 sg13g2_tiehi _22137__1598 (.L_HI(net1598));
 sg13g2_tiehi _22136__1599 (.L_HI(net1599));
 sg13g2_tiehi _22135__1600 (.L_HI(net1600));
 sg13g2_tiehi _22134__1601 (.L_HI(net1601));
 sg13g2_tiehi _22133__1602 (.L_HI(net1602));
 sg13g2_tiehi _22132__1603 (.L_HI(net1603));
 sg13g2_tiehi _22131__1604 (.L_HI(net1604));
 sg13g2_tiehi _22130__1605 (.L_HI(net1605));
 sg13g2_tiehi _22129__1606 (.L_HI(net1606));
 sg13g2_tiehi _22128__1607 (.L_HI(net1607));
 sg13g2_tiehi _22127__1608 (.L_HI(net1608));
 sg13g2_tiehi _22126__1609 (.L_HI(net1609));
 sg13g2_tiehi _22125__1610 (.L_HI(net1610));
 sg13g2_tiehi _22124__1611 (.L_HI(net1611));
 sg13g2_tiehi _22123__1612 (.L_HI(net1612));
 sg13g2_tiehi _22122__1613 (.L_HI(net1613));
 sg13g2_tiehi _22121__1614 (.L_HI(net1614));
 sg13g2_tiehi _22120__1615 (.L_HI(net1615));
 sg13g2_tiehi _22119__1616 (.L_HI(net1616));
 sg13g2_tiehi _22118__1617 (.L_HI(net1617));
 sg13g2_tiehi _22117__1618 (.L_HI(net1618));
 sg13g2_tiehi _22116__1619 (.L_HI(net1619));
 sg13g2_tiehi _22115__1620 (.L_HI(net1620));
 sg13g2_tiehi _22114__1621 (.L_HI(net1621));
 sg13g2_tiehi _22113__1622 (.L_HI(net1622));
 sg13g2_tiehi _22112__1623 (.L_HI(net1623));
 sg13g2_tiehi _22111__1624 (.L_HI(net1624));
 sg13g2_tiehi _22110__1625 (.L_HI(net1625));
 sg13g2_tiehi _22109__1626 (.L_HI(net1626));
 sg13g2_tiehi _22108__1627 (.L_HI(net1627));
 sg13g2_tiehi _22107__1628 (.L_HI(net1628));
 sg13g2_tiehi _22106__1629 (.L_HI(net1629));
 sg13g2_tiehi _22105__1630 (.L_HI(net1630));
 sg13g2_tiehi _22104__1631 (.L_HI(net1631));
 sg13g2_tiehi _22103__1632 (.L_HI(net1632));
 sg13g2_tiehi _22102__1633 (.L_HI(net1633));
 sg13g2_tiehi _22101__1634 (.L_HI(net1634));
 sg13g2_tiehi _22100__1635 (.L_HI(net1635));
 sg13g2_tiehi _22099__1636 (.L_HI(net1636));
 sg13g2_tiehi _22098__1637 (.L_HI(net1637));
 sg13g2_tiehi _22097__1638 (.L_HI(net1638));
 sg13g2_tiehi _22096__1639 (.L_HI(net1639));
 sg13g2_tiehi _22095__1640 (.L_HI(net1640));
 sg13g2_tiehi _22094__1641 (.L_HI(net1641));
 sg13g2_tiehi _22093__1642 (.L_HI(net1642));
 sg13g2_tiehi _22092__1643 (.L_HI(net1643));
 sg13g2_tiehi _22091__1644 (.L_HI(net1644));
 sg13g2_tiehi _22090__1645 (.L_HI(net1645));
 sg13g2_tiehi _22089__1646 (.L_HI(net1646));
 sg13g2_tiehi _22088__1647 (.L_HI(net1647));
 sg13g2_tiehi _22087__1648 (.L_HI(net1648));
 sg13g2_tiehi _22086__1649 (.L_HI(net1649));
 sg13g2_tiehi _22085__1650 (.L_HI(net1650));
 sg13g2_tiehi _22084__1651 (.L_HI(net1651));
 sg13g2_tiehi _22083__1652 (.L_HI(net1652));
 sg13g2_tiehi _22082__1653 (.L_HI(net1653));
 sg13g2_tiehi _22081__1654 (.L_HI(net1654));
 sg13g2_tiehi _22080__1655 (.L_HI(net1655));
 sg13g2_tiehi _22079__1656 (.L_HI(net1656));
 sg13g2_tiehi _22078__1657 (.L_HI(net1657));
 sg13g2_tiehi _22077__1658 (.L_HI(net1658));
 sg13g2_tiehi _22076__1659 (.L_HI(net1659));
 sg13g2_tiehi _22075__1660 (.L_HI(net1660));
 sg13g2_tiehi _22074__1661 (.L_HI(net1661));
 sg13g2_tiehi _22073__1662 (.L_HI(net1662));
 sg13g2_tiehi _22072__1663 (.L_HI(net1663));
 sg13g2_tiehi _22071__1664 (.L_HI(net1664));
 sg13g2_tiehi _22070__1665 (.L_HI(net1665));
 sg13g2_tiehi _22069__1666 (.L_HI(net1666));
 sg13g2_tiehi _22068__1667 (.L_HI(net1667));
 sg13g2_tiehi _22067__1668 (.L_HI(net1668));
 sg13g2_tiehi _22066__1669 (.L_HI(net1669));
 sg13g2_tiehi _22065__1670 (.L_HI(net1670));
 sg13g2_tiehi _22064__1671 (.L_HI(net1671));
 sg13g2_tiehi _22063__1672 (.L_HI(net1672));
 sg13g2_tiehi _22062__1673 (.L_HI(net1673));
 sg13g2_tiehi _22061__1674 (.L_HI(net1674));
 sg13g2_tiehi _22060__1675 (.L_HI(net1675));
 sg13g2_tiehi _22059__1676 (.L_HI(net1676));
 sg13g2_tiehi _22058__1677 (.L_HI(net1677));
 sg13g2_tiehi _22057__1678 (.L_HI(net1678));
 sg13g2_tiehi _22056__1679 (.L_HI(net1679));
 sg13g2_tiehi _22055__1680 (.L_HI(net1680));
 sg13g2_tiehi _22054__1681 (.L_HI(net1681));
 sg13g2_tiehi _22053__1682 (.L_HI(net1682));
 sg13g2_tiehi _22052__1683 (.L_HI(net1683));
 sg13g2_tiehi _22051__1684 (.L_HI(net1684));
 sg13g2_tiehi _22050__1685 (.L_HI(net1685));
 sg13g2_tiehi _22049__1686 (.L_HI(net1686));
 sg13g2_tiehi _22048__1687 (.L_HI(net1687));
 sg13g2_tiehi _22047__1688 (.L_HI(net1688));
 sg13g2_tiehi _22046__1689 (.L_HI(net1689));
 sg13g2_tiehi _22045__1690 (.L_HI(net1690));
 sg13g2_tiehi _22044__1691 (.L_HI(net1691));
 sg13g2_tiehi _22043__1692 (.L_HI(net1692));
 sg13g2_tiehi _22042__1693 (.L_HI(net1693));
 sg13g2_tiehi _22041__1694 (.L_HI(net1694));
 sg13g2_tiehi _22040__1695 (.L_HI(net1695));
 sg13g2_tiehi _22039__1696 (.L_HI(net1696));
 sg13g2_tiehi _22038__1697 (.L_HI(net1697));
 sg13g2_tiehi _22037__1698 (.L_HI(net1698));
 sg13g2_tiehi _22036__1699 (.L_HI(net1699));
 sg13g2_tiehi _22035__1700 (.L_HI(net1700));
 sg13g2_tiehi _22034__1701 (.L_HI(net1701));
 sg13g2_tiehi _22033__1702 (.L_HI(net1702));
 sg13g2_tiehi _22032__1703 (.L_HI(net1703));
 sg13g2_tiehi _22031__1704 (.L_HI(net1704));
 sg13g2_tiehi _22030__1705 (.L_HI(net1705));
 sg13g2_tiehi _22029__1706 (.L_HI(net1706));
 sg13g2_tiehi _22028__1707 (.L_HI(net1707));
 sg13g2_tiehi _22027__1708 (.L_HI(net1708));
 sg13g2_tiehi _22026__1709 (.L_HI(net1709));
 sg13g2_tiehi _22025__1710 (.L_HI(net1710));
 sg13g2_tiehi _22024__1711 (.L_HI(net1711));
 sg13g2_tiehi _22023__1712 (.L_HI(net1712));
 sg13g2_tiehi _22022__1713 (.L_HI(net1713));
 sg13g2_tiehi _22021__1714 (.L_HI(net1714));
 sg13g2_tiehi _22020__1715 (.L_HI(net1715));
 sg13g2_tiehi _22019__1716 (.L_HI(net1716));
 sg13g2_tiehi _22018__1717 (.L_HI(net1717));
 sg13g2_tiehi _22017__1718 (.L_HI(net1718));
 sg13g2_tiehi _22016__1719 (.L_HI(net1719));
 sg13g2_tiehi _22015__1720 (.L_HI(net1720));
 sg13g2_tiehi _22014__1721 (.L_HI(net1721));
 sg13g2_tiehi _22013__1722 (.L_HI(net1722));
 sg13g2_tiehi _22012__1723 (.L_HI(net1723));
 sg13g2_tiehi _22011__1724 (.L_HI(net1724));
 sg13g2_tiehi _22010__1725 (.L_HI(net1725));
 sg13g2_tiehi _22009__1726 (.L_HI(net1726));
 sg13g2_tiehi _22008__1727 (.L_HI(net1727));
 sg13g2_tiehi _22007__1728 (.L_HI(net1728));
 sg13g2_tiehi _22006__1729 (.L_HI(net1729));
 sg13g2_tiehi _22005__1730 (.L_HI(net1730));
 sg13g2_tiehi _22004__1731 (.L_HI(net1731));
 sg13g2_tiehi _22003__1732 (.L_HI(net1732));
 sg13g2_tiehi _22002__1733 (.L_HI(net1733));
 sg13g2_tiehi _22001__1734 (.L_HI(net1734));
 sg13g2_tiehi _22000__1735 (.L_HI(net1735));
 sg13g2_tiehi _21999__1736 (.L_HI(net1736));
 sg13g2_tiehi _21998__1737 (.L_HI(net1737));
 sg13g2_tiehi _21997__1738 (.L_HI(net1738));
 sg13g2_tiehi _21996__1739 (.L_HI(net1739));
 sg13g2_tiehi _21995__1740 (.L_HI(net1740));
 sg13g2_tiehi _21994__1741 (.L_HI(net1741));
 sg13g2_tiehi _21993__1742 (.L_HI(net1742));
 sg13g2_tiehi _21992__1743 (.L_HI(net1743));
 sg13g2_tiehi _21991__1744 (.L_HI(net1744));
 sg13g2_tiehi _21990__1745 (.L_HI(net1745));
 sg13g2_tiehi _21989__1746 (.L_HI(net1746));
 sg13g2_tiehi _21988__1747 (.L_HI(net1747));
 sg13g2_tiehi _21987__1748 (.L_HI(net1748));
 sg13g2_tiehi _21986__1749 (.L_HI(net1749));
 sg13g2_tiehi _21985__1750 (.L_HI(net1750));
 sg13g2_tiehi _21984__1751 (.L_HI(net1751));
 sg13g2_tiehi _21983__1752 (.L_HI(net1752));
 sg13g2_tiehi _21982__1753 (.L_HI(net1753));
 sg13g2_tiehi _21981__1754 (.L_HI(net1754));
 sg13g2_tiehi _21980__1755 (.L_HI(net1755));
 sg13g2_tiehi _21979__1756 (.L_HI(net1756));
 sg13g2_tiehi _21978__1757 (.L_HI(net1757));
 sg13g2_tiehi _21977__1758 (.L_HI(net1758));
 sg13g2_tiehi _21976__1759 (.L_HI(net1759));
 sg13g2_tiehi _21975__1760 (.L_HI(net1760));
 sg13g2_tiehi _21974__1761 (.L_HI(net1761));
 sg13g2_tiehi _21973__1762 (.L_HI(net1762));
 sg13g2_tiehi _21972__1763 (.L_HI(net1763));
 sg13g2_tiehi _21971__1764 (.L_HI(net1764));
 sg13g2_tiehi _21970__1765 (.L_HI(net1765));
 sg13g2_tiehi _21969__1766 (.L_HI(net1766));
 sg13g2_tiehi _21968__1767 (.L_HI(net1767));
 sg13g2_tiehi _21967__1768 (.L_HI(net1768));
 sg13g2_tiehi _21966__1769 (.L_HI(net1769));
 sg13g2_tiehi _21965__1770 (.L_HI(net1770));
 sg13g2_tiehi _21964__1771 (.L_HI(net1771));
 sg13g2_tiehi _21963__1772 (.L_HI(net1772));
 sg13g2_tiehi _21962__1773 (.L_HI(net1773));
 sg13g2_tiehi _21961__1774 (.L_HI(net1774));
 sg13g2_tiehi _21960__1775 (.L_HI(net1775));
 sg13g2_tiehi _21959__1776 (.L_HI(net1776));
 sg13g2_tiehi _21958__1777 (.L_HI(net1777));
 sg13g2_tiehi _21957__1778 (.L_HI(net1778));
 sg13g2_tiehi _21956__1779 (.L_HI(net1779));
 sg13g2_tiehi _21955__1780 (.L_HI(net1780));
 sg13g2_tiehi _21954__1781 (.L_HI(net1781));
 sg13g2_tiehi _21953__1782 (.L_HI(net1782));
 sg13g2_tiehi _21952__1783 (.L_HI(net1783));
 sg13g2_tiehi _21951__1784 (.L_HI(net1784));
 sg13g2_tiehi _21950__1785 (.L_HI(net1785));
 sg13g2_tiehi _21949__1786 (.L_HI(net1786));
 sg13g2_tiehi _21948__1787 (.L_HI(net1787));
 sg13g2_tiehi _21947__1788 (.L_HI(net1788));
 sg13g2_tiehi _21946__1789 (.L_HI(net1789));
 sg13g2_tiehi _21945__1790 (.L_HI(net1790));
 sg13g2_tiehi _21944__1791 (.L_HI(net1791));
 sg13g2_tiehi _21943__1792 (.L_HI(net1792));
 sg13g2_tiehi _21942__1793 (.L_HI(net1793));
 sg13g2_tiehi _21941__1794 (.L_HI(net1794));
 sg13g2_tiehi _21940__1795 (.L_HI(net1795));
 sg13g2_tiehi _21939__1796 (.L_HI(net1796));
 sg13g2_tiehi _21938__1797 (.L_HI(net1797));
 sg13g2_tiehi _21937__1798 (.L_HI(net1798));
 sg13g2_tiehi _21936__1799 (.L_HI(net1799));
 sg13g2_tiehi _21935__1800 (.L_HI(net1800));
 sg13g2_tiehi _21934__1801 (.L_HI(net1801));
 sg13g2_tiehi _21933__1802 (.L_HI(net1802));
 sg13g2_tiehi _21932__1803 (.L_HI(net1803));
 sg13g2_tiehi _21931__1804 (.L_HI(net1804));
 sg13g2_tiehi _21930__1805 (.L_HI(net1805));
 sg13g2_tiehi _21929__1806 (.L_HI(net1806));
 sg13g2_tiehi _21928__1807 (.L_HI(net1807));
 sg13g2_tiehi _21927__1808 (.L_HI(net1808));
 sg13g2_tiehi _21926__1809 (.L_HI(net1809));
 sg13g2_tiehi _21925__1810 (.L_HI(net1810));
 sg13g2_tiehi _21924__1811 (.L_HI(net1811));
 sg13g2_tiehi _21923__1812 (.L_HI(net1812));
 sg13g2_tiehi _21922__1813 (.L_HI(net1813));
 sg13g2_tiehi _21921__1814 (.L_HI(net1814));
 sg13g2_tiehi _21920__1815 (.L_HI(net1815));
 sg13g2_tiehi _21919__1816 (.L_HI(net1816));
 sg13g2_tiehi _21918__1817 (.L_HI(net1817));
 sg13g2_tiehi _21917__1818 (.L_HI(net1818));
 sg13g2_tiehi _21916__1819 (.L_HI(net1819));
 sg13g2_tiehi _21915__1820 (.L_HI(net1820));
 sg13g2_tiehi _21914__1821 (.L_HI(net1821));
 sg13g2_tiehi _21913__1822 (.L_HI(net1822));
 sg13g2_tiehi _21912__1823 (.L_HI(net1823));
 sg13g2_tiehi _21911__1824 (.L_HI(net1824));
 sg13g2_tiehi _21910__1825 (.L_HI(net1825));
 sg13g2_tiehi _21909__1826 (.L_HI(net1826));
 sg13g2_tiehi _21908__1827 (.L_HI(net1827));
 sg13g2_tiehi _21907__1828 (.L_HI(net1828));
 sg13g2_tiehi _21906__1829 (.L_HI(net1829));
 sg13g2_tiehi _21905__1830 (.L_HI(net1830));
 sg13g2_tiehi _21904__1831 (.L_HI(net1831));
 sg13g2_tiehi _21903__1832 (.L_HI(net1832));
 sg13g2_tiehi _21902__1833 (.L_HI(net1833));
 sg13g2_tiehi _21901__1834 (.L_HI(net1834));
 sg13g2_tiehi _21900__1835 (.L_HI(net1835));
 sg13g2_tiehi _21899__1836 (.L_HI(net1836));
 sg13g2_tiehi _21898__1837 (.L_HI(net1837));
 sg13g2_tiehi _21897__1838 (.L_HI(net1838));
 sg13g2_tiehi _21896__1839 (.L_HI(net1839));
 sg13g2_tiehi _21895__1840 (.L_HI(net1840));
 sg13g2_tiehi _21894__1841 (.L_HI(net1841));
 sg13g2_tiehi _21893__1842 (.L_HI(net1842));
 sg13g2_tiehi _21892__1843 (.L_HI(net1843));
 sg13g2_tiehi _21891__1844 (.L_HI(net1844));
 sg13g2_tiehi _21890__1845 (.L_HI(net1845));
 sg13g2_tiehi _21889__1846 (.L_HI(net1846));
 sg13g2_tiehi _21888__1847 (.L_HI(net1847));
 sg13g2_tiehi _21887__1848 (.L_HI(net1848));
 sg13g2_tiehi _21886__1849 (.L_HI(net1849));
 sg13g2_tiehi _21885__1850 (.L_HI(net1850));
 sg13g2_tiehi _21884__1851 (.L_HI(net1851));
 sg13g2_tiehi _21883__1852 (.L_HI(net1852));
 sg13g2_tiehi _21882__1853 (.L_HI(net1853));
 sg13g2_tiehi _21881__1854 (.L_HI(net1854));
 sg13g2_tiehi _21880__1855 (.L_HI(net1855));
 sg13g2_tiehi _21879__1856 (.L_HI(net1856));
 sg13g2_tiehi _21878__1857 (.L_HI(net1857));
 sg13g2_tiehi _21877__1858 (.L_HI(net1858));
 sg13g2_tiehi _21876__1859 (.L_HI(net1859));
 sg13g2_tiehi _21875__1860 (.L_HI(net1860));
 sg13g2_tiehi _21874__1861 (.L_HI(net1861));
 sg13g2_tiehi _21873__1862 (.L_HI(net1862));
 sg13g2_tiehi _21872__1863 (.L_HI(net1863));
 sg13g2_tiehi _21871__1864 (.L_HI(net1864));
 sg13g2_tiehi _21870__1865 (.L_HI(net1865));
 sg13g2_tiehi _21869__1866 (.L_HI(net1866));
 sg13g2_tiehi _21868__1867 (.L_HI(net1867));
 sg13g2_tiehi _21867__1868 (.L_HI(net1868));
 sg13g2_tiehi _21866__1869 (.L_HI(net1869));
 sg13g2_tiehi _21865__1870 (.L_HI(net1870));
 sg13g2_tiehi _21864__1871 (.L_HI(net1871));
 sg13g2_tiehi _21863__1872 (.L_HI(net1872));
 sg13g2_tiehi _21862__1873 (.L_HI(net1873));
 sg13g2_tiehi _21861__1874 (.L_HI(net1874));
 sg13g2_tiehi _21860__1875 (.L_HI(net1875));
 sg13g2_tiehi _21859__1876 (.L_HI(net1876));
 sg13g2_tiehi _21858__1877 (.L_HI(net1877));
 sg13g2_tiehi _21857__1878 (.L_HI(net1878));
 sg13g2_tiehi _21856__1879 (.L_HI(net1879));
 sg13g2_tiehi _21855__1880 (.L_HI(net1880));
 sg13g2_tiehi _21854__1881 (.L_HI(net1881));
 sg13g2_tiehi _21853__1882 (.L_HI(net1882));
 sg13g2_tiehi _21852__1883 (.L_HI(net1883));
 sg13g2_tiehi _21851__1884 (.L_HI(net1884));
 sg13g2_tiehi _21850__1885 (.L_HI(net1885));
 sg13g2_tiehi _21849__1886 (.L_HI(net1886));
 sg13g2_tiehi _21848__1887 (.L_HI(net1887));
 sg13g2_tiehi _21847__1888 (.L_HI(net1888));
 sg13g2_tiehi _21846__1889 (.L_HI(net1889));
 sg13g2_tiehi _21845__1890 (.L_HI(net1890));
 sg13g2_tiehi _21844__1891 (.L_HI(net1891));
 sg13g2_tiehi _21843__1892 (.L_HI(net1892));
 sg13g2_tiehi _21842__1893 (.L_HI(net1893));
 sg13g2_tiehi _21841__1894 (.L_HI(net1894));
 sg13g2_tiehi _21840__1895 (.L_HI(net1895));
 sg13g2_tiehi _21839__1896 (.L_HI(net1896));
 sg13g2_tiehi _21838__1897 (.L_HI(net1897));
 sg13g2_tiehi _21837__1898 (.L_HI(net1898));
 sg13g2_tiehi _21836__1899 (.L_HI(net1899));
 sg13g2_tiehi _21835__1900 (.L_HI(net1900));
 sg13g2_tiehi _21834__1901 (.L_HI(net1901));
 sg13g2_tiehi _21833__1902 (.L_HI(net1902));
 sg13g2_tiehi _21832__1903 (.L_HI(net1903));
 sg13g2_tiehi _21831__1904 (.L_HI(net1904));
 sg13g2_tiehi _21830__1905 (.L_HI(net1905));
 sg13g2_tiehi _21829__1906 (.L_HI(net1906));
 sg13g2_tiehi _21828__1907 (.L_HI(net1907));
 sg13g2_tiehi _21827__1908 (.L_HI(net1908));
 sg13g2_tiehi _21826__1909 (.L_HI(net1909));
 sg13g2_tiehi _21825__1910 (.L_HI(net1910));
 sg13g2_tiehi _21824__1911 (.L_HI(net1911));
 sg13g2_tiehi _21823__1912 (.L_HI(net1912));
 sg13g2_tiehi _21822__1913 (.L_HI(net1913));
 sg13g2_tiehi _21821__1914 (.L_HI(net1914));
 sg13g2_tiehi _21820__1915 (.L_HI(net1915));
 sg13g2_tiehi _21819__1916 (.L_HI(net1916));
 sg13g2_tiehi _21818__1917 (.L_HI(net1917));
 sg13g2_tiehi _21817__1918 (.L_HI(net1918));
 sg13g2_tiehi _21816__1919 (.L_HI(net1919));
 sg13g2_tiehi _21815__1920 (.L_HI(net1920));
 sg13g2_tiehi _21814__1921 (.L_HI(net1921));
 sg13g2_tiehi _21813__1922 (.L_HI(net1922));
 sg13g2_tiehi _21812__1923 (.L_HI(net1923));
 sg13g2_tiehi _21811__1924 (.L_HI(net1924));
 sg13g2_tiehi _21810__1925 (.L_HI(net1925));
 sg13g2_tiehi _21809__1926 (.L_HI(net1926));
 sg13g2_tiehi _21808__1927 (.L_HI(net1927));
 sg13g2_tiehi _21807__1928 (.L_HI(net1928));
 sg13g2_tiehi _21806__1929 (.L_HI(net1929));
 sg13g2_tiehi _21805__1930 (.L_HI(net1930));
 sg13g2_tiehi _21804__1931 (.L_HI(net1931));
 sg13g2_tiehi _21803__1932 (.L_HI(net1932));
 sg13g2_tiehi _21802__1933 (.L_HI(net1933));
 sg13g2_tiehi _21801__1934 (.L_HI(net1934));
 sg13g2_tiehi _21800__1935 (.L_HI(net1935));
 sg13g2_tiehi _21799__1936 (.L_HI(net1936));
 sg13g2_tiehi _21798__1937 (.L_HI(net1937));
 sg13g2_tiehi _21797__1938 (.L_HI(net1938));
 sg13g2_tiehi _21796__1939 (.L_HI(net1939));
 sg13g2_tiehi _21795__1940 (.L_HI(net1940));
 sg13g2_tiehi _21794__1941 (.L_HI(net1941));
 sg13g2_tiehi _21793__1942 (.L_HI(net1942));
 sg13g2_tiehi _21792__1943 (.L_HI(net1943));
 sg13g2_tiehi _21791__1944 (.L_HI(net1944));
 sg13g2_tiehi _21790__1945 (.L_HI(net1945));
 sg13g2_tiehi _21789__1946 (.L_HI(net1946));
 sg13g2_tiehi _21788__1947 (.L_HI(net1947));
 sg13g2_tiehi _21787__1948 (.L_HI(net1948));
 sg13g2_tiehi _21786__1949 (.L_HI(net1949));
 sg13g2_tiehi _21785__1950 (.L_HI(net1950));
 sg13g2_tiehi _21784__1951 (.L_HI(net1951));
 sg13g2_tiehi _21783__1952 (.L_HI(net1952));
 sg13g2_tiehi _21782__1953 (.L_HI(net1953));
 sg13g2_tiehi _21781__1954 (.L_HI(net1954));
 sg13g2_tiehi _21780__1955 (.L_HI(net1955));
 sg13g2_tiehi _21779__1956 (.L_HI(net1956));
 sg13g2_tiehi _21778__1957 (.L_HI(net1957));
 sg13g2_tiehi _21777__1958 (.L_HI(net1958));
 sg13g2_tiehi _21776__1959 (.L_HI(net1959));
 sg13g2_tiehi _21775__1960 (.L_HI(net1960));
 sg13g2_tiehi _21774__1961 (.L_HI(net1961));
 sg13g2_tiehi _21773__1962 (.L_HI(net1962));
 sg13g2_tiehi _21772__1963 (.L_HI(net1963));
 sg13g2_tiehi _21771__1964 (.L_HI(net1964));
 sg13g2_tiehi _21770__1965 (.L_HI(net1965));
 sg13g2_tiehi _21769__1966 (.L_HI(net1966));
 sg13g2_tiehi _21768__1967 (.L_HI(net1967));
 sg13g2_tiehi _21767__1968 (.L_HI(net1968));
 sg13g2_tiehi _21766__1969 (.L_HI(net1969));
 sg13g2_tiehi _21765__1970 (.L_HI(net1970));
 sg13g2_tiehi _21764__1971 (.L_HI(net1971));
 sg13g2_tiehi _21763__1972 (.L_HI(net1972));
 sg13g2_tiehi _21762__1973 (.L_HI(net1973));
 sg13g2_tiehi _21761__1974 (.L_HI(net1974));
 sg13g2_tiehi _21760__1975 (.L_HI(net1975));
 sg13g2_tiehi _21759__1976 (.L_HI(net1976));
 sg13g2_tiehi _21758__1977 (.L_HI(net1977));
 sg13g2_tiehi _21757__1978 (.L_HI(net1978));
 sg13g2_tiehi _21756__1979 (.L_HI(net1979));
 sg13g2_tiehi _21755__1980 (.L_HI(net1980));
 sg13g2_tiehi _21754__1981 (.L_HI(net1981));
 sg13g2_tiehi _21753__1982 (.L_HI(net1982));
 sg13g2_tiehi _21752__1983 (.L_HI(net1983));
 sg13g2_tiehi _21751__1984 (.L_HI(net1984));
 sg13g2_tiehi _21750__1985 (.L_HI(net1985));
 sg13g2_tiehi _21749__1986 (.L_HI(net1986));
 sg13g2_tiehi _21748__1987 (.L_HI(net1987));
 sg13g2_tiehi _21747__1988 (.L_HI(net1988));
 sg13g2_tiehi _21746__1989 (.L_HI(net1989));
 sg13g2_tiehi _21745__1990 (.L_HI(net1990));
 sg13g2_tiehi _21744__1991 (.L_HI(net1991));
 sg13g2_tiehi _21743__1992 (.L_HI(net1992));
 sg13g2_tiehi _21742__1993 (.L_HI(net1993));
 sg13g2_tiehi _21741__1994 (.L_HI(net1994));
 sg13g2_tiehi _21740__1995 (.L_HI(net1995));
 sg13g2_tiehi _21739__1996 (.L_HI(net1996));
 sg13g2_tiehi _21738__1997 (.L_HI(net1997));
 sg13g2_tiehi _21737__1998 (.L_HI(net1998));
 sg13g2_tiehi _21736__1999 (.L_HI(net1999));
 sg13g2_tiehi _21735__2000 (.L_HI(net2000));
 sg13g2_tiehi _21734__2001 (.L_HI(net2001));
 sg13g2_tiehi _21733__2002 (.L_HI(net2002));
 sg13g2_tiehi _21732__2003 (.L_HI(net2003));
 sg13g2_tiehi _21731__2004 (.L_HI(net2004));
 sg13g2_tiehi _21730__2005 (.L_HI(net2005));
 sg13g2_tiehi _21729__2006 (.L_HI(net2006));
 sg13g2_tiehi _21728__2007 (.L_HI(net2007));
 sg13g2_tiehi _21727__2008 (.L_HI(net2008));
 sg13g2_tiehi _21726__2009 (.L_HI(net2009));
 sg13g2_tiehi _21725__2010 (.L_HI(net2010));
 sg13g2_tiehi _21724__2011 (.L_HI(net2011));
 sg13g2_tiehi _21723__2012 (.L_HI(net2012));
 sg13g2_tiehi _21722__2013 (.L_HI(net2013));
 sg13g2_tiehi _21721__2014 (.L_HI(net2014));
 sg13g2_tiehi _21720__2015 (.L_HI(net2015));
 sg13g2_tiehi _21719__2016 (.L_HI(net2016));
 sg13g2_tiehi _21718__2017 (.L_HI(net2017));
 sg13g2_tiehi _21717__2018 (.L_HI(net2018));
 sg13g2_tiehi _21716__2019 (.L_HI(net2019));
 sg13g2_tiehi _21715__2020 (.L_HI(net2020));
 sg13g2_tiehi _21714__2021 (.L_HI(net2021));
 sg13g2_tiehi _21713__2022 (.L_HI(net2022));
 sg13g2_tiehi _21712__2023 (.L_HI(net2023));
 sg13g2_tiehi _21711__2024 (.L_HI(net2024));
 sg13g2_tiehi _21710__2025 (.L_HI(net2025));
 sg13g2_tiehi _21709__2026 (.L_HI(net2026));
 sg13g2_tiehi _21708__2027 (.L_HI(net2027));
 sg13g2_tiehi _21707__2028 (.L_HI(net2028));
 sg13g2_tiehi _21706__2029 (.L_HI(net2029));
 sg13g2_tiehi _21705__2030 (.L_HI(net2030));
 sg13g2_tiehi _21704__2031 (.L_HI(net2031));
 sg13g2_tiehi _21703__2032 (.L_HI(net2032));
 sg13g2_tiehi _21702__2033 (.L_HI(net2033));
 sg13g2_tiehi _21701__2034 (.L_HI(net2034));
 sg13g2_tiehi _21700__2035 (.L_HI(net2035));
 sg13g2_tiehi _21699__2036 (.L_HI(net2036));
 sg13g2_tiehi _21698__2037 (.L_HI(net2037));
 sg13g2_tiehi _21697__2038 (.L_HI(net2038));
 sg13g2_tiehi _21696__2039 (.L_HI(net2039));
 sg13g2_tiehi _21695__2040 (.L_HI(net2040));
 sg13g2_tiehi _21694__2041 (.L_HI(net2041));
 sg13g2_tiehi _21693__2042 (.L_HI(net2042));
 sg13g2_tiehi _21692__2043 (.L_HI(net2043));
 sg13g2_tiehi _21691__2044 (.L_HI(net2044));
 sg13g2_tiehi _21690__2045 (.L_HI(net2045));
 sg13g2_tiehi _21689__2046 (.L_HI(net2046));
 sg13g2_tiehi _21688__2047 (.L_HI(net2047));
 sg13g2_tiehi _21687__2048 (.L_HI(net2048));
 sg13g2_tiehi _21686__2049 (.L_HI(net2049));
 sg13g2_tiehi _21685__2050 (.L_HI(net2050));
 sg13g2_tiehi _21684__2051 (.L_HI(net2051));
 sg13g2_tiehi _21683__2052 (.L_HI(net2052));
 sg13g2_tiehi _21682__2053 (.L_HI(net2053));
 sg13g2_tiehi _21681__2054 (.L_HI(net2054));
 sg13g2_tiehi _21680__2055 (.L_HI(net2055));
 sg13g2_tiehi _21679__2056 (.L_HI(net2056));
 sg13g2_tiehi _21678__2057 (.L_HI(net2057));
 sg13g2_tiehi _21677__2058 (.L_HI(net2058));
 sg13g2_tiehi _21676__2059 (.L_HI(net2059));
 sg13g2_tiehi _21675__2060 (.L_HI(net2060));
 sg13g2_tiehi _21674__2061 (.L_HI(net2061));
 sg13g2_tiehi _21673__2062 (.L_HI(net2062));
 sg13g2_tiehi _21672__2063 (.L_HI(net2063));
 sg13g2_tiehi _21671__2064 (.L_HI(net2064));
 sg13g2_tiehi _21670__2065 (.L_HI(net2065));
 sg13g2_tiehi _21669__2066 (.L_HI(net2066));
 sg13g2_tiehi _21668__2067 (.L_HI(net2067));
 sg13g2_tiehi _21667__2068 (.L_HI(net2068));
 sg13g2_tiehi _21666__2069 (.L_HI(net2069));
 sg13g2_tiehi _21665__2070 (.L_HI(net2070));
 sg13g2_tiehi _21664__2071 (.L_HI(net2071));
 sg13g2_tiehi _21663__2072 (.L_HI(net2072));
 sg13g2_tiehi _21662__2073 (.L_HI(net2073));
 sg13g2_tiehi _21661__2074 (.L_HI(net2074));
 sg13g2_tiehi _21660__2075 (.L_HI(net2075));
 sg13g2_tiehi _21659__2076 (.L_HI(net2076));
 sg13g2_tiehi _21658__2077 (.L_HI(net2077));
 sg13g2_tiehi _21657__2078 (.L_HI(net2078));
 sg13g2_tiehi _21656__2079 (.L_HI(net2079));
 sg13g2_tiehi _21655__2080 (.L_HI(net2080));
 sg13g2_tiehi _21654__2081 (.L_HI(net2081));
 sg13g2_tiehi _21653__2082 (.L_HI(net2082));
 sg13g2_tiehi _21652__2083 (.L_HI(net2083));
 sg13g2_tiehi _21651__2084 (.L_HI(net2084));
 sg13g2_tiehi _21650__2085 (.L_HI(net2085));
 sg13g2_tiehi _21649__2086 (.L_HI(net2086));
 sg13g2_tiehi _21648__2087 (.L_HI(net2087));
 sg13g2_tiehi _21647__2088 (.L_HI(net2088));
 sg13g2_tiehi _21646__2089 (.L_HI(net2089));
 sg13g2_tiehi _21645__2090 (.L_HI(net2090));
 sg13g2_tiehi _21644__2091 (.L_HI(net2091));
 sg13g2_tiehi _21643__2092 (.L_HI(net2092));
 sg13g2_tiehi _21642__2093 (.L_HI(net2093));
 sg13g2_tiehi _21641__2094 (.L_HI(net2094));
 sg13g2_tiehi _21640__2095 (.L_HI(net2095));
 sg13g2_tiehi _21639__2096 (.L_HI(net2096));
 sg13g2_tiehi _21638__2097 (.L_HI(net2097));
 sg13g2_tiehi _21637__2098 (.L_HI(net2098));
 sg13g2_tiehi _21636__2099 (.L_HI(net2099));
 sg13g2_tiehi _21635__2100 (.L_HI(net2100));
 sg13g2_tiehi _21634__2101 (.L_HI(net2101));
 sg13g2_tiehi _21633__2102 (.L_HI(net2102));
 sg13g2_tiehi _21632__2103 (.L_HI(net2103));
 sg13g2_tiehi _21631__2104 (.L_HI(net2104));
 sg13g2_tiehi _21630__2105 (.L_HI(net2105));
 sg13g2_tiehi _21629__2106 (.L_HI(net2106));
 sg13g2_tiehi _21628__2107 (.L_HI(net2107));
 sg13g2_tiehi _21627__2108 (.L_HI(net2108));
 sg13g2_tiehi _21626__2109 (.L_HI(net2109));
 sg13g2_tiehi _21625__2110 (.L_HI(net2110));
 sg13g2_tiehi _21624__2111 (.L_HI(net2111));
 sg13g2_tiehi _21623__2112 (.L_HI(net2112));
 sg13g2_tiehi _21622__2113 (.L_HI(net2113));
 sg13g2_tiehi _21621__2114 (.L_HI(net2114));
 sg13g2_tiehi _21620__2115 (.L_HI(net2115));
 sg13g2_tiehi _21619__2116 (.L_HI(net2116));
 sg13g2_tiehi _21618__2117 (.L_HI(net2117));
 sg13g2_tiehi _21617__2118 (.L_HI(net2118));
 sg13g2_tiehi _21616__2119 (.L_HI(net2119));
 sg13g2_tiehi _21615__2120 (.L_HI(net2120));
 sg13g2_tiehi _21614__2121 (.L_HI(net2121));
 sg13g2_tiehi _21613__2122 (.L_HI(net2122));
 sg13g2_tiehi _21612__2123 (.L_HI(net2123));
 sg13g2_tiehi _21611__2124 (.L_HI(net2124));
 sg13g2_tiehi _21610__2125 (.L_HI(net2125));
 sg13g2_tiehi _21609__2126 (.L_HI(net2126));
 sg13g2_tiehi _21608__2127 (.L_HI(net2127));
 sg13g2_tiehi _21607__2128 (.L_HI(net2128));
 sg13g2_tiehi _21606__2129 (.L_HI(net2129));
 sg13g2_tiehi _21605__2130 (.L_HI(net2130));
 sg13g2_tiehi _21604__2131 (.L_HI(net2131));
 sg13g2_tiehi _21603__2132 (.L_HI(net2132));
 sg13g2_tiehi _21602__2133 (.L_HI(net2133));
 sg13g2_tiehi _21601__2134 (.L_HI(net2134));
 sg13g2_tiehi _21600__2135 (.L_HI(net2135));
 sg13g2_tiehi _21599__2136 (.L_HI(net2136));
 sg13g2_tiehi _21598__2137 (.L_HI(net2137));
 sg13g2_tiehi _21597__2138 (.L_HI(net2138));
 sg13g2_tiehi _21596__2139 (.L_HI(net2139));
 sg13g2_tiehi _21595__2140 (.L_HI(net2140));
 sg13g2_tiehi _21594__2141 (.L_HI(net2141));
 sg13g2_tiehi _21593__2142 (.L_HI(net2142));
 sg13g2_tiehi _21592__2143 (.L_HI(net2143));
 sg13g2_tiehi _21591__2144 (.L_HI(net2144));
 sg13g2_tiehi _21590__2145 (.L_HI(net2145));
 sg13g2_tiehi _21589__2146 (.L_HI(net2146));
 sg13g2_tiehi _21588__2147 (.L_HI(net2147));
 sg13g2_tiehi _21587__2148 (.L_HI(net2148));
 sg13g2_tiehi _21586__2149 (.L_HI(net2149));
 sg13g2_tiehi _21585__2150 (.L_HI(net2150));
 sg13g2_tiehi _21584__2151 (.L_HI(net2151));
 sg13g2_tiehi _21583__2152 (.L_HI(net2152));
 sg13g2_tiehi _21582__2153 (.L_HI(net2153));
 sg13g2_tiehi _21581__2154 (.L_HI(net2154));
 sg13g2_tiehi _21580__2155 (.L_HI(net2155));
 sg13g2_tiehi _21579__2156 (.L_HI(net2156));
 sg13g2_tiehi _21578__2157 (.L_HI(net2157));
 sg13g2_tiehi _21577__2158 (.L_HI(net2158));
 sg13g2_tiehi _21576__2159 (.L_HI(net2159));
 sg13g2_tiehi _21575__2160 (.L_HI(net2160));
 sg13g2_tiehi _21574__2161 (.L_HI(net2161));
 sg13g2_tiehi _21573__2162 (.L_HI(net2162));
 sg13g2_tiehi _21572__2163 (.L_HI(net2163));
 sg13g2_tiehi _21571__2164 (.L_HI(net2164));
 sg13g2_tiehi _21570__2165 (.L_HI(net2165));
 sg13g2_tiehi _21569__2166 (.L_HI(net2166));
 sg13g2_tiehi _21568__2167 (.L_HI(net2167));
 sg13g2_tiehi _21567__2168 (.L_HI(net2168));
 sg13g2_tiehi _21566__2169 (.L_HI(net2169));
 sg13g2_tiehi _21565__2170 (.L_HI(net2170));
 sg13g2_tiehi _21564__2171 (.L_HI(net2171));
 sg13g2_tiehi _21563__2172 (.L_HI(net2172));
 sg13g2_tiehi _21562__2173 (.L_HI(net2173));
 sg13g2_tiehi _21561__2174 (.L_HI(net2174));
 sg13g2_tiehi _21560__2175 (.L_HI(net2175));
 sg13g2_tiehi _21559__2176 (.L_HI(net2176));
 sg13g2_tiehi _21558__2177 (.L_HI(net2177));
 sg13g2_tiehi _21557__2178 (.L_HI(net2178));
 sg13g2_tiehi _21556__2179 (.L_HI(net2179));
 sg13g2_tiehi _21555__2180 (.L_HI(net2180));
 sg13g2_tiehi _21554__2181 (.L_HI(net2181));
 sg13g2_tiehi _21553__2182 (.L_HI(net2182));
 sg13g2_tiehi _21552__2183 (.L_HI(net2183));
 sg13g2_tiehi _21551__2184 (.L_HI(net2184));
 sg13g2_tiehi _21550__2185 (.L_HI(net2185));
 sg13g2_tiehi _21549__2186 (.L_HI(net2186));
 sg13g2_tiehi _21548__2187 (.L_HI(net2187));
 sg13g2_tiehi _21547__2188 (.L_HI(net2188));
 sg13g2_tiehi _21546__2189 (.L_HI(net2189));
 sg13g2_tiehi _21545__2190 (.L_HI(net2190));
 sg13g2_tiehi _21544__2191 (.L_HI(net2191));
 sg13g2_tiehi _21543__2192 (.L_HI(net2192));
 sg13g2_tiehi _21542__2193 (.L_HI(net2193));
 sg13g2_tiehi _21541__2194 (.L_HI(net2194));
 sg13g2_tiehi _21540__2195 (.L_HI(net2195));
 sg13g2_tiehi _21539__2196 (.L_HI(net2196));
 sg13g2_tiehi _21538__2197 (.L_HI(net2197));
 sg13g2_tiehi _21537__2198 (.L_HI(net2198));
 sg13g2_tiehi _21536__2199 (.L_HI(net2199));
 sg13g2_tiehi _21535__2200 (.L_HI(net2200));
 sg13g2_tiehi _21534__2201 (.L_HI(net2201));
 sg13g2_tiehi _21533__2202 (.L_HI(net2202));
 sg13g2_tiehi _21532__2203 (.L_HI(net2203));
 sg13g2_tiehi _21531__2204 (.L_HI(net2204));
 sg13g2_tiehi _21530__2205 (.L_HI(net2205));
 sg13g2_tiehi _21529__2206 (.L_HI(net2206));
 sg13g2_tiehi _21528__2207 (.L_HI(net2207));
 sg13g2_tiehi _21527__2208 (.L_HI(net2208));
 sg13g2_tiehi _21526__2209 (.L_HI(net2209));
 sg13g2_tiehi _21525__2210 (.L_HI(net2210));
 sg13g2_tiehi _21524__2211 (.L_HI(net2211));
 sg13g2_tiehi _21523__2212 (.L_HI(net2212));
 sg13g2_tiehi _21522__2213 (.L_HI(net2213));
 sg13g2_tiehi _21521__2214 (.L_HI(net2214));
 sg13g2_tiehi _21520__2215 (.L_HI(net2215));
 sg13g2_tiehi _21519__2216 (.L_HI(net2216));
 sg13g2_tiehi _21518__2217 (.L_HI(net2217));
 sg13g2_tiehi _21517__2218 (.L_HI(net2218));
 sg13g2_tiehi _21516__2219 (.L_HI(net2219));
 sg13g2_tiehi _21515__2220 (.L_HI(net2220));
 sg13g2_tiehi _21514__2221 (.L_HI(net2221));
 sg13g2_tiehi _21513__2222 (.L_HI(net2222));
 sg13g2_tiehi _21512__2223 (.L_HI(net2223));
 sg13g2_tiehi _21511__2224 (.L_HI(net2224));
 sg13g2_tiehi _21510__2225 (.L_HI(net2225));
 sg13g2_tiehi _21509__2226 (.L_HI(net2226));
 sg13g2_tiehi _21508__2227 (.L_HI(net2227));
 sg13g2_tiehi _21507__2228 (.L_HI(net2228));
 sg13g2_tiehi _21506__2229 (.L_HI(net2229));
 sg13g2_tiehi _21505__2230 (.L_HI(net2230));
 sg13g2_tiehi _21504__2231 (.L_HI(net2231));
 sg13g2_tiehi _21503__2232 (.L_HI(net2232));
 sg13g2_tiehi _21502__2233 (.L_HI(net2233));
 sg13g2_tiehi _21501__2234 (.L_HI(net2234));
 sg13g2_tiehi _21500__2235 (.L_HI(net2235));
 sg13g2_tiehi _21499__2236 (.L_HI(net2236));
 sg13g2_tiehi _21498__2237 (.L_HI(net2237));
 sg13g2_tiehi _21497__2238 (.L_HI(net2238));
 sg13g2_tiehi _21496__2239 (.L_HI(net2239));
 sg13g2_tiehi _21495__2240 (.L_HI(net2240));
 sg13g2_tiehi _21494__2241 (.L_HI(net2241));
 sg13g2_tiehi _21493__2242 (.L_HI(net2242));
 sg13g2_tiehi _21492__2243 (.L_HI(net2243));
 sg13g2_tiehi _21491__2244 (.L_HI(net2244));
 sg13g2_tiehi _21490__2245 (.L_HI(net2245));
 sg13g2_tiehi _21489__2246 (.L_HI(net2246));
 sg13g2_tiehi _21488__2247 (.L_HI(net2247));
 sg13g2_tiehi _21487__2248 (.L_HI(net2248));
 sg13g2_tiehi _21486__2249 (.L_HI(net2249));
 sg13g2_tiehi _21485__2250 (.L_HI(net2250));
 sg13g2_tiehi _21484__2251 (.L_HI(net2251));
 sg13g2_tiehi _21483__2252 (.L_HI(net2252));
 sg13g2_tiehi _21482__2253 (.L_HI(net2253));
 sg13g2_tiehi _21481__2254 (.L_HI(net2254));
 sg13g2_tiehi _21480__2255 (.L_HI(net2255));
 sg13g2_tiehi _21479__2256 (.L_HI(net2256));
 sg13g2_tiehi _21478__2257 (.L_HI(net2257));
 sg13g2_tiehi _21477__2258 (.L_HI(net2258));
 sg13g2_tiehi _21476__2259 (.L_HI(net2259));
 sg13g2_tiehi _21475__2260 (.L_HI(net2260));
 sg13g2_tiehi _21474__2261 (.L_HI(net2261));
 sg13g2_tiehi _21473__2262 (.L_HI(net2262));
 sg13g2_tiehi _21472__2263 (.L_HI(net2263));
 sg13g2_tiehi _21471__2264 (.L_HI(net2264));
 sg13g2_tiehi _21470__2265 (.L_HI(net2265));
 sg13g2_tiehi _21469__2266 (.L_HI(net2266));
 sg13g2_tiehi _21468__2267 (.L_HI(net2267));
 sg13g2_tiehi _21467__2268 (.L_HI(net2268));
 sg13g2_tiehi _21466__2269 (.L_HI(net2269));
 sg13g2_tiehi _21465__2270 (.L_HI(net2270));
 sg13g2_tiehi _21464__2271 (.L_HI(net2271));
 sg13g2_tiehi _21463__2272 (.L_HI(net2272));
 sg13g2_tiehi _21462__2273 (.L_HI(net2273));
 sg13g2_tiehi _21461__2274 (.L_HI(net2274));
 sg13g2_tiehi _21460__2275 (.L_HI(net2275));
 sg13g2_tiehi _21459__2276 (.L_HI(net2276));
 sg13g2_tiehi _21458__2277 (.L_HI(net2277));
 sg13g2_tiehi _21457__2278 (.L_HI(net2278));
 sg13g2_tiehi _21456__2279 (.L_HI(net2279));
 sg13g2_tiehi _21455__2280 (.L_HI(net2280));
 sg13g2_tiehi _21454__2281 (.L_HI(net2281));
 sg13g2_tiehi _21453__2282 (.L_HI(net2282));
 sg13g2_tiehi _21452__2283 (.L_HI(net2283));
 sg13g2_tiehi _21451__2284 (.L_HI(net2284));
 sg13g2_tiehi _21450__2285 (.L_HI(net2285));
 sg13g2_tiehi _21449__2286 (.L_HI(net2286));
 sg13g2_tiehi _21448__2287 (.L_HI(net2287));
 sg13g2_tiehi _21447__2288 (.L_HI(net2288));
 sg13g2_tiehi _21446__2289 (.L_HI(net2289));
 sg13g2_tiehi _21445__2290 (.L_HI(net2290));
 sg13g2_tiehi _21444__2291 (.L_HI(net2291));
 sg13g2_tiehi _21443__2292 (.L_HI(net2292));
 sg13g2_tiehi _21442__2293 (.L_HI(net2293));
 sg13g2_tiehi _21441__2294 (.L_HI(net2294));
 sg13g2_tiehi _21440__2295 (.L_HI(net2295));
 sg13g2_tiehi _21439__2296 (.L_HI(net2296));
 sg13g2_tiehi _21438__2297 (.L_HI(net2297));
 sg13g2_tiehi _21437__2298 (.L_HI(net2298));
 sg13g2_tiehi _21436__2299 (.L_HI(net2299));
 sg13g2_tiehi _21435__2300 (.L_HI(net2300));
 sg13g2_tiehi _21434__2301 (.L_HI(net2301));
 sg13g2_tiehi _21433__2302 (.L_HI(net2302));
 sg13g2_tiehi _21432__2303 (.L_HI(net2303));
 sg13g2_tiehi _21431__2304 (.L_HI(net2304));
 sg13g2_tiehi _21430__2305 (.L_HI(net2305));
 sg13g2_tiehi _21429__2306 (.L_HI(net2306));
 sg13g2_tiehi _21428__2307 (.L_HI(net2307));
 sg13g2_tiehi _21427__2308 (.L_HI(net2308));
 sg13g2_tiehi _21426__2309 (.L_HI(net2309));
 sg13g2_tiehi _21425__2310 (.L_HI(net2310));
 sg13g2_tiehi _21424__2311 (.L_HI(net2311));
 sg13g2_tiehi _21423__2312 (.L_HI(net2312));
 sg13g2_tiehi _21422__2313 (.L_HI(net2313));
 sg13g2_tiehi _21421__2314 (.L_HI(net2314));
 sg13g2_tiehi _21420__2315 (.L_HI(net2315));
 sg13g2_tiehi _21419__2316 (.L_HI(net2316));
 sg13g2_tiehi _21418__2317 (.L_HI(net2317));
 sg13g2_tiehi _21417__2318 (.L_HI(net2318));
 sg13g2_tiehi _21416__2319 (.L_HI(net2319));
 sg13g2_tiehi _21415__2320 (.L_HI(net2320));
 sg13g2_tiehi _21414__2321 (.L_HI(net2321));
 sg13g2_tiehi _21413__2322 (.L_HI(net2322));
 sg13g2_tiehi _21412__2323 (.L_HI(net2323));
 sg13g2_tiehi _21411__2324 (.L_HI(net2324));
 sg13g2_tiehi _21410__2325 (.L_HI(net2325));
 sg13g2_tiehi _21409__2326 (.L_HI(net2326));
 sg13g2_tiehi _21408__2327 (.L_HI(net2327));
 sg13g2_tiehi _21407__2328 (.L_HI(net2328));
 sg13g2_tiehi _21406__2329 (.L_HI(net2329));
 sg13g2_tiehi _21405__2330 (.L_HI(net2330));
 sg13g2_tiehi _21404__2331 (.L_HI(net2331));
 sg13g2_tiehi _21403__2332 (.L_HI(net2332));
 sg13g2_tiehi _21402__2333 (.L_HI(net2333));
 sg13g2_tiehi _21401__2334 (.L_HI(net2334));
 sg13g2_tiehi _21400__2335 (.L_HI(net2335));
 sg13g2_tiehi _21399__2336 (.L_HI(net2336));
 sg13g2_tiehi _21398__2337 (.L_HI(net2337));
 sg13g2_tiehi _21397__2338 (.L_HI(net2338));
 sg13g2_tiehi _21396__2339 (.L_HI(net2339));
 sg13g2_tiehi _21395__2340 (.L_HI(net2340));
 sg13g2_tiehi _21394__2341 (.L_HI(net2341));
 sg13g2_tiehi _21393__2342 (.L_HI(net2342));
 sg13g2_tiehi _21392__2343 (.L_HI(net2343));
 sg13g2_tiehi _21391__2344 (.L_HI(net2344));
 sg13g2_tiehi _21390__2345 (.L_HI(net2345));
 sg13g2_tiehi _21389__2346 (.L_HI(net2346));
 sg13g2_tiehi _21388__2347 (.L_HI(net2347));
 sg13g2_tiehi _21387__2348 (.L_HI(net2348));
 sg13g2_tiehi _21386__2349 (.L_HI(net2349));
 sg13g2_tiehi _21385__2350 (.L_HI(net2350));
 sg13g2_tiehi _21384__2351 (.L_HI(net2351));
 sg13g2_tiehi _21383__2352 (.L_HI(net2352));
 sg13g2_tiehi _21382__2353 (.L_HI(net2353));
 sg13g2_tiehi _21381__2354 (.L_HI(net2354));
 sg13g2_tiehi _21380__2355 (.L_HI(net2355));
 sg13g2_tiehi _21379__2356 (.L_HI(net2356));
 sg13g2_tiehi _21378__2357 (.L_HI(net2357));
 sg13g2_tiehi _21377__2358 (.L_HI(net2358));
 sg13g2_tiehi _21376__2359 (.L_HI(net2359));
 sg13g2_tiehi _21375__2360 (.L_HI(net2360));
 sg13g2_tiehi _21374__2361 (.L_HI(net2361));
 sg13g2_tiehi _21373__2362 (.L_HI(net2362));
 sg13g2_tiehi _21372__2363 (.L_HI(net2363));
 sg13g2_tiehi _21371__2364 (.L_HI(net2364));
 sg13g2_tiehi _21370__2365 (.L_HI(net2365));
 sg13g2_tiehi _21369__2366 (.L_HI(net2366));
 sg13g2_tiehi _21368__2367 (.L_HI(net2367));
 sg13g2_tiehi _21367__2368 (.L_HI(net2368));
 sg13g2_tiehi _21366__2369 (.L_HI(net2369));
 sg13g2_tiehi _21365__2370 (.L_HI(net2370));
 sg13g2_tiehi _21364__2371 (.L_HI(net2371));
 sg13g2_tiehi _21363__2372 (.L_HI(net2372));
 sg13g2_tiehi _21362__2373 (.L_HI(net2373));
 sg13g2_tiehi _21361__2374 (.L_HI(net2374));
 sg13g2_tiehi _21360__2375 (.L_HI(net2375));
 sg13g2_tiehi _21359__2376 (.L_HI(net2376));
 sg13g2_tiehi _21358__2377 (.L_HI(net2377));
 sg13g2_tiehi _21357__2378 (.L_HI(net2378));
 sg13g2_tiehi _21356__2379 (.L_HI(net2379));
 sg13g2_tiehi _21355__2380 (.L_HI(net2380));
 sg13g2_tiehi _21354__2381 (.L_HI(net2381));
 sg13g2_tiehi _21353__2382 (.L_HI(net2382));
 sg13g2_tiehi _21352__2383 (.L_HI(net2383));
 sg13g2_tiehi _21351__2384 (.L_HI(net2384));
 sg13g2_tiehi _21350__2385 (.L_HI(net2385));
 sg13g2_tiehi _21349__2386 (.L_HI(net2386));
 sg13g2_tiehi _21348__2387 (.L_HI(net2387));
 sg13g2_tiehi _21347__2388 (.L_HI(net2388));
 sg13g2_tiehi _21346__2389 (.L_HI(net2389));
 sg13g2_tiehi _21345__2390 (.L_HI(net2390));
 sg13g2_tiehi _21344__2391 (.L_HI(net2391));
 sg13g2_tiehi _21343__2392 (.L_HI(net2392));
 sg13g2_tiehi _21342__2393 (.L_HI(net2393));
 sg13g2_tiehi _21341__2394 (.L_HI(net2394));
 sg13g2_tiehi _21340__2395 (.L_HI(net2395));
 sg13g2_tiehi _21339__2396 (.L_HI(net2396));
 sg13g2_tiehi _21338__2397 (.L_HI(net2397));
 sg13g2_tiehi _21337__2398 (.L_HI(net2398));
 sg13g2_tiehi _21336__2399 (.L_HI(net2399));
 sg13g2_tiehi _21335__2400 (.L_HI(net2400));
 sg13g2_tiehi _21334__2401 (.L_HI(net2401));
 sg13g2_tiehi _21333__2402 (.L_HI(net2402));
 sg13g2_tiehi _21332__2403 (.L_HI(net2403));
 sg13g2_tiehi _21331__2404 (.L_HI(net2404));
 sg13g2_tiehi _21330__2405 (.L_HI(net2405));
 sg13g2_tiehi _21329__2406 (.L_HI(net2406));
 sg13g2_tiehi _21328__2407 (.L_HI(net2407));
 sg13g2_tiehi _21327__2408 (.L_HI(net2408));
 sg13g2_tiehi _21326__2409 (.L_HI(net2409));
 sg13g2_tiehi _21325__2410 (.L_HI(net2410));
 sg13g2_tiehi _21324__2411 (.L_HI(net2411));
 sg13g2_tiehi _21323__2412 (.L_HI(net2412));
 sg13g2_tiehi _21322__2413 (.L_HI(net2413));
 sg13g2_tiehi _21321__2414 (.L_HI(net2414));
 sg13g2_tiehi _21320__2415 (.L_HI(net2415));
 sg13g2_tiehi _21319__2416 (.L_HI(net2416));
 sg13g2_tiehi _21318__2417 (.L_HI(net2417));
 sg13g2_tiehi _21317__2418 (.L_HI(net2418));
 sg13g2_tiehi _21316__2419 (.L_HI(net2419));
 sg13g2_tiehi _21315__2420 (.L_HI(net2420));
 sg13g2_tiehi _21314__2421 (.L_HI(net2421));
 sg13g2_tiehi _21313__2422 (.L_HI(net2422));
 sg13g2_tiehi _21312__2423 (.L_HI(net2423));
 sg13g2_tiehi _21311__2424 (.L_HI(net2424));
 sg13g2_tiehi _21310__2425 (.L_HI(net2425));
 sg13g2_tiehi _21309__2426 (.L_HI(net2426));
 sg13g2_tiehi _21308__2427 (.L_HI(net2427));
 sg13g2_tiehi _21307__2428 (.L_HI(net2428));
 sg13g2_tiehi _21306__2429 (.L_HI(net2429));
 sg13g2_tiehi _21305__2430 (.L_HI(net2430));
 sg13g2_tiehi _21304__2431 (.L_HI(net2431));
 sg13g2_tiehi _21303__2432 (.L_HI(net2432));
 sg13g2_tiehi _21302__2433 (.L_HI(net2433));
 sg13g2_tiehi _21301__2434 (.L_HI(net2434));
 sg13g2_tiehi _21300__2435 (.L_HI(net2435));
 sg13g2_tiehi _21299__2436 (.L_HI(net2436));
 sg13g2_tiehi _21298__2437 (.L_HI(net2437));
 sg13g2_tiehi _21297__2438 (.L_HI(net2438));
 sg13g2_buf_2 \clkbuf_leaf_0_top1.acquisition_clk  (.A(\clknet_6_0_0_top1.acquisition_clk ),
    .X(\clknet_leaf_0_top1.acquisition_clk ));
 sg13g2_tielo tt_um_Coline3003_spect_top_18 (.L_LO(net18));
 sg13g2_tielo tt_um_Coline3003_spect_top_19 (.L_LO(net19));
 sg13g2_tielo tt_um_Coline3003_spect_top_20 (.L_LO(net20));
 sg13g2_tielo tt_um_Coline3003_spect_top_21 (.L_LO(net21));
 sg13g2_tielo tt_um_Coline3003_spect_top_22 (.L_LO(net22));
 sg13g2_tielo tt_um_Coline3003_spect_top_23 (.L_LO(net23));
 sg13g2_tielo tt_um_Coline3003_spect_top_24 (.L_LO(net24));
 sg13g2_tielo tt_um_Coline3003_spect_top_25 (.L_LO(net25));
 sg13g2_tielo tt_um_Coline3003_spect_top_26 (.L_LO(net26));
 sg13g2_tielo tt_um_Coline3003_spect_top_27 (.L_LO(net27));
 sg13g2_tielo tt_um_Coline3003_spect_top_28 (.L_LO(net28));
 sg13g2_tielo tt_um_Coline3003_spect_top_29 (.L_LO(net29));
 sg13g2_tielo tt_um_Coline3003_spect_top_30 (.L_LO(net30));
 sg13g2_tielo tt_um_Coline3003_spect_top_31 (.L_LO(net31));
 sg13g2_tielo tt_um_Coline3003_spect_top_32 (.L_LO(net32));
 sg13g2_tiehi _21296__33 (.L_HI(net33));
 sg13g2_buf_4 _24853_ (.X(uo_out[0]),
    .A(\top1.mux.data_out ));
 sg13g2_buf_2 _24854_ (.A(\top1.reg2.serial_out ),
    .X(uo_out[1]));
 sg13g2_buf_2 _24855_ (.A(net5826),
    .X(uo_out[2]));
 sg13g2_buf_8 _24856_ (.A(net5823),
    .X(uo_out[3]));
 sg13g2_buf_2 _24857_ (.A(net7567),
    .X(uo_out[4]));
 sg13g2_buf_4 _24858_ (.X(uo_out[5]),
    .A(net7560));
 sg13g2_buf_4 _24859_ (.X(uo_out[6]),
    .A(\top1.fsm.serial_readout ));
 sg13g2_buf_4 _24860_ (.X(uo_out[7]),
    .A(\top1.fsm.sending_data ));
 sg13g2_buf_2 fanout5822 (.A(net5823),
    .X(net5822));
 sg13g2_buf_4 fanout5823 (.X(net5823),
    .A(\top1.SL_ch ));
 sg13g2_buf_4 fanout5824 (.X(net5824),
    .A(_07321_));
 sg13g2_buf_4 fanout5825 (.X(net5825),
    .A(net5826));
 sg13g2_buf_4 fanout5826 (.X(net5826),
    .A(net5830));
 sg13g2_buf_4 fanout5827 (.X(net5827),
    .A(net5828));
 sg13g2_buf_2 fanout5828 (.A(net5829),
    .X(net5828));
 sg13g2_buf_2 fanout5829 (.A(net5830),
    .X(net5829));
 sg13g2_buf_2 fanout5830 (.A(\top1.SL_time ),
    .X(net5830));
 sg13g2_buf_4 fanout5831 (.X(net5831),
    .A(_05515_));
 sg13g2_buf_4 fanout5832 (.X(net5832),
    .A(net5833));
 sg13g2_buf_2 fanout5833 (.A(net5834),
    .X(net5833));
 sg13g2_buf_2 fanout5834 (.A(net5835),
    .X(net5834));
 sg13g2_buf_4 fanout5835 (.X(net5835),
    .A(_05444_));
 sg13g2_buf_8 fanout5836 (.A(_05444_),
    .X(net5836));
 sg13g2_buf_4 fanout5837 (.X(net5837),
    .A(_05453_));
 sg13g2_buf_4 fanout5838 (.X(net5838),
    .A(net5841));
 sg13g2_buf_2 fanout5839 (.A(net5841),
    .X(net5839));
 sg13g2_buf_4 fanout5840 (.X(net5840),
    .A(net5841));
 sg13g2_buf_4 fanout5841 (.X(net5841),
    .A(_05453_));
 sg13g2_buf_4 fanout5842 (.X(net5842),
    .A(net5844));
 sg13g2_buf_2 fanout5843 (.A(net5844),
    .X(net5843));
 sg13g2_buf_4 fanout5844 (.X(net5844),
    .A(net5846));
 sg13g2_buf_8 fanout5845 (.A(net5846),
    .X(net5845));
 sg13g2_buf_4 fanout5846 (.X(net5846),
    .A(net5849));
 sg13g2_buf_8 fanout5847 (.A(net5848),
    .X(net5847));
 sg13g2_buf_8 fanout5848 (.A(net5849),
    .X(net5848));
 sg13g2_buf_8 fanout5849 (.A(_05422_),
    .X(net5849));
 sg13g2_buf_4 fanout5850 (.X(net5850),
    .A(net5852));
 sg13g2_buf_4 fanout5851 (.X(net5851),
    .A(net5852));
 sg13g2_buf_8 fanout5852 (.A(net5866),
    .X(net5852));
 sg13g2_buf_4 fanout5853 (.X(net5853),
    .A(net5855));
 sg13g2_buf_4 fanout5854 (.X(net5854),
    .A(net5855));
 sg13g2_buf_4 fanout5855 (.X(net5855),
    .A(net5866));
 sg13g2_buf_4 fanout5856 (.X(net5856),
    .A(net5858));
 sg13g2_buf_4 fanout5857 (.X(net5857),
    .A(net5858));
 sg13g2_buf_8 fanout5858 (.A(net5866),
    .X(net5858));
 sg13g2_buf_4 fanout5859 (.X(net5859),
    .A(net5860));
 sg13g2_buf_4 fanout5860 (.X(net5860),
    .A(net5861));
 sg13g2_buf_4 fanout5861 (.X(net5861),
    .A(net5866));
 sg13g2_buf_4 fanout5862 (.X(net5862),
    .A(net5863));
 sg13g2_buf_2 fanout5863 (.A(net5865),
    .X(net5863));
 sg13g2_buf_4 fanout5864 (.X(net5864),
    .A(net5865));
 sg13g2_buf_2 fanout5865 (.A(net5866),
    .X(net5865));
 sg13g2_buf_8 fanout5866 (.A(_05421_),
    .X(net5866));
 sg13g2_buf_4 fanout5867 (.X(net5867),
    .A(net5868));
 sg13g2_buf_8 fanout5868 (.A(net5869),
    .X(net5868));
 sg13g2_buf_8 fanout5869 (.A(net5872),
    .X(net5869));
 sg13g2_buf_4 fanout5870 (.X(net5870),
    .A(net5871));
 sg13g2_buf_8 fanout5871 (.A(net5872),
    .X(net5871));
 sg13g2_buf_8 fanout5872 (.A(_05419_),
    .X(net5872));
 sg13g2_buf_4 fanout5873 (.X(net5873),
    .A(net5874));
 sg13g2_buf_4 fanout5874 (.X(net5874),
    .A(net5876));
 sg13g2_buf_4 fanout5875 (.X(net5875),
    .A(net5876));
 sg13g2_buf_2 fanout5876 (.A(_05418_),
    .X(net5876));
 sg13g2_buf_4 fanout5877 (.X(net5877),
    .A(net5879));
 sg13g2_buf_1 fanout5878 (.A(net5879),
    .X(net5878));
 sg13g2_buf_8 fanout5879 (.A(_05418_),
    .X(net5879));
 sg13g2_buf_4 fanout5880 (.X(net5880),
    .A(net5881));
 sg13g2_buf_4 fanout5881 (.X(net5881),
    .A(net5889));
 sg13g2_buf_4 fanout5882 (.X(net5882),
    .A(net5883));
 sg13g2_buf_8 fanout5883 (.A(net5889),
    .X(net5883));
 sg13g2_buf_4 fanout5884 (.X(net5884),
    .A(net5885));
 sg13g2_buf_4 fanout5885 (.X(net5885),
    .A(net5889));
 sg13g2_buf_4 fanout5886 (.X(net5886),
    .A(net5888));
 sg13g2_buf_2 fanout5887 (.A(net5888),
    .X(net5887));
 sg13g2_buf_4 fanout5888 (.X(net5888),
    .A(net5889));
 sg13g2_buf_8 fanout5889 (.A(_05418_),
    .X(net5889));
 sg13g2_buf_4 fanout5890 (.X(net5890),
    .A(net5893));
 sg13g2_buf_4 fanout5891 (.X(net5891),
    .A(net5892));
 sg13g2_buf_4 fanout5892 (.X(net5892),
    .A(net5893));
 sg13g2_buf_2 fanout5893 (.A(net5900),
    .X(net5893));
 sg13g2_buf_4 fanout5894 (.X(net5894),
    .A(net5895));
 sg13g2_buf_4 fanout5895 (.X(net5895),
    .A(net5896));
 sg13g2_buf_4 fanout5896 (.X(net5896),
    .A(net5900));
 sg13g2_buf_2 fanout5897 (.A(net5898),
    .X(net5897));
 sg13g2_buf_4 fanout5898 (.X(net5898),
    .A(net5899));
 sg13g2_buf_8 fanout5899 (.A(net5900),
    .X(net5899));
 sg13g2_buf_8 fanout5900 (.A(_05411_),
    .X(net5900));
 sg13g2_buf_4 fanout5901 (.X(net5901),
    .A(net5902));
 sg13g2_buf_4 fanout5902 (.X(net5902),
    .A(net5910));
 sg13g2_buf_4 fanout5903 (.X(net5903),
    .A(net5904));
 sg13g2_buf_4 fanout5904 (.X(net5904),
    .A(net5910));
 sg13g2_buf_4 fanout5905 (.X(net5905),
    .A(net5907));
 sg13g2_buf_2 fanout5906 (.A(net5907),
    .X(net5906));
 sg13g2_buf_4 fanout5907 (.X(net5907),
    .A(net5910));
 sg13g2_buf_4 fanout5908 (.X(net5908),
    .A(net5910));
 sg13g2_buf_2 fanout5909 (.A(net5910),
    .X(net5909));
 sg13g2_buf_4 fanout5910 (.X(net5910),
    .A(net5917));
 sg13g2_buf_4 fanout5911 (.X(net5911),
    .A(net5917));
 sg13g2_buf_4 fanout5912 (.X(net5912),
    .A(net5917));
 sg13g2_buf_4 fanout5913 (.X(net5913),
    .A(net5914));
 sg13g2_buf_4 fanout5914 (.X(net5914),
    .A(net5916));
 sg13g2_buf_4 fanout5915 (.X(net5915),
    .A(net5916));
 sg13g2_buf_2 fanout5916 (.A(net5917),
    .X(net5916));
 sg13g2_buf_4 fanout5917 (.X(net5917),
    .A(_05410_));
 sg13g2_buf_4 fanout5918 (.X(net5918),
    .A(net5920));
 sg13g2_buf_4 fanout5919 (.X(net5919),
    .A(net5920));
 sg13g2_buf_2 fanout5920 (.A(net5925),
    .X(net5920));
 sg13g2_buf_4 fanout5921 (.X(net5921),
    .A(net5922));
 sg13g2_buf_4 fanout5922 (.X(net5922),
    .A(net5925));
 sg13g2_buf_4 fanout5923 (.X(net5923),
    .A(net5924));
 sg13g2_buf_2 fanout5924 (.A(net5925),
    .X(net5924));
 sg13g2_buf_2 fanout5925 (.A(_05410_),
    .X(net5925));
 sg13g2_buf_4 fanout5926 (.X(net5926),
    .A(net5929));
 sg13g2_buf_4 fanout5927 (.X(net5927),
    .A(net5928));
 sg13g2_buf_4 fanout5928 (.X(net5928),
    .A(net5929));
 sg13g2_buf_8 fanout5929 (.A(_05410_),
    .X(net5929));
 sg13g2_buf_4 fanout5930 (.X(net5930),
    .A(net5931));
 sg13g2_buf_4 fanout5931 (.X(net5931),
    .A(net5932));
 sg13g2_buf_4 fanout5932 (.X(net5932),
    .A(net5941));
 sg13g2_buf_4 fanout5933 (.X(net5933),
    .A(net5936));
 sg13g2_buf_4 fanout5934 (.X(net5934),
    .A(net5936));
 sg13g2_buf_4 fanout5935 (.X(net5935),
    .A(net5936));
 sg13g2_buf_4 fanout5936 (.X(net5936),
    .A(net5941));
 sg13g2_buf_4 fanout5937 (.X(net5937),
    .A(net5938));
 sg13g2_buf_4 fanout5938 (.X(net5938),
    .A(net5939));
 sg13g2_buf_4 fanout5939 (.X(net5939),
    .A(net5940));
 sg13g2_buf_8 fanout5940 (.A(net5941),
    .X(net5940));
 sg13g2_buf_4 fanout5941 (.X(net5941),
    .A(_05409_));
 sg13g2_buf_4 fanout5942 (.X(net5942),
    .A(net5943));
 sg13g2_buf_4 fanout5943 (.X(net5943),
    .A(net5957));
 sg13g2_buf_4 fanout5944 (.X(net5944),
    .A(net5945));
 sg13g2_buf_4 fanout5945 (.X(net5945),
    .A(net5957));
 sg13g2_buf_4 fanout5946 (.X(net5946),
    .A(net5947));
 sg13g2_buf_4 fanout5947 (.X(net5947),
    .A(net5950));
 sg13g2_buf_4 fanout5948 (.X(net5948),
    .A(net5949));
 sg13g2_buf_4 fanout5949 (.X(net5949),
    .A(net5950));
 sg13g2_buf_2 fanout5950 (.A(net5957),
    .X(net5950));
 sg13g2_buf_4 fanout5951 (.X(net5951),
    .A(net5957));
 sg13g2_buf_4 fanout5952 (.X(net5952),
    .A(net5957));
 sg13g2_buf_4 fanout5953 (.X(net5953),
    .A(net5954));
 sg13g2_buf_2 fanout5954 (.A(net5956),
    .X(net5954));
 sg13g2_buf_4 fanout5955 (.X(net5955),
    .A(net5956));
 sg13g2_buf_2 fanout5956 (.A(net5957),
    .X(net5956));
 sg13g2_buf_8 fanout5957 (.A(_05408_),
    .X(net5957));
 sg13g2_buf_4 fanout5958 (.X(net5958),
    .A(net5960));
 sg13g2_buf_4 fanout5959 (.X(net5959),
    .A(net5960));
 sg13g2_buf_2 fanout5960 (.A(net5965),
    .X(net5960));
 sg13g2_buf_4 fanout5961 (.X(net5961),
    .A(net5962));
 sg13g2_buf_4 fanout5962 (.X(net5962),
    .A(net5965));
 sg13g2_buf_4 fanout5963 (.X(net5963),
    .A(net5964));
 sg13g2_buf_2 fanout5964 (.A(net5965),
    .X(net5964));
 sg13g2_buf_2 fanout5965 (.A(_05408_),
    .X(net5965));
 sg13g2_buf_4 fanout5966 (.X(net5966),
    .A(net5969));
 sg13g2_buf_4 fanout5967 (.X(net5967),
    .A(net5968));
 sg13g2_buf_4 fanout5968 (.X(net5968),
    .A(net5969));
 sg13g2_buf_8 fanout5969 (.A(_05408_),
    .X(net5969));
 sg13g2_buf_4 fanout5970 (.X(net5970),
    .A(net5971));
 sg13g2_buf_4 fanout5971 (.X(net5971),
    .A(net5972));
 sg13g2_buf_4 fanout5972 (.X(net5972),
    .A(net5976));
 sg13g2_buf_4 fanout5973 (.X(net5973),
    .A(net5974));
 sg13g2_buf_4 fanout5974 (.X(net5974),
    .A(net5975));
 sg13g2_buf_4 fanout5975 (.X(net5975),
    .A(net5976));
 sg13g2_buf_2 fanout5976 (.A(net5980),
    .X(net5976));
 sg13g2_buf_4 fanout5977 (.X(net5977),
    .A(net5978));
 sg13g2_buf_4 fanout5978 (.X(net5978),
    .A(net5979));
 sg13g2_buf_8 fanout5979 (.A(net5980),
    .X(net5979));
 sg13g2_buf_8 fanout5980 (.A(_05406_),
    .X(net5980));
 sg13g2_buf_4 fanout5981 (.X(net5981),
    .A(net5982));
 sg13g2_buf_4 fanout5982 (.X(net5982),
    .A(net5985));
 sg13g2_buf_4 fanout5983 (.X(net5983),
    .A(net5984));
 sg13g2_buf_4 fanout5984 (.X(net5984),
    .A(net5985));
 sg13g2_buf_4 fanout5985 (.X(net5985),
    .A(net5991));
 sg13g2_buf_4 fanout5986 (.X(net5986),
    .A(net5988));
 sg13g2_buf_2 fanout5987 (.A(net5988),
    .X(net5987));
 sg13g2_buf_2 fanout5988 (.A(net5991),
    .X(net5988));
 sg13g2_buf_4 fanout5989 (.X(net5989),
    .A(net5991));
 sg13g2_buf_2 fanout5990 (.A(net5991),
    .X(net5990));
 sg13g2_buf_2 fanout5991 (.A(_05405_),
    .X(net5991));
 sg13g2_buf_4 fanout5992 (.X(net5992),
    .A(net5993));
 sg13g2_buf_4 fanout5993 (.X(net5993),
    .A(net5998));
 sg13g2_buf_4 fanout5994 (.X(net5994),
    .A(net5997));
 sg13g2_buf_4 fanout5995 (.X(net5995),
    .A(net5996));
 sg13g2_buf_4 fanout5996 (.X(net5996),
    .A(net5997));
 sg13g2_buf_2 fanout5997 (.A(net5998),
    .X(net5997));
 sg13g2_buf_4 fanout5998 (.X(net5998),
    .A(_05405_));
 sg13g2_buf_4 fanout5999 (.X(net5999),
    .A(net6001));
 sg13g2_buf_4 fanout6000 (.X(net6000),
    .A(net6001));
 sg13g2_buf_2 fanout6001 (.A(net6010),
    .X(net6001));
 sg13g2_buf_4 fanout6002 (.X(net6002),
    .A(net6003));
 sg13g2_buf_2 fanout6003 (.A(net6010),
    .X(net6003));
 sg13g2_buf_4 fanout6004 (.X(net6004),
    .A(net6005));
 sg13g2_buf_2 fanout6005 (.A(net6010),
    .X(net6005));
 sg13g2_buf_4 fanout6006 (.X(net6006),
    .A(net6009));
 sg13g2_buf_4 fanout6007 (.X(net6007),
    .A(net6009));
 sg13g2_buf_4 fanout6008 (.X(net6008),
    .A(net6009));
 sg13g2_buf_4 fanout6009 (.X(net6009),
    .A(net6010));
 sg13g2_buf_4 fanout6010 (.X(net6010),
    .A(_05405_));
 sg13g2_buf_8 fanout6011 (.A(net6015),
    .X(net6011));
 sg13g2_buf_4 fanout6012 (.X(net6012),
    .A(net6014));
 sg13g2_buf_2 fanout6013 (.A(net6014),
    .X(net6013));
 sg13g2_buf_8 fanout6014 (.A(net6015),
    .X(net6014));
 sg13g2_buf_8 fanout6015 (.A(_05403_),
    .X(net6015));
 sg13g2_buf_4 fanout6016 (.X(net6016),
    .A(net6017));
 sg13g2_buf_2 fanout6017 (.A(net6018),
    .X(net6017));
 sg13g2_buf_2 fanout6018 (.A(net6024),
    .X(net6018));
 sg13g2_buf_4 fanout6019 (.X(net6019),
    .A(net6020));
 sg13g2_buf_4 fanout6020 (.X(net6020),
    .A(net6024));
 sg13g2_buf_4 fanout6021 (.X(net6021),
    .A(net6023));
 sg13g2_buf_2 fanout6022 (.A(net6023),
    .X(net6022));
 sg13g2_buf_8 fanout6023 (.A(net6024),
    .X(net6023));
 sg13g2_buf_4 fanout6024 (.X(net6024),
    .A(_05402_));
 sg13g2_buf_4 fanout6025 (.X(net6025),
    .A(net6026));
 sg13g2_buf_4 fanout6026 (.X(net6026),
    .A(net6029));
 sg13g2_buf_4 fanout6027 (.X(net6027),
    .A(net6029));
 sg13g2_buf_2 fanout6028 (.A(net6029),
    .X(net6028));
 sg13g2_buf_2 fanout6029 (.A(_05402_),
    .X(net6029));
 sg13g2_buf_4 fanout6030 (.X(net6030),
    .A(net6032));
 sg13g2_buf_4 fanout6031 (.X(net6031),
    .A(net6035));
 sg13g2_buf_2 fanout6032 (.A(net6035),
    .X(net6032));
 sg13g2_buf_4 fanout6033 (.X(net6033),
    .A(net6034));
 sg13g2_buf_4 fanout6034 (.X(net6034),
    .A(net6035));
 sg13g2_buf_4 fanout6035 (.X(net6035),
    .A(_05402_));
 sg13g2_buf_4 fanout6036 (.X(net6036),
    .A(net6038));
 sg13g2_buf_2 fanout6037 (.A(net6038),
    .X(net6037));
 sg13g2_buf_4 fanout6038 (.X(net6038),
    .A(net6042));
 sg13g2_buf_4 fanout6039 (.X(net6039),
    .A(net6040));
 sg13g2_buf_4 fanout6040 (.X(net6040),
    .A(net6041));
 sg13g2_buf_4 fanout6041 (.X(net6041),
    .A(net6042));
 sg13g2_buf_4 fanout6042 (.X(net6042),
    .A(_03984_));
 sg13g2_buf_4 fanout6043 (.X(net6043),
    .A(net6044));
 sg13g2_buf_4 fanout6044 (.X(net6044),
    .A(net6045));
 sg13g2_buf_8 fanout6045 (.A(_03984_),
    .X(net6045));
 sg13g2_buf_4 fanout6046 (.X(net6046),
    .A(net6047));
 sg13g2_buf_4 fanout6047 (.X(net6047),
    .A(net6049));
 sg13g2_buf_4 fanout6048 (.X(net6048),
    .A(net6049));
 sg13g2_buf_4 fanout6049 (.X(net6049),
    .A(net6055));
 sg13g2_buf_4 fanout6050 (.X(net6050),
    .A(net6051));
 sg13g2_buf_2 fanout6051 (.A(net6052),
    .X(net6051));
 sg13g2_buf_2 fanout6052 (.A(net6055),
    .X(net6052));
 sg13g2_buf_4 fanout6053 (.X(net6053),
    .A(net6055));
 sg13g2_buf_2 fanout6054 (.A(net6055),
    .X(net6054));
 sg13g2_buf_4 fanout6055 (.X(net6055),
    .A(net6074));
 sg13g2_buf_4 fanout6056 (.X(net6056),
    .A(net6062));
 sg13g2_buf_4 fanout6057 (.X(net6057),
    .A(net6062));
 sg13g2_buf_4 fanout6058 (.X(net6058),
    .A(net6059));
 sg13g2_buf_2 fanout6059 (.A(net6062),
    .X(net6059));
 sg13g2_buf_4 fanout6060 (.X(net6060),
    .A(net6061));
 sg13g2_buf_4 fanout6061 (.X(net6061),
    .A(net6062));
 sg13g2_buf_2 fanout6062 (.A(net6074),
    .X(net6062));
 sg13g2_buf_4 fanout6063 (.X(net6063),
    .A(net6064));
 sg13g2_buf_4 fanout6064 (.X(net6064),
    .A(net6069));
 sg13g2_buf_4 fanout6065 (.X(net6065),
    .A(net6068));
 sg13g2_buf_4 fanout6066 (.X(net6066),
    .A(net6067));
 sg13g2_buf_2 fanout6067 (.A(net6068),
    .X(net6067));
 sg13g2_buf_4 fanout6068 (.X(net6068),
    .A(net6069));
 sg13g2_buf_2 fanout6069 (.A(net6074),
    .X(net6069));
 sg13g2_buf_4 fanout6070 (.X(net6070),
    .A(net6073));
 sg13g2_buf_4 fanout6071 (.X(net6071),
    .A(net6073));
 sg13g2_buf_4 fanout6072 (.X(net6072),
    .A(net6073));
 sg13g2_buf_4 fanout6073 (.X(net6073),
    .A(net6074));
 sg13g2_buf_4 fanout6074 (.X(net6074),
    .A(_03983_));
 sg13g2_buf_4 fanout6075 (.X(net6075),
    .A(net6076));
 sg13g2_buf_8 fanout6076 (.A(net6079),
    .X(net6076));
 sg13g2_buf_8 fanout6077 (.A(net6079),
    .X(net6077));
 sg13g2_buf_2 fanout6078 (.A(net6079),
    .X(net6078));
 sg13g2_buf_4 fanout6079 (.X(net6079),
    .A(_03982_));
 sg13g2_buf_4 fanout6080 (.X(net6080),
    .A(net6081));
 sg13g2_buf_4 fanout6081 (.X(net6081),
    .A(net6082));
 sg13g2_buf_8 fanout6082 (.A(_03982_),
    .X(net6082));
 sg13g2_buf_4 fanout6083 (.X(net6083),
    .A(net6086));
 sg13g2_buf_8 fanout6084 (.A(net6086),
    .X(net6084));
 sg13g2_buf_2 fanout6085 (.A(net6086),
    .X(net6085));
 sg13g2_buf_4 fanout6086 (.X(net6086),
    .A(net6088));
 sg13g2_buf_8 fanout6087 (.A(net6088),
    .X(net6087));
 sg13g2_buf_4 fanout6088 (.X(net6088),
    .A(net6100));
 sg13g2_buf_8 fanout6089 (.A(net6090),
    .X(net6089));
 sg13g2_buf_4 fanout6090 (.X(net6090),
    .A(net6092));
 sg13g2_buf_4 fanout6091 (.X(net6091),
    .A(net6092));
 sg13g2_buf_2 fanout6092 (.A(net6100),
    .X(net6092));
 sg13g2_buf_4 fanout6093 (.X(net6093),
    .A(net6096));
 sg13g2_buf_4 fanout6094 (.X(net6094),
    .A(net6095));
 sg13g2_buf_4 fanout6095 (.X(net6095),
    .A(net6096));
 sg13g2_buf_2 fanout6096 (.A(net6100),
    .X(net6096));
 sg13g2_buf_4 fanout6097 (.X(net6097),
    .A(net6099));
 sg13g2_buf_2 fanout6098 (.A(net6099),
    .X(net6098));
 sg13g2_buf_4 fanout6099 (.X(net6099),
    .A(net6100));
 sg13g2_buf_8 fanout6100 (.A(_03981_),
    .X(net6100));
 sg13g2_buf_2 fanout6101 (.A(_03832_),
    .X(net6101));
 sg13g2_buf_8 fanout6102 (.A(_03830_),
    .X(net6102));
 sg13g2_buf_8 fanout6103 (.A(_03829_),
    .X(net6103));
 sg13g2_buf_4 fanout6104 (.X(net6104),
    .A(net6105));
 sg13g2_buf_8 fanout6105 (.A(net6107),
    .X(net6105));
 sg13g2_buf_8 fanout6106 (.A(net6107),
    .X(net6106));
 sg13g2_buf_8 fanout6107 (.A(_03828_),
    .X(net6107));
 sg13g2_buf_2 fanout6108 (.A(\top1.addr_out[8] ),
    .X(net6108));
 sg13g2_buf_1 fanout6109 (.A(\top1.addr_out[8] ),
    .X(net6109));
 sg13g2_buf_2 fanout6110 (.A(\top1.fsm.state_reg[0] ),
    .X(net6110));
 sg13g2_buf_4 fanout6111 (.X(net6111),
    .A(\top1.addr_out[7] ));
 sg13g2_buf_4 fanout6112 (.X(net6112),
    .A(\top1.addr_out[7] ));
 sg13g2_buf_4 fanout6113 (.X(net6113),
    .A(net6115));
 sg13g2_buf_2 fanout6114 (.A(net6115),
    .X(net6114));
 sg13g2_buf_2 fanout6115 (.A(net6116),
    .X(net6115));
 sg13g2_buf_8 fanout6116 (.A(\top1.addr_out[6] ),
    .X(net6116));
 sg13g2_buf_8 fanout6117 (.A(net6119),
    .X(net6117));
 sg13g2_buf_4 fanout6118 (.X(net6118),
    .A(net6119));
 sg13g2_buf_8 fanout6119 (.A(\top1.addr_out[5] ),
    .X(net6119));
 sg13g2_buf_4 fanout6120 (.X(net6120),
    .A(net6121));
 sg13g2_buf_4 fanout6121 (.X(net6121),
    .A(net6126));
 sg13g2_buf_8 fanout6122 (.A(net6123),
    .X(net6122));
 sg13g2_buf_2 fanout6123 (.A(net6126),
    .X(net6123));
 sg13g2_buf_8 fanout6124 (.A(net6126),
    .X(net6124));
 sg13g2_buf_2 fanout6125 (.A(net6126),
    .X(net6125));
 sg13g2_buf_8 fanout6126 (.A(\top1.addr_out[4] ),
    .X(net6126));
 sg13g2_buf_4 fanout6127 (.X(net6127),
    .A(\top1.addr_out[3] ));
 sg13g2_buf_2 fanout6128 (.A(net6129),
    .X(net6128));
 sg13g2_buf_2 fanout6129 (.A(net6130),
    .X(net6129));
 sg13g2_buf_2 fanout6130 (.A(net6132),
    .X(net6130));
 sg13g2_buf_4 fanout6131 (.X(net6131),
    .A(net6132));
 sg13g2_buf_2 fanout6132 (.A(\top1.addr_out[2] ),
    .X(net6132));
 sg13g2_buf_4 fanout6133 (.X(net6133),
    .A(net6134));
 sg13g2_buf_4 fanout6134 (.X(net6134),
    .A(net6135));
 sg13g2_buf_4 fanout6135 (.X(net6135),
    .A(net6143));
 sg13g2_buf_4 fanout6136 (.X(net6136),
    .A(net6137));
 sg13g2_buf_4 fanout6137 (.X(net6137),
    .A(net6138));
 sg13g2_buf_4 fanout6138 (.X(net6138),
    .A(net6143));
 sg13g2_buf_8 fanout6139 (.A(net6142),
    .X(net6139));
 sg13g2_buf_4 fanout6140 (.X(net6140),
    .A(net6142));
 sg13g2_buf_4 fanout6141 (.X(net6141),
    .A(net6142));
 sg13g2_buf_4 fanout6142 (.X(net6142),
    .A(net6143));
 sg13g2_buf_4 fanout6143 (.X(net6143),
    .A(net6154));
 sg13g2_buf_4 fanout6144 (.X(net6144),
    .A(net6145));
 sg13g2_buf_2 fanout6145 (.A(net6154),
    .X(net6145));
 sg13g2_buf_4 fanout6146 (.X(net6146),
    .A(net6148));
 sg13g2_buf_4 fanout6147 (.X(net6147),
    .A(net6148));
 sg13g2_buf_4 fanout6148 (.X(net6148),
    .A(net6149));
 sg13g2_buf_4 fanout6149 (.X(net6149),
    .A(net6154));
 sg13g2_buf_4 fanout6150 (.X(net6150),
    .A(net6153));
 sg13g2_buf_4 fanout6151 (.X(net6151),
    .A(net6152));
 sg13g2_buf_4 fanout6152 (.X(net6152),
    .A(net6153));
 sg13g2_buf_4 fanout6153 (.X(net6153),
    .A(net6154));
 sg13g2_buf_4 fanout6154 (.X(net6154),
    .A(\top1.addr_out[1] ));
 sg13g2_buf_4 fanout6155 (.X(net6155),
    .A(net6156));
 sg13g2_buf_4 fanout6156 (.X(net6156),
    .A(net6157));
 sg13g2_buf_4 fanout6157 (.X(net6157),
    .A(net6163));
 sg13g2_buf_4 fanout6158 (.X(net6158),
    .A(net6159));
 sg13g2_buf_4 fanout6159 (.X(net6159),
    .A(net6162));
 sg13g2_buf_4 fanout6160 (.X(net6160),
    .A(net6162));
 sg13g2_buf_4 fanout6161 (.X(net6161),
    .A(net6162));
 sg13g2_buf_4 fanout6162 (.X(net6162),
    .A(net6163));
 sg13g2_buf_2 fanout6163 (.A(net6196),
    .X(net6163));
 sg13g2_buf_4 fanout6164 (.X(net6164),
    .A(net6166));
 sg13g2_buf_4 fanout6165 (.X(net6165),
    .A(net6166));
 sg13g2_buf_4 fanout6166 (.X(net6166),
    .A(net6196));
 sg13g2_buf_4 fanout6167 (.X(net6167),
    .A(net6170));
 sg13g2_buf_2 fanout6168 (.A(net6170),
    .X(net6168));
 sg13g2_buf_4 fanout6169 (.X(net6169),
    .A(net6170));
 sg13g2_buf_2 fanout6170 (.A(net6196),
    .X(net6170));
 sg13g2_buf_4 fanout6171 (.X(net6171),
    .A(net6173));
 sg13g2_buf_4 fanout6172 (.X(net6172),
    .A(net6173));
 sg13g2_buf_4 fanout6173 (.X(net6173),
    .A(net6183));
 sg13g2_buf_4 fanout6174 (.X(net6174),
    .A(net6183));
 sg13g2_buf_4 fanout6175 (.X(net6175),
    .A(net6183));
 sg13g2_buf_4 fanout6176 (.X(net6176),
    .A(net6179));
 sg13g2_buf_2 fanout6177 (.A(net6179),
    .X(net6177));
 sg13g2_buf_4 fanout6178 (.X(net6178),
    .A(net6179));
 sg13g2_buf_2 fanout6179 (.A(net6182),
    .X(net6179));
 sg13g2_buf_4 fanout6180 (.X(net6180),
    .A(net6181));
 sg13g2_buf_4 fanout6181 (.X(net6181),
    .A(net6182));
 sg13g2_buf_4 fanout6182 (.X(net6182),
    .A(net6183));
 sg13g2_buf_2 fanout6183 (.A(net6196),
    .X(net6183));
 sg13g2_buf_4 fanout6184 (.X(net6184),
    .A(net6195));
 sg13g2_buf_4 fanout6185 (.X(net6185),
    .A(net6195));
 sg13g2_buf_4 fanout6186 (.X(net6186),
    .A(net6188));
 sg13g2_buf_4 fanout6187 (.X(net6187),
    .A(net6188));
 sg13g2_buf_4 fanout6188 (.X(net6188),
    .A(net6195));
 sg13g2_buf_4 fanout6189 (.X(net6189),
    .A(net6191));
 sg13g2_buf_4 fanout6190 (.X(net6190),
    .A(net6191));
 sg13g2_buf_2 fanout6191 (.A(net6194),
    .X(net6191));
 sg13g2_buf_4 fanout6192 (.X(net6192),
    .A(net6193));
 sg13g2_buf_4 fanout6193 (.X(net6193),
    .A(net6194));
 sg13g2_buf_2 fanout6194 (.A(net6195),
    .X(net6194));
 sg13g2_buf_2 fanout6195 (.A(net6196),
    .X(net6195));
 sg13g2_buf_4 fanout6196 (.X(net6196),
    .A(\top1.addr_out[1] ));
 sg13g2_buf_8 fanout6197 (.A(net6198),
    .X(net6197));
 sg13g2_buf_8 fanout6198 (.A(net6199),
    .X(net6198));
 sg13g2_buf_8 fanout6199 (.A(net6208),
    .X(net6199));
 sg13g2_buf_8 fanout6200 (.A(net6201),
    .X(net6200));
 sg13g2_buf_8 fanout6201 (.A(net6202),
    .X(net6201));
 sg13g2_buf_8 fanout6202 (.A(net6208),
    .X(net6202));
 sg13g2_buf_8 fanout6203 (.A(net6207),
    .X(net6203));
 sg13g2_buf_4 fanout6204 (.X(net6204),
    .A(net6207));
 sg13g2_buf_8 fanout6205 (.A(net6207),
    .X(net6205));
 sg13g2_buf_4 fanout6206 (.X(net6206),
    .A(net6207));
 sg13g2_buf_4 fanout6207 (.X(net6207),
    .A(net6208));
 sg13g2_buf_4 fanout6208 (.X(net6208),
    .A(net6219));
 sg13g2_buf_8 fanout6209 (.A(net6210),
    .X(net6209));
 sg13g2_buf_4 fanout6210 (.X(net6210),
    .A(net6219));
 sg13g2_buf_4 fanout6211 (.X(net6211),
    .A(net6213));
 sg13g2_buf_8 fanout6212 (.A(net6213),
    .X(net6212));
 sg13g2_buf_4 fanout6213 (.X(net6213),
    .A(net6214));
 sg13g2_buf_8 fanout6214 (.A(net6219),
    .X(net6214));
 sg13g2_buf_8 fanout6215 (.A(net6218),
    .X(net6215));
 sg13g2_buf_8 fanout6216 (.A(net6217),
    .X(net6216));
 sg13g2_buf_8 fanout6217 (.A(net6218),
    .X(net6217));
 sg13g2_buf_4 fanout6218 (.X(net6218),
    .A(net6219));
 sg13g2_buf_4 fanout6219 (.X(net6219),
    .A(\top1.addr_out[0] ));
 sg13g2_buf_8 fanout6220 (.A(net6221),
    .X(net6220));
 sg13g2_buf_8 fanout6221 (.A(net6222),
    .X(net6221));
 sg13g2_buf_8 fanout6222 (.A(net6228),
    .X(net6222));
 sg13g2_buf_8 fanout6223 (.A(net6224),
    .X(net6223));
 sg13g2_buf_8 fanout6224 (.A(net6227),
    .X(net6224));
 sg13g2_buf_8 fanout6225 (.A(net6227),
    .X(net6225));
 sg13g2_buf_4 fanout6226 (.X(net6226),
    .A(net6227));
 sg13g2_buf_8 fanout6227 (.A(net6228),
    .X(net6227));
 sg13g2_buf_2 fanout6228 (.A(net6261),
    .X(net6228));
 sg13g2_buf_8 fanout6229 (.A(net6231),
    .X(net6229));
 sg13g2_buf_8 fanout6230 (.A(net6231),
    .X(net6230));
 sg13g2_buf_8 fanout6231 (.A(net6261),
    .X(net6231));
 sg13g2_buf_8 fanout6232 (.A(net6235),
    .X(net6232));
 sg13g2_buf_4 fanout6233 (.X(net6233),
    .A(net6235));
 sg13g2_buf_8 fanout6234 (.A(net6235),
    .X(net6234));
 sg13g2_buf_4 fanout6235 (.X(net6235),
    .A(net6261));
 sg13g2_buf_8 fanout6236 (.A(net6238),
    .X(net6236));
 sg13g2_buf_8 fanout6237 (.A(net6238),
    .X(net6237));
 sg13g2_buf_8 fanout6238 (.A(net6248),
    .X(net6238));
 sg13g2_buf_8 fanout6239 (.A(net6248),
    .X(net6239));
 sg13g2_buf_8 fanout6240 (.A(net6248),
    .X(net6240));
 sg13g2_buf_8 fanout6241 (.A(net6244),
    .X(net6241));
 sg13g2_buf_4 fanout6242 (.X(net6242),
    .A(net6244));
 sg13g2_buf_8 fanout6243 (.A(net6244),
    .X(net6243));
 sg13g2_buf_4 fanout6244 (.X(net6244),
    .A(net6247));
 sg13g2_buf_8 fanout6245 (.A(net6246),
    .X(net6245));
 sg13g2_buf_8 fanout6246 (.A(net6247),
    .X(net6246));
 sg13g2_buf_4 fanout6247 (.X(net6247),
    .A(net6248));
 sg13g2_buf_2 fanout6248 (.A(net6261),
    .X(net6248));
 sg13g2_buf_8 fanout6249 (.A(net6260),
    .X(net6249));
 sg13g2_buf_8 fanout6250 (.A(net6260),
    .X(net6250));
 sg13g2_buf_8 fanout6251 (.A(net6253),
    .X(net6251));
 sg13g2_buf_8 fanout6252 (.A(net6253),
    .X(net6252));
 sg13g2_buf_8 fanout6253 (.A(net6260),
    .X(net6253));
 sg13g2_buf_8 fanout6254 (.A(net6256),
    .X(net6254));
 sg13g2_buf_8 fanout6255 (.A(net6256),
    .X(net6255));
 sg13g2_buf_4 fanout6256 (.X(net6256),
    .A(net6259));
 sg13g2_buf_8 fanout6257 (.A(net6258),
    .X(net6257));
 sg13g2_buf_8 fanout6258 (.A(net6259),
    .X(net6258));
 sg13g2_buf_4 fanout6259 (.X(net6259),
    .A(net6260));
 sg13g2_buf_4 fanout6260 (.X(net6260),
    .A(net6261));
 sg13g2_buf_8 fanout6261 (.A(\top1.addr_out[0] ),
    .X(net6261));
 sg13g2_buf_2 fanout6262 (.A(_02611_),
    .X(net6262));
 sg13g2_buf_2 fanout6263 (.A(_02611_),
    .X(net6263));
 sg13g2_buf_2 fanout6264 (.A(_02603_),
    .X(net6264));
 sg13g2_buf_1 fanout6265 (.A(_02603_),
    .X(net6265));
 sg13g2_buf_2 fanout6266 (.A(_02579_),
    .X(net6266));
 sg13g2_buf_1 fanout6267 (.A(_02579_),
    .X(net6267));
 sg13g2_buf_2 fanout6268 (.A(_02564_),
    .X(net6268));
 sg13g2_buf_1 fanout6269 (.A(_02564_),
    .X(net6269));
 sg13g2_buf_2 fanout6270 (.A(_02556_),
    .X(net6270));
 sg13g2_buf_1 fanout6271 (.A(_02556_),
    .X(net6271));
 sg13g2_buf_2 fanout6272 (.A(_07454_),
    .X(net6272));
 sg13g2_buf_2 fanout6273 (.A(_07454_),
    .X(net6273));
 sg13g2_buf_2 fanout6274 (.A(_07450_),
    .X(net6274));
 sg13g2_buf_1 fanout6275 (.A(_07450_),
    .X(net6275));
 sg13g2_buf_2 fanout6276 (.A(_07402_),
    .X(net6276));
 sg13g2_buf_1 fanout6277 (.A(_07402_),
    .X(net6277));
 sg13g2_buf_2 fanout6278 (.A(_07398_),
    .X(net6278));
 sg13g2_buf_1 fanout6279 (.A(_07398_),
    .X(net6279));
 sg13g2_buf_2 fanout6280 (.A(_07394_),
    .X(net6280));
 sg13g2_buf_1 fanout6281 (.A(_07394_),
    .X(net6281));
 sg13g2_buf_2 fanout6282 (.A(_07390_),
    .X(net6282));
 sg13g2_buf_1 fanout6283 (.A(_07390_),
    .X(net6283));
 sg13g2_buf_2 fanout6284 (.A(_07382_),
    .X(net6284));
 sg13g2_buf_1 fanout6285 (.A(_07382_),
    .X(net6285));
 sg13g2_buf_2 fanout6286 (.A(_07374_),
    .X(net6286));
 sg13g2_buf_1 fanout6287 (.A(_07374_),
    .X(net6287));
 sg13g2_buf_2 fanout6288 (.A(_07370_),
    .X(net6288));
 sg13g2_buf_1 fanout6289 (.A(_07370_),
    .X(net6289));
 sg13g2_buf_2 fanout6290 (.A(_07366_),
    .X(net6290));
 sg13g2_buf_1 fanout6291 (.A(_07366_),
    .X(net6291));
 sg13g2_buf_2 fanout6292 (.A(_07354_),
    .X(net6292));
 sg13g2_buf_1 fanout6293 (.A(_07354_),
    .X(net6293));
 sg13g2_buf_2 fanout6294 (.A(_07350_),
    .X(net6294));
 sg13g2_buf_1 fanout6295 (.A(_07350_),
    .X(net6295));
 sg13g2_buf_2 fanout6296 (.A(_07346_),
    .X(net6296));
 sg13g2_buf_1 fanout6297 (.A(_07346_),
    .X(net6297));
 sg13g2_buf_2 fanout6298 (.A(_07342_),
    .X(net6298));
 sg13g2_buf_1 fanout6299 (.A(_07342_),
    .X(net6299));
 sg13g2_buf_2 fanout6300 (.A(_07314_),
    .X(net6300));
 sg13g2_buf_2 fanout6301 (.A(_07314_),
    .X(net6301));
 sg13g2_buf_4 fanout6302 (.X(net6302),
    .A(_07310_));
 sg13g2_buf_1 fanout6303 (.A(_07310_),
    .X(net6303));
 sg13g2_buf_2 fanout6304 (.A(_07306_),
    .X(net6304));
 sg13g2_buf_1 fanout6305 (.A(_07306_),
    .X(net6305));
 sg13g2_buf_4 fanout6306 (.X(net6306),
    .A(_07267_));
 sg13g2_buf_1 fanout6307 (.A(_07267_),
    .X(net6307));
 sg13g2_buf_2 fanout6308 (.A(_07263_),
    .X(net6308));
 sg13g2_buf_1 fanout6309 (.A(_07263_),
    .X(net6309));
 sg13g2_buf_4 fanout6310 (.X(net6310),
    .A(_07259_));
 sg13g2_buf_1 fanout6311 (.A(_07259_),
    .X(net6311));
 sg13g2_buf_2 fanout6312 (.A(_07255_),
    .X(net6312));
 sg13g2_buf_1 fanout6313 (.A(_07255_),
    .X(net6313));
 sg13g2_buf_2 fanout6314 (.A(_07251_),
    .X(net6314));
 sg13g2_buf_1 fanout6315 (.A(_07251_),
    .X(net6315));
 sg13g2_buf_2 fanout6316 (.A(_07247_),
    .X(net6316));
 sg13g2_buf_1 fanout6317 (.A(_07247_),
    .X(net6317));
 sg13g2_buf_2 fanout6318 (.A(_07243_),
    .X(net6318));
 sg13g2_buf_1 fanout6319 (.A(_07243_),
    .X(net6319));
 sg13g2_buf_2 fanout6320 (.A(_07239_),
    .X(net6320));
 sg13g2_buf_1 fanout6321 (.A(_07239_),
    .X(net6321));
 sg13g2_buf_2 fanout6322 (.A(_07235_),
    .X(net6322));
 sg13g2_buf_1 fanout6323 (.A(_07235_),
    .X(net6323));
 sg13g2_buf_2 fanout6324 (.A(_07231_),
    .X(net6324));
 sg13g2_buf_1 fanout6325 (.A(_07231_),
    .X(net6325));
 sg13g2_buf_2 fanout6326 (.A(_07227_),
    .X(net6326));
 sg13g2_buf_1 fanout6327 (.A(_07227_),
    .X(net6327));
 sg13g2_buf_2 fanout6328 (.A(_07223_),
    .X(net6328));
 sg13g2_buf_1 fanout6329 (.A(_07223_),
    .X(net6329));
 sg13g2_buf_2 fanout6330 (.A(_07215_),
    .X(net6330));
 sg13g2_buf_1 fanout6331 (.A(_07215_),
    .X(net6331));
 sg13g2_buf_2 fanout6332 (.A(_07211_),
    .X(net6332));
 sg13g2_buf_1 fanout6333 (.A(_07211_),
    .X(net6333));
 sg13g2_buf_2 fanout6334 (.A(_07207_),
    .X(net6334));
 sg13g2_buf_1 fanout6335 (.A(_07207_),
    .X(net6335));
 sg13g2_buf_2 fanout6336 (.A(_07203_),
    .X(net6336));
 sg13g2_buf_1 fanout6337 (.A(_07203_),
    .X(net6337));
 sg13g2_buf_4 fanout6338 (.X(net6338),
    .A(_07198_));
 sg13g2_buf_1 fanout6339 (.A(_07198_),
    .X(net6339));
 sg13g2_buf_2 fanout6340 (.A(_07194_),
    .X(net6340));
 sg13g2_buf_1 fanout6341 (.A(_07194_),
    .X(net6341));
 sg13g2_buf_2 fanout6342 (.A(_07190_),
    .X(net6342));
 sg13g2_buf_1 fanout6343 (.A(_07190_),
    .X(net6343));
 sg13g2_buf_2 fanout6344 (.A(_07182_),
    .X(net6344));
 sg13g2_buf_1 fanout6345 (.A(_07182_),
    .X(net6345));
 sg13g2_buf_2 fanout6346 (.A(_07178_),
    .X(net6346));
 sg13g2_buf_1 fanout6347 (.A(_07178_),
    .X(net6347));
 sg13g2_buf_2 fanout6348 (.A(_07174_),
    .X(net6348));
 sg13g2_buf_1 fanout6349 (.A(_07174_),
    .X(net6349));
 sg13g2_buf_4 fanout6350 (.X(net6350),
    .A(_07170_));
 sg13g2_buf_2 fanout6351 (.A(_07170_),
    .X(net6351));
 sg13g2_buf_2 fanout6352 (.A(_06307_),
    .X(net6352));
 sg13g2_buf_1 fanout6353 (.A(_06307_),
    .X(net6353));
 sg13g2_buf_2 fanout6354 (.A(_06303_),
    .X(net6354));
 sg13g2_buf_1 fanout6355 (.A(_06303_),
    .X(net6355));
 sg13g2_buf_2 fanout6356 (.A(_06295_),
    .X(net6356));
 sg13g2_buf_1 fanout6357 (.A(_06295_),
    .X(net6357));
 sg13g2_buf_4 fanout6358 (.X(net6358),
    .A(_06287_));
 sg13g2_buf_2 fanout6359 (.A(_06287_),
    .X(net6359));
 sg13g2_buf_2 fanout6360 (.A(_06283_),
    .X(net6360));
 sg13g2_buf_2 fanout6361 (.A(_06283_),
    .X(net6361));
 sg13g2_buf_2 fanout6362 (.A(_05386_),
    .X(net6362));
 sg13g2_buf_1 fanout6363 (.A(_05386_),
    .X(net6363));
 sg13g2_buf_2 fanout6364 (.A(_05382_),
    .X(net6364));
 sg13g2_buf_1 fanout6365 (.A(_05382_),
    .X(net6365));
 sg13g2_buf_2 fanout6366 (.A(_05378_),
    .X(net6366));
 sg13g2_buf_1 fanout6367 (.A(_05378_),
    .X(net6367));
 sg13g2_buf_4 fanout6368 (.X(net6368),
    .A(_05370_));
 sg13g2_buf_1 fanout6369 (.A(_05370_),
    .X(net6369));
 sg13g2_buf_4 fanout6370 (.X(net6370),
    .A(_05366_));
 sg13g2_buf_2 fanout6371 (.A(_05366_),
    .X(net6371));
 sg13g2_buf_4 fanout6372 (.X(net6372),
    .A(_05362_));
 sg13g2_buf_2 fanout6373 (.A(_05362_),
    .X(net6373));
 sg13g2_buf_4 fanout6374 (.X(net6374),
    .A(_05354_));
 sg13g2_buf_1 fanout6375 (.A(_05354_),
    .X(net6375));
 sg13g2_buf_2 fanout6376 (.A(_05350_),
    .X(net6376));
 sg13g2_buf_2 fanout6377 (.A(_05350_),
    .X(net6377));
 sg13g2_buf_2 fanout6378 (.A(_05346_),
    .X(net6378));
 sg13g2_buf_1 fanout6379 (.A(_05346_),
    .X(net6379));
 sg13g2_buf_2 fanout6380 (.A(_05342_),
    .X(net6380));
 sg13g2_buf_1 fanout6381 (.A(_05342_),
    .X(net6381));
 sg13g2_buf_2 fanout6382 (.A(_05338_),
    .X(net6382));
 sg13g2_buf_1 fanout6383 (.A(_05338_),
    .X(net6383));
 sg13g2_buf_2 fanout6384 (.A(_05334_),
    .X(net6384));
 sg13g2_buf_1 fanout6385 (.A(_05334_),
    .X(net6385));
 sg13g2_buf_2 fanout6386 (.A(_05326_),
    .X(net6386));
 sg13g2_buf_1 fanout6387 (.A(_05326_),
    .X(net6387));
 sg13g2_buf_2 fanout6388 (.A(_05314_),
    .X(net6388));
 sg13g2_buf_2 fanout6389 (.A(_05314_),
    .X(net6389));
 sg13g2_buf_2 fanout6390 (.A(_05290_),
    .X(net6390));
 sg13g2_buf_1 fanout6391 (.A(_05290_),
    .X(net6391));
 sg13g2_buf_2 fanout6392 (.A(_05286_),
    .X(net6392));
 sg13g2_buf_1 fanout6393 (.A(_05286_),
    .X(net6393));
 sg13g2_buf_2 fanout6394 (.A(_05282_),
    .X(net6394));
 sg13g2_buf_1 fanout6395 (.A(_05282_),
    .X(net6395));
 sg13g2_buf_2 fanout6396 (.A(_05278_),
    .X(net6396));
 sg13g2_buf_1 fanout6397 (.A(_05278_),
    .X(net6397));
 sg13g2_buf_2 fanout6398 (.A(_05274_),
    .X(net6398));
 sg13g2_buf_1 fanout6399 (.A(_05274_),
    .X(net6399));
 sg13g2_buf_2 fanout6400 (.A(_05270_),
    .X(net6400));
 sg13g2_buf_1 fanout6401 (.A(_05270_),
    .X(net6401));
 sg13g2_buf_2 fanout6402 (.A(_05266_),
    .X(net6402));
 sg13g2_buf_1 fanout6403 (.A(_05266_),
    .X(net6403));
 sg13g2_buf_2 fanout6404 (.A(_05258_),
    .X(net6404));
 sg13g2_buf_1 fanout6405 (.A(_05258_),
    .X(net6405));
 sg13g2_buf_2 fanout6406 (.A(_05254_),
    .X(net6406));
 sg13g2_buf_1 fanout6407 (.A(_05254_),
    .X(net6407));
 sg13g2_buf_2 fanout6408 (.A(_05234_),
    .X(net6408));
 sg13g2_buf_1 fanout6409 (.A(_05234_),
    .X(net6409));
 sg13g2_buf_2 fanout6410 (.A(_05230_),
    .X(net6410));
 sg13g2_buf_1 fanout6411 (.A(_05230_),
    .X(net6411));
 sg13g2_buf_2 fanout6412 (.A(_05226_),
    .X(net6412));
 sg13g2_buf_1 fanout6413 (.A(_05226_),
    .X(net6413));
 sg13g2_buf_2 fanout6414 (.A(_05218_),
    .X(net6414));
 sg13g2_buf_1 fanout6415 (.A(_05218_),
    .X(net6415));
 sg13g2_buf_2 fanout6416 (.A(_05214_),
    .X(net6416));
 sg13g2_buf_1 fanout6417 (.A(_05214_),
    .X(net6417));
 sg13g2_buf_2 fanout6418 (.A(_05206_),
    .X(net6418));
 sg13g2_buf_1 fanout6419 (.A(_05206_),
    .X(net6419));
 sg13g2_buf_2 fanout6420 (.A(_05202_),
    .X(net6420));
 sg13g2_buf_1 fanout6421 (.A(_05202_),
    .X(net6421));
 sg13g2_buf_2 fanout6422 (.A(_05194_),
    .X(net6422));
 sg13g2_buf_1 fanout6423 (.A(_05194_),
    .X(net6423));
 sg13g2_buf_2 fanout6424 (.A(_05190_),
    .X(net6424));
 sg13g2_buf_1 fanout6425 (.A(_05190_),
    .X(net6425));
 sg13g2_buf_2 fanout6426 (.A(_05182_),
    .X(net6426));
 sg13g2_buf_1 fanout6427 (.A(_05182_),
    .X(net6427));
 sg13g2_buf_2 fanout6428 (.A(_05178_),
    .X(net6428));
 sg13g2_buf_1 fanout6429 (.A(_05178_),
    .X(net6429));
 sg13g2_buf_2 fanout6430 (.A(_05146_),
    .X(net6430));
 sg13g2_buf_1 fanout6431 (.A(_05146_),
    .X(net6431));
 sg13g2_buf_2 fanout6432 (.A(_05142_),
    .X(net6432));
 sg13g2_buf_1 fanout6433 (.A(_05142_),
    .X(net6433));
 sg13g2_buf_4 fanout6434 (.X(net6434),
    .A(_05138_));
 sg13g2_buf_1 fanout6435 (.A(_05138_),
    .X(net6435));
 sg13g2_buf_2 fanout6436 (.A(_05134_),
    .X(net6436));
 sg13g2_buf_1 fanout6437 (.A(_05134_),
    .X(net6437));
 sg13g2_buf_2 fanout6438 (.A(_05106_),
    .X(net6438));
 sg13g2_buf_1 fanout6439 (.A(_05106_),
    .X(net6439));
 sg13g2_buf_2 fanout6440 (.A(_05098_),
    .X(net6440));
 sg13g2_buf_1 fanout6441 (.A(_05098_),
    .X(net6441));
 sg13g2_buf_2 fanout6442 (.A(_05094_),
    .X(net6442));
 sg13g2_buf_1 fanout6443 (.A(_05094_),
    .X(net6443));
 sg13g2_buf_2 fanout6444 (.A(_05090_),
    .X(net6444));
 sg13g2_buf_1 fanout6445 (.A(_05090_),
    .X(net6445));
 sg13g2_buf_2 fanout6446 (.A(_05086_),
    .X(net6446));
 sg13g2_buf_1 fanout6447 (.A(_05086_),
    .X(net6447));
 sg13g2_buf_2 fanout6448 (.A(_05082_),
    .X(net6448));
 sg13g2_buf_1 fanout6449 (.A(_05082_),
    .X(net6449));
 sg13g2_buf_2 fanout6450 (.A(_05078_),
    .X(net6450));
 sg13g2_buf_1 fanout6451 (.A(_05078_),
    .X(net6451));
 sg13g2_buf_2 fanout6452 (.A(_05074_),
    .X(net6452));
 sg13g2_buf_1 fanout6453 (.A(_05074_),
    .X(net6453));
 sg13g2_buf_2 fanout6454 (.A(_05070_),
    .X(net6454));
 sg13g2_buf_1 fanout6455 (.A(_05070_),
    .X(net6455));
 sg13g2_buf_2 fanout6456 (.A(_05062_),
    .X(net6456));
 sg13g2_buf_1 fanout6457 (.A(_05062_),
    .X(net6457));
 sg13g2_buf_2 fanout6458 (.A(_05058_),
    .X(net6458));
 sg13g2_buf_1 fanout6459 (.A(_05058_),
    .X(net6459));
 sg13g2_buf_2 fanout6460 (.A(_05027_),
    .X(net6460));
 sg13g2_buf_1 fanout6461 (.A(_05027_),
    .X(net6461));
 sg13g2_buf_2 fanout6462 (.A(_05023_),
    .X(net6462));
 sg13g2_buf_1 fanout6463 (.A(_05023_),
    .X(net6463));
 sg13g2_buf_2 fanout6464 (.A(_05015_),
    .X(net6464));
 sg13g2_buf_1 fanout6465 (.A(_05015_),
    .X(net6465));
 sg13g2_buf_2 fanout6466 (.A(_05011_),
    .X(net6466));
 sg13g2_buf_1 fanout6467 (.A(_05011_),
    .X(net6467));
 sg13g2_buf_2 fanout6468 (.A(_05007_),
    .X(net6468));
 sg13g2_buf_1 fanout6469 (.A(_05007_),
    .X(net6469));
 sg13g2_buf_2 fanout6470 (.A(_04995_),
    .X(net6470));
 sg13g2_buf_1 fanout6471 (.A(_04995_),
    .X(net6471));
 sg13g2_buf_2 fanout6472 (.A(_04987_),
    .X(net6472));
 sg13g2_buf_1 fanout6473 (.A(_04987_),
    .X(net6473));
 sg13g2_buf_2 fanout6474 (.A(_04983_),
    .X(net6474));
 sg13g2_buf_1 fanout6475 (.A(_04983_),
    .X(net6475));
 sg13g2_buf_2 fanout6476 (.A(_04979_),
    .X(net6476));
 sg13g2_buf_1 fanout6477 (.A(_04979_),
    .X(net6477));
 sg13g2_buf_2 fanout6478 (.A(_04975_),
    .X(net6478));
 sg13g2_buf_1 fanout6479 (.A(_04975_),
    .X(net6479));
 sg13g2_buf_2 fanout6480 (.A(_04971_),
    .X(net6480));
 sg13g2_buf_1 fanout6481 (.A(_04971_),
    .X(net6481));
 sg13g2_buf_2 fanout6482 (.A(_04963_),
    .X(net6482));
 sg13g2_buf_1 fanout6483 (.A(_04963_),
    .X(net6483));
 sg13g2_buf_2 fanout6484 (.A(_04959_),
    .X(net6484));
 sg13g2_buf_1 fanout6485 (.A(_04959_),
    .X(net6485));
 sg13g2_buf_2 fanout6486 (.A(_04951_),
    .X(net6486));
 sg13g2_buf_1 fanout6487 (.A(_04951_),
    .X(net6487));
 sg13g2_buf_2 fanout6488 (.A(_04947_),
    .X(net6488));
 sg13g2_buf_1 fanout6489 (.A(_04947_),
    .X(net6489));
 sg13g2_buf_4 fanout6490 (.X(net6490),
    .A(_04943_));
 sg13g2_buf_1 fanout6491 (.A(_04943_),
    .X(net6491));
 sg13g2_buf_2 fanout6492 (.A(_04939_),
    .X(net6492));
 sg13g2_buf_1 fanout6493 (.A(_04939_),
    .X(net6493));
 sg13g2_buf_2 fanout6494 (.A(_04935_),
    .X(net6494));
 sg13g2_buf_1 fanout6495 (.A(_04935_),
    .X(net6495));
 sg13g2_buf_2 fanout6496 (.A(_04931_),
    .X(net6496));
 sg13g2_buf_1 fanout6497 (.A(_04931_),
    .X(net6497));
 sg13g2_buf_2 fanout6498 (.A(_04927_),
    .X(net6498));
 sg13g2_buf_1 fanout6499 (.A(_04927_),
    .X(net6499));
 sg13g2_buf_4 fanout6500 (.X(net6500),
    .A(_04923_));
 sg13g2_buf_1 fanout6501 (.A(_04923_),
    .X(net6501));
 sg13g2_buf_2 fanout6502 (.A(_04911_),
    .X(net6502));
 sg13g2_buf_1 fanout6503 (.A(_04911_),
    .X(net6503));
 sg13g2_buf_2 fanout6504 (.A(_04907_),
    .X(net6504));
 sg13g2_buf_1 fanout6505 (.A(_04907_),
    .X(net6505));
 sg13g2_buf_2 fanout6506 (.A(_04903_),
    .X(net6506));
 sg13g2_buf_1 fanout6507 (.A(_04903_),
    .X(net6507));
 sg13g2_buf_2 fanout6508 (.A(_04899_),
    .X(net6508));
 sg13g2_buf_1 fanout6509 (.A(_04899_),
    .X(net6509));
 sg13g2_buf_2 fanout6510 (.A(_04895_),
    .X(net6510));
 sg13g2_buf_1 fanout6511 (.A(_04895_),
    .X(net6511));
 sg13g2_buf_2 fanout6512 (.A(_04891_),
    .X(net6512));
 sg13g2_buf_1 fanout6513 (.A(_04891_),
    .X(net6513));
 sg13g2_buf_2 fanout6514 (.A(_04887_),
    .X(net6514));
 sg13g2_buf_1 fanout6515 (.A(_04887_),
    .X(net6515));
 sg13g2_buf_2 fanout6516 (.A(_04865_),
    .X(net6516));
 sg13g2_buf_1 fanout6517 (.A(_04865_),
    .X(net6517));
 sg13g2_buf_2 fanout6518 (.A(_04853_),
    .X(net6518));
 sg13g2_buf_1 fanout6519 (.A(_04853_),
    .X(net6519));
 sg13g2_buf_4 fanout6520 (.X(net6520),
    .A(_04849_));
 sg13g2_buf_1 fanout6521 (.A(_04849_),
    .X(net6521));
 sg13g2_buf_2 fanout6522 (.A(_04841_),
    .X(net6522));
 sg13g2_buf_1 fanout6523 (.A(_04841_),
    .X(net6523));
 sg13g2_buf_2 fanout6524 (.A(_04837_),
    .X(net6524));
 sg13g2_buf_1 fanout6525 (.A(_04837_),
    .X(net6525));
 sg13g2_buf_2 fanout6526 (.A(_04833_),
    .X(net6526));
 sg13g2_buf_1 fanout6527 (.A(_04833_),
    .X(net6527));
 sg13g2_buf_2 fanout6528 (.A(_04829_),
    .X(net6528));
 sg13g2_buf_1 fanout6529 (.A(_04829_),
    .X(net6529));
 sg13g2_buf_4 fanout6530 (.X(net6530),
    .A(_04825_));
 sg13g2_buf_1 fanout6531 (.A(_04825_),
    .X(net6531));
 sg13g2_buf_2 fanout6532 (.A(_04821_),
    .X(net6532));
 sg13g2_buf_1 fanout6533 (.A(_04821_),
    .X(net6533));
 sg13g2_buf_2 fanout6534 (.A(_04817_),
    .X(net6534));
 sg13g2_buf_1 fanout6535 (.A(_04817_),
    .X(net6535));
 sg13g2_buf_2 fanout6536 (.A(_04813_),
    .X(net6536));
 sg13g2_buf_1 fanout6537 (.A(_04813_),
    .X(net6537));
 sg13g2_buf_2 fanout6538 (.A(_04809_),
    .X(net6538));
 sg13g2_buf_1 fanout6539 (.A(_04809_),
    .X(net6539));
 sg13g2_buf_2 fanout6540 (.A(_04805_),
    .X(net6540));
 sg13g2_buf_1 fanout6541 (.A(_04805_),
    .X(net6541));
 sg13g2_buf_2 fanout6542 (.A(_04801_),
    .X(net6542));
 sg13g2_buf_1 fanout6543 (.A(_04801_),
    .X(net6543));
 sg13g2_buf_2 fanout6544 (.A(_04793_),
    .X(net6544));
 sg13g2_buf_1 fanout6545 (.A(_04793_),
    .X(net6545));
 sg13g2_buf_2 fanout6546 (.A(_04781_),
    .X(net6546));
 sg13g2_buf_1 fanout6547 (.A(_04781_),
    .X(net6547));
 sg13g2_buf_2 fanout6548 (.A(_04769_),
    .X(net6548));
 sg13g2_buf_1 fanout6549 (.A(_04769_),
    .X(net6549));
 sg13g2_buf_2 fanout6550 (.A(_04761_),
    .X(net6550));
 sg13g2_buf_1 fanout6551 (.A(_04761_),
    .X(net6551));
 sg13g2_buf_2 fanout6552 (.A(_04753_),
    .X(net6552));
 sg13g2_buf_1 fanout6553 (.A(_04753_),
    .X(net6553));
 sg13g2_buf_2 fanout6554 (.A(_04749_),
    .X(net6554));
 sg13g2_buf_1 fanout6555 (.A(_04749_),
    .X(net6555));
 sg13g2_buf_2 fanout6556 (.A(_04745_),
    .X(net6556));
 sg13g2_buf_1 fanout6557 (.A(_04745_),
    .X(net6557));
 sg13g2_buf_2 fanout6558 (.A(_04741_),
    .X(net6558));
 sg13g2_buf_1 fanout6559 (.A(_04741_),
    .X(net6559));
 sg13g2_buf_2 fanout6560 (.A(_04733_),
    .X(net6560));
 sg13g2_buf_1 fanout6561 (.A(_04733_),
    .X(net6561));
 sg13g2_buf_2 fanout6562 (.A(_04721_),
    .X(net6562));
 sg13g2_buf_1 fanout6563 (.A(_04721_),
    .X(net6563));
 sg13g2_buf_2 fanout6564 (.A(_04712_),
    .X(net6564));
 sg13g2_buf_1 fanout6565 (.A(_04712_),
    .X(net6565));
 sg13g2_buf_2 fanout6566 (.A(_04708_),
    .X(net6566));
 sg13g2_buf_1 fanout6567 (.A(_04708_),
    .X(net6567));
 sg13g2_buf_2 fanout6568 (.A(_04704_),
    .X(net6568));
 sg13g2_buf_1 fanout6569 (.A(_04704_),
    .X(net6569));
 sg13g2_buf_2 fanout6570 (.A(_04700_),
    .X(net6570));
 sg13g2_buf_1 fanout6571 (.A(_04700_),
    .X(net6571));
 sg13g2_buf_2 fanout6572 (.A(_04696_),
    .X(net6572));
 sg13g2_buf_1 fanout6573 (.A(_04696_),
    .X(net6573));
 sg13g2_buf_2 fanout6574 (.A(_04692_),
    .X(net6574));
 sg13g2_buf_1 fanout6575 (.A(_04692_),
    .X(net6575));
 sg13g2_buf_2 fanout6576 (.A(_04688_),
    .X(net6576));
 sg13g2_buf_1 fanout6577 (.A(_04688_),
    .X(net6577));
 sg13g2_buf_2 fanout6578 (.A(_04684_),
    .X(net6578));
 sg13g2_buf_1 fanout6579 (.A(_04684_),
    .X(net6579));
 sg13g2_buf_2 fanout6580 (.A(_04672_),
    .X(net6580));
 sg13g2_buf_1 fanout6581 (.A(_04672_),
    .X(net6581));
 sg13g2_buf_2 fanout6582 (.A(_04664_),
    .X(net6582));
 sg13g2_buf_1 fanout6583 (.A(_04664_),
    .X(net6583));
 sg13g2_buf_4 fanout6584 (.X(net6584),
    .A(_04660_));
 sg13g2_buf_1 fanout6585 (.A(_04660_),
    .X(net6585));
 sg13g2_buf_2 fanout6586 (.A(_04656_),
    .X(net6586));
 sg13g2_buf_1 fanout6587 (.A(_04656_),
    .X(net6587));
 sg13g2_buf_2 fanout6588 (.A(_04652_),
    .X(net6588));
 sg13g2_buf_1 fanout6589 (.A(_04652_),
    .X(net6589));
 sg13g2_buf_2 fanout6590 (.A(_04648_),
    .X(net6590));
 sg13g2_buf_1 fanout6591 (.A(_04648_),
    .X(net6591));
 sg13g2_buf_2 fanout6592 (.A(_04644_),
    .X(net6592));
 sg13g2_buf_1 fanout6593 (.A(_04644_),
    .X(net6593));
 sg13g2_buf_2 fanout6594 (.A(_04640_),
    .X(net6594));
 sg13g2_buf_1 fanout6595 (.A(_04640_),
    .X(net6595));
 sg13g2_buf_4 fanout6596 (.X(net6596),
    .A(_04636_));
 sg13g2_buf_1 fanout6597 (.A(_04636_),
    .X(net6597));
 sg13g2_buf_2 fanout6598 (.A(_04632_),
    .X(net6598));
 sg13g2_buf_1 fanout6599 (.A(_04632_),
    .X(net6599));
 sg13g2_buf_2 fanout6600 (.A(_04628_),
    .X(net6600));
 sg13g2_buf_1 fanout6601 (.A(_04628_),
    .X(net6601));
 sg13g2_buf_2 fanout6602 (.A(_04624_),
    .X(net6602));
 sg13g2_buf_1 fanout6603 (.A(_04624_),
    .X(net6603));
 sg13g2_buf_2 fanout6604 (.A(_04616_),
    .X(net6604));
 sg13g2_buf_1 fanout6605 (.A(_04616_),
    .X(net6605));
 sg13g2_buf_2 fanout6606 (.A(_04612_),
    .X(net6606));
 sg13g2_buf_1 fanout6607 (.A(_04612_),
    .X(net6607));
 sg13g2_buf_4 fanout6608 (.X(net6608),
    .A(_04608_));
 sg13g2_buf_1 fanout6609 (.A(_04608_),
    .X(net6609));
 sg13g2_buf_2 fanout6610 (.A(_04604_),
    .X(net6610));
 sg13g2_buf_1 fanout6611 (.A(_04604_),
    .X(net6611));
 sg13g2_buf_2 fanout6612 (.A(_04600_),
    .X(net6612));
 sg13g2_buf_1 fanout6613 (.A(_04600_),
    .X(net6613));
 sg13g2_buf_4 fanout6614 (.X(net6614),
    .A(_04596_));
 sg13g2_buf_1 fanout6615 (.A(_04596_),
    .X(net6615));
 sg13g2_buf_2 fanout6616 (.A(_04588_),
    .X(net6616));
 sg13g2_buf_1 fanout6617 (.A(_04588_),
    .X(net6617));
 sg13g2_buf_2 fanout6618 (.A(_04584_),
    .X(net6618));
 sg13g2_buf_1 fanout6619 (.A(_04584_),
    .X(net6619));
 sg13g2_buf_2 fanout6620 (.A(_04576_),
    .X(net6620));
 sg13g2_buf_2 fanout6621 (.A(_04576_),
    .X(net6621));
 sg13g2_buf_2 fanout6622 (.A(_04572_),
    .X(net6622));
 sg13g2_buf_1 fanout6623 (.A(_04572_),
    .X(net6623));
 sg13g2_buf_2 fanout6624 (.A(_04504_),
    .X(net6624));
 sg13g2_buf_1 fanout6625 (.A(_04504_),
    .X(net6625));
 sg13g2_buf_2 fanout6626 (.A(_04500_),
    .X(net6626));
 sg13g2_buf_1 fanout6627 (.A(_04500_),
    .X(net6627));
 sg13g2_buf_2 fanout6628 (.A(_04496_),
    .X(net6628));
 sg13g2_buf_1 fanout6629 (.A(_04496_),
    .X(net6629));
 sg13g2_buf_2 fanout6630 (.A(_04492_),
    .X(net6630));
 sg13g2_buf_1 fanout6631 (.A(_04492_),
    .X(net6631));
 sg13g2_buf_2 fanout6632 (.A(_04460_),
    .X(net6632));
 sg13g2_buf_1 fanout6633 (.A(_04460_),
    .X(net6633));
 sg13g2_buf_2 fanout6634 (.A(_04456_),
    .X(net6634));
 sg13g2_buf_1 fanout6635 (.A(_04456_),
    .X(net6635));
 sg13g2_buf_2 fanout6636 (.A(_04452_),
    .X(net6636));
 sg13g2_buf_1 fanout6637 (.A(_04452_),
    .X(net6637));
 sg13g2_buf_2 fanout6638 (.A(_04448_),
    .X(net6638));
 sg13g2_buf_1 fanout6639 (.A(_04448_),
    .X(net6639));
 sg13g2_buf_2 fanout6640 (.A(_04444_),
    .X(net6640));
 sg13g2_buf_1 fanout6641 (.A(_04444_),
    .X(net6641));
 sg13g2_buf_2 fanout6642 (.A(_04440_),
    .X(net6642));
 sg13g2_buf_2 fanout6643 (.A(_04440_),
    .X(net6643));
 sg13g2_buf_2 fanout6644 (.A(_04432_),
    .X(net6644));
 sg13g2_buf_1 fanout6645 (.A(_04432_),
    .X(net6645));
 sg13g2_buf_2 fanout6646 (.A(_04428_),
    .X(net6646));
 sg13g2_buf_1 fanout6647 (.A(_04428_),
    .X(net6647));
 sg13g2_buf_2 fanout6648 (.A(_04424_),
    .X(net6648));
 sg13g2_buf_1 fanout6649 (.A(_04424_),
    .X(net6649));
 sg13g2_buf_2 fanout6650 (.A(_04420_),
    .X(net6650));
 sg13g2_buf_1 fanout6651 (.A(_04420_),
    .X(net6651));
 sg13g2_buf_2 fanout6652 (.A(_04416_),
    .X(net6652));
 sg13g2_buf_1 fanout6653 (.A(_04416_),
    .X(net6653));
 sg13g2_buf_2 fanout6654 (.A(_04412_),
    .X(net6654));
 sg13g2_buf_1 fanout6655 (.A(_04412_),
    .X(net6655));
 sg13g2_buf_2 fanout6656 (.A(_04376_),
    .X(net6656));
 sg13g2_buf_1 fanout6657 (.A(_04376_),
    .X(net6657));
 sg13g2_buf_2 fanout6658 (.A(_04372_),
    .X(net6658));
 sg13g2_buf_1 fanout6659 (.A(_04372_),
    .X(net6659));
 sg13g2_buf_2 fanout6660 (.A(_04368_),
    .X(net6660));
 sg13g2_buf_1 fanout6661 (.A(_04368_),
    .X(net6661));
 sg13g2_buf_2 fanout6662 (.A(_04364_),
    .X(net6662));
 sg13g2_buf_2 fanout6663 (.A(_04364_),
    .X(net6663));
 sg13g2_buf_2 fanout6664 (.A(_04332_),
    .X(net6664));
 sg13g2_buf_1 fanout6665 (.A(_04332_),
    .X(net6665));
 sg13g2_buf_2 fanout6666 (.A(_04328_),
    .X(net6666));
 sg13g2_buf_1 fanout6667 (.A(_04328_),
    .X(net6667));
 sg13g2_buf_4 fanout6668 (.X(net6668),
    .A(_04324_));
 sg13g2_buf_1 fanout6669 (.A(_04324_),
    .X(net6669));
 sg13g2_buf_2 fanout6670 (.A(_04320_),
    .X(net6670));
 sg13g2_buf_1 fanout6671 (.A(_04320_),
    .X(net6671));
 sg13g2_buf_2 fanout6672 (.A(_04316_),
    .X(net6672));
 sg13g2_buf_1 fanout6673 (.A(_04316_),
    .X(net6673));
 sg13g2_buf_2 fanout6674 (.A(_04312_),
    .X(net6674));
 sg13g2_buf_1 fanout6675 (.A(_04312_),
    .X(net6675));
 sg13g2_buf_2 fanout6676 (.A(_04308_),
    .X(net6676));
 sg13g2_buf_1 fanout6677 (.A(_04308_),
    .X(net6677));
 sg13g2_buf_2 fanout6678 (.A(_04304_),
    .X(net6678));
 sg13g2_buf_1 fanout6679 (.A(_04304_),
    .X(net6679));
 sg13g2_buf_2 fanout6680 (.A(_04300_),
    .X(net6680));
 sg13g2_buf_1 fanout6681 (.A(_04300_),
    .X(net6681));
 sg13g2_buf_2 fanout6682 (.A(_04296_),
    .X(net6682));
 sg13g2_buf_1 fanout6683 (.A(_04296_),
    .X(net6683));
 sg13g2_buf_2 fanout6684 (.A(_04292_),
    .X(net6684));
 sg13g2_buf_1 fanout6685 (.A(_04292_),
    .X(net6685));
 sg13g2_buf_2 fanout6686 (.A(_04286_),
    .X(net6686));
 sg13g2_buf_1 fanout6687 (.A(_04286_),
    .X(net6687));
 sg13g2_buf_2 fanout6688 (.A(_04282_),
    .X(net6688));
 sg13g2_buf_1 fanout6689 (.A(_04282_),
    .X(net6689));
 sg13g2_buf_2 fanout6690 (.A(_04278_),
    .X(net6690));
 sg13g2_buf_1 fanout6691 (.A(_04278_),
    .X(net6691));
 sg13g2_buf_2 fanout6692 (.A(_04274_),
    .X(net6692));
 sg13g2_buf_1 fanout6693 (.A(_04274_),
    .X(net6693));
 sg13g2_buf_2 fanout6694 (.A(_04270_),
    .X(net6694));
 sg13g2_buf_1 fanout6695 (.A(_04270_),
    .X(net6695));
 sg13g2_buf_2 fanout6696 (.A(_04266_),
    .X(net6696));
 sg13g2_buf_1 fanout6697 (.A(_04266_),
    .X(net6697));
 sg13g2_buf_2 fanout6698 (.A(_04258_),
    .X(net6698));
 sg13g2_buf_1 fanout6699 (.A(_04258_),
    .X(net6699));
 sg13g2_buf_2 fanout6700 (.A(_04254_),
    .X(net6700));
 sg13g2_buf_1 fanout6701 (.A(_04254_),
    .X(net6701));
 sg13g2_buf_2 fanout6702 (.A(_04246_),
    .X(net6702));
 sg13g2_buf_1 fanout6703 (.A(_04246_),
    .X(net6703));
 sg13g2_buf_2 fanout6704 (.A(_04242_),
    .X(net6704));
 sg13g2_buf_1 fanout6705 (.A(_04242_),
    .X(net6705));
 sg13g2_buf_2 fanout6706 (.A(_04230_),
    .X(net6706));
 sg13g2_buf_1 fanout6707 (.A(_04230_),
    .X(net6707));
 sg13g2_buf_2 fanout6708 (.A(_04222_),
    .X(net6708));
 sg13g2_buf_1 fanout6709 (.A(_04222_),
    .X(net6709));
 sg13g2_buf_2 fanout6710 (.A(_04212_),
    .X(net6710));
 sg13g2_buf_1 fanout6711 (.A(_04212_),
    .X(net6711));
 sg13g2_buf_2 fanout6712 (.A(_04203_),
    .X(net6712));
 sg13g2_buf_1 fanout6713 (.A(_04203_),
    .X(net6713));
 sg13g2_buf_2 fanout6714 (.A(_04199_),
    .X(net6714));
 sg13g2_buf_1 fanout6715 (.A(_04199_),
    .X(net6715));
 sg13g2_buf_2 fanout6716 (.A(_04189_),
    .X(net6716));
 sg13g2_buf_1 fanout6717 (.A(_04189_),
    .X(net6717));
 sg13g2_buf_2 fanout6718 (.A(_04178_),
    .X(net6718));
 sg13g2_buf_1 fanout6719 (.A(_04178_),
    .X(net6719));
 sg13g2_buf_2 fanout6720 (.A(_04170_),
    .X(net6720));
 sg13g2_buf_1 fanout6721 (.A(_04170_),
    .X(net6721));
 sg13g2_buf_4 fanout6722 (.X(net6722),
    .A(_04160_));
 sg13g2_buf_1 fanout6723 (.A(_04160_),
    .X(net6723));
 sg13g2_buf_2 fanout6724 (.A(_04155_),
    .X(net6724));
 sg13g2_buf_1 fanout6725 (.A(_04155_),
    .X(net6725));
 sg13g2_buf_2 fanout6726 (.A(_04136_),
    .X(net6726));
 sg13g2_buf_1 fanout6727 (.A(_04136_),
    .X(net6727));
 sg13g2_buf_2 fanout6728 (.A(_04124_),
    .X(net6728));
 sg13g2_buf_1 fanout6729 (.A(_04124_),
    .X(net6729));
 sg13g2_buf_2 fanout6730 (.A(_04120_),
    .X(net6730));
 sg13g2_buf_1 fanout6731 (.A(_04120_),
    .X(net6731));
 sg13g2_buf_2 fanout6732 (.A(_04111_),
    .X(net6732));
 sg13g2_buf_1 fanout6733 (.A(_04111_),
    .X(net6733));
 sg13g2_buf_2 fanout6734 (.A(_04102_),
    .X(net6734));
 sg13g2_buf_1 fanout6735 (.A(_04102_),
    .X(net6735));
 sg13g2_buf_2 fanout6736 (.A(net6737),
    .X(net6736));
 sg13g2_buf_4 fanout6737 (.X(net6737),
    .A(net6738));
 sg13g2_buf_2 fanout6738 (.A(net6743),
    .X(net6738));
 sg13g2_buf_2 fanout6739 (.A(net6743),
    .X(net6739));
 sg13g2_buf_2 fanout6740 (.A(net6742),
    .X(net6740));
 sg13g2_buf_2 fanout6741 (.A(net6742),
    .X(net6741));
 sg13g2_buf_2 fanout6742 (.A(net6743),
    .X(net6742));
 sg13g2_buf_2 fanout6743 (.A(\top1.fsm.clk ),
    .X(net6743));
 sg13g2_buf_2 fanout6744 (.A(net6745),
    .X(net6744));
 sg13g2_buf_2 fanout6745 (.A(net6746),
    .X(net6745));
 sg13g2_buf_4 fanout6746 (.X(net6746),
    .A(\top1.fsm.clk ));
 sg13g2_buf_2 fanout6747 (.A(_02622_),
    .X(net6747));
 sg13g2_buf_1 fanout6748 (.A(_02622_),
    .X(net6748));
 sg13g2_buf_2 fanout6749 (.A(_02599_),
    .X(net6749));
 sg13g2_buf_1 fanout6750 (.A(_02599_),
    .X(net6750));
 sg13g2_buf_2 fanout6751 (.A(_02595_),
    .X(net6751));
 sg13g2_buf_1 fanout6752 (.A(_02595_),
    .X(net6752));
 sg13g2_buf_2 fanout6753 (.A(net6754),
    .X(net6753));
 sg13g2_buf_2 fanout6754 (.A(_02591_),
    .X(net6754));
 sg13g2_buf_2 fanout6755 (.A(_02587_),
    .X(net6755));
 sg13g2_buf_1 fanout6756 (.A(_02587_),
    .X(net6756));
 sg13g2_buf_2 fanout6757 (.A(_02583_),
    .X(net6757));
 sg13g2_buf_1 fanout6758 (.A(_02583_),
    .X(net6758));
 sg13g2_buf_2 fanout6759 (.A(_02568_),
    .X(net6759));
 sg13g2_buf_1 fanout6760 (.A(_02568_),
    .X(net6760));
 sg13g2_buf_2 fanout6761 (.A(_02560_),
    .X(net6761));
 sg13g2_buf_1 fanout6762 (.A(_02560_),
    .X(net6762));
 sg13g2_buf_2 fanout6763 (.A(_02552_),
    .X(net6763));
 sg13g2_buf_1 fanout6764 (.A(_02552_),
    .X(net6764));
 sg13g2_buf_2 fanout6765 (.A(_02548_),
    .X(net6765));
 sg13g2_buf_1 fanout6766 (.A(_02548_),
    .X(net6766));
 sg13g2_buf_2 fanout6767 (.A(_02544_),
    .X(net6767));
 sg13g2_buf_1 fanout6768 (.A(_02544_),
    .X(net6768));
 sg13g2_buf_2 fanout6769 (.A(_02540_),
    .X(net6769));
 sg13g2_buf_1 fanout6770 (.A(_02540_),
    .X(net6770));
 sg13g2_buf_2 fanout6771 (.A(_02536_),
    .X(net6771));
 sg13g2_buf_1 fanout6772 (.A(_02536_),
    .X(net6772));
 sg13g2_buf_2 fanout6773 (.A(_02532_),
    .X(net6773));
 sg13g2_buf_1 fanout6774 (.A(_02532_),
    .X(net6774));
 sg13g2_buf_2 fanout6775 (.A(_02528_),
    .X(net6775));
 sg13g2_buf_1 fanout6776 (.A(_02528_),
    .X(net6776));
 sg13g2_buf_2 fanout6777 (.A(_07458_),
    .X(net6777));
 sg13g2_buf_1 fanout6778 (.A(_07458_),
    .X(net6778));
 sg13g2_buf_2 fanout6779 (.A(_07446_),
    .X(net6779));
 sg13g2_buf_1 fanout6780 (.A(_07446_),
    .X(net6780));
 sg13g2_buf_2 fanout6781 (.A(_07442_),
    .X(net6781));
 sg13g2_buf_1 fanout6782 (.A(_07442_),
    .X(net6782));
 sg13g2_buf_2 fanout6783 (.A(_07438_),
    .X(net6783));
 sg13g2_buf_1 fanout6784 (.A(_07438_),
    .X(net6784));
 sg13g2_buf_2 fanout6785 (.A(_07434_),
    .X(net6785));
 sg13g2_buf_1 fanout6786 (.A(_07434_),
    .X(net6786));
 sg13g2_buf_2 fanout6787 (.A(_07430_),
    .X(net6787));
 sg13g2_buf_1 fanout6788 (.A(_07430_),
    .X(net6788));
 sg13g2_buf_2 fanout6789 (.A(_07426_),
    .X(net6789));
 sg13g2_buf_1 fanout6790 (.A(_07426_),
    .X(net6790));
 sg13g2_buf_2 fanout6791 (.A(_07422_),
    .X(net6791));
 sg13g2_buf_1 fanout6792 (.A(_07422_),
    .X(net6792));
 sg13g2_buf_2 fanout6793 (.A(_07418_),
    .X(net6793));
 sg13g2_buf_1 fanout6794 (.A(_07418_),
    .X(net6794));
 sg13g2_buf_2 fanout6795 (.A(_07414_),
    .X(net6795));
 sg13g2_buf_1 fanout6796 (.A(_07414_),
    .X(net6796));
 sg13g2_buf_2 fanout6797 (.A(_07410_),
    .X(net6797));
 sg13g2_buf_1 fanout6798 (.A(_07410_),
    .X(net6798));
 sg13g2_buf_2 fanout6799 (.A(_07406_),
    .X(net6799));
 sg13g2_buf_1 fanout6800 (.A(_07406_),
    .X(net6800));
 sg13g2_buf_2 fanout6801 (.A(_07386_),
    .X(net6801));
 sg13g2_buf_1 fanout6802 (.A(_07386_),
    .X(net6802));
 sg13g2_buf_2 fanout6803 (.A(_07378_),
    .X(net6803));
 sg13g2_buf_1 fanout6804 (.A(_07378_),
    .X(net6804));
 sg13g2_buf_2 fanout6805 (.A(_07362_),
    .X(net6805));
 sg13g2_buf_1 fanout6806 (.A(_07362_),
    .X(net6806));
 sg13g2_buf_2 fanout6807 (.A(_07358_),
    .X(net6807));
 sg13g2_buf_1 fanout6808 (.A(_07358_),
    .X(net6808));
 sg13g2_buf_2 fanout6809 (.A(_07289_),
    .X(net6809));
 sg13g2_buf_1 fanout6810 (.A(_07289_),
    .X(net6810));
 sg13g2_buf_2 fanout6811 (.A(_07275_),
    .X(net6811));
 sg13g2_buf_1 fanout6812 (.A(_07275_),
    .X(net6812));
 sg13g2_buf_2 fanout6813 (.A(_07271_),
    .X(net6813));
 sg13g2_buf_1 fanout6814 (.A(_07271_),
    .X(net6814));
 sg13g2_buf_2 fanout6815 (.A(_07219_),
    .X(net6815));
 sg13g2_buf_1 fanout6816 (.A(_07219_),
    .X(net6816));
 sg13g2_buf_2 fanout6817 (.A(_07186_),
    .X(net6817));
 sg13g2_buf_1 fanout6818 (.A(_07186_),
    .X(net6818));
 sg13g2_buf_2 fanout6819 (.A(_06311_),
    .X(net6819));
 sg13g2_buf_1 fanout6820 (.A(_06311_),
    .X(net6820));
 sg13g2_buf_2 fanout6821 (.A(_06299_),
    .X(net6821));
 sg13g2_buf_1 fanout6822 (.A(_06299_),
    .X(net6822));
 sg13g2_buf_4 fanout6823 (.X(net6823),
    .A(_06291_));
 sg13g2_buf_1 fanout6824 (.A(_06291_),
    .X(net6824));
 sg13g2_buf_2 fanout6825 (.A(_06279_),
    .X(net6825));
 sg13g2_buf_1 fanout6826 (.A(_06279_),
    .X(net6826));
 sg13g2_buf_2 fanout6827 (.A(_05390_),
    .X(net6827));
 sg13g2_buf_1 fanout6828 (.A(_05390_),
    .X(net6828));
 sg13g2_buf_2 fanout6829 (.A(_05374_),
    .X(net6829));
 sg13g2_buf_1 fanout6830 (.A(_05374_),
    .X(net6830));
 sg13g2_buf_2 fanout6831 (.A(_05358_),
    .X(net6831));
 sg13g2_buf_1 fanout6832 (.A(_05358_),
    .X(net6832));
 sg13g2_buf_2 fanout6833 (.A(_05330_),
    .X(net6833));
 sg13g2_buf_1 fanout6834 (.A(_05330_),
    .X(net6834));
 sg13g2_buf_2 fanout6835 (.A(_05322_),
    .X(net6835));
 sg13g2_buf_1 fanout6836 (.A(_05322_),
    .X(net6836));
 sg13g2_buf_2 fanout6837 (.A(_05318_),
    .X(net6837));
 sg13g2_buf_1 fanout6838 (.A(_05318_),
    .X(net6838));
 sg13g2_buf_2 fanout6839 (.A(_05310_),
    .X(net6839));
 sg13g2_buf_1 fanout6840 (.A(_05310_),
    .X(net6840));
 sg13g2_buf_2 fanout6841 (.A(_05306_),
    .X(net6841));
 sg13g2_buf_1 fanout6842 (.A(_05306_),
    .X(net6842));
 sg13g2_buf_2 fanout6843 (.A(_05302_),
    .X(net6843));
 sg13g2_buf_1 fanout6844 (.A(_05302_),
    .X(net6844));
 sg13g2_buf_2 fanout6845 (.A(_05298_),
    .X(net6845));
 sg13g2_buf_1 fanout6846 (.A(_05298_),
    .X(net6846));
 sg13g2_buf_2 fanout6847 (.A(_05294_),
    .X(net6847));
 sg13g2_buf_1 fanout6848 (.A(_05294_),
    .X(net6848));
 sg13g2_buf_2 fanout6849 (.A(_05262_),
    .X(net6849));
 sg13g2_buf_1 fanout6850 (.A(_05262_),
    .X(net6850));
 sg13g2_buf_4 fanout6851 (.X(net6851),
    .A(_05250_));
 sg13g2_buf_1 fanout6852 (.A(_05250_),
    .X(net6852));
 sg13g2_buf_2 fanout6853 (.A(_05246_),
    .X(net6853));
 sg13g2_buf_1 fanout6854 (.A(_05246_),
    .X(net6854));
 sg13g2_buf_2 fanout6855 (.A(_05242_),
    .X(net6855));
 sg13g2_buf_1 fanout6856 (.A(_05242_),
    .X(net6856));
 sg13g2_buf_2 fanout6857 (.A(_05238_),
    .X(net6857));
 sg13g2_buf_1 fanout6858 (.A(_05238_),
    .X(net6858));
 sg13g2_buf_2 fanout6859 (.A(_05222_),
    .X(net6859));
 sg13g2_buf_1 fanout6860 (.A(_05222_),
    .X(net6860));
 sg13g2_buf_2 fanout6861 (.A(_05210_),
    .X(net6861));
 sg13g2_buf_1 fanout6862 (.A(_05210_),
    .X(net6862));
 sg13g2_buf_2 fanout6863 (.A(_05198_),
    .X(net6863));
 sg13g2_buf_1 fanout6864 (.A(_05198_),
    .X(net6864));
 sg13g2_buf_2 fanout6865 (.A(_05186_),
    .X(net6865));
 sg13g2_buf_1 fanout6866 (.A(_05186_),
    .X(net6866));
 sg13g2_buf_2 fanout6867 (.A(_05174_),
    .X(net6867));
 sg13g2_buf_1 fanout6868 (.A(_05174_),
    .X(net6868));
 sg13g2_buf_2 fanout6869 (.A(_05170_),
    .X(net6869));
 sg13g2_buf_1 fanout6870 (.A(_05170_),
    .X(net6870));
 sg13g2_buf_2 fanout6871 (.A(_05166_),
    .X(net6871));
 sg13g2_buf_1 fanout6872 (.A(_05166_),
    .X(net6872));
 sg13g2_buf_2 fanout6873 (.A(_05162_),
    .X(net6873));
 sg13g2_buf_1 fanout6874 (.A(_05162_),
    .X(net6874));
 sg13g2_buf_2 fanout6875 (.A(_05158_),
    .X(net6875));
 sg13g2_buf_1 fanout6876 (.A(_05158_),
    .X(net6876));
 sg13g2_buf_2 fanout6877 (.A(_05154_),
    .X(net6877));
 sg13g2_buf_1 fanout6878 (.A(_05154_),
    .X(net6878));
 sg13g2_buf_2 fanout6879 (.A(_05150_),
    .X(net6879));
 sg13g2_buf_1 fanout6880 (.A(_05150_),
    .X(net6880));
 sg13g2_buf_2 fanout6881 (.A(_05130_),
    .X(net6881));
 sg13g2_buf_1 fanout6882 (.A(_05130_),
    .X(net6882));
 sg13g2_buf_2 fanout6883 (.A(_05126_),
    .X(net6883));
 sg13g2_buf_1 fanout6884 (.A(_05126_),
    .X(net6884));
 sg13g2_buf_2 fanout6885 (.A(_05122_),
    .X(net6885));
 sg13g2_buf_1 fanout6886 (.A(_05122_),
    .X(net6886));
 sg13g2_buf_2 fanout6887 (.A(_05118_),
    .X(net6887));
 sg13g2_buf_1 fanout6888 (.A(_05118_),
    .X(net6888));
 sg13g2_buf_2 fanout6889 (.A(_05114_),
    .X(net6889));
 sg13g2_buf_1 fanout6890 (.A(_05114_),
    .X(net6890));
 sg13g2_buf_2 fanout6891 (.A(_05110_),
    .X(net6891));
 sg13g2_buf_1 fanout6892 (.A(_05110_),
    .X(net6892));
 sg13g2_buf_2 fanout6893 (.A(_05102_),
    .X(net6893));
 sg13g2_buf_1 fanout6894 (.A(_05102_),
    .X(net6894));
 sg13g2_buf_2 fanout6895 (.A(_05066_),
    .X(net6895));
 sg13g2_buf_1 fanout6896 (.A(_05066_),
    .X(net6896));
 sg13g2_buf_2 fanout6897 (.A(_05043_),
    .X(net6897));
 sg13g2_buf_2 fanout6898 (.A(_05031_),
    .X(net6898));
 sg13g2_buf_1 fanout6899 (.A(_05031_),
    .X(net6899));
 sg13g2_buf_4 fanout6900 (.X(net6900),
    .A(_05019_));
 sg13g2_buf_1 fanout6901 (.A(_05019_),
    .X(net6901));
 sg13g2_buf_2 fanout6902 (.A(_05003_),
    .X(net6902));
 sg13g2_buf_1 fanout6903 (.A(_05003_),
    .X(net6903));
 sg13g2_buf_2 fanout6904 (.A(_04999_),
    .X(net6904));
 sg13g2_buf_1 fanout6905 (.A(_04999_),
    .X(net6905));
 sg13g2_buf_2 fanout6906 (.A(_04991_),
    .X(net6906));
 sg13g2_buf_1 fanout6907 (.A(_04991_),
    .X(net6907));
 sg13g2_buf_2 fanout6908 (.A(_04967_),
    .X(net6908));
 sg13g2_buf_1 fanout6909 (.A(_04967_),
    .X(net6909));
 sg13g2_buf_2 fanout6910 (.A(_04955_),
    .X(net6910));
 sg13g2_buf_1 fanout6911 (.A(_04955_),
    .X(net6911));
 sg13g2_buf_2 fanout6912 (.A(_04919_),
    .X(net6912));
 sg13g2_buf_1 fanout6913 (.A(_04919_),
    .X(net6913));
 sg13g2_buf_2 fanout6914 (.A(_04915_),
    .X(net6914));
 sg13g2_buf_1 fanout6915 (.A(_04915_),
    .X(net6915));
 sg13g2_buf_2 fanout6916 (.A(_04883_),
    .X(net6916));
 sg13g2_buf_1 fanout6917 (.A(_04883_),
    .X(net6917));
 sg13g2_buf_2 fanout6918 (.A(_04879_),
    .X(net6918));
 sg13g2_buf_1 fanout6919 (.A(_04879_),
    .X(net6919));
 sg13g2_buf_2 fanout6920 (.A(_04875_),
    .X(net6920));
 sg13g2_buf_1 fanout6921 (.A(_04875_),
    .X(net6921));
 sg13g2_buf_2 fanout6922 (.A(_04871_),
    .X(net6922));
 sg13g2_buf_1 fanout6923 (.A(_04871_),
    .X(net6923));
 sg13g2_buf_2 fanout6924 (.A(_04861_),
    .X(net6924));
 sg13g2_buf_1 fanout6925 (.A(_04861_),
    .X(net6925));
 sg13g2_buf_2 fanout6926 (.A(_04857_),
    .X(net6926));
 sg13g2_buf_1 fanout6927 (.A(_04857_),
    .X(net6927));
 sg13g2_buf_2 fanout6928 (.A(_04845_),
    .X(net6928));
 sg13g2_buf_1 fanout6929 (.A(_04845_),
    .X(net6929));
 sg13g2_buf_2 fanout6930 (.A(_04797_),
    .X(net6930));
 sg13g2_buf_1 fanout6931 (.A(_04797_),
    .X(net6931));
 sg13g2_buf_2 fanout6932 (.A(_04789_),
    .X(net6932));
 sg13g2_buf_1 fanout6933 (.A(_04789_),
    .X(net6933));
 sg13g2_buf_2 fanout6934 (.A(_04785_),
    .X(net6934));
 sg13g2_buf_1 fanout6935 (.A(_04785_),
    .X(net6935));
 sg13g2_buf_2 fanout6936 (.A(_04777_),
    .X(net6936));
 sg13g2_buf_1 fanout6937 (.A(_04777_),
    .X(net6937));
 sg13g2_buf_2 fanout6938 (.A(_04773_),
    .X(net6938));
 sg13g2_buf_1 fanout6939 (.A(_04773_),
    .X(net6939));
 sg13g2_buf_2 fanout6940 (.A(_04765_),
    .X(net6940));
 sg13g2_buf_1 fanout6941 (.A(_04765_),
    .X(net6941));
 sg13g2_buf_2 fanout6942 (.A(_04757_),
    .X(net6942));
 sg13g2_buf_1 fanout6943 (.A(_04757_),
    .X(net6943));
 sg13g2_buf_2 fanout6944 (.A(_04737_),
    .X(net6944));
 sg13g2_buf_1 fanout6945 (.A(_04737_),
    .X(net6945));
 sg13g2_buf_2 fanout6946 (.A(_04729_),
    .X(net6946));
 sg13g2_buf_1 fanout6947 (.A(_04729_),
    .X(net6947));
 sg13g2_buf_2 fanout6948 (.A(_04725_),
    .X(net6948));
 sg13g2_buf_1 fanout6949 (.A(_04725_),
    .X(net6949));
 sg13g2_buf_2 fanout6950 (.A(_04717_),
    .X(net6950));
 sg13g2_buf_1 fanout6951 (.A(_04717_),
    .X(net6951));
 sg13g2_buf_2 fanout6952 (.A(_04680_),
    .X(net6952));
 sg13g2_buf_1 fanout6953 (.A(_04680_),
    .X(net6953));
 sg13g2_buf_2 fanout6954 (.A(_04676_),
    .X(net6954));
 sg13g2_buf_1 fanout6955 (.A(_04676_),
    .X(net6955));
 sg13g2_buf_2 fanout6956 (.A(_04668_),
    .X(net6956));
 sg13g2_buf_1 fanout6957 (.A(_04668_),
    .X(net6957));
 sg13g2_buf_2 fanout6958 (.A(_04620_),
    .X(net6958));
 sg13g2_buf_1 fanout6959 (.A(_04620_),
    .X(net6959));
 sg13g2_buf_2 fanout6960 (.A(net6961),
    .X(net6960));
 sg13g2_buf_1 fanout6961 (.A(_04592_),
    .X(net6961));
 sg13g2_buf_2 fanout6962 (.A(_04580_),
    .X(net6962));
 sg13g2_buf_1 fanout6963 (.A(_04580_),
    .X(net6963));
 sg13g2_buf_2 fanout6964 (.A(_04568_),
    .X(net6964));
 sg13g2_buf_1 fanout6965 (.A(_04568_),
    .X(net6965));
 sg13g2_buf_2 fanout6966 (.A(_04564_),
    .X(net6966));
 sg13g2_buf_1 fanout6967 (.A(_04564_),
    .X(net6967));
 sg13g2_buf_2 fanout6968 (.A(_04560_),
    .X(net6968));
 sg13g2_buf_1 fanout6969 (.A(_04560_),
    .X(net6969));
 sg13g2_buf_2 fanout6970 (.A(_04556_),
    .X(net6970));
 sg13g2_buf_1 fanout6971 (.A(_04556_),
    .X(net6971));
 sg13g2_buf_2 fanout6972 (.A(_04552_),
    .X(net6972));
 sg13g2_buf_1 fanout6973 (.A(_04552_),
    .X(net6973));
 sg13g2_buf_2 fanout6974 (.A(_04548_),
    .X(net6974));
 sg13g2_buf_1 fanout6975 (.A(_04548_),
    .X(net6975));
 sg13g2_buf_2 fanout6976 (.A(_04544_),
    .X(net6976));
 sg13g2_buf_1 fanout6977 (.A(_04544_),
    .X(net6977));
 sg13g2_buf_2 fanout6978 (.A(_04540_),
    .X(net6978));
 sg13g2_buf_1 fanout6979 (.A(_04540_),
    .X(net6979));
 sg13g2_buf_4 fanout6980 (.X(net6980),
    .A(_04536_));
 sg13g2_buf_1 fanout6981 (.A(_04536_),
    .X(net6981));
 sg13g2_buf_4 fanout6982 (.X(net6982),
    .A(_04532_));
 sg13g2_buf_1 fanout6983 (.A(_04532_),
    .X(net6983));
 sg13g2_buf_2 fanout6984 (.A(_04528_),
    .X(net6984));
 sg13g2_buf_1 fanout6985 (.A(_04528_),
    .X(net6985));
 sg13g2_buf_2 fanout6986 (.A(_04524_),
    .X(net6986));
 sg13g2_buf_1 fanout6987 (.A(_04524_),
    .X(net6987));
 sg13g2_buf_2 fanout6988 (.A(_04520_),
    .X(net6988));
 sg13g2_buf_1 fanout6989 (.A(_04520_),
    .X(net6989));
 sg13g2_buf_2 fanout6990 (.A(_04516_),
    .X(net6990));
 sg13g2_buf_1 fanout6991 (.A(_04516_),
    .X(net6991));
 sg13g2_buf_2 fanout6992 (.A(_04512_),
    .X(net6992));
 sg13g2_buf_1 fanout6993 (.A(_04512_),
    .X(net6993));
 sg13g2_buf_2 fanout6994 (.A(_04508_),
    .X(net6994));
 sg13g2_buf_1 fanout6995 (.A(_04508_),
    .X(net6995));
 sg13g2_buf_2 fanout6996 (.A(_04488_),
    .X(net6996));
 sg13g2_buf_1 fanout6997 (.A(_04488_),
    .X(net6997));
 sg13g2_buf_2 fanout6998 (.A(_04484_),
    .X(net6998));
 sg13g2_buf_1 fanout6999 (.A(_04484_),
    .X(net6999));
 sg13g2_buf_2 fanout7000 (.A(_04480_),
    .X(net7000));
 sg13g2_buf_1 fanout7001 (.A(_04480_),
    .X(net7001));
 sg13g2_buf_2 fanout7002 (.A(_04476_),
    .X(net7002));
 sg13g2_buf_1 fanout7003 (.A(_04476_),
    .X(net7003));
 sg13g2_buf_2 fanout7004 (.A(_04472_),
    .X(net7004));
 sg13g2_buf_1 fanout7005 (.A(_04472_),
    .X(net7005));
 sg13g2_buf_2 fanout7006 (.A(_04468_),
    .X(net7006));
 sg13g2_buf_1 fanout7007 (.A(_04468_),
    .X(net7007));
 sg13g2_buf_2 fanout7008 (.A(_04464_),
    .X(net7008));
 sg13g2_buf_1 fanout7009 (.A(_04464_),
    .X(net7009));
 sg13g2_buf_2 fanout7010 (.A(_04436_),
    .X(net7010));
 sg13g2_buf_1 fanout7011 (.A(_04436_),
    .X(net7011));
 sg13g2_buf_2 fanout7012 (.A(_04408_),
    .X(net7012));
 sg13g2_buf_1 fanout7013 (.A(_04408_),
    .X(net7013));
 sg13g2_buf_2 fanout7014 (.A(_04404_),
    .X(net7014));
 sg13g2_buf_1 fanout7015 (.A(_04404_),
    .X(net7015));
 sg13g2_buf_2 fanout7016 (.A(_04400_),
    .X(net7016));
 sg13g2_buf_1 fanout7017 (.A(_04400_),
    .X(net7017));
 sg13g2_buf_2 fanout7018 (.A(_04396_),
    .X(net7018));
 sg13g2_buf_1 fanout7019 (.A(_04396_),
    .X(net7019));
 sg13g2_buf_2 fanout7020 (.A(_04392_),
    .X(net7020));
 sg13g2_buf_1 fanout7021 (.A(_04392_),
    .X(net7021));
 sg13g2_buf_2 fanout7022 (.A(_04388_),
    .X(net7022));
 sg13g2_buf_1 fanout7023 (.A(_04388_),
    .X(net7023));
 sg13g2_buf_2 fanout7024 (.A(_04384_),
    .X(net7024));
 sg13g2_buf_1 fanout7025 (.A(_04384_),
    .X(net7025));
 sg13g2_buf_2 fanout7026 (.A(_04380_),
    .X(net7026));
 sg13g2_buf_1 fanout7027 (.A(_04380_),
    .X(net7027));
 sg13g2_buf_2 fanout7028 (.A(_04360_),
    .X(net7028));
 sg13g2_buf_1 fanout7029 (.A(_04360_),
    .X(net7029));
 sg13g2_buf_2 fanout7030 (.A(_04356_),
    .X(net7030));
 sg13g2_buf_1 fanout7031 (.A(_04356_),
    .X(net7031));
 sg13g2_buf_2 fanout7032 (.A(_04352_),
    .X(net7032));
 sg13g2_buf_1 fanout7033 (.A(_04352_),
    .X(net7033));
 sg13g2_buf_4 fanout7034 (.X(net7034),
    .A(_04348_));
 sg13g2_buf_1 fanout7035 (.A(_04348_),
    .X(net7035));
 sg13g2_buf_2 fanout7036 (.A(net7037),
    .X(net7036));
 sg13g2_buf_1 fanout7037 (.A(_04344_),
    .X(net7037));
 sg13g2_buf_2 fanout7038 (.A(net7039),
    .X(net7038));
 sg13g2_buf_1 fanout7039 (.A(_04340_),
    .X(net7039));
 sg13g2_buf_2 fanout7040 (.A(_04336_),
    .X(net7040));
 sg13g2_buf_1 fanout7041 (.A(_04336_),
    .X(net7041));
 sg13g2_buf_8 fanout7042 (.A(net7043),
    .X(net7042));
 sg13g2_buf_8 fanout7043 (.A(_04290_),
    .X(net7043));
 sg13g2_buf_2 fanout7044 (.A(_04262_),
    .X(net7044));
 sg13g2_buf_1 fanout7045 (.A(_04262_),
    .X(net7045));
 sg13g2_buf_2 fanout7046 (.A(_04250_),
    .X(net7046));
 sg13g2_buf_1 fanout7047 (.A(_04250_),
    .X(net7047));
 sg13g2_buf_2 fanout7048 (.A(net7050),
    .X(net7048));
 sg13g2_buf_2 fanout7049 (.A(net7050),
    .X(net7049));
 sg13g2_buf_2 fanout7050 (.A(net7052),
    .X(net7050));
 sg13g2_buf_4 fanout7051 (.X(net7051),
    .A(net7052));
 sg13g2_buf_4 fanout7052 (.X(net7052),
    .A(_04241_));
 sg13g2_buf_2 fanout7053 (.A(_04236_),
    .X(net7053));
 sg13g2_buf_1 fanout7054 (.A(_04236_),
    .X(net7054));
 sg13g2_buf_2 fanout7055 (.A(_04226_),
    .X(net7055));
 sg13g2_buf_1 fanout7056 (.A(_04226_),
    .X(net7056));
 sg13g2_buf_2 fanout7057 (.A(_04218_),
    .X(net7057));
 sg13g2_buf_1 fanout7058 (.A(_04218_),
    .X(net7058));
 sg13g2_buf_2 fanout7059 (.A(_04208_),
    .X(net7059));
 sg13g2_buf_1 fanout7060 (.A(_04208_),
    .X(net7060));
 sg13g2_buf_2 fanout7061 (.A(_04193_),
    .X(net7061));
 sg13g2_buf_1 fanout7062 (.A(_04193_),
    .X(net7062));
 sg13g2_buf_2 fanout7063 (.A(_04185_),
    .X(net7063));
 sg13g2_buf_1 fanout7064 (.A(_04185_),
    .X(net7064));
 sg13g2_buf_8 fanout7065 (.A(net7067),
    .X(net7065));
 sg13g2_buf_8 fanout7066 (.A(net7067),
    .X(net7066));
 sg13g2_buf_8 fanout7067 (.A(_04183_),
    .X(net7067));
 sg13g2_buf_2 fanout7068 (.A(_04174_),
    .X(net7068));
 sg13g2_buf_1 fanout7069 (.A(_04174_),
    .X(net7069));
 sg13g2_buf_2 fanout7070 (.A(_04166_),
    .X(net7070));
 sg13g2_buf_2 fanout7071 (.A(_04166_),
    .X(net7071));
 sg13g2_buf_2 fanout7072 (.A(net7073),
    .X(net7072));
 sg13g2_buf_2 fanout7073 (.A(net7077),
    .X(net7073));
 sg13g2_buf_2 fanout7074 (.A(net7076),
    .X(net7074));
 sg13g2_buf_1 fanout7075 (.A(net7076),
    .X(net7075));
 sg13g2_buf_2 fanout7076 (.A(net7077),
    .X(net7076));
 sg13g2_buf_4 fanout7077 (.X(net7077),
    .A(_04159_));
 sg13g2_buf_2 fanout7078 (.A(net7079),
    .X(net7078));
 sg13g2_buf_2 fanout7079 (.A(_04153_),
    .X(net7079));
 sg13g2_buf_2 fanout7080 (.A(net7082),
    .X(net7080));
 sg13g2_buf_1 fanout7081 (.A(net7082),
    .X(net7081));
 sg13g2_buf_2 fanout7082 (.A(_04153_),
    .X(net7082));
 sg13g2_buf_8 fanout7083 (.A(net7085),
    .X(net7083));
 sg13g2_buf_4 fanout7084 (.X(net7084),
    .A(net7085));
 sg13g2_buf_8 fanout7085 (.A(_04151_),
    .X(net7085));
 sg13g2_buf_2 fanout7086 (.A(_04147_),
    .X(net7086));
 sg13g2_buf_1 fanout7087 (.A(_04147_),
    .X(net7087));
 sg13g2_buf_2 fanout7088 (.A(_04143_),
    .X(net7088));
 sg13g2_buf_1 fanout7089 (.A(_04143_),
    .X(net7089));
 sg13g2_buf_2 fanout7090 (.A(_04131_),
    .X(net7090));
 sg13g2_buf_1 fanout7091 (.A(_04131_),
    .X(net7091));
 sg13g2_buf_4 fanout7092 (.X(net7092),
    .A(_04119_));
 sg13g2_buf_2 fanout7093 (.A(_04119_),
    .X(net7093));
 sg13g2_buf_2 fanout7094 (.A(net7095),
    .X(net7094));
 sg13g2_buf_1 fanout7095 (.A(_04118_),
    .X(net7095));
 sg13g2_buf_2 fanout7096 (.A(_04118_),
    .X(net7096));
 sg13g2_buf_4 fanout7097 (.X(net7097),
    .A(_04110_));
 sg13g2_buf_1 fanout7098 (.A(_04110_),
    .X(net7098));
 sg13g2_buf_2 fanout7099 (.A(net7101),
    .X(net7099));
 sg13g2_buf_2 fanout7100 (.A(net7101),
    .X(net7100));
 sg13g2_buf_2 fanout7101 (.A(_04109_),
    .X(net7101));
 sg13g2_buf_8 fanout7102 (.A(net7104),
    .X(net7102));
 sg13g2_buf_4 fanout7103 (.X(net7103),
    .A(net7104));
 sg13g2_buf_8 fanout7104 (.A(_04100_),
    .X(net7104));
 sg13g2_buf_2 fanout7105 (.A(_04094_),
    .X(net7105));
 sg13g2_buf_1 fanout7106 (.A(_04094_),
    .X(net7106));
 sg13g2_buf_8 fanout7107 (.A(_04093_),
    .X(net7107));
 sg13g2_buf_4 fanout7108 (.X(net7108),
    .A(_04088_));
 sg13g2_buf_1 fanout7109 (.A(_04088_),
    .X(net7109));
 sg13g2_buf_2 fanout7110 (.A(_04080_),
    .X(net7110));
 sg13g2_buf_1 fanout7111 (.A(_04080_),
    .X(net7111));
 sg13g2_buf_2 fanout7112 (.A(_04066_),
    .X(net7112));
 sg13g2_buf_1 fanout7113 (.A(_04066_),
    .X(net7113));
 sg13g2_buf_2 fanout7114 (.A(_04057_),
    .X(net7114));
 sg13g2_buf_2 fanout7115 (.A(_04057_),
    .X(net7115));
 sg13g2_buf_2 fanout7116 (.A(net7117),
    .X(net7116));
 sg13g2_buf_2 fanout7117 (.A(_04057_),
    .X(net7117));
 sg13g2_buf_2 fanout7118 (.A(net7119),
    .X(net7118));
 sg13g2_buf_2 fanout7119 (.A(net7135),
    .X(net7119));
 sg13g2_buf_2 fanout7120 (.A(net7122),
    .X(net7120));
 sg13g2_buf_1 fanout7121 (.A(net7122),
    .X(net7121));
 sg13g2_buf_2 fanout7122 (.A(net7135),
    .X(net7122));
 sg13g2_buf_2 fanout7123 (.A(net7126),
    .X(net7123));
 sg13g2_buf_2 fanout7124 (.A(net7126),
    .X(net7124));
 sg13g2_buf_4 fanout7125 (.X(net7125),
    .A(net7126));
 sg13g2_buf_4 fanout7126 (.X(net7126),
    .A(net7135));
 sg13g2_buf_2 fanout7127 (.A(net7131),
    .X(net7127));
 sg13g2_buf_1 fanout7128 (.A(net7131),
    .X(net7128));
 sg13g2_buf_2 fanout7129 (.A(net7131),
    .X(net7129));
 sg13g2_buf_2 fanout7130 (.A(net7131),
    .X(net7130));
 sg13g2_buf_2 fanout7131 (.A(net7135),
    .X(net7131));
 sg13g2_buf_2 fanout7132 (.A(net7133),
    .X(net7132));
 sg13g2_buf_2 fanout7133 (.A(net7135),
    .X(net7133));
 sg13g2_buf_2 fanout7134 (.A(net7135),
    .X(net7134));
 sg13g2_buf_8 fanout7135 (.A(net7191),
    .X(net7135));
 sg13g2_buf_4 fanout7136 (.X(net7136),
    .A(net7139));
 sg13g2_buf_2 fanout7137 (.A(net7139),
    .X(net7137));
 sg13g2_buf_4 fanout7138 (.X(net7138),
    .A(net7139));
 sg13g2_buf_2 fanout7139 (.A(net7144),
    .X(net7139));
 sg13g2_buf_4 fanout7140 (.X(net7140),
    .A(net7141));
 sg13g2_buf_2 fanout7141 (.A(net7144),
    .X(net7141));
 sg13g2_buf_4 fanout7142 (.X(net7142),
    .A(net7144));
 sg13g2_buf_2 fanout7143 (.A(net7144),
    .X(net7143));
 sg13g2_buf_2 fanout7144 (.A(net7191),
    .X(net7144));
 sg13g2_buf_4 fanout7145 (.X(net7145),
    .A(net7147));
 sg13g2_buf_4 fanout7146 (.X(net7146),
    .A(net7147));
 sg13g2_buf_2 fanout7147 (.A(net7152),
    .X(net7147));
 sg13g2_buf_4 fanout7148 (.X(net7148),
    .A(net7152));
 sg13g2_buf_4 fanout7149 (.X(net7149),
    .A(net7151));
 sg13g2_buf_1 fanout7150 (.A(net7151),
    .X(net7150));
 sg13g2_buf_2 fanout7151 (.A(net7152),
    .X(net7151));
 sg13g2_buf_2 fanout7152 (.A(net7191),
    .X(net7152));
 sg13g2_buf_4 fanout7153 (.X(net7153),
    .A(net7162));
 sg13g2_buf_2 fanout7154 (.A(net7162),
    .X(net7154));
 sg13g2_buf_2 fanout7155 (.A(net7156),
    .X(net7155));
 sg13g2_buf_2 fanout7156 (.A(net7162),
    .X(net7156));
 sg13g2_buf_2 fanout7157 (.A(net7161),
    .X(net7157));
 sg13g2_buf_1 fanout7158 (.A(net7161),
    .X(net7158));
 sg13g2_buf_4 fanout7159 (.X(net7159),
    .A(net7161));
 sg13g2_buf_2 fanout7160 (.A(net7161),
    .X(net7160));
 sg13g2_buf_2 fanout7161 (.A(net7162),
    .X(net7161));
 sg13g2_buf_4 fanout7162 (.X(net7162),
    .A(net7190));
 sg13g2_buf_4 fanout7163 (.X(net7163),
    .A(net7170));
 sg13g2_buf_2 fanout7164 (.A(net7165),
    .X(net7164));
 sg13g2_buf_4 fanout7165 (.X(net7165),
    .A(net7170));
 sg13g2_buf_4 fanout7166 (.X(net7166),
    .A(net7170));
 sg13g2_buf_2 fanout7167 (.A(net7170),
    .X(net7167));
 sg13g2_buf_2 fanout7168 (.A(net7170),
    .X(net7168));
 sg13g2_buf_2 fanout7169 (.A(net7170),
    .X(net7169));
 sg13g2_buf_4 fanout7170 (.X(net7170),
    .A(net7190));
 sg13g2_buf_4 fanout7171 (.X(net7171),
    .A(net7174));
 sg13g2_buf_1 fanout7172 (.A(net7174),
    .X(net7172));
 sg13g2_buf_4 fanout7173 (.X(net7173),
    .A(net7174));
 sg13g2_buf_2 fanout7174 (.A(net7180),
    .X(net7174));
 sg13g2_buf_2 fanout7175 (.A(net7178),
    .X(net7175));
 sg13g2_buf_2 fanout7176 (.A(net7178),
    .X(net7176));
 sg13g2_buf_1 fanout7177 (.A(net7178),
    .X(net7177));
 sg13g2_buf_4 fanout7178 (.X(net7178),
    .A(net7180));
 sg13g2_buf_4 fanout7179 (.X(net7179),
    .A(net7180));
 sg13g2_buf_2 fanout7180 (.A(net7190),
    .X(net7180));
 sg13g2_buf_2 fanout7181 (.A(net7185),
    .X(net7181));
 sg13g2_buf_1 fanout7182 (.A(net7185),
    .X(net7182));
 sg13g2_buf_4 fanout7183 (.X(net7183),
    .A(net7185));
 sg13g2_buf_1 fanout7184 (.A(net7185),
    .X(net7184));
 sg13g2_buf_2 fanout7185 (.A(net7189),
    .X(net7185));
 sg13g2_buf_4 fanout7186 (.X(net7186),
    .A(net7189));
 sg13g2_buf_1 fanout7187 (.A(net7189),
    .X(net7187));
 sg13g2_buf_2 fanout7188 (.A(net7189),
    .X(net7188));
 sg13g2_buf_2 fanout7189 (.A(net7190),
    .X(net7189));
 sg13g2_buf_8 fanout7190 (.A(net7191),
    .X(net7190));
 sg13g2_buf_8 fanout7191 (.A(_02571_),
    .X(net7191));
 sg13g2_buf_2 fanout7192 (.A(net7196),
    .X(net7192));
 sg13g2_buf_1 fanout7193 (.A(net7196),
    .X(net7193));
 sg13g2_buf_2 fanout7194 (.A(net7196),
    .X(net7194));
 sg13g2_buf_2 fanout7195 (.A(net7196),
    .X(net7195));
 sg13g2_buf_2 fanout7196 (.A(net7197),
    .X(net7196));
 sg13g2_buf_4 fanout7197 (.X(net7197),
    .A(net7199));
 sg13g2_buf_4 fanout7198 (.X(net7198),
    .A(net7199));
 sg13g2_buf_8 fanout7199 (.A(_04870_),
    .X(net7199));
 sg13g2_buf_4 fanout7200 (.X(net7200),
    .A(net7201));
 sg13g2_buf_2 fanout7201 (.A(net7202),
    .X(net7201));
 sg13g2_buf_8 fanout7202 (.A(_04870_),
    .X(net7202));
 sg13g2_buf_4 fanout7203 (.X(net7203),
    .A(net7207));
 sg13g2_buf_2 fanout7204 (.A(net7205),
    .X(net7204));
 sg13g2_buf_2 fanout7205 (.A(net7207),
    .X(net7205));
 sg13g2_buf_4 fanout7206 (.X(net7206),
    .A(net7207));
 sg13g2_buf_4 fanout7207 (.X(net7207),
    .A(_04869_));
 sg13g2_buf_4 fanout7208 (.X(net7208),
    .A(net7210));
 sg13g2_buf_2 fanout7209 (.A(net7210),
    .X(net7209));
 sg13g2_buf_2 fanout7210 (.A(net7211),
    .X(net7210));
 sg13g2_buf_4 fanout7211 (.X(net7211),
    .A(net7212));
 sg13g2_buf_1 fanout7212 (.A(_04869_),
    .X(net7212));
 sg13g2_buf_2 fanout7213 (.A(net7216),
    .X(net7213));
 sg13g2_buf_2 fanout7214 (.A(net7216),
    .X(net7214));
 sg13g2_buf_2 fanout7215 (.A(net7216),
    .X(net7215));
 sg13g2_buf_4 fanout7216 (.X(net7216),
    .A(net7227));
 sg13g2_buf_2 fanout7217 (.A(net7219),
    .X(net7217));
 sg13g2_buf_2 fanout7218 (.A(net7219),
    .X(net7218));
 sg13g2_buf_4 fanout7219 (.X(net7219),
    .A(net7220));
 sg13g2_buf_2 fanout7220 (.A(net7227),
    .X(net7220));
 sg13g2_buf_2 fanout7221 (.A(net7225),
    .X(net7221));
 sg13g2_buf_2 fanout7222 (.A(net7224),
    .X(net7222));
 sg13g2_buf_1 fanout7223 (.A(net7224),
    .X(net7223));
 sg13g2_buf_2 fanout7224 (.A(net7225),
    .X(net7224));
 sg13g2_buf_2 fanout7225 (.A(net7226),
    .X(net7225));
 sg13g2_buf_1 fanout7226 (.A(net7227),
    .X(net7226));
 sg13g2_buf_4 fanout7227 (.X(net7227),
    .A(_04869_));
 sg13g2_buf_2 fanout7228 (.A(net7230),
    .X(net7228));
 sg13g2_buf_1 fanout7229 (.A(net7230),
    .X(net7229));
 sg13g2_buf_2 fanout7230 (.A(_04716_),
    .X(net7230));
 sg13g2_buf_2 fanout7231 (.A(net7232),
    .X(net7231));
 sg13g2_buf_1 fanout7232 (.A(net7233),
    .X(net7232));
 sg13g2_buf_2 fanout7233 (.A(_04716_),
    .X(net7233));
 sg13g2_buf_16 fanout7234 (.X(net7234),
    .A(_04291_));
 sg13g2_buf_8 fanout7235 (.A(_04234_),
    .X(net7235));
 sg13g2_buf_8 fanout7236 (.A(_04234_),
    .X(net7236));
 sg13g2_buf_8 fanout7237 (.A(net7239),
    .X(net7237));
 sg13g2_buf_8 fanout7238 (.A(net7239),
    .X(net7238));
 sg13g2_buf_8 fanout7239 (.A(_04216_),
    .X(net7239));
 sg13g2_buf_2 fanout7240 (.A(net7242),
    .X(net7240));
 sg13g2_buf_1 fanout7241 (.A(net7242),
    .X(net7241));
 sg13g2_buf_2 fanout7242 (.A(_04207_),
    .X(net7242));
 sg13g2_buf_2 fanout7243 (.A(net7244),
    .X(net7243));
 sg13g2_buf_2 fanout7244 (.A(_04207_),
    .X(net7244));
 sg13g2_buf_8 fanout7245 (.A(_04198_),
    .X(net7245));
 sg13g2_buf_8 fanout7246 (.A(_04198_),
    .X(net7246));
 sg13g2_buf_16 fanout7247 (.X(net7247),
    .A(_04197_));
 sg13g2_buf_4 fanout7248 (.X(net7248),
    .A(_04197_));
 sg13g2_buf_2 fanout7249 (.A(net7253),
    .X(net7249));
 sg13g2_buf_2 fanout7250 (.A(net7253),
    .X(net7250));
 sg13g2_buf_4 fanout7251 (.X(net7251),
    .A(net7253));
 sg13g2_buf_2 fanout7252 (.A(net7253),
    .X(net7252));
 sg13g2_buf_4 fanout7253 (.X(net7253),
    .A(_04182_));
 sg13g2_buf_2 fanout7254 (.A(net7255),
    .X(net7254));
 sg13g2_buf_2 fanout7255 (.A(net7256),
    .X(net7255));
 sg13g2_buf_4 fanout7256 (.X(net7256),
    .A(_04164_));
 sg13g2_buf_2 fanout7257 (.A(_04164_),
    .X(net7257));
 sg13g2_buf_4 fanout7258 (.X(net7258),
    .A(net7260));
 sg13g2_buf_1 fanout7259 (.A(net7260),
    .X(net7259));
 sg13g2_buf_2 fanout7260 (.A(_04142_),
    .X(net7260));
 sg13g2_buf_2 fanout7261 (.A(net7263),
    .X(net7261));
 sg13g2_buf_1 fanout7262 (.A(net7263),
    .X(net7262));
 sg13g2_buf_2 fanout7263 (.A(_04142_),
    .X(net7263));
 sg13g2_buf_8 fanout7264 (.A(net7266),
    .X(net7264));
 sg13g2_buf_8 fanout7265 (.A(net7266),
    .X(net7265));
 sg13g2_buf_8 fanout7266 (.A(_04140_),
    .X(net7266));
 sg13g2_buf_4 fanout7267 (.X(net7267),
    .A(net7268));
 sg13g2_buf_2 fanout7268 (.A(_04130_),
    .X(net7268));
 sg13g2_buf_4 fanout7269 (.X(net7269),
    .A(_04130_));
 sg13g2_buf_2 fanout7270 (.A(_04130_),
    .X(net7270));
 sg13g2_buf_8 fanout7271 (.A(_04116_),
    .X(net7271));
 sg13g2_buf_8 fanout7272 (.A(_04116_),
    .X(net7272));
 sg13g2_buf_16 fanout7273 (.X(net7273),
    .A(_04115_));
 sg13g2_buf_4 fanout7274 (.X(net7274),
    .A(_04115_));
 sg13g2_buf_8 fanout7275 (.A(_04107_),
    .X(net7275));
 sg13g2_buf_8 fanout7276 (.A(_04107_),
    .X(net7276));
 sg13g2_buf_16 fanout7277 (.X(net7277),
    .A(_04106_));
 sg13g2_buf_4 fanout7278 (.X(net7278),
    .A(_04106_));
 sg13g2_buf_8 fanout7279 (.A(net7280),
    .X(net7279));
 sg13g2_buf_8 fanout7280 (.A(_04092_),
    .X(net7280));
 sg13g2_buf_8 fanout7281 (.A(net7283),
    .X(net7281));
 sg13g2_buf_8 fanout7282 (.A(net7283),
    .X(net7282));
 sg13g2_buf_8 fanout7283 (.A(_04086_),
    .X(net7283));
 sg13g2_buf_8 fanout7284 (.A(_04079_),
    .X(net7284));
 sg13g2_buf_8 fanout7285 (.A(_04078_),
    .X(net7285));
 sg13g2_buf_16 fanout7286 (.X(net7286),
    .A(_04078_));
 sg13g2_buf_2 fanout7287 (.A(net7291),
    .X(net7287));
 sg13g2_buf_1 fanout7288 (.A(net7291),
    .X(net7288));
 sg13g2_buf_2 fanout7289 (.A(net7291),
    .X(net7289));
 sg13g2_buf_2 fanout7290 (.A(net7291),
    .X(net7290));
 sg13g2_buf_2 fanout7291 (.A(net7296),
    .X(net7291));
 sg13g2_buf_2 fanout7292 (.A(net7295),
    .X(net7292));
 sg13g2_buf_1 fanout7293 (.A(net7295),
    .X(net7293));
 sg13g2_buf_2 fanout7294 (.A(net7295),
    .X(net7294));
 sg13g2_buf_4 fanout7295 (.X(net7295),
    .A(net7296));
 sg13g2_buf_2 fanout7296 (.A(net7323),
    .X(net7296));
 sg13g2_buf_2 fanout7297 (.A(net7300),
    .X(net7297));
 sg13g2_buf_4 fanout7298 (.X(net7298),
    .A(net7300));
 sg13g2_buf_1 fanout7299 (.A(net7300),
    .X(net7299));
 sg13g2_buf_2 fanout7300 (.A(net7323),
    .X(net7300));
 sg13g2_buf_2 fanout7301 (.A(net7302),
    .X(net7301));
 sg13g2_buf_2 fanout7302 (.A(net7305),
    .X(net7302));
 sg13g2_buf_4 fanout7303 (.X(net7303),
    .A(net7305));
 sg13g2_buf_2 fanout7304 (.A(net7305),
    .X(net7304));
 sg13g2_buf_2 fanout7305 (.A(net7323),
    .X(net7305));
 sg13g2_buf_4 fanout7306 (.X(net7306),
    .A(net7308));
 sg13g2_buf_1 fanout7307 (.A(net7308),
    .X(net7307));
 sg13g2_buf_4 fanout7308 (.X(net7308),
    .A(net7314));
 sg13g2_buf_2 fanout7309 (.A(net7310),
    .X(net7309));
 sg13g2_buf_2 fanout7310 (.A(net7311),
    .X(net7310));
 sg13g2_buf_2 fanout7311 (.A(net7314),
    .X(net7311));
 sg13g2_buf_4 fanout7312 (.X(net7312),
    .A(net7314));
 sg13g2_buf_1 fanout7313 (.A(net7314),
    .X(net7313));
 sg13g2_buf_4 fanout7314 (.X(net7314),
    .A(net7323));
 sg13g2_buf_4 fanout7315 (.X(net7315),
    .A(net7322));
 sg13g2_buf_4 fanout7316 (.X(net7316),
    .A(net7322));
 sg13g2_buf_4 fanout7317 (.X(net7317),
    .A(net7321));
 sg13g2_buf_1 fanout7318 (.A(net7321),
    .X(net7318));
 sg13g2_buf_2 fanout7319 (.A(net7321),
    .X(net7319));
 sg13g2_buf_1 fanout7320 (.A(net7321),
    .X(net7320));
 sg13g2_buf_2 fanout7321 (.A(net7322),
    .X(net7321));
 sg13g2_buf_2 fanout7322 (.A(net7323),
    .X(net7322));
 sg13g2_buf_8 fanout7323 (.A(_04069_),
    .X(net7323));
 sg13g2_buf_2 fanout7324 (.A(net7326),
    .X(net7324));
 sg13g2_buf_2 fanout7325 (.A(net7326),
    .X(net7325));
 sg13g2_buf_4 fanout7326 (.X(net7326),
    .A(net7332));
 sg13g2_buf_4 fanout7327 (.X(net7327),
    .A(net7331));
 sg13g2_buf_2 fanout7328 (.A(net7331),
    .X(net7328));
 sg13g2_buf_2 fanout7329 (.A(net7331),
    .X(net7329));
 sg13g2_buf_1 fanout7330 (.A(net7331),
    .X(net7330));
 sg13g2_buf_2 fanout7331 (.A(net7332),
    .X(net7331));
 sg13g2_buf_2 fanout7332 (.A(net7360),
    .X(net7332));
 sg13g2_buf_4 fanout7333 (.X(net7333),
    .A(net7336));
 sg13g2_buf_4 fanout7334 (.X(net7334),
    .A(net7336));
 sg13g2_buf_2 fanout7335 (.A(net7336),
    .X(net7335));
 sg13g2_buf_4 fanout7336 (.X(net7336),
    .A(net7360));
 sg13g2_buf_4 fanout7337 (.X(net7337),
    .A(net7340));
 sg13g2_buf_4 fanout7338 (.X(net7338),
    .A(net7340));
 sg13g2_buf_1 fanout7339 (.A(net7340),
    .X(net7339));
 sg13g2_buf_2 fanout7340 (.A(net7360),
    .X(net7340));
 sg13g2_buf_2 fanout7341 (.A(net7345),
    .X(net7341));
 sg13g2_buf_1 fanout7342 (.A(net7345),
    .X(net7342));
 sg13g2_buf_2 fanout7343 (.A(net7345),
    .X(net7343));
 sg13g2_buf_1 fanout7344 (.A(net7345),
    .X(net7344));
 sg13g2_buf_2 fanout7345 (.A(net7360),
    .X(net7345));
 sg13g2_buf_2 fanout7346 (.A(net7350),
    .X(net7346));
 sg13g2_buf_2 fanout7347 (.A(net7350),
    .X(net7347));
 sg13g2_buf_2 fanout7348 (.A(net7350),
    .X(net7348));
 sg13g2_buf_1 fanout7349 (.A(net7350),
    .X(net7349));
 sg13g2_buf_2 fanout7350 (.A(net7360),
    .X(net7350));
 sg13g2_buf_2 fanout7351 (.A(net7353),
    .X(net7351));
 sg13g2_buf_2 fanout7352 (.A(net7359),
    .X(net7352));
 sg13g2_buf_1 fanout7353 (.A(net7359),
    .X(net7353));
 sg13g2_buf_2 fanout7354 (.A(net7359),
    .X(net7354));
 sg13g2_buf_4 fanout7355 (.X(net7355),
    .A(net7356));
 sg13g2_buf_2 fanout7356 (.A(net7359),
    .X(net7356));
 sg13g2_buf_2 fanout7357 (.A(net7358),
    .X(net7357));
 sg13g2_buf_2 fanout7358 (.A(net7359),
    .X(net7358));
 sg13g2_buf_4 fanout7359 (.X(net7359),
    .A(net7360));
 sg13g2_buf_8 fanout7360 (.A(_04069_),
    .X(net7360));
 sg13g2_buf_8 fanout7361 (.A(net7363),
    .X(net7361));
 sg13g2_buf_8 fanout7362 (.A(net7363),
    .X(net7362));
 sg13g2_buf_8 fanout7363 (.A(_04064_),
    .X(net7363));
 sg13g2_buf_4 fanout7364 (.X(net7364),
    .A(net7371));
 sg13g2_buf_2 fanout7365 (.A(net7371),
    .X(net7365));
 sg13g2_buf_4 fanout7366 (.X(net7366),
    .A(net7368));
 sg13g2_buf_2 fanout7367 (.A(net7368),
    .X(net7367));
 sg13g2_buf_2 fanout7368 (.A(net7371),
    .X(net7368));
 sg13g2_buf_8 fanout7369 (.A(net7371),
    .X(net7369));
 sg13g2_buf_4 fanout7370 (.X(net7370),
    .A(net7371));
 sg13g2_buf_8 fanout7371 (.A(_04061_),
    .X(net7371));
 sg13g2_buf_2 fanout7372 (.A(net7373),
    .X(net7372));
 sg13g2_buf_2 fanout7373 (.A(net7374),
    .X(net7373));
 sg13g2_buf_8 fanout7374 (.A(_04061_),
    .X(net7374));
 sg13g2_buf_2 fanout7375 (.A(net7376),
    .X(net7375));
 sg13g2_buf_1 fanout7376 (.A(net7380),
    .X(net7376));
 sg13g2_buf_2 fanout7377 (.A(net7378),
    .X(net7377));
 sg13g2_buf_2 fanout7378 (.A(net7379),
    .X(net7378));
 sg13g2_buf_4 fanout7379 (.X(net7379),
    .A(net7380));
 sg13g2_buf_2 fanout7380 (.A(net7401),
    .X(net7380));
 sg13g2_buf_2 fanout7381 (.A(net7383),
    .X(net7381));
 sg13g2_buf_2 fanout7382 (.A(net7383),
    .X(net7382));
 sg13g2_buf_4 fanout7383 (.X(net7383),
    .A(net7384));
 sg13g2_buf_2 fanout7384 (.A(net7401),
    .X(net7384));
 sg13g2_buf_2 fanout7385 (.A(net7389),
    .X(net7385));
 sg13g2_buf_2 fanout7386 (.A(net7388),
    .X(net7386));
 sg13g2_buf_1 fanout7387 (.A(net7388),
    .X(net7387));
 sg13g2_buf_2 fanout7388 (.A(net7389),
    .X(net7388));
 sg13g2_buf_2 fanout7389 (.A(net7401),
    .X(net7389));
 sg13g2_buf_2 fanout7390 (.A(net7394),
    .X(net7390));
 sg13g2_buf_2 fanout7391 (.A(net7392),
    .X(net7391));
 sg13g2_buf_2 fanout7392 (.A(net7393),
    .X(net7392));
 sg13g2_buf_1 fanout7393 (.A(net7394),
    .X(net7393));
 sg13g2_buf_4 fanout7394 (.X(net7394),
    .A(net7400));
 sg13g2_buf_2 fanout7395 (.A(net7400),
    .X(net7395));
 sg13g2_buf_1 fanout7396 (.A(net7400),
    .X(net7396));
 sg13g2_buf_2 fanout7397 (.A(net7399),
    .X(net7397));
 sg13g2_buf_1 fanout7398 (.A(net7399),
    .X(net7398));
 sg13g2_buf_2 fanout7399 (.A(net7400),
    .X(net7399));
 sg13g2_buf_2 fanout7400 (.A(net7401),
    .X(net7400));
 sg13g2_buf_4 fanout7401 (.X(net7401),
    .A(_04060_));
 sg13g2_buf_8 fanout7402 (.A(_04045_),
    .X(net7402));
 sg13g2_buf_8 fanout7403 (.A(net7404),
    .X(net7403));
 sg13g2_buf_8 fanout7404 (.A(_04044_),
    .X(net7404));
 sg13g2_buf_8 fanout7405 (.A(_04044_),
    .X(net7405));
 sg13g2_buf_4 fanout7406 (.X(net7406),
    .A(net7409));
 sg13g2_buf_8 fanout7407 (.A(net7409),
    .X(net7407));
 sg13g2_buf_8 fanout7408 (.A(net7409),
    .X(net7408));
 sg13g2_buf_8 fanout7409 (.A(_04039_),
    .X(net7409));
 sg13g2_buf_4 fanout7410 (.X(net7410),
    .A(net7412));
 sg13g2_buf_2 fanout7411 (.A(net7412),
    .X(net7411));
 sg13g2_buf_2 fanout7412 (.A(_04036_),
    .X(net7412));
 sg13g2_buf_2 fanout7413 (.A(net7414),
    .X(net7413));
 sg13g2_buf_2 fanout7414 (.A(net7421),
    .X(net7414));
 sg13g2_buf_2 fanout7415 (.A(net7421),
    .X(net7415));
 sg13g2_buf_1 fanout7416 (.A(net7421),
    .X(net7416));
 sg13g2_buf_2 fanout7417 (.A(net7418),
    .X(net7417));
 sg13g2_buf_2 fanout7418 (.A(net7421),
    .X(net7418));
 sg13g2_buf_2 fanout7419 (.A(net7420),
    .X(net7419));
 sg13g2_buf_2 fanout7420 (.A(net7421),
    .X(net7420));
 sg13g2_buf_8 fanout7421 (.A(net7429),
    .X(net7421));
 sg13g2_buf_4 fanout7422 (.X(net7422),
    .A(net7426));
 sg13g2_buf_1 fanout7423 (.A(net7426),
    .X(net7423));
 sg13g2_buf_4 fanout7424 (.X(net7424),
    .A(net7426));
 sg13g2_buf_2 fanout7425 (.A(net7426),
    .X(net7425));
 sg13g2_buf_2 fanout7426 (.A(net7429),
    .X(net7426));
 sg13g2_buf_4 fanout7427 (.X(net7427),
    .A(net7429));
 sg13g2_buf_2 fanout7428 (.A(net7429),
    .X(net7428));
 sg13g2_buf_4 fanout7429 (.X(net7429),
    .A(net7448));
 sg13g2_buf_2 fanout7430 (.A(net7433),
    .X(net7430));
 sg13g2_buf_1 fanout7431 (.A(net7433),
    .X(net7431));
 sg13g2_buf_4 fanout7432 (.X(net7432),
    .A(net7433));
 sg13g2_buf_2 fanout7433 (.A(net7448),
    .X(net7433));
 sg13g2_buf_2 fanout7434 (.A(net7435),
    .X(net7434));
 sg13g2_buf_2 fanout7435 (.A(net7437),
    .X(net7435));
 sg13g2_buf_4 fanout7436 (.X(net7436),
    .A(net7437));
 sg13g2_buf_2 fanout7437 (.A(net7448),
    .X(net7437));
 sg13g2_buf_4 fanout7438 (.X(net7438),
    .A(net7447));
 sg13g2_buf_2 fanout7439 (.A(net7441),
    .X(net7439));
 sg13g2_buf_1 fanout7440 (.A(net7441),
    .X(net7440));
 sg13g2_buf_2 fanout7441 (.A(net7442),
    .X(net7441));
 sg13g2_buf_2 fanout7442 (.A(net7447),
    .X(net7442));
 sg13g2_buf_4 fanout7443 (.X(net7443),
    .A(net7446));
 sg13g2_buf_4 fanout7444 (.X(net7444),
    .A(net7445));
 sg13g2_buf_2 fanout7445 (.A(net7446),
    .X(net7445));
 sg13g2_buf_2 fanout7446 (.A(net7447),
    .X(net7446));
 sg13g2_buf_4 fanout7447 (.X(net7447),
    .A(net7448));
 sg13g2_buf_8 fanout7448 (.A(_02575_),
    .X(net7448));
 sg13g2_buf_2 fanout7449 (.A(net7452),
    .X(net7449));
 sg13g2_buf_1 fanout7450 (.A(net7452),
    .X(net7450));
 sg13g2_buf_4 fanout7451 (.X(net7451),
    .A(net7452));
 sg13g2_buf_2 fanout7452 (.A(net7466),
    .X(net7452));
 sg13g2_buf_2 fanout7453 (.A(net7454),
    .X(net7453));
 sg13g2_buf_2 fanout7454 (.A(net7457),
    .X(net7454));
 sg13g2_buf_1 fanout7455 (.A(net7457),
    .X(net7455));
 sg13g2_buf_4 fanout7456 (.X(net7456),
    .A(net7457));
 sg13g2_buf_4 fanout7457 (.X(net7457),
    .A(net7466));
 sg13g2_buf_2 fanout7458 (.A(net7460),
    .X(net7458));
 sg13g2_buf_1 fanout7459 (.A(net7460),
    .X(net7459));
 sg13g2_buf_2 fanout7460 (.A(net7461),
    .X(net7460));
 sg13g2_buf_2 fanout7461 (.A(net7466),
    .X(net7461));
 sg13g2_buf_2 fanout7462 (.A(net7464),
    .X(net7462));
 sg13g2_buf_1 fanout7463 (.A(net7464),
    .X(net7463));
 sg13g2_buf_2 fanout7464 (.A(net7465),
    .X(net7464));
 sg13g2_buf_4 fanout7465 (.X(net7465),
    .A(net7466));
 sg13g2_buf_8 fanout7466 (.A(net7487),
    .X(net7466));
 sg13g2_buf_4 fanout7467 (.X(net7467),
    .A(net7470));
 sg13g2_buf_1 fanout7468 (.A(net7470),
    .X(net7468));
 sg13g2_buf_4 fanout7469 (.X(net7469),
    .A(net7470));
 sg13g2_buf_2 fanout7470 (.A(net7487),
    .X(net7470));
 sg13g2_buf_2 fanout7471 (.A(net7476),
    .X(net7471));
 sg13g2_buf_1 fanout7472 (.A(net7476),
    .X(net7472));
 sg13g2_buf_2 fanout7473 (.A(net7474),
    .X(net7473));
 sg13g2_buf_4 fanout7474 (.X(net7474),
    .A(net7476));
 sg13g2_buf_1 fanout7475 (.A(net7476),
    .X(net7475));
 sg13g2_buf_2 fanout7476 (.A(net7487),
    .X(net7476));
 sg13g2_buf_2 fanout7477 (.A(net7478),
    .X(net7477));
 sg13g2_buf_4 fanout7478 (.X(net7478),
    .A(net7482));
 sg13g2_buf_1 fanout7479 (.A(net7482),
    .X(net7479));
 sg13g2_buf_4 fanout7480 (.X(net7480),
    .A(net7482));
 sg13g2_buf_2 fanout7481 (.A(net7482),
    .X(net7481));
 sg13g2_buf_1 fanout7482 (.A(net7486),
    .X(net7482));
 sg13g2_buf_2 fanout7483 (.A(net7486),
    .X(net7483));
 sg13g2_buf_1 fanout7484 (.A(net7486),
    .X(net7484));
 sg13g2_buf_4 fanout7485 (.X(net7485),
    .A(net7486));
 sg13g2_buf_2 fanout7486 (.A(net7487),
    .X(net7486));
 sg13g2_buf_4 fanout7487 (.X(net7487),
    .A(_02575_));
 sg13g2_buf_2 fanout7488 (.A(net7490),
    .X(net7488));
 sg13g2_buf_2 fanout7489 (.A(net7490),
    .X(net7489));
 sg13g2_buf_4 fanout7490 (.X(net7490),
    .A(net7494));
 sg13g2_buf_2 fanout7491 (.A(net7492),
    .X(net7491));
 sg13g2_buf_4 fanout7492 (.X(net7492),
    .A(net7494));
 sg13g2_buf_4 fanout7493 (.X(net7493),
    .A(net7494));
 sg13g2_buf_2 fanout7494 (.A(net7522),
    .X(net7494));
 sg13g2_buf_2 fanout7495 (.A(net7499),
    .X(net7495));
 sg13g2_buf_2 fanout7496 (.A(net7499),
    .X(net7496));
 sg13g2_buf_4 fanout7497 (.X(net7497),
    .A(net7499));
 sg13g2_buf_2 fanout7498 (.A(net7499),
    .X(net7498));
 sg13g2_buf_4 fanout7499 (.X(net7499),
    .A(net7522));
 sg13g2_buf_2 fanout7500 (.A(net7503),
    .X(net7500));
 sg13g2_buf_2 fanout7501 (.A(net7503),
    .X(net7501));
 sg13g2_buf_4 fanout7502 (.X(net7502),
    .A(net7503));
 sg13g2_buf_2 fanout7503 (.A(net7522),
    .X(net7503));
 sg13g2_buf_2 fanout7504 (.A(net7508),
    .X(net7504));
 sg13g2_buf_2 fanout7505 (.A(net7508),
    .X(net7505));
 sg13g2_buf_4 fanout7506 (.X(net7506),
    .A(net7507));
 sg13g2_buf_4 fanout7507 (.X(net7507),
    .A(net7508));
 sg13g2_buf_2 fanout7508 (.A(net7513),
    .X(net7508));
 sg13g2_buf_2 fanout7509 (.A(net7513),
    .X(net7509));
 sg13g2_buf_4 fanout7510 (.X(net7510),
    .A(net7512));
 sg13g2_buf_2 fanout7511 (.A(net7512),
    .X(net7511));
 sg13g2_buf_2 fanout7512 (.A(net7513),
    .X(net7512));
 sg13g2_buf_4 fanout7513 (.X(net7513),
    .A(net7522));
 sg13g2_buf_4 fanout7514 (.X(net7514),
    .A(net7521));
 sg13g2_buf_1 fanout7515 (.A(net7521),
    .X(net7515));
 sg13g2_buf_4 fanout7516 (.X(net7516),
    .A(net7521));
 sg13g2_buf_2 fanout7517 (.A(net7518),
    .X(net7517));
 sg13g2_buf_2 fanout7518 (.A(net7521),
    .X(net7518));
 sg13g2_buf_4 fanout7519 (.X(net7519),
    .A(net7520));
 sg13g2_buf_2 fanout7520 (.A(net7521),
    .X(net7520));
 sg13g2_buf_2 fanout7521 (.A(net7522),
    .X(net7521));
 sg13g2_buf_8 fanout7522 (.A(_04073_),
    .X(net7522));
 sg13g2_buf_2 fanout7523 (.A(net7525),
    .X(net7523));
 sg13g2_buf_2 fanout7524 (.A(net7525),
    .X(net7524));
 sg13g2_buf_4 fanout7525 (.X(net7525),
    .A(net7529));
 sg13g2_buf_4 fanout7526 (.X(net7526),
    .A(net7528));
 sg13g2_buf_1 fanout7527 (.A(net7528),
    .X(net7527));
 sg13g2_buf_4 fanout7528 (.X(net7528),
    .A(net7529));
 sg13g2_buf_2 fanout7529 (.A(net7558),
    .X(net7529));
 sg13g2_buf_4 fanout7530 (.X(net7530),
    .A(net7532));
 sg13g2_buf_2 fanout7531 (.A(net7532),
    .X(net7531));
 sg13g2_buf_2 fanout7532 (.A(net7533),
    .X(net7532));
 sg13g2_buf_4 fanout7533 (.X(net7533),
    .A(net7538));
 sg13g2_buf_4 fanout7534 (.X(net7534),
    .A(net7538));
 sg13g2_buf_2 fanout7535 (.A(net7538),
    .X(net7535));
 sg13g2_buf_2 fanout7536 (.A(net7537),
    .X(net7536));
 sg13g2_buf_4 fanout7537 (.X(net7537),
    .A(net7538));
 sg13g2_buf_2 fanout7538 (.A(net7558),
    .X(net7538));
 sg13g2_buf_2 fanout7539 (.A(net7543),
    .X(net7539));
 sg13g2_buf_2 fanout7540 (.A(net7543),
    .X(net7540));
 sg13g2_buf_2 fanout7541 (.A(net7543),
    .X(net7541));
 sg13g2_buf_1 fanout7542 (.A(net7543),
    .X(net7542));
 sg13g2_buf_2 fanout7543 (.A(net7558),
    .X(net7543));
 sg13g2_buf_2 fanout7544 (.A(net7548),
    .X(net7544));
 sg13g2_buf_2 fanout7545 (.A(net7548),
    .X(net7545));
 sg13g2_buf_4 fanout7546 (.X(net7546),
    .A(net7548));
 sg13g2_buf_4 fanout7547 (.X(net7547),
    .A(net7548));
 sg13g2_buf_2 fanout7548 (.A(net7558),
    .X(net7548));
 sg13g2_buf_2 fanout7549 (.A(net7557),
    .X(net7549));
 sg13g2_buf_2 fanout7550 (.A(net7557),
    .X(net7550));
 sg13g2_buf_2 fanout7551 (.A(net7557),
    .X(net7551));
 sg13g2_buf_2 fanout7552 (.A(net7556),
    .X(net7552));
 sg13g2_buf_2 fanout7553 (.A(net7556),
    .X(net7553));
 sg13g2_buf_2 fanout7554 (.A(net7556),
    .X(net7554));
 sg13g2_buf_1 fanout7555 (.A(net7556),
    .X(net7555));
 sg13g2_buf_2 fanout7556 (.A(net7557),
    .X(net7556));
 sg13g2_buf_4 fanout7557 (.X(net7557),
    .A(net7558));
 sg13g2_buf_8 fanout7558 (.A(_04073_),
    .X(net7558));
 sg13g2_buf_2 fanout7559 (.A(net7560),
    .X(net7559));
 sg13g2_buf_4 fanout7560 (.X(net7560),
    .A(\top1.fsm.memorization_completed ));
 sg13g2_buf_4 fanout7561 (.X(net7561),
    .A(net4869));
 sg13g2_buf_4 fanout7562 (.X(net7562),
    .A(\top1.addr_in[6] ));
 sg13g2_buf_2 fanout7563 (.A(net4868),
    .X(net7563));
 sg13g2_buf_4 fanout7564 (.X(net7564),
    .A(\top1.addr_in[1] ));
 sg13g2_buf_4 fanout7565 (.X(net7565),
    .A(net4863));
 sg13g2_buf_4 fanout7566 (.X(net7566),
    .A(net4625));
 sg13g2_buf_2 fanout7567 (.A(net7569),
    .X(net7567));
 sg13g2_buf_1 fanout7568 (.A(net7569),
    .X(net7568));
 sg13g2_buf_4 fanout7569 (.X(net7569),
    .A(net7570));
 sg13g2_buf_2 fanout7570 (.A(net7572),
    .X(net7570));
 sg13g2_buf_2 fanout7571 (.A(net7572),
    .X(net7571));
 sg13g2_buf_2 fanout7572 (.A(\top1.mem_ctl.signal_detected ),
    .X(net7572));
 sg13g2_buf_2 fanout7573 (.A(net7574),
    .X(net7573));
 sg13g2_buf_4 fanout7574 (.X(net7574),
    .A(net7576));
 sg13g2_buf_2 fanout7575 (.A(net7576),
    .X(net7575));
 sg13g2_buf_2 fanout7576 (.A(net7607),
    .X(net7576));
 sg13g2_buf_4 fanout7577 (.X(net7577),
    .A(net7580));
 sg13g2_buf_4 fanout7578 (.X(net7578),
    .A(net7580));
 sg13g2_buf_2 fanout7579 (.A(net7580),
    .X(net7579));
 sg13g2_buf_2 fanout7580 (.A(net7607),
    .X(net7580));
 sg13g2_buf_2 fanout7581 (.A(net7585),
    .X(net7581));
 sg13g2_buf_2 fanout7582 (.A(net7585),
    .X(net7582));
 sg13g2_buf_4 fanout7583 (.X(net7583),
    .A(net7585));
 sg13g2_buf_2 fanout7584 (.A(net7585),
    .X(net7584));
 sg13g2_buf_4 fanout7585 (.X(net7585),
    .A(net7589));
 sg13g2_buf_2 fanout7586 (.A(net7589),
    .X(net7586));
 sg13g2_buf_4 fanout7587 (.X(net7587),
    .A(net7588));
 sg13g2_buf_4 fanout7588 (.X(net7588),
    .A(net7589));
 sg13g2_buf_2 fanout7589 (.A(net7607),
    .X(net7589));
 sg13g2_buf_4 fanout7590 (.X(net7590),
    .A(net7594));
 sg13g2_buf_2 fanout7591 (.A(net7594),
    .X(net7591));
 sg13g2_buf_4 fanout7592 (.X(net7592),
    .A(net7594));
 sg13g2_buf_1 fanout7593 (.A(net7594),
    .X(net7593));
 sg13g2_buf_2 fanout7594 (.A(net7598),
    .X(net7594));
 sg13g2_buf_2 fanout7595 (.A(net7596),
    .X(net7595));
 sg13g2_buf_2 fanout7596 (.A(net7597),
    .X(net7596));
 sg13g2_buf_4 fanout7597 (.X(net7597),
    .A(net7598));
 sg13g2_buf_2 fanout7598 (.A(net7607),
    .X(net7598));
 sg13g2_buf_2 fanout7599 (.A(net7606),
    .X(net7599));
 sg13g2_buf_4 fanout7600 (.X(net7600),
    .A(net7606));
 sg13g2_buf_4 fanout7601 (.X(net7601),
    .A(net7605));
 sg13g2_buf_1 fanout7602 (.A(net7605),
    .X(net7602));
 sg13g2_buf_2 fanout7603 (.A(net7605),
    .X(net7603));
 sg13g2_buf_1 fanout7604 (.A(net7605),
    .X(net7604));
 sg13g2_buf_2 fanout7605 (.A(net7606),
    .X(net7605));
 sg13g2_buf_2 fanout7606 (.A(net7607),
    .X(net7606));
 sg13g2_buf_8 fanout7607 (.A(_02577_),
    .X(net7607));
 sg13g2_buf_2 fanout7608 (.A(net7611),
    .X(net7608));
 sg13g2_buf_1 fanout7609 (.A(net7611),
    .X(net7609));
 sg13g2_buf_4 fanout7610 (.X(net7610),
    .A(net7611));
 sg13g2_buf_4 fanout7611 (.X(net7611),
    .A(net7644));
 sg13g2_buf_2 fanout7612 (.A(net7615),
    .X(net7612));
 sg13g2_buf_4 fanout7613 (.X(net7613),
    .A(net7615));
 sg13g2_buf_2 fanout7614 (.A(net7615),
    .X(net7614));
 sg13g2_buf_4 fanout7615 (.X(net7615),
    .A(net7644));
 sg13g2_buf_2 fanout7616 (.A(net7617),
    .X(net7616));
 sg13g2_buf_2 fanout7617 (.A(net7625),
    .X(net7617));
 sg13g2_buf_2 fanout7618 (.A(net7625),
    .X(net7618));
 sg13g2_buf_1 fanout7619 (.A(net7625),
    .X(net7619));
 sg13g2_buf_4 fanout7620 (.X(net7620),
    .A(net7622));
 sg13g2_buf_2 fanout7621 (.A(net7622),
    .X(net7621));
 sg13g2_buf_2 fanout7622 (.A(net7625),
    .X(net7622));
 sg13g2_buf_2 fanout7623 (.A(net7625),
    .X(net7623));
 sg13g2_buf_4 fanout7624 (.X(net7624),
    .A(net7625));
 sg13g2_buf_4 fanout7625 (.X(net7625),
    .A(net7644));
 sg13g2_buf_4 fanout7626 (.X(net7626),
    .A(net7630));
 sg13g2_buf_2 fanout7627 (.A(net7630),
    .X(net7627));
 sg13g2_buf_4 fanout7628 (.X(net7628),
    .A(net7630));
 sg13g2_buf_1 fanout7629 (.A(net7630),
    .X(net7629));
 sg13g2_buf_2 fanout7630 (.A(net7635),
    .X(net7630));
 sg13g2_buf_2 fanout7631 (.A(net7635),
    .X(net7631));
 sg13g2_buf_1 fanout7632 (.A(net7635),
    .X(net7632));
 sg13g2_buf_2 fanout7633 (.A(net7634),
    .X(net7633));
 sg13g2_buf_2 fanout7634 (.A(net7635),
    .X(net7634));
 sg13g2_buf_2 fanout7635 (.A(net7643),
    .X(net7635));
 sg13g2_buf_4 fanout7636 (.X(net7636),
    .A(net7638));
 sg13g2_buf_4 fanout7637 (.X(net7637),
    .A(net7638));
 sg13g2_buf_2 fanout7638 (.A(net7643),
    .X(net7638));
 sg13g2_buf_2 fanout7639 (.A(net7640),
    .X(net7639));
 sg13g2_buf_4 fanout7640 (.X(net7640),
    .A(net7641));
 sg13g2_buf_4 fanout7641 (.X(net7641),
    .A(net7643));
 sg13g2_buf_1 fanout7642 (.A(net7643),
    .X(net7642));
 sg13g2_buf_4 fanout7643 (.X(net7643),
    .A(net7644));
 sg13g2_buf_2 fanout7644 (.A(_02577_),
    .X(net7644));
 sg13g2_buf_4 fanout7645 (.X(net7645),
    .A(net7646));
 sg13g2_buf_4 fanout7646 (.X(net7646),
    .A(net7654));
 sg13g2_buf_2 fanout7647 (.A(net7654),
    .X(net7647));
 sg13g2_buf_2 fanout7648 (.A(net7654),
    .X(net7648));
 sg13g2_buf_4 fanout7649 (.X(net7649),
    .A(net7653));
 sg13g2_buf_2 fanout7650 (.A(net7653),
    .X(net7650));
 sg13g2_buf_2 fanout7651 (.A(net7653),
    .X(net7651));
 sg13g2_buf_1 fanout7652 (.A(net7653),
    .X(net7652));
 sg13g2_buf_4 fanout7653 (.X(net7653),
    .A(net7654));
 sg13g2_buf_2 fanout7654 (.A(net7662),
    .X(net7654));
 sg13g2_buf_2 fanout7655 (.A(net7659),
    .X(net7655));
 sg13g2_buf_1 fanout7656 (.A(net7659),
    .X(net7656));
 sg13g2_buf_2 fanout7657 (.A(net7659),
    .X(net7657));
 sg13g2_buf_2 fanout7658 (.A(net7659),
    .X(net7658));
 sg13g2_buf_2 fanout7659 (.A(net7662),
    .X(net7659));
 sg13g2_buf_2 fanout7660 (.A(net7662),
    .X(net7660));
 sg13g2_buf_4 fanout7661 (.X(net7661),
    .A(net7662));
 sg13g2_buf_4 fanout7662 (.X(net7662),
    .A(net7717));
 sg13g2_buf_2 fanout7663 (.A(net7664),
    .X(net7663));
 sg13g2_buf_2 fanout7664 (.A(net7665),
    .X(net7664));
 sg13g2_buf_4 fanout7665 (.X(net7665),
    .A(net7679));
 sg13g2_buf_2 fanout7666 (.A(net7668),
    .X(net7666));
 sg13g2_buf_1 fanout7667 (.A(net7668),
    .X(net7667));
 sg13g2_buf_2 fanout7668 (.A(net7669),
    .X(net7668));
 sg13g2_buf_4 fanout7669 (.X(net7669),
    .A(net7679));
 sg13g2_buf_4 fanout7670 (.X(net7670),
    .A(net7674));
 sg13g2_buf_4 fanout7671 (.X(net7671),
    .A(net7672));
 sg13g2_buf_2 fanout7672 (.A(net7673),
    .X(net7672));
 sg13g2_buf_2 fanout7673 (.A(net7674),
    .X(net7673));
 sg13g2_buf_2 fanout7674 (.A(net7678),
    .X(net7674));
 sg13g2_buf_2 fanout7675 (.A(net7678),
    .X(net7675));
 sg13g2_buf_2 fanout7676 (.A(net7678),
    .X(net7676));
 sg13g2_buf_2 fanout7677 (.A(net7678),
    .X(net7677));
 sg13g2_buf_2 fanout7678 (.A(net7679),
    .X(net7678));
 sg13g2_buf_2 fanout7679 (.A(net7717),
    .X(net7679));
 sg13g2_buf_2 fanout7680 (.A(net7683),
    .X(net7680));
 sg13g2_buf_2 fanout7681 (.A(net7683),
    .X(net7681));
 sg13g2_buf_2 fanout7682 (.A(net7683),
    .X(net7682));
 sg13g2_buf_2 fanout7683 (.A(net7699),
    .X(net7683));
 sg13g2_buf_2 fanout7684 (.A(net7688),
    .X(net7684));
 sg13g2_buf_1 fanout7685 (.A(net7688),
    .X(net7685));
 sg13g2_buf_2 fanout7686 (.A(net7687),
    .X(net7686));
 sg13g2_buf_2 fanout7687 (.A(net7688),
    .X(net7687));
 sg13g2_buf_2 fanout7688 (.A(net7699),
    .X(net7688));
 sg13g2_buf_2 fanout7689 (.A(net7693),
    .X(net7689));
 sg13g2_buf_1 fanout7690 (.A(net7693),
    .X(net7690));
 sg13g2_buf_4 fanout7691 (.X(net7691),
    .A(net7692));
 sg13g2_buf_4 fanout7692 (.X(net7692),
    .A(net7693));
 sg13g2_buf_2 fanout7693 (.A(net7699),
    .X(net7693));
 sg13g2_buf_4 fanout7694 (.X(net7694),
    .A(net7698));
 sg13g2_buf_1 fanout7695 (.A(net7698),
    .X(net7695));
 sg13g2_buf_2 fanout7696 (.A(net7698),
    .X(net7696));
 sg13g2_buf_1 fanout7697 (.A(net7698),
    .X(net7697));
 sg13g2_buf_2 fanout7698 (.A(net7699),
    .X(net7698));
 sg13g2_buf_4 fanout7699 (.X(net7699),
    .A(net7717));
 sg13g2_buf_4 fanout7700 (.X(net7700),
    .A(net7702));
 sg13g2_buf_1 fanout7701 (.A(net7702),
    .X(net7701));
 sg13g2_buf_4 fanout7702 (.X(net7702),
    .A(net7708));
 sg13g2_buf_2 fanout7703 (.A(net7708),
    .X(net7703));
 sg13g2_buf_1 fanout7704 (.A(net7708),
    .X(net7704));
 sg13g2_buf_2 fanout7705 (.A(net7707),
    .X(net7705));
 sg13g2_buf_2 fanout7706 (.A(net7707),
    .X(net7706));
 sg13g2_buf_2 fanout7707 (.A(net7708),
    .X(net7707));
 sg13g2_buf_4 fanout7708 (.X(net7708),
    .A(net7717));
 sg13g2_buf_4 fanout7709 (.X(net7709),
    .A(net7712));
 sg13g2_buf_2 fanout7710 (.A(net7712),
    .X(net7710));
 sg13g2_buf_2 fanout7711 (.A(net7712),
    .X(net7711));
 sg13g2_buf_2 fanout7712 (.A(net7716),
    .X(net7712));
 sg13g2_buf_4 fanout7713 (.X(net7713),
    .A(net7716));
 sg13g2_buf_4 fanout7714 (.X(net7714),
    .A(net7715));
 sg13g2_buf_2 fanout7715 (.A(net7716),
    .X(net7715));
 sg13g2_buf_4 fanout7716 (.X(net7716),
    .A(net7717));
 sg13g2_buf_8 fanout7717 (.A(_04075_),
    .X(net7717));
 sg13g2_buf_2 fanout7718 (.A(net7719),
    .X(net7718));
 sg13g2_buf_2 fanout7719 (.A(net8),
    .X(net7719));
 sg13g2_buf_2 fanout7720 (.A(net7721),
    .X(net7720));
 sg13g2_buf_1 fanout7721 (.A(net7722),
    .X(net7721));
 sg13g2_buf_2 fanout7722 (.A(net8),
    .X(net7722));
 sg13g2_buf_4 fanout7723 (.X(net7723),
    .A(net7724));
 sg13g2_buf_4 fanout7724 (.X(net7724),
    .A(net7725));
 sg13g2_buf_4 fanout7725 (.X(net7725),
    .A(net7731));
 sg13g2_buf_4 fanout7726 (.X(net7726),
    .A(net7728));
 sg13g2_buf_2 fanout7727 (.A(net7728),
    .X(net7727));
 sg13g2_buf_4 fanout7728 (.X(net7728),
    .A(net7731));
 sg13g2_buf_4 fanout7729 (.X(net7729),
    .A(net7730));
 sg13g2_buf_2 fanout7730 (.A(net7731),
    .X(net7730));
 sg13g2_buf_2 fanout7731 (.A(net7741),
    .X(net7731));
 sg13g2_buf_4 fanout7732 (.X(net7732),
    .A(net7733));
 sg13g2_buf_2 fanout7733 (.A(net7740),
    .X(net7733));
 sg13g2_buf_4 fanout7734 (.X(net7734),
    .A(net7740));
 sg13g2_buf_4 fanout7735 (.X(net7735),
    .A(net7736));
 sg13g2_buf_4 fanout7736 (.X(net7736),
    .A(net7739));
 sg13g2_buf_4 fanout7737 (.X(net7737),
    .A(net7739));
 sg13g2_buf_2 fanout7738 (.A(net7739),
    .X(net7738));
 sg13g2_buf_2 fanout7739 (.A(net7740),
    .X(net7739));
 sg13g2_buf_2 fanout7740 (.A(net7741),
    .X(net7740));
 sg13g2_buf_4 fanout7741 (.X(net7741),
    .A(net7750));
 sg13g2_buf_4 fanout7742 (.X(net7742),
    .A(net7743));
 sg13g2_buf_2 fanout7743 (.A(net7749),
    .X(net7743));
 sg13g2_buf_4 fanout7744 (.X(net7744),
    .A(net7747));
 sg13g2_buf_4 fanout7745 (.X(net7745),
    .A(net7747));
 sg13g2_buf_4 fanout7746 (.X(net7746),
    .A(net7747));
 sg13g2_buf_4 fanout7747 (.X(net7747),
    .A(net7748));
 sg13g2_buf_2 fanout7748 (.A(net7749),
    .X(net7748));
 sg13g2_buf_4 fanout7749 (.X(net7749),
    .A(net7750));
 sg13g2_buf_4 fanout7750 (.X(net7750),
    .A(rst_n));
 sg13g2_buf_8 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_8 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_8 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_8 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_8 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_8 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_8 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_8 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_8 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_8 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_8 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_8 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_8 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_8 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_2 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tielo tt_um_Coline3003_spect_top_17 (.L_LO(net17));
 sg13g2_buf_2 \clkbuf_leaf_1_top1.acquisition_clk  (.A(\clknet_6_0_0_top1.acquisition_clk ),
    .X(\clknet_leaf_1_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_2_top1.acquisition_clk  (.A(\clknet_6_1_0_top1.acquisition_clk ),
    .X(\clknet_leaf_2_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_3_top1.acquisition_clk  (.A(\clknet_6_1_0_top1.acquisition_clk ),
    .X(\clknet_leaf_3_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_4_top1.acquisition_clk  (.A(\clknet_6_1_0_top1.acquisition_clk ),
    .X(\clknet_leaf_4_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_5_top1.acquisition_clk  (.A(\clknet_6_1_0_top1.acquisition_clk ),
    .X(\clknet_leaf_5_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_6_top1.acquisition_clk  (.A(\clknet_6_3_0_top1.acquisition_clk ),
    .X(\clknet_leaf_6_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_7_top1.acquisition_clk  (.A(\clknet_6_3_0_top1.acquisition_clk ),
    .X(\clknet_leaf_7_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_8_top1.acquisition_clk  (.A(\clknet_6_3_0_top1.acquisition_clk ),
    .X(\clknet_leaf_8_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_9_top1.acquisition_clk  (.A(\clknet_6_6_0_top1.acquisition_clk ),
    .X(\clknet_leaf_9_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_10_top1.acquisition_clk  (.A(\clknet_6_6_0_top1.acquisition_clk ),
    .X(\clknet_leaf_10_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_11_top1.acquisition_clk  (.A(\clknet_6_4_0_top1.acquisition_clk ),
    .X(\clknet_leaf_11_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_12_top1.acquisition_clk  (.A(\clknet_6_4_0_top1.acquisition_clk ),
    .X(\clknet_leaf_12_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_13_top1.acquisition_clk  (.A(\clknet_6_1_0_top1.acquisition_clk ),
    .X(\clknet_leaf_13_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_14_top1.acquisition_clk  (.A(\clknet_6_4_0_top1.acquisition_clk ),
    .X(\clknet_leaf_14_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_15_top1.acquisition_clk  (.A(\clknet_6_4_0_top1.acquisition_clk ),
    .X(\clknet_leaf_15_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_16_top1.acquisition_clk  (.A(\clknet_6_4_0_top1.acquisition_clk ),
    .X(\clknet_leaf_16_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_17_top1.acquisition_clk  (.A(\clknet_6_5_0_top1.acquisition_clk ),
    .X(\clknet_leaf_17_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_18_top1.acquisition_clk  (.A(\clknet_6_5_0_top1.acquisition_clk ),
    .X(\clknet_leaf_18_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_19_top1.acquisition_clk  (.A(\clknet_6_5_0_top1.acquisition_clk ),
    .X(\clknet_leaf_19_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_20_top1.acquisition_clk  (.A(\clknet_6_5_0_top1.acquisition_clk ),
    .X(\clknet_leaf_20_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_21_top1.acquisition_clk  (.A(\clknet_6_5_0_top1.acquisition_clk ),
    .X(\clknet_leaf_21_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_22_top1.acquisition_clk  (.A(\clknet_6_7_0_top1.acquisition_clk ),
    .X(\clknet_leaf_22_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_23_top1.acquisition_clk  (.A(\clknet_6_7_0_top1.acquisition_clk ),
    .X(\clknet_leaf_23_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_24_top1.acquisition_clk  (.A(\clknet_6_7_0_top1.acquisition_clk ),
    .X(\clknet_leaf_24_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_25_top1.acquisition_clk  (.A(\clknet_6_7_0_top1.acquisition_clk ),
    .X(\clknet_leaf_25_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_26_top1.acquisition_clk  (.A(\clknet_6_6_0_top1.acquisition_clk ),
    .X(\clknet_leaf_26_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_27_top1.acquisition_clk  (.A(\clknet_6_6_0_top1.acquisition_clk ),
    .X(\clknet_leaf_27_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_28_top1.acquisition_clk  (.A(\clknet_6_6_0_top1.acquisition_clk ),
    .X(\clknet_leaf_28_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_29_top1.acquisition_clk  (.A(\clknet_6_12_0_top1.acquisition_clk ),
    .X(\clknet_leaf_29_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_30_top1.acquisition_clk  (.A(\clknet_6_12_0_top1.acquisition_clk ),
    .X(\clknet_leaf_30_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_31_top1.acquisition_clk  (.A(\clknet_6_13_0_top1.acquisition_clk ),
    .X(\clknet_leaf_31_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_32_top1.acquisition_clk  (.A(\clknet_6_12_0_top1.acquisition_clk ),
    .X(\clknet_leaf_32_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_33_top1.acquisition_clk  (.A(\clknet_6_24_0_top1.acquisition_clk ),
    .X(\clknet_leaf_33_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_34_top1.acquisition_clk  (.A(\clknet_6_24_0_top1.acquisition_clk ),
    .X(\clknet_leaf_34_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_35_top1.acquisition_clk  (.A(\clknet_6_24_0_top1.acquisition_clk ),
    .X(\clknet_leaf_35_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_36_top1.acquisition_clk  (.A(\clknet_6_24_0_top1.acquisition_clk ),
    .X(\clknet_leaf_36_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_37_top1.acquisition_clk  (.A(\clknet_6_26_0_top1.acquisition_clk ),
    .X(\clknet_leaf_37_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_38_top1.acquisition_clk  (.A(\clknet_6_25_0_top1.acquisition_clk ),
    .X(\clknet_leaf_38_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_39_top1.acquisition_clk  (.A(\clknet_6_24_0_top1.acquisition_clk ),
    .X(\clknet_leaf_39_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_40_top1.acquisition_clk  (.A(\clknet_6_25_0_top1.acquisition_clk ),
    .X(\clknet_leaf_40_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_41_top1.acquisition_clk  (.A(\clknet_6_25_0_top1.acquisition_clk ),
    .X(\clknet_leaf_41_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_42_top1.acquisition_clk  (.A(\clknet_6_19_0_top1.acquisition_clk ),
    .X(\clknet_leaf_42_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_43_top1.acquisition_clk  (.A(\clknet_6_18_0_top1.acquisition_clk ),
    .X(\clknet_leaf_43_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_44_top1.acquisition_clk  (.A(\clknet_6_17_0_top1.acquisition_clk ),
    .X(\clknet_leaf_44_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_45_top1.acquisition_clk  (.A(\clknet_6_18_0_top1.acquisition_clk ),
    .X(\clknet_leaf_45_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_46_top1.acquisition_clk  (.A(\clknet_6_18_0_top1.acquisition_clk ),
    .X(\clknet_leaf_46_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_47_top1.acquisition_clk  (.A(\clknet_6_18_0_top1.acquisition_clk ),
    .X(\clknet_leaf_47_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_48_top1.acquisition_clk  (.A(\clknet_6_18_0_top1.acquisition_clk ),
    .X(\clknet_leaf_48_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_49_top1.acquisition_clk  (.A(\clknet_6_16_0_top1.acquisition_clk ),
    .X(\clknet_leaf_49_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_50_top1.acquisition_clk  (.A(\clknet_6_16_0_top1.acquisition_clk ),
    .X(\clknet_leaf_50_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_51_top1.acquisition_clk  (.A(\clknet_6_16_0_top1.acquisition_clk ),
    .X(\clknet_leaf_51_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_52_top1.acquisition_clk  (.A(\clknet_6_16_0_top1.acquisition_clk ),
    .X(\clknet_leaf_52_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_53_top1.acquisition_clk  (.A(\clknet_6_16_0_top1.acquisition_clk ),
    .X(\clknet_leaf_53_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_54_top1.acquisition_clk  (.A(\clknet_6_17_0_top1.acquisition_clk ),
    .X(\clknet_leaf_54_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_55_top1.acquisition_clk  (.A(\clknet_6_17_0_top1.acquisition_clk ),
    .X(\clknet_leaf_55_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_56_top1.acquisition_clk  (.A(\clknet_6_17_0_top1.acquisition_clk ),
    .X(\clknet_leaf_56_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_57_top1.acquisition_clk  (.A(\clknet_6_17_0_top1.acquisition_clk ),
    .X(\clknet_leaf_57_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_58_top1.acquisition_clk  (.A(\clknet_6_19_0_top1.acquisition_clk ),
    .X(\clknet_leaf_58_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_59_top1.acquisition_clk  (.A(\clknet_6_19_0_top1.acquisition_clk ),
    .X(\clknet_leaf_59_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_60_top1.acquisition_clk  (.A(\clknet_6_20_0_top1.acquisition_clk ),
    .X(\clknet_leaf_60_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_61_top1.acquisition_clk  (.A(\clknet_6_20_0_top1.acquisition_clk ),
    .X(\clknet_leaf_61_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_62_top1.acquisition_clk  (.A(\clknet_6_20_0_top1.acquisition_clk ),
    .X(\clknet_leaf_62_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_63_top1.acquisition_clk  (.A(\clknet_6_20_0_top1.acquisition_clk ),
    .X(\clknet_leaf_63_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_64_top1.acquisition_clk  (.A(\clknet_6_20_0_top1.acquisition_clk ),
    .X(\clknet_leaf_64_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_65_top1.acquisition_clk  (.A(\clknet_6_21_0_top1.acquisition_clk ),
    .X(\clknet_leaf_65_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_66_top1.acquisition_clk  (.A(\clknet_6_21_0_top1.acquisition_clk ),
    .X(\clknet_leaf_66_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_67_top1.acquisition_clk  (.A(\clknet_6_21_0_top1.acquisition_clk ),
    .X(\clknet_leaf_67_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_68_top1.acquisition_clk  (.A(\clknet_6_21_0_top1.acquisition_clk ),
    .X(\clknet_leaf_68_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_69_top1.acquisition_clk  (.A(\clknet_6_21_0_top1.acquisition_clk ),
    .X(\clknet_leaf_69_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_70_top1.acquisition_clk  (.A(\clknet_6_23_0_top1.acquisition_clk ),
    .X(\clknet_leaf_70_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_71_top1.acquisition_clk  (.A(\clknet_6_23_0_top1.acquisition_clk ),
    .X(\clknet_leaf_71_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_72_top1.acquisition_clk  (.A(\clknet_6_23_0_top1.acquisition_clk ),
    .X(\clknet_leaf_72_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_73_top1.acquisition_clk  (.A(\clknet_6_22_0_top1.acquisition_clk ),
    .X(\clknet_leaf_73_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_74_top1.acquisition_clk  (.A(\clknet_6_22_0_top1.acquisition_clk ),
    .X(\clknet_leaf_74_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_75_top1.acquisition_clk  (.A(\clknet_6_22_0_top1.acquisition_clk ),
    .X(\clknet_leaf_75_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_76_top1.acquisition_clk  (.A(\clknet_6_22_0_top1.acquisition_clk ),
    .X(\clknet_leaf_76_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_77_top1.acquisition_clk  (.A(\clknet_6_22_0_top1.acquisition_clk ),
    .X(\clknet_leaf_77_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_78_top1.acquisition_clk  (.A(\clknet_6_29_0_top1.acquisition_clk ),
    .X(\clknet_leaf_78_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_79_top1.acquisition_clk  (.A(\clknet_6_29_0_top1.acquisition_clk ),
    .X(\clknet_leaf_79_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_80_top1.acquisition_clk  (.A(\clknet_6_29_0_top1.acquisition_clk ),
    .X(\clknet_leaf_80_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_81_top1.acquisition_clk  (.A(\clknet_6_23_0_top1.acquisition_clk ),
    .X(\clknet_leaf_81_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_82_top1.acquisition_clk  (.A(\clknet_6_29_0_top1.acquisition_clk ),
    .X(\clknet_leaf_82_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_83_top1.acquisition_clk  (.A(\clknet_6_28_0_top1.acquisition_clk ),
    .X(\clknet_leaf_83_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_84_top1.acquisition_clk  (.A(\clknet_6_28_0_top1.acquisition_clk ),
    .X(\clknet_leaf_84_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_85_top1.acquisition_clk  (.A(\clknet_6_31_0_top1.acquisition_clk ),
    .X(\clknet_leaf_85_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_86_top1.acquisition_clk  (.A(\clknet_6_31_0_top1.acquisition_clk ),
    .X(\clknet_leaf_86_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_87_top1.acquisition_clk  (.A(\clknet_6_31_0_top1.acquisition_clk ),
    .X(\clknet_leaf_87_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_88_top1.acquisition_clk  (.A(\clknet_6_31_0_top1.acquisition_clk ),
    .X(\clknet_leaf_88_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_89_top1.acquisition_clk  (.A(\clknet_6_30_0_top1.acquisition_clk ),
    .X(\clknet_leaf_89_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_90_top1.acquisition_clk  (.A(\clknet_6_28_0_top1.acquisition_clk ),
    .X(\clknet_leaf_90_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_91_top1.acquisition_clk  (.A(\clknet_6_30_0_top1.acquisition_clk ),
    .X(\clknet_leaf_91_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_92_top1.acquisition_clk  (.A(\clknet_6_30_0_top1.acquisition_clk ),
    .X(\clknet_leaf_92_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_93_top1.acquisition_clk  (.A(\clknet_6_30_0_top1.acquisition_clk ),
    .X(\clknet_leaf_93_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_94_top1.acquisition_clk  (.A(\clknet_6_28_0_top1.acquisition_clk ),
    .X(\clknet_leaf_94_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_95_top1.acquisition_clk  (.A(\clknet_6_28_0_top1.acquisition_clk ),
    .X(\clknet_leaf_95_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_96_top1.acquisition_clk  (.A(\clknet_6_29_0_top1.acquisition_clk ),
    .X(\clknet_leaf_96_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_97_top1.acquisition_clk  (.A(\clknet_6_19_0_top1.acquisition_clk ),
    .X(\clknet_leaf_97_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_98_top1.acquisition_clk  (.A(\clknet_6_25_0_top1.acquisition_clk ),
    .X(\clknet_leaf_98_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_99_top1.acquisition_clk  (.A(\clknet_6_25_0_top1.acquisition_clk ),
    .X(\clknet_leaf_99_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_100_top1.acquisition_clk  (.A(\clknet_6_27_0_top1.acquisition_clk ),
    .X(\clknet_leaf_100_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_101_top1.acquisition_clk  (.A(\clknet_6_30_0_top1.acquisition_clk ),
    .X(\clknet_leaf_101_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_102_top1.acquisition_clk  (.A(\clknet_6_27_0_top1.acquisition_clk ),
    .X(\clknet_leaf_102_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_103_top1.acquisition_clk  (.A(\clknet_6_27_0_top1.acquisition_clk ),
    .X(\clknet_leaf_103_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_104_top1.acquisition_clk  (.A(\clknet_6_27_0_top1.acquisition_clk ),
    .X(\clknet_leaf_104_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_105_top1.acquisition_clk  (.A(\clknet_6_26_0_top1.acquisition_clk ),
    .X(\clknet_leaf_105_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_106_top1.acquisition_clk  (.A(\clknet_6_26_0_top1.acquisition_clk ),
    .X(\clknet_leaf_106_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_107_top1.acquisition_clk  (.A(\clknet_6_26_0_top1.acquisition_clk ),
    .X(\clknet_leaf_107_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_108_top1.acquisition_clk  (.A(\clknet_6_49_0_top1.acquisition_clk ),
    .X(\clknet_leaf_108_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_109_top1.acquisition_clk  (.A(\clknet_6_49_0_top1.acquisition_clk ),
    .X(\clknet_leaf_109_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_110_top1.acquisition_clk  (.A(\clknet_6_49_0_top1.acquisition_clk ),
    .X(\clknet_leaf_110_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_111_top1.acquisition_clk  (.A(\clknet_6_49_0_top1.acquisition_clk ),
    .X(\clknet_leaf_111_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_112_top1.acquisition_clk  (.A(\clknet_6_49_0_top1.acquisition_clk ),
    .X(\clknet_leaf_112_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_113_top1.acquisition_clk  (.A(\clknet_6_48_0_top1.acquisition_clk ),
    .X(\clknet_leaf_113_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_114_top1.acquisition_clk  (.A(\clknet_6_48_0_top1.acquisition_clk ),
    .X(\clknet_leaf_114_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_115_top1.acquisition_clk  (.A(\clknet_6_48_0_top1.acquisition_clk ),
    .X(\clknet_leaf_115_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_116_top1.acquisition_clk  (.A(\clknet_6_51_0_top1.acquisition_clk ),
    .X(\clknet_leaf_116_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_117_top1.acquisition_clk  (.A(\clknet_6_51_0_top1.acquisition_clk ),
    .X(\clknet_leaf_117_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_118_top1.acquisition_clk  (.A(\clknet_6_51_0_top1.acquisition_clk ),
    .X(\clknet_leaf_118_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_119_top1.acquisition_clk  (.A(\clknet_6_52_0_top1.acquisition_clk ),
    .X(\clknet_leaf_119_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_120_top1.acquisition_clk  (.A(\clknet_6_52_0_top1.acquisition_clk ),
    .X(\clknet_leaf_120_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_121_top1.acquisition_clk  (.A(\clknet_6_52_0_top1.acquisition_clk ),
    .X(\clknet_leaf_121_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_122_top1.acquisition_clk  (.A(\clknet_6_52_0_top1.acquisition_clk ),
    .X(\clknet_leaf_122_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_123_top1.acquisition_clk  (.A(\clknet_6_52_0_top1.acquisition_clk ),
    .X(\clknet_leaf_123_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_124_top1.acquisition_clk  (.A(\clknet_6_53_0_top1.acquisition_clk ),
    .X(\clknet_leaf_124_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_125_top1.acquisition_clk  (.A(\clknet_6_53_0_top1.acquisition_clk ),
    .X(\clknet_leaf_125_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_126_top1.acquisition_clk  (.A(\clknet_6_53_0_top1.acquisition_clk ),
    .X(\clknet_leaf_126_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_127_top1.acquisition_clk  (.A(\clknet_6_53_0_top1.acquisition_clk ),
    .X(\clknet_leaf_127_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_128_top1.acquisition_clk  (.A(\clknet_6_53_0_top1.acquisition_clk ),
    .X(\clknet_leaf_128_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_129_top1.acquisition_clk  (.A(\clknet_6_55_0_top1.acquisition_clk ),
    .X(\clknet_leaf_129_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_130_top1.acquisition_clk  (.A(\clknet_6_55_0_top1.acquisition_clk ),
    .X(\clknet_leaf_130_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_131_top1.acquisition_clk  (.A(\clknet_6_55_0_top1.acquisition_clk ),
    .X(\clknet_leaf_131_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_132_top1.acquisition_clk  (.A(\clknet_6_55_0_top1.acquisition_clk ),
    .X(\clknet_leaf_132_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_133_top1.acquisition_clk  (.A(\clknet_6_54_0_top1.acquisition_clk ),
    .X(\clknet_leaf_133_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_134_top1.acquisition_clk  (.A(\clknet_6_54_0_top1.acquisition_clk ),
    .X(\clknet_leaf_134_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_135_top1.acquisition_clk  (.A(\clknet_6_54_0_top1.acquisition_clk ),
    .X(\clknet_leaf_135_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_136_top1.acquisition_clk  (.A(\clknet_6_54_0_top1.acquisition_clk ),
    .X(\clknet_leaf_136_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_137_top1.acquisition_clk  (.A(\clknet_6_54_0_top1.acquisition_clk ),
    .X(\clknet_leaf_137_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_138_top1.acquisition_clk  (.A(\clknet_6_60_0_top1.acquisition_clk ),
    .X(\clknet_leaf_138_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_139_top1.acquisition_clk  (.A(\clknet_6_60_0_top1.acquisition_clk ),
    .X(\clknet_leaf_139_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_140_top1.acquisition_clk  (.A(\clknet_6_60_0_top1.acquisition_clk ),
    .X(\clknet_leaf_140_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_141_top1.acquisition_clk  (.A(\clknet_6_61_0_top1.acquisition_clk ),
    .X(\clknet_leaf_141_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_142_top1.acquisition_clk  (.A(\clknet_6_61_0_top1.acquisition_clk ),
    .X(\clknet_leaf_142_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_143_top1.acquisition_clk  (.A(\clknet_6_61_0_top1.acquisition_clk ),
    .X(\clknet_leaf_143_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_144_top1.acquisition_clk  (.A(\clknet_6_61_0_top1.acquisition_clk ),
    .X(\clknet_leaf_144_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_145_top1.acquisition_clk  (.A(\clknet_6_63_0_top1.acquisition_clk ),
    .X(\clknet_leaf_145_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_146_top1.acquisition_clk  (.A(\clknet_6_63_0_top1.acquisition_clk ),
    .X(\clknet_leaf_146_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_147_top1.acquisition_clk  (.A(\clknet_6_63_0_top1.acquisition_clk ),
    .X(\clknet_leaf_147_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_148_top1.acquisition_clk  (.A(\clknet_6_63_0_top1.acquisition_clk ),
    .X(\clknet_leaf_148_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_149_top1.acquisition_clk  (.A(\clknet_6_62_0_top1.acquisition_clk ),
    .X(\clknet_leaf_149_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_150_top1.acquisition_clk  (.A(\clknet_6_62_0_top1.acquisition_clk ),
    .X(\clknet_leaf_150_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_151_top1.acquisition_clk  (.A(\clknet_6_62_0_top1.acquisition_clk ),
    .X(\clknet_leaf_151_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_152_top1.acquisition_clk  (.A(\clknet_6_62_0_top1.acquisition_clk ),
    .X(\clknet_leaf_152_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_153_top1.acquisition_clk  (.A(\clknet_6_62_0_top1.acquisition_clk ),
    .X(\clknet_leaf_153_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_154_top1.acquisition_clk  (.A(\clknet_6_60_0_top1.acquisition_clk ),
    .X(\clknet_leaf_154_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_155_top1.acquisition_clk  (.A(\clknet_6_57_0_top1.acquisition_clk ),
    .X(\clknet_leaf_155_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_156_top1.acquisition_clk  (.A(\clknet_6_60_0_top1.acquisition_clk ),
    .X(\clknet_leaf_156_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_157_top1.acquisition_clk  (.A(\clknet_6_57_0_top1.acquisition_clk ),
    .X(\clknet_leaf_157_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_158_top1.acquisition_clk  (.A(\clknet_6_57_0_top1.acquisition_clk ),
    .X(\clknet_leaf_158_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_159_top1.acquisition_clk  (.A(\clknet_6_59_0_top1.acquisition_clk ),
    .X(\clknet_leaf_159_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_160_top1.acquisition_clk  (.A(\clknet_6_59_0_top1.acquisition_clk ),
    .X(\clknet_leaf_160_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_161_top1.acquisition_clk  (.A(\clknet_6_59_0_top1.acquisition_clk ),
    .X(\clknet_leaf_161_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_162_top1.acquisition_clk  (.A(\clknet_6_59_0_top1.acquisition_clk ),
    .X(\clknet_leaf_162_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_163_top1.acquisition_clk  (.A(\clknet_6_58_0_top1.acquisition_clk ),
    .X(\clknet_leaf_163_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_164_top1.acquisition_clk  (.A(\clknet_6_58_0_top1.acquisition_clk ),
    .X(\clknet_leaf_164_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_165_top1.acquisition_clk  (.A(\clknet_6_58_0_top1.acquisition_clk ),
    .X(\clknet_leaf_165_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_166_top1.acquisition_clk  (.A(\clknet_6_58_0_top1.acquisition_clk ),
    .X(\clknet_leaf_166_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_167_top1.acquisition_clk  (.A(\clknet_6_58_0_top1.acquisition_clk ),
    .X(\clknet_leaf_167_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_168_top1.acquisition_clk  (.A(\clknet_6_56_0_top1.acquisition_clk ),
    .X(\clknet_leaf_168_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_169_top1.acquisition_clk  (.A(\clknet_6_56_0_top1.acquisition_clk ),
    .X(\clknet_leaf_169_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_170_top1.acquisition_clk  (.A(\clknet_6_56_0_top1.acquisition_clk ),
    .X(\clknet_leaf_170_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_171_top1.acquisition_clk  (.A(\clknet_6_56_0_top1.acquisition_clk ),
    .X(\clknet_leaf_171_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_172_top1.acquisition_clk  (.A(\clknet_6_56_0_top1.acquisition_clk ),
    .X(\clknet_leaf_172_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_173_top1.acquisition_clk  (.A(\clknet_6_57_0_top1.acquisition_clk ),
    .X(\clknet_leaf_173_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_174_top1.acquisition_clk  (.A(\clknet_6_57_0_top1.acquisition_clk ),
    .X(\clknet_leaf_174_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_175_top1.acquisition_clk  (.A(\clknet_6_51_0_top1.acquisition_clk ),
    .X(\clknet_leaf_175_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_176_top1.acquisition_clk  (.A(\clknet_6_50_0_top1.acquisition_clk ),
    .X(\clknet_leaf_176_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_177_top1.acquisition_clk  (.A(\clknet_6_50_0_top1.acquisition_clk ),
    .X(\clknet_leaf_177_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_178_top1.acquisition_clk  (.A(\clknet_6_50_0_top1.acquisition_clk ),
    .X(\clknet_leaf_178_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_179_top1.acquisition_clk  (.A(\clknet_6_50_0_top1.acquisition_clk ),
    .X(\clknet_leaf_179_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_180_top1.acquisition_clk  (.A(\clknet_6_50_0_top1.acquisition_clk ),
    .X(\clknet_leaf_180_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_181_top1.acquisition_clk  (.A(\clknet_6_48_0_top1.acquisition_clk ),
    .X(\clknet_leaf_181_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_182_top1.acquisition_clk  (.A(\clknet_6_48_0_top1.acquisition_clk ),
    .X(\clknet_leaf_182_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_183_top1.acquisition_clk  (.A(\clknet_6_37_0_top1.acquisition_clk ),
    .X(\clknet_leaf_183_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_184_top1.acquisition_clk  (.A(\clknet_6_37_0_top1.acquisition_clk ),
    .X(\clknet_leaf_184_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_185_top1.acquisition_clk  (.A(\clknet_6_37_0_top1.acquisition_clk ),
    .X(\clknet_leaf_185_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_186_top1.acquisition_clk  (.A(\clknet_6_39_0_top1.acquisition_clk ),
    .X(\clknet_leaf_186_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_187_top1.acquisition_clk  (.A(\clknet_6_39_0_top1.acquisition_clk ),
    .X(\clknet_leaf_187_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_188_top1.acquisition_clk  (.A(\clknet_6_39_0_top1.acquisition_clk ),
    .X(\clknet_leaf_188_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_189_top1.acquisition_clk  (.A(\clknet_6_39_0_top1.acquisition_clk ),
    .X(\clknet_leaf_189_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_190_top1.acquisition_clk  (.A(\clknet_6_38_0_top1.acquisition_clk ),
    .X(\clknet_leaf_190_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_191_top1.acquisition_clk  (.A(\clknet_6_38_0_top1.acquisition_clk ),
    .X(\clknet_leaf_191_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_192_top1.acquisition_clk  (.A(\clknet_6_38_0_top1.acquisition_clk ),
    .X(\clknet_leaf_192_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_193_top1.acquisition_clk  (.A(\clknet_6_44_0_top1.acquisition_clk ),
    .X(\clknet_leaf_193_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_194_top1.acquisition_clk  (.A(\clknet_6_44_0_top1.acquisition_clk ),
    .X(\clknet_leaf_194_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_195_top1.acquisition_clk  (.A(\clknet_6_44_0_top1.acquisition_clk ),
    .X(\clknet_leaf_195_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_196_top1.acquisition_clk  (.A(\clknet_6_45_0_top1.acquisition_clk ),
    .X(\clknet_leaf_196_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_197_top1.acquisition_clk  (.A(\clknet_6_45_0_top1.acquisition_clk ),
    .X(\clknet_leaf_197_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_198_top1.acquisition_clk  (.A(\clknet_6_45_0_top1.acquisition_clk ),
    .X(\clknet_leaf_198_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_199_top1.acquisition_clk  (.A(\clknet_6_45_0_top1.acquisition_clk ),
    .X(\clknet_leaf_199_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_200_top1.acquisition_clk  (.A(\clknet_6_45_0_top1.acquisition_clk ),
    .X(\clknet_leaf_200_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_201_top1.acquisition_clk  (.A(\clknet_6_47_0_top1.acquisition_clk ),
    .X(\clknet_leaf_201_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_202_top1.acquisition_clk  (.A(\clknet_6_47_0_top1.acquisition_clk ),
    .X(\clknet_leaf_202_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_203_top1.acquisition_clk  (.A(\clknet_6_47_0_top1.acquisition_clk ),
    .X(\clknet_leaf_203_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_204_top1.acquisition_clk  (.A(\clknet_6_46_0_top1.acquisition_clk ),
    .X(\clknet_leaf_204_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_205_top1.acquisition_clk  (.A(\clknet_6_47_0_top1.acquisition_clk ),
    .X(\clknet_leaf_205_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_206_top1.acquisition_clk  (.A(\clknet_6_46_0_top1.acquisition_clk ),
    .X(\clknet_leaf_206_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_207_top1.acquisition_clk  (.A(\clknet_6_46_0_top1.acquisition_clk ),
    .X(\clknet_leaf_207_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_208_top1.acquisition_clk  (.A(\clknet_6_44_0_top1.acquisition_clk ),
    .X(\clknet_leaf_208_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_209_top1.acquisition_clk  (.A(\clknet_6_44_0_top1.acquisition_clk ),
    .X(\clknet_leaf_209_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_210_top1.acquisition_clk  (.A(\clknet_6_41_0_top1.acquisition_clk ),
    .X(\clknet_leaf_210_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_211_top1.acquisition_clk  (.A(\clknet_6_41_0_top1.acquisition_clk ),
    .X(\clknet_leaf_211_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_212_top1.acquisition_clk  (.A(\clknet_6_41_0_top1.acquisition_clk ),
    .X(\clknet_leaf_212_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_213_top1.acquisition_clk  (.A(\clknet_6_42_0_top1.acquisition_clk ),
    .X(\clknet_leaf_213_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_214_top1.acquisition_clk  (.A(\clknet_6_43_0_top1.acquisition_clk ),
    .X(\clknet_leaf_214_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_215_top1.acquisition_clk  (.A(\clknet_6_46_0_top1.acquisition_clk ),
    .X(\clknet_leaf_215_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_216_top1.acquisition_clk  (.A(\clknet_6_46_0_top1.acquisition_clk ),
    .X(\clknet_leaf_216_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_217_top1.acquisition_clk  (.A(\clknet_6_43_0_top1.acquisition_clk ),
    .X(\clknet_leaf_217_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_218_top1.acquisition_clk  (.A(\clknet_6_43_0_top1.acquisition_clk ),
    .X(\clknet_leaf_218_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_219_top1.acquisition_clk  (.A(\clknet_6_43_0_top1.acquisition_clk ),
    .X(\clknet_leaf_219_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_220_top1.acquisition_clk  (.A(\clknet_6_42_0_top1.acquisition_clk ),
    .X(\clknet_leaf_220_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_221_top1.acquisition_clk  (.A(\clknet_6_42_0_top1.acquisition_clk ),
    .X(\clknet_leaf_221_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_222_top1.acquisition_clk  (.A(\clknet_6_42_0_top1.acquisition_clk ),
    .X(\clknet_leaf_222_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_223_top1.acquisition_clk  (.A(\clknet_6_42_0_top1.acquisition_clk ),
    .X(\clknet_leaf_223_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_224_top1.acquisition_clk  (.A(\clknet_6_40_0_top1.acquisition_clk ),
    .X(\clknet_leaf_224_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_225_top1.acquisition_clk  (.A(\clknet_6_40_0_top1.acquisition_clk ),
    .X(\clknet_leaf_225_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_226_top1.acquisition_clk  (.A(\clknet_6_40_0_top1.acquisition_clk ),
    .X(\clknet_leaf_226_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_227_top1.acquisition_clk  (.A(\clknet_6_40_0_top1.acquisition_clk ),
    .X(\clknet_leaf_227_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_228_top1.acquisition_clk  (.A(\clknet_6_40_0_top1.acquisition_clk ),
    .X(\clknet_leaf_228_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_229_top1.acquisition_clk  (.A(\clknet_6_41_0_top1.acquisition_clk ),
    .X(\clknet_leaf_229_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_230_top1.acquisition_clk  (.A(\clknet_6_41_0_top1.acquisition_clk ),
    .X(\clknet_leaf_230_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_231_top1.acquisition_clk  (.A(\clknet_6_35_0_top1.acquisition_clk ),
    .X(\clknet_leaf_231_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_232_top1.acquisition_clk  (.A(\clknet_6_35_0_top1.acquisition_clk ),
    .X(\clknet_leaf_232_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_233_top1.acquisition_clk  (.A(\clknet_6_34_0_top1.acquisition_clk ),
    .X(\clknet_leaf_233_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_234_top1.acquisition_clk  (.A(\clknet_6_34_0_top1.acquisition_clk ),
    .X(\clknet_leaf_234_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_235_top1.acquisition_clk  (.A(\clknet_6_34_0_top1.acquisition_clk ),
    .X(\clknet_leaf_235_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_236_top1.acquisition_clk  (.A(\clknet_6_34_0_top1.acquisition_clk ),
    .X(\clknet_leaf_236_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_237_top1.acquisition_clk  (.A(\clknet_6_34_0_top1.acquisition_clk ),
    .X(\clknet_leaf_237_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_238_top1.acquisition_clk  (.A(\clknet_6_32_0_top1.acquisition_clk ),
    .X(\clknet_leaf_238_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_239_top1.acquisition_clk  (.A(\clknet_6_32_0_top1.acquisition_clk ),
    .X(\clknet_leaf_239_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_240_top1.acquisition_clk  (.A(\clknet_6_32_0_top1.acquisition_clk ),
    .X(\clknet_leaf_240_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_241_top1.acquisition_clk  (.A(\clknet_6_32_0_top1.acquisition_clk ),
    .X(\clknet_leaf_241_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_242_top1.acquisition_clk  (.A(\clknet_6_32_0_top1.acquisition_clk ),
    .X(\clknet_leaf_242_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_243_top1.acquisition_clk  (.A(\clknet_6_33_0_top1.acquisition_clk ),
    .X(\clknet_leaf_243_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_244_top1.acquisition_clk  (.A(\clknet_6_33_0_top1.acquisition_clk ),
    .X(\clknet_leaf_244_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_245_top1.acquisition_clk  (.A(\clknet_6_33_0_top1.acquisition_clk ),
    .X(\clknet_leaf_245_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_246_top1.acquisition_clk  (.A(\clknet_6_14_0_top1.acquisition_clk ),
    .X(\clknet_leaf_246_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_247_top1.acquisition_clk  (.A(\clknet_6_33_0_top1.acquisition_clk ),
    .X(\clknet_leaf_247_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_248_top1.acquisition_clk  (.A(\clknet_6_36_0_top1.acquisition_clk ),
    .X(\clknet_leaf_248_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_249_top1.acquisition_clk  (.A(\clknet_6_33_0_top1.acquisition_clk ),
    .X(\clknet_leaf_249_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_250_top1.acquisition_clk  (.A(\clknet_6_35_0_top1.acquisition_clk ),
    .X(\clknet_leaf_250_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_251_top1.acquisition_clk  (.A(\clknet_6_35_0_top1.acquisition_clk ),
    .X(\clknet_leaf_251_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_252_top1.acquisition_clk  (.A(\clknet_6_38_0_top1.acquisition_clk ),
    .X(\clknet_leaf_252_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_253_top1.acquisition_clk  (.A(\clknet_6_38_0_top1.acquisition_clk ),
    .X(\clknet_leaf_253_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_254_top1.acquisition_clk  (.A(\clknet_6_36_0_top1.acquisition_clk ),
    .X(\clknet_leaf_254_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_255_top1.acquisition_clk  (.A(\clknet_6_36_0_top1.acquisition_clk ),
    .X(\clknet_leaf_255_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_256_top1.acquisition_clk  (.A(\clknet_6_36_0_top1.acquisition_clk ),
    .X(\clknet_leaf_256_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_257_top1.acquisition_clk  (.A(\clknet_6_36_0_top1.acquisition_clk ),
    .X(\clknet_leaf_257_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_258_top1.acquisition_clk  (.A(\clknet_6_37_0_top1.acquisition_clk ),
    .X(\clknet_leaf_258_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_259_top1.acquisition_clk  (.A(\clknet_6_37_0_top1.acquisition_clk ),
    .X(\clknet_leaf_259_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_260_top1.acquisition_clk  (.A(\clknet_6_26_0_top1.acquisition_clk ),
    .X(\clknet_leaf_260_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_261_top1.acquisition_clk  (.A(\clknet_6_15_0_top1.acquisition_clk ),
    .X(\clknet_leaf_261_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_262_top1.acquisition_clk  (.A(\clknet_6_15_0_top1.acquisition_clk ),
    .X(\clknet_leaf_262_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_263_top1.acquisition_clk  (.A(\clknet_6_15_0_top1.acquisition_clk ),
    .X(\clknet_leaf_263_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_264_top1.acquisition_clk  (.A(\clknet_6_15_0_top1.acquisition_clk ),
    .X(\clknet_leaf_264_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_265_top1.acquisition_clk  (.A(\clknet_6_14_0_top1.acquisition_clk ),
    .X(\clknet_leaf_265_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_266_top1.acquisition_clk  (.A(\clknet_6_13_0_top1.acquisition_clk ),
    .X(\clknet_leaf_266_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_267_top1.acquisition_clk  (.A(\clknet_6_13_0_top1.acquisition_clk ),
    .X(\clknet_leaf_267_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_268_top1.acquisition_clk  (.A(\clknet_6_13_0_top1.acquisition_clk ),
    .X(\clknet_leaf_268_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_269_top1.acquisition_clk  (.A(\clknet_6_12_0_top1.acquisition_clk ),
    .X(\clknet_leaf_269_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_270_top1.acquisition_clk  (.A(\clknet_6_13_0_top1.acquisition_clk ),
    .X(\clknet_leaf_270_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_271_top1.acquisition_clk  (.A(\clknet_6_11_0_top1.acquisition_clk ),
    .X(\clknet_leaf_271_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_272_top1.acquisition_clk  (.A(\clknet_6_14_0_top1.acquisition_clk ),
    .X(\clknet_leaf_272_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_273_top1.acquisition_clk  (.A(\clknet_6_14_0_top1.acquisition_clk ),
    .X(\clknet_leaf_273_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_274_top1.acquisition_clk  (.A(\clknet_6_14_0_top1.acquisition_clk ),
    .X(\clknet_leaf_274_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_275_top1.acquisition_clk  (.A(\clknet_6_11_0_top1.acquisition_clk ),
    .X(\clknet_leaf_275_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_276_top1.acquisition_clk  (.A(\clknet_6_11_0_top1.acquisition_clk ),
    .X(\clknet_leaf_276_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_277_top1.acquisition_clk  (.A(\clknet_6_11_0_top1.acquisition_clk ),
    .X(\clknet_leaf_277_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_278_top1.acquisition_clk  (.A(\clknet_6_10_0_top1.acquisition_clk ),
    .X(\clknet_leaf_278_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_279_top1.acquisition_clk  (.A(\clknet_6_10_0_top1.acquisition_clk ),
    .X(\clknet_leaf_279_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_280_top1.acquisition_clk  (.A(\clknet_6_10_0_top1.acquisition_clk ),
    .X(\clknet_leaf_280_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_281_top1.acquisition_clk  (.A(\clknet_6_10_0_top1.acquisition_clk ),
    .X(\clknet_leaf_281_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_282_top1.acquisition_clk  (.A(\clknet_6_10_0_top1.acquisition_clk ),
    .X(\clknet_leaf_282_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_283_top1.acquisition_clk  (.A(\clknet_6_8_0_top1.acquisition_clk ),
    .X(\clknet_leaf_283_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_284_top1.acquisition_clk  (.A(\clknet_6_8_0_top1.acquisition_clk ),
    .X(\clknet_leaf_284_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_285_top1.acquisition_clk  (.A(\clknet_6_8_0_top1.acquisition_clk ),
    .X(\clknet_leaf_285_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_286_top1.acquisition_clk  (.A(\clknet_6_9_0_top1.acquisition_clk ),
    .X(\clknet_leaf_286_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_287_top1.acquisition_clk  (.A(\clknet_6_9_0_top1.acquisition_clk ),
    .X(\clknet_leaf_287_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_288_top1.acquisition_clk  (.A(\clknet_6_9_0_top1.acquisition_clk ),
    .X(\clknet_leaf_288_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_289_top1.acquisition_clk  (.A(\clknet_6_9_0_top1.acquisition_clk ),
    .X(\clknet_leaf_289_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_290_top1.acquisition_clk  (.A(\clknet_6_12_0_top1.acquisition_clk ),
    .X(\clknet_leaf_290_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_291_top1.acquisition_clk  (.A(\clknet_6_9_0_top1.acquisition_clk ),
    .X(\clknet_leaf_291_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_292_top1.acquisition_clk  (.A(\clknet_6_3_0_top1.acquisition_clk ),
    .X(\clknet_leaf_292_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_293_top1.acquisition_clk  (.A(\clknet_6_2_0_top1.acquisition_clk ),
    .X(\clknet_leaf_293_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_294_top1.acquisition_clk  (.A(\clknet_6_8_0_top1.acquisition_clk ),
    .X(\clknet_leaf_294_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_295_top1.acquisition_clk  (.A(\clknet_6_8_0_top1.acquisition_clk ),
    .X(\clknet_leaf_295_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_296_top1.acquisition_clk  (.A(\clknet_6_2_0_top1.acquisition_clk ),
    .X(\clknet_leaf_296_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_297_top1.acquisition_clk  (.A(\clknet_6_2_0_top1.acquisition_clk ),
    .X(\clknet_leaf_297_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_298_top1.acquisition_clk  (.A(\clknet_6_2_0_top1.acquisition_clk ),
    .X(\clknet_leaf_298_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_299_top1.acquisition_clk  (.A(\clknet_6_2_0_top1.acquisition_clk ),
    .X(\clknet_leaf_299_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_300_top1.acquisition_clk  (.A(\clknet_6_0_0_top1.acquisition_clk ),
    .X(\clknet_leaf_300_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_301_top1.acquisition_clk  (.A(\clknet_6_0_0_top1.acquisition_clk ),
    .X(\clknet_leaf_301_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_leaf_302_top1.acquisition_clk  (.A(\clknet_6_0_0_top1.acquisition_clk ),
    .X(\clknet_leaf_302_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_0_top1.acquisition_clk  (.A(\top1.acquisition_clk ),
    .X(\clknet_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_3_0_0_top1.acquisition_clk  (.A(\clknet_0_top1.acquisition_clk ),
    .X(\clknet_3_0_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_3_1_0_top1.acquisition_clk  (.A(\clknet_0_top1.acquisition_clk ),
    .X(\clknet_3_1_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_3_2_0_top1.acquisition_clk  (.A(\clknet_0_top1.acquisition_clk ),
    .X(\clknet_3_2_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_3_3_0_top1.acquisition_clk  (.A(\clknet_0_top1.acquisition_clk ),
    .X(\clknet_3_3_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_3_4_0_top1.acquisition_clk  (.A(\clknet_0_top1.acquisition_clk ),
    .X(\clknet_3_4_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_3_5_0_top1.acquisition_clk  (.A(\clknet_0_top1.acquisition_clk ),
    .X(\clknet_3_5_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_3_6_0_top1.acquisition_clk  (.A(\clknet_0_top1.acquisition_clk ),
    .X(\clknet_3_6_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_3_7_0_top1.acquisition_clk  (.A(\clknet_0_top1.acquisition_clk ),
    .X(\clknet_3_7_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_0_0_top1.acquisition_clk  (.A(\clknet_3_0_0_top1.acquisition_clk ),
    .X(\clknet_6_0_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_1_0_top1.acquisition_clk  (.A(\clknet_3_0_0_top1.acquisition_clk ),
    .X(\clknet_6_1_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_2_0_top1.acquisition_clk  (.A(\clknet_3_0_0_top1.acquisition_clk ),
    .X(\clknet_6_2_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_3_0_top1.acquisition_clk  (.A(\clknet_3_0_0_top1.acquisition_clk ),
    .X(\clknet_6_3_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_4_0_top1.acquisition_clk  (.A(\clknet_3_0_0_top1.acquisition_clk ),
    .X(\clknet_6_4_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_5_0_top1.acquisition_clk  (.A(\clknet_3_0_0_top1.acquisition_clk ),
    .X(\clknet_6_5_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_6_0_top1.acquisition_clk  (.A(\clknet_3_0_0_top1.acquisition_clk ),
    .X(\clknet_6_6_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_7_0_top1.acquisition_clk  (.A(\clknet_3_0_0_top1.acquisition_clk ),
    .X(\clknet_6_7_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_8_0_top1.acquisition_clk  (.A(\clknet_3_1_0_top1.acquisition_clk ),
    .X(\clknet_6_8_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_9_0_top1.acquisition_clk  (.A(\clknet_3_1_0_top1.acquisition_clk ),
    .X(\clknet_6_9_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_10_0_top1.acquisition_clk  (.A(\clknet_3_1_0_top1.acquisition_clk ),
    .X(\clknet_6_10_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_11_0_top1.acquisition_clk  (.A(\clknet_3_1_0_top1.acquisition_clk ),
    .X(\clknet_6_11_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_12_0_top1.acquisition_clk  (.A(\clknet_3_1_0_top1.acquisition_clk ),
    .X(\clknet_6_12_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_13_0_top1.acquisition_clk  (.A(\clknet_3_1_0_top1.acquisition_clk ),
    .X(\clknet_6_13_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_14_0_top1.acquisition_clk  (.A(\clknet_3_1_0_top1.acquisition_clk ),
    .X(\clknet_6_14_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_15_0_top1.acquisition_clk  (.A(\clknet_3_1_0_top1.acquisition_clk ),
    .X(\clknet_6_15_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_16_0_top1.acquisition_clk  (.A(\clknet_3_2_0_top1.acquisition_clk ),
    .X(\clknet_6_16_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_17_0_top1.acquisition_clk  (.A(\clknet_3_2_0_top1.acquisition_clk ),
    .X(\clknet_6_17_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_18_0_top1.acquisition_clk  (.A(\clknet_3_2_0_top1.acquisition_clk ),
    .X(\clknet_6_18_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_19_0_top1.acquisition_clk  (.A(\clknet_3_2_0_top1.acquisition_clk ),
    .X(\clknet_6_19_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_20_0_top1.acquisition_clk  (.A(\clknet_3_2_0_top1.acquisition_clk ),
    .X(\clknet_6_20_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_21_0_top1.acquisition_clk  (.A(\clknet_3_2_0_top1.acquisition_clk ),
    .X(\clknet_6_21_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_22_0_top1.acquisition_clk  (.A(\clknet_3_2_0_top1.acquisition_clk ),
    .X(\clknet_6_22_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_23_0_top1.acquisition_clk  (.A(\clknet_3_2_0_top1.acquisition_clk ),
    .X(\clknet_6_23_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_24_0_top1.acquisition_clk  (.A(\clknet_3_3_0_top1.acquisition_clk ),
    .X(\clknet_6_24_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_25_0_top1.acquisition_clk  (.A(\clknet_3_3_0_top1.acquisition_clk ),
    .X(\clknet_6_25_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_26_0_top1.acquisition_clk  (.A(\clknet_3_3_0_top1.acquisition_clk ),
    .X(\clknet_6_26_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_27_0_top1.acquisition_clk  (.A(\clknet_3_3_0_top1.acquisition_clk ),
    .X(\clknet_6_27_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_28_0_top1.acquisition_clk  (.A(\clknet_3_3_0_top1.acquisition_clk ),
    .X(\clknet_6_28_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_29_0_top1.acquisition_clk  (.A(\clknet_3_3_0_top1.acquisition_clk ),
    .X(\clknet_6_29_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_30_0_top1.acquisition_clk  (.A(\clknet_3_3_0_top1.acquisition_clk ),
    .X(\clknet_6_30_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_31_0_top1.acquisition_clk  (.A(\clknet_3_3_0_top1.acquisition_clk ),
    .X(\clknet_6_31_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_32_0_top1.acquisition_clk  (.A(\clknet_3_4_0_top1.acquisition_clk ),
    .X(\clknet_6_32_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_33_0_top1.acquisition_clk  (.A(\clknet_3_4_0_top1.acquisition_clk ),
    .X(\clknet_6_33_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_34_0_top1.acquisition_clk  (.A(\clknet_3_4_0_top1.acquisition_clk ),
    .X(\clknet_6_34_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_35_0_top1.acquisition_clk  (.A(\clknet_3_4_0_top1.acquisition_clk ),
    .X(\clknet_6_35_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_36_0_top1.acquisition_clk  (.A(\clknet_3_4_0_top1.acquisition_clk ),
    .X(\clknet_6_36_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_37_0_top1.acquisition_clk  (.A(\clknet_3_4_0_top1.acquisition_clk ),
    .X(\clknet_6_37_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_38_0_top1.acquisition_clk  (.A(\clknet_3_4_0_top1.acquisition_clk ),
    .X(\clknet_6_38_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_39_0_top1.acquisition_clk  (.A(\clknet_3_4_0_top1.acquisition_clk ),
    .X(\clknet_6_39_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_40_0_top1.acquisition_clk  (.A(\clknet_3_5_0_top1.acquisition_clk ),
    .X(\clknet_6_40_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_41_0_top1.acquisition_clk  (.A(\clknet_3_5_0_top1.acquisition_clk ),
    .X(\clknet_6_41_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_42_0_top1.acquisition_clk  (.A(\clknet_3_5_0_top1.acquisition_clk ),
    .X(\clknet_6_42_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_43_0_top1.acquisition_clk  (.A(\clknet_3_5_0_top1.acquisition_clk ),
    .X(\clknet_6_43_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_44_0_top1.acquisition_clk  (.A(\clknet_3_5_0_top1.acquisition_clk ),
    .X(\clknet_6_44_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_45_0_top1.acquisition_clk  (.A(\clknet_3_5_0_top1.acquisition_clk ),
    .X(\clknet_6_45_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_46_0_top1.acquisition_clk  (.A(\clknet_3_5_0_top1.acquisition_clk ),
    .X(\clknet_6_46_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_47_0_top1.acquisition_clk  (.A(\clknet_3_5_0_top1.acquisition_clk ),
    .X(\clknet_6_47_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_48_0_top1.acquisition_clk  (.A(\clknet_3_6_0_top1.acquisition_clk ),
    .X(\clknet_6_48_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_49_0_top1.acquisition_clk  (.A(\clknet_3_6_0_top1.acquisition_clk ),
    .X(\clknet_6_49_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_50_0_top1.acquisition_clk  (.A(\clknet_3_6_0_top1.acquisition_clk ),
    .X(\clknet_6_50_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_51_0_top1.acquisition_clk  (.A(\clknet_3_6_0_top1.acquisition_clk ),
    .X(\clknet_6_51_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_52_0_top1.acquisition_clk  (.A(\clknet_3_6_0_top1.acquisition_clk ),
    .X(\clknet_6_52_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_53_0_top1.acquisition_clk  (.A(\clknet_3_6_0_top1.acquisition_clk ),
    .X(\clknet_6_53_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_54_0_top1.acquisition_clk  (.A(\clknet_3_6_0_top1.acquisition_clk ),
    .X(\clknet_6_54_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_55_0_top1.acquisition_clk  (.A(\clknet_3_6_0_top1.acquisition_clk ),
    .X(\clknet_6_55_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_56_0_top1.acquisition_clk  (.A(\clknet_3_7_0_top1.acquisition_clk ),
    .X(\clknet_6_56_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_57_0_top1.acquisition_clk  (.A(\clknet_3_7_0_top1.acquisition_clk ),
    .X(\clknet_6_57_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_58_0_top1.acquisition_clk  (.A(\clknet_3_7_0_top1.acquisition_clk ),
    .X(\clknet_6_58_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_59_0_top1.acquisition_clk  (.A(\clknet_3_7_0_top1.acquisition_clk ),
    .X(\clknet_6_59_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_60_0_top1.acquisition_clk  (.A(\clknet_3_7_0_top1.acquisition_clk ),
    .X(\clknet_6_60_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_61_0_top1.acquisition_clk  (.A(\clknet_3_7_0_top1.acquisition_clk ),
    .X(\clknet_6_61_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_62_0_top1.acquisition_clk  (.A(\clknet_3_7_0_top1.acquisition_clk ),
    .X(\clknet_6_62_0_top1.acquisition_clk ));
 sg13g2_buf_2 \clkbuf_6_63_0_top1.acquisition_clk  (.A(\clknet_3_7_0_top1.acquisition_clk ),
    .X(\clknet_6_63_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload0 (.A(\clknet_6_3_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload1 (.A(\clknet_6_7_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload2 (.A(\clknet_6_11_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload3 (.A(\clknet_6_15_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload4 (.A(\clknet_6_19_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload5 (.A(\clknet_6_23_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload6 (.A(\clknet_6_27_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload7 (.A(\clknet_6_31_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload8 (.A(\clknet_6_35_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload9 (.A(\clknet_6_39_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload10 (.A(\clknet_6_43_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload11 (.A(\clknet_6_47_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload12 (.A(\clknet_6_51_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload13 (.A(\clknet_6_55_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload14 (.A(\clknet_6_59_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload15 (.A(\clknet_6_61_0_top1.acquisition_clk ));
 sg13g2_buf_2 clkload16 (.A(\clknet_6_63_0_top1.acquisition_clk ));
 sg13g2_inv_4 clkload17 (.A(\clknet_leaf_302_top1.acquisition_clk ));
 sg13g2_dlygate4sd3_1 hold1 (.A(\top1.memory2.mem2[159][1] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold2 (.A(\top1.memory2.mem1[156][0] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold3 (.A(\top1.memory1.mem2[151][2] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold4 (.A(\top1.memory2.mem2[168][1] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold5 (.A(\top1.memory2.mem2[93][2] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold6 (.A(\top1.memory1.mem2[28][1] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold7 (.A(\top1.memory1.mem2[191][0] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold8 (.A(\top1.memory2.mem1[147][2] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold9 (.A(\top1.memory1.mem2[184][0] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold10 (.A(\top1.memory1.mem2[28][0] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold11 (.A(\top1.memory2.mem1[180][2] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold12 (.A(\top1.memory2.mem1[122][0] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold13 (.A(\top1.memory1.mem2[195][2] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold14 (.A(\top1.memory2.mem2[147][1] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold15 (.A(\top1.memory2.mem2[195][0] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold16 (.A(\top1.memory2.mem2[125][2] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold17 (.A(\top1.memory1.mem1[180][2] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold18 (.A(\top1.memory1.mem2[172][1] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold19 (.A(\top1.memory1.mem1[91][1] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold20 (.A(\top1.memory2.mem1[61][1] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold21 (.A(\top1.memory2.mem2[40][2] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold22 (.A(\top1.memory1.mem1[14][0] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold23 (.A(\top1.memory1.mem1[183][2] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold24 (.A(\top1.memory2.mem2[11][2] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold25 (.A(\top1.memory2.mem1[44][2] ),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold26 (.A(\top1.memory1.mem1[44][0] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold27 (.A(\top1.memory2.mem2[55][0] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold28 (.A(\top1.memory2.mem2[17][0] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold29 (.A(\top1.memory1.mem1[51][2] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold30 (.A(\top1.memory2.mem2[40][0] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold31 (.A(\top1.memory1.mem2[91][0] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold32 (.A(\top1.memory1.mem2[61][1] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold33 (.A(\top1.memory1.mem2[175][1] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold34 (.A(\top1.memory2.mem1[159][0] ),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold35 (.A(\top1.memory2.mem1[95][2] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold36 (.A(\top1.memory2.mem2[31][0] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold37 (.A(\top1.memory1.mem1[185][1] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold38 (.A(\top1.memory2.mem1[171][0] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold39 (.A(\top1.memory2.mem2[24][0] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold40 (.A(\top1.memory2.mem2[169][1] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold41 (.A(\top1.memory1.mem1[93][0] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold42 (.A(\top1.memory2.mem2[56][2] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold43 (.A(\top1.memory2.mem2[157][1] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold44 (.A(\top1.memory2.mem2[95][1] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold45 (.A(\top1.memory2.mem2[37][1] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold46 (.A(\top1.memory2.mem2[44][2] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold47 (.A(\top1.memory1.mem1[158][0] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold48 (.A(\top1.memory2.mem2[28][0] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold49 (.A(\top1.memory2.mem1[16][1] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold50 (.A(\top1.memory1.mem1[159][0] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold51 (.A(\top1.memory2.mem1[89][0] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold52 (.A(\top1.memory1.mem2[158][2] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold53 (.A(\top1.memory1.mem1[36][0] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold54 (.A(\top1.memory1.mem1[165][2] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold55 (.A(\top1.memory1.mem1[89][0] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold56 (.A(\top1.memory1.mem1[182][0] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold57 (.A(\top1.memory2.mem1[191][1] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold58 (.A(\top1.memory2.mem2[13][0] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold59 (.A(\top1.memory1.mem2[34][0] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold60 (.A(\top1.memory1.mem1[16][2] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold61 (.A(\top1.memory2.mem1[114][2] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold62 (.A(\top1.memory2.mem1[193][1] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold63 (.A(\top1.memory1.mem2[187][1] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold64 (.A(\top1.memory2.mem2[168][0] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold65 (.A(\top1.memory2.mem1[35][2] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold66 (.A(\top1.memory2.mem1[187][0] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold67 (.A(\top1.memory2.mem2[116][0] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold68 (.A(\top1.memory1.mem2[157][2] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold69 (.A(\top1.memory1.mem2[172][2] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold70 (.A(\top1.memory1.mem1[152][1] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold71 (.A(\top1.memory1.mem1[33][1] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold72 (.A(\top1.memory1.mem2[53][0] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold73 (.A(\top1.memory2.mem2[164][1] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold74 (.A(\top1.memory2.mem1[60][2] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold75 (.A(\top1.memory2.mem1[62][1] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold76 (.A(\top1.memory2.mem1[56][2] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold77 (.A(\top1.memory1.mem2[159][1] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold78 (.A(\top1.memory2.mem1[52][0] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold79 (.A(\top1.memory1.mem2[108][0] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold80 (.A(\top1.memory2.mem2[89][2] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold81 (.A(\top1.memory1.mem1[165][1] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold82 (.A(\top1.memory2.mem2[39][2] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold83 (.A(\top1.memory2.mem1[150][0] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold84 (.A(\top1.memory2.mem1[32][2] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold85 (.A(\top1.memory1.mem2[156][1] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold86 (.A(\top1.memory1.mem2[103][1] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold87 (.A(\top1.memory2.mem1[191][0] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold88 (.A(\top1.memory2.mem2[164][0] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold89 (.A(\top1.memory1.mem2[108][2] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold90 (.A(\top1.memory1.mem1[153][1] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold91 (.A(\top1.memory2.mem1[47][1] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold92 (.A(\top1.memory1.mem1[91][2] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold93 (.A(\top1.memory2.mem2[18][0] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold94 (.A(\top1.memory1.mem2[38][1] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold95 (.A(\top1.memory1.mem1[13][0] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold96 (.A(\top1.memory2.mem2[177][1] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold97 (.A(\top1.memory1.mem1[93][1] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold98 (.A(\top1.memory1.mem1[157][1] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold99 (.A(\top1.memory1.mem2[170][2] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold100 (.A(\top1.memory2.mem2[36][2] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold101 (.A(\top1.memory1.mem1[18][2] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold102 (.A(\top1.memory2.mem2[180][0] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold103 (.A(\top1.memory2.mem1[196][1] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold104 (.A(\top1.memory2.mem1[21][2] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold105 (.A(\top1.memory2.mem2[55][2] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold106 (.A(\top1.memory2.mem2[89][1] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold107 (.A(\top1.memory2.mem2[56][1] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold108 (.A(\top1.memory1.mem2[16][1] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold109 (.A(\top1.memory1.mem2[149][2] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold110 (.A(\top1.memory2.mem2[32][2] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold111 (.A(\top1.memory1.mem1[92][0] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold112 (.A(\top1.memory1.mem1[90][2] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold113 (.A(\top1.memory2.mem1[170][1] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold114 (.A(\top1.memory2.mem2[51][1] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold115 (.A(\top1.memory2.mem2[44][0] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold116 (.A(\top1.memory2.mem2[36][1] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold117 (.A(\top1.memory2.mem2[28][2] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold118 (.A(\top1.memory2.mem1[22][0] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold119 (.A(\top1.memory1.mem2[92][2] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold120 (.A(\top1.memory2.mem1[148][0] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold121 (.A(\top1.memory1.mem2[13][1] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold122 (.A(\top1.memory2.mem2[184][0] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold123 (.A(\top1.memory1.mem2[158][0] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold124 (.A(\top1.memory1.mem2[51][2] ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold125 (.A(\top1.memory1.mem2[192][0] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold126 (.A(\top1.memory1.mem1[28][1] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold127 (.A(\top1.memory2.mem2[49][0] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold128 (.A(\top1.memory2.mem1[20][0] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold129 (.A(\top1.memory2.mem1[92][0] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold130 (.A(\top1.memory1.mem1[17][0] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold131 (.A(\top1.memory2.mem1[71][1] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold132 (.A(\top1.memory2.mem2[180][1] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold133 (.A(\top1.memory1.mem1[193][1] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold134 (.A(\top1.memory2.mem2[71][1] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold135 (.A(\top1.memory1.mem1[155][1] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold136 (.A(\top1.memory2.mem1[179][2] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold137 (.A(\top1.memory2.mem1[24][0] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold138 (.A(\top1.memory1.mem1[147][1] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold139 (.A(\top1.memory2.mem2[175][2] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold140 (.A(\top1.memory2.mem2[87][1] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold141 (.A(\top1.memory2.mem2[188][0] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold142 (.A(\top1.memory2.mem2[120][0] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold143 (.A(\top1.memory1.mem2[38][0] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold144 (.A(\top1.memory1.mem1[120][0] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold145 (.A(\top1.memory1.mem1[71][1] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold146 (.A(\top1.memory1.mem2[30][0] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold147 (.A(\top1.memory1.mem1[155][0] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold148 (.A(\top1.memory1.mem1[49][0] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold149 (.A(\top1.memory1.mem2[121][0] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold150 (.A(\top1.memory2.mem1[169][2] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold151 (.A(\top1.memory1.mem1[193][2] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold152 (.A(\top1.memory1.mem2[44][1] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold153 (.A(\top1.memory2.mem1[198][0] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold154 (.A(\top1.memory1.mem1[112][1] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold155 (.A(\top1.memory2.mem2[183][2] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold156 (.A(\top1.memory1.mem1[62][1] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold157 (.A(\top1.memory2.mem1[175][2] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold158 (.A(\top1.memory2.mem1[103][0] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold159 (.A(\top1.memory1.mem1[179][2] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold160 (.A(\top1.memory2.mem2[181][0] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold161 (.A(\top1.memory1.mem1[184][1] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold162 (.A(\top1.memory1.mem1[176][0] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold163 (.A(\top1.memory1.mem2[194][0] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold164 (.A(\top1.memory1.mem2[164][1] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold165 (.A(\top1.memory1.mem1[7][1] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold166 (.A(\top1.memory2.mem1[90][0] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold167 (.A(\top1.memory2.mem1[89][1] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold168 (.A(\top1.memory2.mem2[27][0] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold169 (.A(\top1.memory1.mem2[155][2] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold170 (.A(\top1.memory1.mem2[154][0] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold171 (.A(\top1.memory2.mem2[30][2] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold172 (.A(\top1.memory2.mem1[177][2] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold173 (.A(\top1.memory1.mem2[93][0] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold174 (.A(\top1.memory1.mem1[164][0] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold175 (.A(\top1.memory1.mem2[19][0] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold176 (.A(\top1.memory1.mem1[171][1] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold177 (.A(\top1.memory2.mem1[32][1] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold178 (.A(\top1.memory2.mem1[89][2] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold179 (.A(\top1.memory1.mem2[32][0] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold180 (.A(\top1.memory1.mem1[24][2] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold181 (.A(\top1.memory2.mem2[27][2] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold182 (.A(\top1.memory1.mem1[184][0] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold183 (.A(\top1.memory1.mem1[150][1] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold184 (.A(\top1.memory2.mem2[171][1] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold185 (.A(\top1.memory2.mem1[117][1] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold186 (.A(\top1.memory2.mem2[174][1] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold187 (.A(\top1.memory1.mem1[103][0] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold188 (.A(\top1.memory2.mem2[36][0] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold189 (.A(\top1.memory1.mem2[177][0] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold190 (.A(\top1.memory2.mem2[48][2] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold191 (.A(\top1.memory2.mem1[60][0] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold192 (.A(\top1.memory2.mem2[24][1] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold193 (.A(\top1.memory2.mem2[11][0] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold194 (.A(\top1.memory1.mem2[95][2] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold195 (.A(\top1.memory1.mem1[44][2] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold196 (.A(\top1.memory2.mem1[163][0] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold197 (.A(\top1.memory1.mem2[155][0] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold198 (.A(\top1.memory1.mem1[20][1] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold199 (.A(\top1.memory1.mem1[48][1] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold200 (.A(\top1.memory1.mem2[52][0] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold201 (.A(\top1.memory2.mem2[159][0] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold202 (.A(\top1.memory2.mem1[86][2] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold203 (.A(\top1.memory2.mem1[85][0] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold204 (.A(\top1.memory2.mem2[90][0] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold205 (.A(\top1.memory1.mem1[28][0] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold206 (.A(\top1.memory1.mem1[195][2] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold207 (.A(\top1.memory1.mem1[105][1] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold208 (.A(\top1.memory2.mem2[43][0] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold209 (.A(\top1.memory1.mem1[147][2] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold210 (.A(\top1.memory1.mem1[35][0] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold211 (.A(\top1.memory1.mem2[123][1] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold212 (.A(\top1.memory2.mem2[46][2] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold213 (.A(\top1.memory1.mem2[150][2] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold214 (.A(\top1.memory2.mem2[52][1] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold215 (.A(\top1.memory2.mem2[47][2] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold216 (.A(\top1.memory1.mem1[175][0] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold217 (.A(\top1.memory2.mem1[90][1] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold218 (.A(\top1.memory1.mem2[95][0] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold219 (.A(\top1.memory1.mem1[124][0] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold220 (.A(\top1.memory1.mem2[197][0] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold221 (.A(\top1.memory2.mem1[190][1] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold222 (.A(\top1.memory2.mem1[59][1] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold223 (.A(\top1.memory1.mem1[23][0] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold224 (.A(\top1.memory2.mem1[91][2] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold225 (.A(\top1.memory2.mem1[187][2] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold226 (.A(\top1.memory2.mem2[102][0] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold227 (.A(\top1.memory1.mem1[125][0] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold228 (.A(\top1.memory1.mem1[57][2] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold229 (.A(\top1.memory1.mem2[164][0] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold230 (.A(\top1.memory1.mem1[22][2] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold231 (.A(\top1.memory1.mem1[11][2] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold232 (.A(\top1.memory2.mem1[182][0] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold233 (.A(\top1.memory2.mem1[155][0] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold234 (.A(\top1.memory1.mem1[41][2] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold235 (.A(\top1.memory2.mem2[26][1] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold236 (.A(\top1.memory1.mem2[124][2] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold237 (.A(\top1.memory2.mem2[85][2] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold238 (.A(\top1.memory1.mem2[183][2] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold239 (.A(\top1.memory1.mem1[165][0] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold240 (.A(\top1.memory2.mem1[71][2] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold241 (.A(\top1.memory1.mem2[54][1] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold242 (.A(\top1.memory2.mem1[155][2] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold243 (.A(\top1.memory2.mem2[117][2] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold244 (.A(\top1.memory2.mem2[34][2] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold245 (.A(\top1.memory2.mem2[180][2] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold246 (.A(\top1.memory1.mem1[111][2] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold247 (.A(\top1.memory2.mem2[25][2] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold248 (.A(\top1.memory1.mem2[92][1] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold249 (.A(\top1.memory2.mem2[48][0] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold250 (.A(\top1.memory2.mem2[149][1] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold251 (.A(\top1.memory2.mem2[177][2] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold252 (.A(\top1.memory1.mem1[26][1] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold253 (.A(\top1.memory1.mem1[198][1] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold254 (.A(\top1.memory1.mem1[173][2] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold255 (.A(\top1.memory1.mem2[193][1] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold256 (.A(\top1.memory2.mem2[111][2] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold257 (.A(\top1.memory2.mem2[19][0] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold258 (.A(\top1.memory1.mem1[152][0] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold259 (.A(\top1.memory1.mem1[56][2] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold260 (.A(\top1.memory2.mem2[22][0] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold261 (.A(\top1.memory2.mem2[152][2] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold262 (.A(\top1.memory1.mem1[44][1] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold263 (.A(\top1.memory2.mem1[102][1] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold264 (.A(\top1.memory1.mem2[42][2] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold265 (.A(\top1.memory1.mem2[107][0] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold266 (.A(\top1.memory2.mem1[14][2] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold267 (.A(\top1.memory2.mem1[91][0] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold268 (.A(\top1.memory1.mem2[56][1] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold269 (.A(\top1.memory1.mem2[122][1] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold270 (.A(\top1.memory1.mem2[22][0] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold271 (.A(\top1.memory2.mem1[196][0] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold272 (.A(\top1.memory1.mem1[190][0] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold273 (.A(\top1.memory2.mem1[195][2] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold274 (.A(\top1.memory2.mem2[87][2] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold275 (.A(\top1.memory2.mem1[194][0] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold276 (.A(\top1.memory2.mem2[166][1] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold277 (.A(\top1.memory2.mem1[180][1] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold278 (.A(\top1.memory2.mem2[182][2] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold279 (.A(\top1.memory1.mem2[168][2] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold280 (.A(\top1.memory1.mem2[184][1] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold281 (.A(\top1.memory1.mem1[56][0] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold282 (.A(\top1.memory2.mem1[126][0] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold283 (.A(\top1.memory1.mem2[90][1] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold284 (.A(\top1.memory2.mem1[53][0] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold285 (.A(\top1.memory1.mem2[111][0] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold286 (.A(\top1.memory2.mem2[193][0] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold287 (.A(\top1.memory2.mem2[91][0] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold288 (.A(\top1.memory1.mem2[152][1] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold289 (.A(\top1.memory2.mem2[109][0] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold290 (.A(\top1.memory2.mem2[113][1] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold291 (.A(\top1.memory1.mem2[114][2] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold292 (.A(\top1.memory1.mem1[32][1] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold293 (.A(\top1.memory2.mem1[102][0] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold294 (.A(\top1.memory2.mem1[47][0] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold295 (.A(\top1.memory2.mem2[57][1] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold296 (.A(\top1.memory2.mem1[55][1] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold297 (.A(\top1.memory1.mem2[110][2] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold298 (.A(\top1.memory2.mem1[194][2] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold299 (.A(\top1.memory1.mem1[111][0] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold300 (.A(\top1.memory1.mem1[32][2] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold301 (.A(\top1.memory1.mem2[113][0] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold302 (.A(\top1.memory1.mem2[55][2] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold303 (.A(\top1.memory2.mem1[196][2] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold304 (.A(\top1.memory1.mem2[150][0] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold305 (.A(\top1.memory2.mem1[11][0] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold306 (.A(\top1.memory1.mem2[176][0] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold307 (.A(\top1.memory2.mem2[43][2] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold308 (.A(\top1.memory2.mem2[191][0] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold309 (.A(\top1.memory2.mem2[119][1] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold310 (.A(\top1.memory1.mem2[168][1] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold311 (.A(\top1.memory2.mem1[181][0] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold312 (.A(\top1.memory2.mem2[184][1] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold313 (.A(\top1.memory2.mem1[119][1] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold314 (.A(\top1.memory2.mem2[87][0] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold315 (.A(\top1.memory2.mem2[43][1] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold316 (.A(\top1.memory2.mem2[193][2] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold317 (.A(\top1.memory1.mem2[198][2] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold318 (.A(\top1.memory2.mem1[192][2] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold319 (.A(\top1.memory1.mem2[31][2] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold320 (.A(\top1.memory2.mem1[163][1] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold321 (.A(\top1.memory2.mem1[28][0] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold322 (.A(\top1.memory2.mem1[92][1] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold323 (.A(\top1.memory1.mem2[60][2] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold324 (.A(\top1.memory1.mem1[186][1] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold325 (.A(\top1.memory2.mem1[27][0] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold326 (.A(\top1.memory1.mem2[159][0] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold327 (.A(\top1.memory2.mem2[41][1] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold328 (.A(\top1.memory1.mem2[177][2] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold329 (.A(\top1.memory1.mem1[147][0] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold330 (.A(\top1.memory2.mem1[170][2] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold331 (.A(\top1.memory1.mem2[179][1] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold332 (.A(\top1.memory1.mem1[95][2] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold333 (.A(\top1.memory1.mem1[113][2] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold334 (.A(\top1.memory2.mem1[48][0] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold335 (.A(\top1.memory1.mem1[148][1] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold336 (.A(\top1.memory1.mem1[59][2] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold337 (.A(\top1.memory1.mem2[16][2] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold338 (.A(\top1.memory2.mem2[173][1] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold339 (.A(\top1.memory1.mem1[63][2] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold340 (.A(\top1.memory1.mem2[23][2] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold341 (.A(\top1.memory1.mem2[87][2] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold342 (.A(\top1.memory1.mem2[182][1] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold343 (.A(\top1.memory2.mem2[61][1] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold344 (.A(\top1.memory1.mem2[158][1] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold345 (.A(\top1.memory1.mem2[56][0] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold346 (.A(\top1.memory1.mem1[32][0] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold347 (.A(\top1.memory1.mem1[121][1] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold348 (.A(\top1.memory2.mem2[154][0] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold349 (.A(\top1.memory1.mem2[61][2] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold350 (.A(\top1.memory1.mem2[7][0] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold351 (.A(\top1.memory1.mem1[120][2] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold352 (.A(\top1.memory2.mem1[176][2] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold353 (.A(\top1.memory2.mem1[121][1] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold354 (.A(\top1.memory1.mem1[87][0] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold355 (.A(\top1.memory1.mem2[122][0] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold356 (.A(\top1.memory1.mem2[57][2] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold357 (.A(\top1.memory2.mem1[175][1] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold358 (.A(\top1.memory2.mem1[181][1] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold359 (.A(\top1.memory1.mem1[94][0] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold360 (.A(\top1.memory2.mem2[190][0] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold361 (.A(\top1.memory2.mem2[171][2] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold362 (.A(\top1.memory1.mem2[167][0] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold363 (.A(\top1.memory1.mem2[56][2] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold364 (.A(\top1.memory2.mem2[62][2] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold365 (.A(\top1.memory1.mem2[198][0] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold366 (.A(\top1.memory1.mem1[58][2] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold367 (.A(\top1.memory1.mem2[51][1] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold368 (.A(\top1.memory1.mem1[47][1] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold369 (.A(\top1.memory1.mem1[87][2] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold370 (.A(\top1.memory2.mem1[112][1] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold371 (.A(\top1.memory2.mem1[14][0] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold372 (.A(\top1.memory1.mem2[186][0] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold373 (.A(\top1.memory2.mem1[101][0] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold374 (.A(\top1.memory1.mem1[20][0] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold375 (.A(\top1.memory1.mem2[169][0] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold376 (.A(\top1.memory2.mem1[183][0] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold377 (.A(\top1.memory1.mem2[86][1] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold378 (.A(\top1.memory1.mem2[105][0] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold379 (.A(\top1.memory2.mem1[13][0] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold380 (.A(\top1.memory1.mem2[124][1] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold381 (.A(\top1.memory2.mem1[147][1] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold382 (.A(\top1.memory1.mem2[17][2] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold383 (.A(\top1.memory2.mem2[153][2] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold384 (.A(\top1.memory2.mem1[17][0] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold385 (.A(\top1.memory2.mem1[34][0] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold386 (.A(\top1.memory1.mem2[35][0] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold387 (.A(\top1.memory1.mem1[18][1] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold388 (.A(\top1.memory2.mem1[31][1] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold389 (.A(\top1.memory2.mem1[33][2] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold390 (.A(\top1.memory2.mem2[51][0] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold391 (.A(\top1.memory1.mem2[93][1] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold392 (.A(\top1.memory1.mem1[62][0] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold393 (.A(\top1.memory2.mem1[87][2] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold394 (.A(\top1.memory1.mem2[7][2] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold395 (.A(\top1.memory1.mem2[183][0] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold396 (.A(\top1.memory2.mem1[123][1] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold397 (.A(\top1.memory1.mem1[46][2] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold398 (.A(\top1.memory2.mem1[90][2] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold399 (.A(\top1.memory2.mem2[13][1] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold400 (.A(\top1.memory2.mem1[86][1] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold401 (.A(\top1.memory1.mem1[188][0] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold402 (.A(\top1.memory1.mem2[157][0] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold403 (.A(\top1.memory2.mem2[158][0] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold404 (.A(\top1.memory2.mem2[108][2] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold405 (.A(\top1.memory2.mem2[186][2] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold406 (.A(\top1.memory1.mem1[108][2] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold407 (.A(\top1.memory2.mem1[103][2] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold408 (.A(\top1.memory2.mem2[192][1] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold409 (.A(\top1.memory2.mem2[163][2] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold410 (.A(\top1.memory1.mem2[42][0] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold411 (.A(\top1.memory1.mem2[47][0] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold412 (.A(\top1.memory1.mem2[101][0] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold413 (.A(\top1.memory2.mem2[101][2] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold414 (.A(\top1.memory1.mem2[122][2] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold415 (.A(\top1.memory1.mem2[71][2] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold416 (.A(\top1.memory2.mem1[95][1] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold417 (.A(\top1.memory1.mem2[166][1] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold418 (.A(\top1.memory1.mem1[50][1] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold419 (.A(\top1.memory1.mem2[60][1] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold420 (.A(\top1.memory1.mem1[174][0] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold421 (.A(\top1.memory2.mem1[111][1] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold422 (.A(\top1.memory1.mem2[43][2] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold423 (.A(\top1.memory2.mem1[56][0] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold424 (.A(\top1.memory2.mem2[152][1] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold425 (.A(\top1.memory2.mem1[46][2] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold426 (.A(\top1.memory2.mem1[147][0] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold427 (.A(\top1.memory2.mem1[115][1] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold428 (.A(\top1.memory2.mem1[115][2] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold429 (.A(\top1.memory1.mem1[116][2] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold430 (.A(\top1.memory1.mem2[154][1] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold431 (.A(\top1.memory1.mem2[125][2] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold432 (.A(\top1.memory1.mem2[191][1] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold433 (.A(\top1.memory1.mem2[102][0] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold434 (.A(\top1.memory2.mem2[172][0] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold435 (.A(\top1.memory1.mem2[23][1] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold436 (.A(\top1.memory2.mem2[155][2] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold437 (.A(\top1.memory1.mem2[116][1] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold438 (.A(\top1.memory1.mem2[106][0] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold439 (.A(\top1.memory1.mem1[31][0] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold440 (.A(\top1.memory2.mem2[108][0] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold441 (.A(\top1.memory2.mem1[22][2] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold442 (.A(\top1.memory1.mem1[41][1] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold443 (.A(\top1.memory1.mem1[101][2] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold444 (.A(\top1.memory1.mem2[178][0] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold445 (.A(\top1.memory1.mem2[21][1] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold446 (.A(\top1.memory2.mem1[11][1] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold447 (.A(\top1.memory2.mem1[165][0] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold448 (.A(\top1.memory2.mem1[171][2] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold449 (.A(\top1.memory2.mem1[105][1] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold450 (.A(\top1.memory2.mem2[35][0] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold451 (.A(\top1.memory2.mem1[180][0] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold452 (.A(\top1.memory1.mem1[60][1] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold453 (.A(\top1.memory1.mem1[43][2] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold454 (.A(\top1.memory2.mem1[169][0] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold455 (.A(\top1.memory1.mem2[44][0] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold456 (.A(\top1.memory2.mem2[86][1] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold457 (.A(\top1.memory1.mem2[105][2] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold458 (.A(\top1.memory2.mem1[176][0] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold459 (.A(\top1.memory2.mem2[191][1] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold460 (.A(\top1.memory1.mem1[85][1] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold461 (.A(\top1.memory2.mem1[21][1] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold462 (.A(\top1.memory2.mem2[56][0] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold463 (.A(\top1.memory1.mem2[14][1] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold464 (.A(\top1.memory2.mem2[34][1] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold465 (.A(\top1.memory1.mem1[168][1] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold466 (.A(\top1.memory2.mem1[47][2] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold467 (.A(\top1.memory1.mem2[33][1] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold468 (.A(\top1.memory2.mem1[56][1] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold469 (.A(\top1.memory2.mem2[117][1] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold470 (.A(\top1.memory1.mem1[125][1] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold471 (.A(\top1.memory2.mem1[57][2] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold472 (.A(\top1.memory1.mem1[23][1] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold473 (.A(\top1.memory1.mem1[157][0] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold474 (.A(\top1.memory1.mem2[176][2] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold475 (.A(\top1.memory2.mem2[151][2] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold476 (.A(\top1.memory2.mem2[39][1] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold477 (.A(\top1.memory2.mem2[183][0] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold478 (.A(\top1.memory1.mem2[32][2] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold479 (.A(\top1.memory2.mem2[112][0] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold480 (.A(\top1.memory2.mem2[189][0] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold481 (.A(\top1.memory2.mem2[71][0] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold482 (.A(\top1.memory1.mem2[163][2] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold483 (.A(\top1.memory1.mem1[155][2] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold484 (.A(\top1.memory2.mem2[61][0] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold485 (.A(\top1.memory1.mem2[35][1] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold486 (.A(\top1.memory2.mem2[48][1] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold487 (.A(\top1.memory2.mem1[92][2] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold488 (.A(\top1.memory1.mem2[108][1] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold489 (.A(\top1.memory2.mem1[29][0] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold490 (.A(\top1.memory1.mem1[178][0] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold491 (.A(\top1.memory2.mem1[35][1] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold492 (.A(\top1.memory1.mem1[87][1] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold493 (.A(\top1.memory1.mem2[40][2] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold494 (.A(\top1.memory2.mem2[165][1] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold495 (.A(\top1.memory1.mem1[22][1] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold496 (.A(\top1.memory2.mem1[167][2] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold497 (.A(\top1.memory2.mem1[46][1] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold498 (.A(\top1.memory1.mem2[28][2] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold499 (.A(\top1.memory2.mem1[34][1] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold500 (.A(\top1.memory2.mem1[125][1] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold501 (.A(\top1.memory1.mem2[89][2] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold502 (.A(\top1.memory1.mem1[192][2] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold503 (.A(\top1.memory1.mem2[150][1] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold504 (.A(\top1.memory1.mem1[48][2] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold505 (.A(\top1.memory2.mem2[16][2] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold506 (.A(\top1.memory1.mem1[185][0] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold507 (.A(\top1.memory1.mem2[118][1] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold508 (.A(\top1.memory2.mem1[109][0] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold509 (.A(\top1.memory1.mem1[105][2] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold510 (.A(\top1.memory1.mem1[71][2] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold511 (.A(\top1.memory2.mem2[91][2] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold512 (.A(\top1.memory1.mem2[27][2] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold513 (.A(\top1.memory1.mem2[119][1] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold514 (.A(\top1.memory2.mem1[7][1] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold515 (.A(\top1.memory2.mem2[183][1] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold516 (.A(\top1.memory1.mem1[164][1] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold517 (.A(\top1.memory1.mem2[50][1] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold518 (.A(\top1.memory2.mem1[61][2] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold519 (.A(\top1.memory1.mem1[122][0] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold520 (.A(\top1.memory1.mem2[20][1] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold521 (.A(\top1.memory1.mem2[193][0] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold522 (.A(\top1.memory1.mem2[110][0] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold523 (.A(\top1.memory2.mem1[169][1] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold524 (.A(\top1.memory2.mem1[17][1] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold525 (.A(\top1.memory1.mem1[61][0] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold526 (.A(\top1.memory1.mem1[192][1] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold527 (.A(\top1.memory2.mem1[45][1] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold528 (.A(\top1.memory1.mem2[85][0] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold529 (.A(\top1.memory2.mem2[126][2] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold530 (.A(\top1.memory2.mem2[95][2] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold531 (.A(\top1.memory1.mem2[61][0] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold532 (.A(\top1.memory2.mem1[120][0] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold533 (.A(\top1.memory2.mem2[147][0] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold534 (.A(\top1.memory1.mem1[149][1] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold535 (.A(\top1.memory2.mem1[93][1] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold536 (.A(\top1.memory1.mem2[37][2] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold537 (.A(\top1.memory2.mem1[119][2] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold538 (.A(\top1.memory2.mem1[185][2] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold539 (.A(\top1.memory1.mem1[16][1] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold540 (.A(\top1.memory2.mem1[195][1] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold541 (.A(\top1.memory2.mem2[33][2] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold542 (.A(\top1.memory1.mem2[170][0] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold543 (.A(\top1.memory2.mem2[31][1] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold544 (.A(\top1.memory2.mem1[57][1] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold545 (.A(\top1.memory1.mem1[169][0] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold546 (.A(\top1.memory2.mem2[192][2] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold547 (.A(\top1.memory2.mem1[120][2] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold548 (.A(\top1.memory1.mem1[169][1] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold549 (.A(\top1.memory1.mem1[14][2] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold550 (.A(\top1.memory2.mem1[55][0] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold551 (.A(\top1.memory1.mem1[19][2] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold552 (.A(\top1.memory2.mem2[167][0] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold553 (.A(\top1.memory1.mem1[95][0] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold554 (.A(\top1.memory1.mem2[180][1] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold555 (.A(\top1.memory1.mem2[17][1] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold556 (.A(\top1.memory2.mem2[29][1] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold557 (.A(\top1.memory1.mem1[25][0] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold558 (.A(\top1.memory1.mem2[103][0] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold559 (.A(\top1.memory1.mem2[63][1] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold560 (.A(\top1.memory2.mem2[45][2] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold561 (.A(\top1.memory2.mem2[197][2] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold562 (.A(\top1.memory1.mem1[17][2] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold563 (.A(\top1.memory2.mem2[44][1] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold564 (.A(\top1.memory2.mem2[20][1] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold565 (.A(\top1.memory2.mem1[154][0] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold566 (.A(\top1.memory2.mem2[58][2] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold567 (.A(\top1.memory2.mem1[192][1] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold568 (.A(\top1.memory2.mem2[54][1] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold569 (.A(\top1.memory1.mem1[191][2] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold570 (.A(\top1.memory1.mem2[193][2] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold571 (.A(\top1.memory2.mem1[185][1] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold572 (.A(\top1.memory2.mem2[120][2] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold573 (.A(\top1.memory1.mem1[114][0] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold574 (.A(\top1.memory2.mem2[169][0] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold575 (.A(\top1.memory1.mem2[168][0] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold576 (.A(\top1.memory1.mem2[197][2] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold577 (.A(\top1.memory2.mem1[152][2] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold578 (.A(\top1.memory2.mem1[115][0] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold579 (.A(\top1.memory1.mem2[89][0] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold580 (.A(\top1.memory2.mem1[26][0] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold581 (.A(\top1.memory1.mem1[120][1] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold582 (.A(\top1.memory2.mem2[14][2] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold583 (.A(\top1.memory2.mem1[87][0] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold584 (.A(\top1.memory2.mem2[92][2] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold585 (.A(\top1.memory2.mem2[173][2] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold586 (.A(\top1.memory2.mem2[14][1] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold587 (.A(\top1.memory1.mem1[95][1] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold588 (.A(\top1.memory2.mem2[164][2] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold589 (.A(\top1.memory2.mem2[163][1] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold590 (.A(\top1.memory2.mem2[120][1] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold591 (.A(\top1.memory1.mem2[36][2] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold592 (.A(\top1.memory1.mem2[169][1] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold593 (.A(\top1.memory1.mem2[155][1] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold594 (.A(\top1.memory1.mem2[187][2] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold595 (.A(\top1.memory1.mem1[193][0] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold596 (.A(\top1.memory1.mem2[171][0] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold597 (.A(\top1.memory1.mem2[46][1] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold598 (.A(\top1.memory1.mem1[184][2] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold599 (.A(\top1.memory1.mem2[149][1] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold600 (.A(\top1.memory1.mem1[39][1] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold601 (.A(\top1.memory2.mem2[168][2] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold602 (.A(\top1.memory2.mem2[158][1] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold603 (.A(\top1.memory1.mem2[91][2] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold604 (.A(\top1.memory1.mem1[113][0] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold605 (.A(\top1.memory1.mem2[184][2] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold606 (.A(\top1.memory1.mem1[151][1] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold607 (.A(\top1.memory1.mem1[90][0] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold608 (.A(\top1.memory2.mem2[188][2] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold609 (.A(\top1.memory1.mem2[45][1] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold610 (.A(\top1.memory2.mem2[111][1] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold611 (.A(\top1.memory1.mem1[40][1] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold612 (.A(\top1.memory2.mem1[151][1] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold613 (.A(\top1.memory1.mem1[163][2] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold614 (.A(\top1.memory2.mem1[164][0] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold615 (.A(\top1.memory1.mem1[176][2] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold616 (.A(\top1.memory1.mem1[182][2] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold617 (.A(\top1.memory2.mem2[40][1] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold618 (.A(\top1.memory1.mem2[95][1] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold619 (.A(\top1.memory1.mem1[176][1] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold620 (.A(\top1.memory1.mem2[194][1] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold621 (.A(\top1.memory2.mem1[178][0] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold622 (.A(\top1.memory1.mem1[33][0] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold623 (.A(\top1.memory2.mem1[52][2] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold624 (.A(\top1.memory2.mem2[19][1] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold625 (.A(\top1.memory1.mem2[151][0] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold626 (.A(\top1.memory2.mem1[125][2] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold627 (.A(\top1.memory1.mem1[121][2] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold628 (.A(\top1.memory2.mem2[103][0] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold629 (.A(\top1.memory1.mem1[197][2] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold630 (.A(\top1.memory2.mem1[34][2] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold631 (.A(\top1.memory1.mem2[121][2] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold632 (.A(\top1.memory1.mem2[156][0] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold633 (.A(\top1.memory1.mem2[54][0] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold634 (.A(\top1.memory1.mem1[163][0] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold635 (.A(\top1.memory1.mem1[27][0] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold636 (.A(\top1.memory2.mem2[176][1] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold637 (.A(\top1.memory2.mem2[71][2] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold638 (.A(\top1.memory1.mem1[158][1] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold639 (.A(\top1.memory1.mem1[183][1] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold640 (.A(\top1.memory2.mem2[174][2] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold641 (.A(\top1.memory2.mem1[94][0] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold642 (.A(\top1.memory2.mem2[189][1] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold643 (.A(\top1.memory2.mem1[44][0] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold644 (.A(\top1.memory2.mem1[58][2] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold645 (.A(\top1.memory2.mem2[16][1] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold646 (.A(\top1.memory1.mem2[30][1] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold647 (.A(\top1.memory2.mem2[191][2] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold648 (.A(\top1.memory1.mem2[93][2] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold649 (.A(\top1.memory1.mem2[171][1] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold650 (.A(\top1.memory1.mem1[187][1] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold651 (.A(\top1.memory2.mem2[154][1] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold652 (.A(\top1.memory1.mem1[154][1] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold653 (.A(\top1.memory2.mem1[53][1] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold654 (.A(\top1.memory1.mem1[185][2] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold655 (.A(\top1.memory2.mem1[27][1] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold656 (.A(\top1.memory2.mem2[38][1] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold657 (.A(\top1.memory2.mem1[108][2] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold658 (.A(\top1.memory2.mem2[107][2] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold659 (.A(\top1.memory1.mem2[60][0] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold660 (.A(\top1.memory2.mem2[118][2] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold661 (.A(\top1.memory2.mem2[23][2] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold662 (.A(\top1.memory2.mem1[150][2] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold663 (.A(\top1.memory1.mem1[49][2] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold664 (.A(\top1.memory1.mem1[27][1] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold665 (.A(\top1.memory2.mem1[20][2] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold666 (.A(\top1.memory1.mem1[24][0] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold667 (.A(\top1.memory1.mem2[17][0] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold668 (.A(\top1.memory2.mem2[181][1] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold669 (.A(\top1.memory1.mem2[117][1] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold670 (.A(\top1.memory1.mem1[7][0] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold671 (.A(\top1.memory2.mem2[194][2] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold672 (.A(\top1.memory1.mem2[181][2] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold673 (.A(\top1.memory1.mem1[37][0] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold674 (.A(\top1.memory1.mem1[119][0] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold675 (.A(\top1.memory2.mem1[152][0] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold676 (.A(\top1.memory1.mem1[101][0] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold677 (.A(\top1.memory2.mem2[124][2] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold678 (.A(\top1.memory2.mem1[20][1] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold679 (.A(\top1.memory1.mem1[103][2] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold680 (.A(\top1.memory2.mem2[165][0] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold681 (.A(\top1.memory1.mem2[153][1] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold682 (.A(\top1.memory1.mem2[29][2] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold683 (.A(\top1.memory2.mem1[49][1] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold684 (.A(\top1.memory1.mem2[111][1] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold685 (.A(\top1.memory1.mem1[21][2] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold686 (.A(\top1.memory1.mem1[108][1] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold687 (.A(\top1.memory2.mem1[119][0] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold688 (.A(\top1.memory2.mem1[94][2] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold689 (.A(\top1.memory2.mem1[45][0] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold690 (.A(\top1.memory1.mem2[26][0] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold691 (.A(\top1.memory1.mem2[25][2] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold692 (.A(\top1.memory2.mem2[188][1] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold693 (.A(\top1.memory2.mem2[21][0] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold694 (.A(\top1.memory1.mem2[36][0] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold695 (.A(\top1.memory1.mem2[163][0] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold696 (.A(\top1.memory2.mem2[153][0] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold697 (.A(\top1.memory2.mem2[21][1] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold698 (.A(\top1.memory1.mem1[121][0] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold699 (.A(\top1.memory2.mem2[182][0] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold700 (.A(\top1.memory2.mem1[172][2] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold701 (.A(\top1.memory1.mem2[147][2] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold702 (.A(\top1.memory1.mem2[173][1] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold703 (.A(\top1.memory1.mem1[35][1] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold704 (.A(\top1.memory1.mem2[48][0] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold705 (.A(\top1.memory2.mem1[11][2] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold706 (.A(\top1.memory2.mem1[195][0] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold707 (.A(\top1.memory2.mem2[187][0] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold708 (.A(\top1.memory1.mem1[196][1] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold709 (.A(\top1.memory1.mem2[196][1] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold710 (.A(\top1.memory1.mem2[105][1] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold711 (.A(\top1.memory2.mem1[124][2] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold712 (.A(\top1.memory2.mem2[86][2] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold713 (.A(\top1.memory2.mem2[92][1] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold714 (.A(\top1.memory2.mem2[108][1] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold715 (.A(\top1.memory2.mem1[36][0] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold716 (.A(\top1.memory2.mem1[57][0] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold717 (.A(\top1.memory2.mem1[173][1] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold718 (.A(\top1.memory2.mem2[174][0] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold719 (.A(\top1.memory1.mem1[181][2] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold720 (.A(\top1.memory2.mem1[153][2] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold721 (.A(\top1.memory1.mem2[175][2] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold722 (.A(\top1.memory2.mem1[148][1] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold723 (.A(\top1.memory1.mem1[110][2] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold724 (.A(\top1.memory1.mem1[166][1] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold725 (.A(\top1.memory2.mem2[31][2] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold726 (.A(\top1.memory2.mem1[108][0] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold727 (.A(\top1.memory2.mem2[122][1] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold728 (.A(\top1.memory2.mem1[165][2] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold729 (.A(\top1.memory2.mem2[190][2] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold730 (.A(\top1.memory1.mem1[164][2] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold731 (.A(\top1.memory1.mem1[39][0] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold732 (.A(\top1.memory1.mem1[101][1] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold733 (.A(\top1.memory2.mem1[39][0] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold734 (.A(\top1.memory1.mem1[17][1] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold735 (.A(\top1.memory2.mem2[166][2] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold736 (.A(\top1.memory2.mem1[110][1] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold737 (.A(\top1.memory1.mem1[167][1] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold738 (.A(\top1.memory1.mem2[20][0] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold739 (.A(\top1.memory1.mem1[124][1] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold740 (.A(\top1.memory1.mem1[191][0] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold741 (.A(\top1.memory1.mem2[183][1] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold742 (.A(\top1.memory2.mem2[185][1] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold743 (.A(\top1.memory2.mem2[152][0] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold744 (.A(\top1.memory1.mem1[30][1] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold745 (.A(\top1.memory1.mem2[103][2] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold746 (.A(\top1.memory1.mem2[156][2] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold747 (.A(\top1.memory2.mem2[34][0] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold748 (.A(\top1.memory1.mem1[91][0] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold749 (.A(\top1.memory1.mem1[89][2] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold750 (.A(\top1.memory2.mem2[16][0] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold751 (.A(\top1.memory1.mem1[149][2] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold752 (.A(\top1.memory1.mem1[86][2] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold753 (.A(\top1.memory2.mem2[7][2] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold754 (.A(\top1.memory1.mem2[94][2] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold755 (.A(\top1.memory2.mem1[30][0] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold756 (.A(\top1.memory1.mem2[172][0] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold757 (.A(\top1.memory2.mem2[35][2] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold758 (.A(\top1.memory2.mem2[60][0] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold759 (.A(\top1.memory1.mem2[53][1] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold760 (.A(\top1.memory2.mem2[32][1] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold761 (.A(\top1.memory1.mem2[47][2] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold762 (.A(\top1.memory1.mem1[170][0] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold763 (.A(\top1.memory1.mem1[190][2] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold764 (.A(\top1.memory2.mem1[41][0] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold765 (.A(\top1.memory1.mem2[86][2] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold766 (.A(\top1.memory2.mem2[149][0] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold767 (.A(\top1.memory1.mem1[31][1] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold768 (.A(\top1.memory1.mem1[178][1] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold769 (.A(\top1.memory2.mem1[40][2] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold770 (.A(\top1.memory2.mem2[113][2] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold771 (.A(\top1.memory1.mem1[150][0] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold772 (.A(\top1.memory1.mem2[188][0] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold773 (.A(\top1.memory2.mem1[171][1] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold774 (.A(\top1.memory2.mem2[11][1] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold775 (.A(\top1.memory2.mem2[114][2] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold776 (.A(\top1.memory2.mem1[86][0] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold777 (.A(\top1.memory2.mem2[13][2] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold778 (.A(\top1.memory2.mem1[186][0] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold779 (.A(\top1.memory2.mem1[42][1] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold780 (.A(\top1.memory2.mem1[112][2] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold781 (.A(\top1.memory1.mem1[52][0] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold782 (.A(\top1.memory2.mem2[7][0] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold783 (.A(\top1.memory1.mem2[26][1] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold784 (.A(\top1.memory2.mem2[89][0] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold785 (.A(\top1.memory2.mem2[187][2] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold786 (.A(\top1.memory2.mem2[116][1] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold787 (.A(\top1.memory2.mem1[37][1] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold788 (.A(\top1.memory1.mem2[126][2] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold789 (.A(\top1.memory1.mem2[167][2] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold790 (.A(\top1.memory1.mem2[120][1] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold791 (.A(\top1.memory2.mem1[40][1] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold792 (.A(\top1.memory2.mem1[159][1] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold793 (.A(\top1.memory1.mem2[180][0] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold794 (.A(\top1.memory1.mem1[59][1] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold795 (.A(\top1.memory2.mem1[111][2] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold796 (.A(\top1.memory1.mem2[53][2] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold797 (.A(\top1.memory1.mem2[176][1] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold798 (.A(\top1.memory2.mem2[159][2] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold799 (.A(\top1.memory1.mem1[151][2] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold800 (.A(\top1.memory1.mem1[92][2] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold801 (.A(\top1.memory1.mem2[62][0] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold802 (.A(\top1.memory1.mem2[192][1] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold803 (.A(\top1.memory2.mem2[179][1] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold804 (.A(\top1.memory2.mem2[187][1] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold805 (.A(\top1.memory2.mem2[30][1] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold806 (.A(\top1.memory1.mem1[50][0] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold807 (.A(\top1.memory1.mem1[54][2] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold808 (.A(\top1.memory1.mem2[114][0] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold809 (.A(\top1.memory1.mem2[13][2] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold810 (.A(\top1.memory2.mem2[179][2] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold811 (.A(\top1.memory1.mem1[34][0] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold812 (.A(\top1.memory2.mem1[118][1] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold813 (.A(\top1.memory1.mem1[198][0] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold814 (.A(\top1.memory1.mem2[180][2] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold815 (.A(\top1.memory2.mem2[41][0] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold816 (.A(\top1.memory2.mem1[19][0] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold817 (.A(\top1.memory1.mem2[58][2] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold818 (.A(\top1.memory2.mem1[48][2] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold819 (.A(\top1.memory2.mem2[19][2] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold820 (.A(\top1.memory1.mem2[31][0] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold821 (.A(\top1.memory2.mem2[176][0] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold822 (.A(\top1.memory2.mem2[195][2] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold823 (.A(\top1.memory2.mem1[107][2] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold824 (.A(\top1.memory1.mem1[179][0] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold825 (.A(\top1.memory1.mem2[164][2] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold826 (.A(\top1.memory1.mem2[182][2] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold827 (.A(\top1.memory1.mem1[21][1] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold828 (.A(\top1.memory1.mem1[46][1] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold829 (.A(\top1.memory1.mem1[125][2] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold830 (.A(\top1.memory1.mem1[86][1] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold831 (.A(\top1.memory1.mem1[175][1] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold832 (.A(\top1.memory2.mem2[166][0] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold833 (.A(\top1.memory2.mem1[110][0] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold834 (.A(\top1.memory2.mem2[198][2] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold835 (.A(\top1.memory2.mem1[198][1] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold836 (.A(\top1.memory2.mem1[181][2] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold837 (.A(\top1.memory2.mem1[126][1] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold838 (.A(\top1.memory1.mem1[186][0] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold839 (.A(\top1.memory2.mem2[53][2] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold840 (.A(\top1.memory2.mem1[182][2] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold841 (.A(\top1.memory1.mem2[174][0] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold842 (.A(\top1.memory2.mem1[177][0] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold843 (.A(\top1.memory2.mem1[29][1] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold844 (.A(\top1.memory1.mem1[180][0] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold845 (.A(\top1.memory2.mem2[114][0] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold846 (.A(\top1.memory2.mem1[158][2] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold847 (.A(\top1.memory2.mem2[121][2] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold848 (.A(\top1.memory2.mem1[149][0] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold849 (.A(\top1.memory2.mem2[112][2] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold850 (.A(\top1.memory1.mem1[152][2] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold851 (.A(\top1.memory2.mem1[113][2] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold852 (.A(\top1.memory1.mem2[107][1] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold853 (.A(\top1.memory1.mem2[187][0] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold854 (.A(\top1.memory2.mem1[198][2] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold855 (.A(\top1.memory1.mem1[116][0] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold856 (.A(\top1.memory1.mem1[168][2] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold857 (.A(\top1.memory1.mem1[54][1] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold858 (.A(\top1.memory2.mem2[49][2] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold859 (.A(\top1.memory2.mem2[194][0] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold860 (.A(\top1.memory1.mem1[117][0] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold861 (.A(\top1.memory1.mem2[71][1] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold862 (.A(\top1.memory1.mem1[105][0] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold863 (.A(\top1.memory2.mem2[155][0] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold864 (.A(\top1.memory1.mem2[165][0] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold865 (.A(\top1.memory1.mem1[21][0] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold866 (.A(\top1.memory1.mem1[106][1] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold867 (.A(\top1.memory2.mem2[163][0] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold868 (.A(\top1.memory2.mem2[113][0] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold869 (.A(\top1.memory2.mem1[149][2] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold870 (.A(\top1.memory2.mem1[41][1] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold871 (.A(\top1.memory2.mem1[91][1] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold872 (.A(\top1.memory1.mem2[173][0] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold873 (.A(\top1.memory1.mem1[153][0] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold874 (.A(\top1.memory2.mem1[164][2] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold875 (.A(\top1.memory1.mem2[157][1] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold876 (.A(\top1.memory2.mem2[103][2] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold877 (.A(\top1.memory2.mem1[155][1] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold878 (.A(\top1.memory1.mem1[108][0] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold879 (.A(\top1.memory2.mem1[175][0] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold880 (.A(\top1.memory2.mem2[38][2] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold881 (.A(\top1.memory2.mem2[112][1] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold882 (.A(\top1.memory2.mem2[176][2] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold883 (.A(\top1.memory2.mem1[18][2] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold884 (.A(\top1.memory2.mem1[50][2] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold885 (.A(\top1.memory2.mem2[110][2] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold886 (.A(\top1.memory2.mem2[47][0] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold887 (.A(\top1.memory2.mem2[197][0] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold888 (.A(\top1.memory1.mem2[195][1] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold889 (.A(\top1.memory2.mem1[140][0] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold890 (.A(\top1.memory2.mem1[18][1] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold891 (.A(\top1.memory1.mem1[25][2] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold892 (.A(\top1.memory2.mem2[95][0] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold893 (.A(\top1.memory1.mem2[62][1] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold894 (.A(\top1.memory2.mem1[32][0] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold895 (.A(\top1.memory2.mem1[26][1] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold896 (.A(\top1.memory1.mem2[106][1] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold897 (.A(\top1.memory2.mem1[42][0] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold898 (.A(\top1.memory1.mem1[38][2] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold899 (.A(\top1.memory2.mem2[185][2] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold900 (.A(\top1.memory1.mem1[124][2] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold901 (.A(\top1.memory2.mem2[86][0] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold902 (.A(\top1.memory2.mem2[192][0] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold903 (.A(\top1.memory1.mem2[188][1] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold904 (.A(\top1.memory1.mem2[16][0] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold905 (.A(\top1.memory1.mem2[118][2] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold906 (.A(\top1.memory2.mem2[156][2] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold907 (.A(\top1.memory2.mem2[189][2] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold908 (.A(\top1.memory2.mem1[150][1] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold909 (.A(\top1.memory2.mem1[41][2] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold910 (.A(\top1.memory1.mem2[112][1] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold911 (.A(\top1.memory1.mem2[118][0] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold912 (.A(\top1.memory2.mem1[62][2] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold913 (.A(\top1.memory2.mem1[168][2] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold914 (.A(\top1.memory2.mem1[63][1] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold915 (.A(\top1.memory1.mem2[11][1] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold916 (.A(\top1.memory1.mem1[157][2] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold917 (.A(\top1.memory2.mem1[188][1] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold918 (.A(\top1.memory2.mem1[149][1] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold919 (.A(\top1.memory2.mem2[158][2] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold920 (.A(\top1.memory1.mem2[31][1] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold921 (.A(\top1.memory2.mem1[187][1] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold922 (.A(\top1.memory1.mem1[35][2] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold923 (.A(\top1.memory1.mem1[11][1] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold924 (.A(\top1.memory2.mem2[182][1] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold925 (.A(\top1.memory2.mem2[171][0] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold926 (.A(\top1.memory2.mem1[28][1] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold927 (.A(\top1.memory1.mem1[52][1] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold928 (.A(\top1.memory1.mem1[115][1] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold929 (.A(\top1.memory1.mem2[120][2] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold930 (.A(\top1.memory2.mem2[58][1] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold931 (.A(\top1.memory1.mem2[126][0] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold932 (.A(\top1.memory1.mem2[39][1] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold933 (.A(\top1.memory1.mem1[170][1] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold934 (.A(\top1.memory1.mem1[48][0] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold935 (.A(\top1.memory2.mem1[179][0] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold936 (.A(\top1.memory1.mem2[186][1] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold937 (.A(\top1.memory2.mem2[194][1] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold938 (.A(\top1.memory1.mem2[179][0] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold939 (.A(\top1.memory2.mem1[197][0] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold940 (.A(\top1.memory1.mem2[174][1] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold941 (.A(\top1.memory2.mem1[168][1] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold942 (.A(\top1.memory2.mem2[106][2] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold943 (.A(\top1.memory1.mem1[85][2] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold944 (.A(\top1.memory1.mem1[33][2] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold945 (.A(\top1.memory1.mem1[49][1] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold946 (.A(\top1.memory1.mem1[114][1] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold947 (.A(\top1.memory2.mem1[112][0] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold948 (.A(\top1.memory1.mem2[36][1] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold949 (.A(\top1.memory2.mem1[53][2] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold950 (.A(\top1.memory2.mem2[116][2] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold951 (.A(\top1.memory1.mem2[112][0] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold952 (.A(\top1.memory1.mem2[0][2] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold953 (.A(\top1.memory2.mem2[109][1] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold954 (.A(\top1.memory1.mem1[106][0] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold955 (.A(\top1.memory2.mem2[93][1] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold956 (.A(\top1.memory2.mem1[118][2] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold957 (.A(\top1.memory2.mem1[114][0] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold958 (.A(\top1.memory1.mem1[71][0] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold959 (.A(\top1.memory2.mem2[37][2] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold960 (.A(\top1.memory2.mem1[157][2] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold961 (.A(\top1.memory1.mem2[30][2] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold962 (.A(\top1.memory1.mem2[44][2] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold963 (.A(\top1.memory2.mem2[124][0] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold964 (.A(\top1.memory2.mem1[19][1] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold965 (.A(\top1.memory1.mem2[115][0] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold966 (.A(\top1.memory1.mem1[117][2] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold967 (.A(\top1.memory1.mem1[183][0] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold968 (.A(\top1.memory1.mem1[174][1] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold969 (.A(\top1.memory1.mem1[115][0] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold970 (.A(\top1.memory1.mem2[40][0] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold971 (.A(\top1.memory1.mem1[113][1] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold972 (.A(\top1.memory1.mem2[39][0] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold973 (.A(\top1.memory1.mem2[50][2] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold974 (.A(\top1.memory2.mem2[22][2] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold975 (.A(\top1.memory2.mem2[63][2] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold976 (.A(\top1.memory1.mem1[159][1] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold977 (.A(\top1.memory2.mem1[48][1] ),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold978 (.A(\top1.memory1.mem1[40][2] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold979 (.A(\top1.memory1.mem2[121][1] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold980 (.A(\top1.memory2.mem1[25][0] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold981 (.A(\top1.memory2.mem2[94][2] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold982 (.A(\top1.memory1.mem1[45][0] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold983 (.A(\top1.memory2.mem1[116][2] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold984 (.A(\top1.memory1.mem1[31][2] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold985 (.A(\top1.memory1.mem2[27][0] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold986 (.A(\top1.memory1.mem1[51][1] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold987 (.A(\top1.memory1.mem1[94][2] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold988 (.A(\top1.memory1.mem2[43][0] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold989 (.A(\top1.memory1.mem2[167][1] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold990 (.A(\top1.memory1.mem2[189][0] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold991 (.A(\top1.memory2.mem2[85][1] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold992 (.A(\top1.memory1.mem1[19][0] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold993 (.A(\top1.memory1.mem1[194][1] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold994 (.A(\top1.memory1.mem1[188][2] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold995 (.A(\top1.memory2.mem1[18][0] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold996 (.A(\top1.memory1.mem1[47][2] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold997 (.A(\top1.memory1.mem2[148][2] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold998 (.A(\top1.memory1.mem2[140][1] ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold999 (.A(\top1.memory1.mem2[52][1] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\top1.memory2.mem1[26][2] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\top1.memory2.mem1[170][0] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\top1.memory2.mem1[188][0] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\top1.memory2.mem1[128][0] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\top1.memory2.mem1[93][2] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\top1.memory2.mem2[21][2] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\top1.memory1.mem1[154][0] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\top1.memory2.mem2[60][1] ),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\top1.memory1.mem2[154][2] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\top1.memory2.mem2[124][1] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\top1.memory2.mem1[27][2] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\top1.memory2.mem1[75][0] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\top1.memory1.mem1[11][0] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\top1.memory1.mem1[29][2] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\top1.memory2.mem2[185][0] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\top1.memory2.mem1[120][1] ),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\top1.memory2.mem2[18][1] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\top1.memory2.mem2[23][1] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\top1.memory1.mem2[94][1] ),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\top1.memory1.mem1[167][2] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\top1.memory2.mem1[151][2] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\top1.memory1.mem1[38][1] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\top1.memory1.mem2[13][0] ),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\top1.memory1.mem2[49][2] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\top1.memory2.mem1[176][1] ),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\top1.memory2.mem2[15][2] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\top1.memory2.mem2[106][0] ),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\top1.memory2.mem2[150][2] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\top1.memory1.mem1[173][0] ),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\top1.memory2.mem1[33][0] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\top1.memory1.mem1[194][2] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\top1.memory1.mem1[47][0] ),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\top1.memory2.mem1[136][2] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\top1.memory2.mem2[45][0] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\top1.memory2.mem2[42][1] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\top1.memory1.mem1[59][0] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\top1.memory1.mem2[41][2] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\top1.memory1.mem2[85][2] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\top1.memory1.mem2[143][2] ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\top1.memory2.mem1[49][2] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\top1.memory2.mem1[16][2] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\top1.memory2.mem2[198][0] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\top1.memory1.mem2[45][2] ),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\top1.memory1.mem1[36][2] ),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\top1.memory2.mem1[59][2] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\top1.memory1.mem2[198][1] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\top1.memory2.mem2[17][2] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\top1.memory2.mem1[165][1] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\top1.memory1.mem1[58][1] ),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\top1.memory1.mem2[101][1] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\top1.memory1.mem1[179][1] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\top1.memory2.mem2[54][2] ),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\top1.memory1.mem1[172][2] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\top1.memory2.mem1[168][0] ),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\top1.memory2.mem1[24][2] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\top1.memory2.mem2[29][2] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\top1.memory1.mem1[149][0] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\top1.memory1.mem1[18][0] ),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\top1.memory2.mem1[58][0] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\top1.memory1.mem1[58][0] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\top1.memory1.mem1[117][1] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\top1.memory2.mem2[151][0] ),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\top1.memory1.mem2[181][1] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\top1.memory2.mem1[158][1] ),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\top1.memory1.mem2[116][0] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\top1.memory2.mem1[36][1] ),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\top1.memory2.mem2[172][1] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\top1.memory2.mem2[90][1] ),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\top1.memory1.mem2[101][2] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\top1.memory2.mem2[151][1] ),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\top1.memory1.mem2[48][2] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\top1.memory2.mem2[91][1] ),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\top1.memory2.mem1[7][0] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\top1.memory2.mem1[25][1] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\top1.memory2.mem2[149][2] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\top1.memory2.mem2[150][0] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\top1.memory2.mem2[178][0] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\top1.memory1.mem2[46][0] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\top1.memory1.mem1[148][0] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\top1.memory1.mem2[186][2] ),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\top1.memory1.mem2[147][0] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\top1.memory2.mem2[115][2] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\top1.memory2.mem2[63][0] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\top1.memory2.mem1[116][1] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\top1.memory1.mem2[190][0] ),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\top1.memory1.mem2[139][0] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\top1.memory1.mem1[62][2] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\top1.memory1.mem2[109][2] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\top1.memory2.mem2[148][2] ),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\top1.memory2.mem2[147][2] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\top1.memory1.mem1[90][1] ),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\top1.memory2.mem1[106][1] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\top1.memory1.mem2[63][0] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\top1.memory2.mem2[181][2] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\top1.memory2.mem1[35][0] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\top1.memory1.mem2[14][2] ),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\top1.memory2.mem1[111][0] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\top1.memory2.mem1[45][2] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\top1.memory2.mem1[113][0] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\top1.memory1.mem2[57][0] ),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\top1.memory1.mem1[86][0] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\top1.memory1.mem2[55][1] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\top1.memory2.mem2[29][0] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\top1.memory2.mem2[175][0] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\top1.memory1.mem2[160][0] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\top1.memory2.mem1[54][0] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\top1.memory2.mem2[22][1] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\top1.memory1.mem2[159][2] ),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\top1.memory1.mem1[126][0] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\top1.memory2.mem2[169][2] ),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\top1.memory1.mem2[163][1] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\top1.memory2.mem2[105][1] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\top1.memory1.mem1[122][2] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\top1.memory2.mem1[28][2] ),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\top1.memory2.mem2[51][2] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\top1.memory1.mem1[156][2] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\top1.memory1.mem1[173][1] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\top1.memory1.mem1[88][1] ),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\top1.memory2.mem2[165][2] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\top1.memory1.mem2[117][2] ),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\top1.memory1.mem1[148][2] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\top1.memory2.mem1[44][1] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\top1.memory1.mem1[61][2] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\top1.memory1.mem1[189][2] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\top1.memory2.mem2[45][1] ),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\top1.memory1.mem1[109][1] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\top1.memory2.mem2[157][2] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\top1.memory1.mem1[194][0] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\top1.memory1.mem2[120][0] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\top1.memory1.mem1[123][1] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\top1.memory2.mem2[148][0] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\top1.memory2.mem1[7][2] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\top1.memory2.mem1[143][2] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\top1.memory2.mem2[196][1] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\top1.memory1.mem2[113][2] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\top1.memory1.mem1[172][1] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\top1.memory2.mem2[50][0] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\top1.memory2.mem2[186][1] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\top1.memory1.mem1[196][0] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\top1.memory1.mem1[180][1] ),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\top1.memory2.mem1[95][0] ),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\top1.memory2.mem2[156][1] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\top1.memory1.mem2[21][0] ),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\top1.memory2.mem2[50][2] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\top1.memory2.mem2[26][2] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\top1.memory2.mem2[177][0] ),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\top1.memory1.mem1[60][2] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\top1.memory2.mem1[94][1] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\top1.memory1.mem2[194][2] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\top1.memory2.mem2[57][0] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\top1.memory1.mem1[38][0] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\top1.memory1.mem2[34][1] ),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\top1.memory1.mem2[195][0] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\top1.memory2.mem1[148][2] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\top1.memory1.mem1[129][1] ),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\top1.memory2.mem1[19][2] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\top1.memory2.mem1[193][0] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\top1.memory2.mem1[159][2] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\top1.memory2.mem2[107][1] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\top1.memory2.mem2[94][1] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\top1.memory2.mem2[111][0] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\top1.memory1.mem2[165][1] ),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\top1.memory1.mem1[55][2] ),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\top1.memory2.mem1[154][1] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\top1.memory2.mem2[195][1] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\top1.memory2.mem2[25][0] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\top1.memory1.mem2[59][2] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\top1.memory1.mem1[45][1] ),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\top1.memory1.mem1[14][1] ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\top1.memory1.mem1[111][1] ),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\top1.memory2.mem1[107][0] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\top1.memory2.mem2[41][2] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\top1.memory2.mem1[38][0] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\top1.memory2.mem2[59][0] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\top1.memory2.mem1[76][0] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\top1.memory2.mem1[156][2] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\top1.memory1.mem1[30][0] ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\top1.memory1.mem2[169][2] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\top1.memory1.mem1[126][1] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\top1.memory2.mem1[101][2] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\top1.memory2.mem2[62][1] ),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\top1.memory2.mem2[157][0] ),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\top1.memory1.mem1[110][0] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\top1.memory1.mem2[62][2] ),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\top1.memory2.mem1[23][1] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\top1.memory1.mem1[45][2] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\top1.memory2.mem1[197][1] ),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\top1.memory1.mem2[7][1] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\top1.memory1.mem1[118][0] ),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\top1.memory2.mem2[144][1] ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\top1.memory1.mem1[55][0] ),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\top1.memory2.mem1[43][1] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\top1.memory2.mem1[61][0] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\top1.memory1.mem2[85][1] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\top1.memory1.mem2[104][0] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\top1.memory2.mem1[13][2] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\top1.memory1.mem2[173][2] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\top1.memory2.mem1[124][0] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\top1.memory2.mem2[32][0] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\top1.memory2.mem1[177][1] ),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\top1.memory1.mem1[63][0] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\top1.memory1.mem1[112][0] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\top1.memory1.mem2[90][2] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\top1.memory2.mem1[174][0] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\top1.memory2.mem1[197][2] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\top1.memory1.mem1[181][0] ),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\top1.memory1.mem2[69][0] ),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\top1.memory2.mem2[30][0] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\top1.memory1.mem1[93][2] ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\top1.memory1.mem1[64][0] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\top1.memory1.mem1[167][0] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\top1.memory1.mem2[71][0] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\top1.memory2.mem2[107][0] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\top1.memory2.mem1[172][0] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\top1.memory2.mem2[131][1] ),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\top1.memory1.mem1[106][2] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\top1.memory2.mem2[126][1] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\top1.memory1.mem1[136][1] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\top1.memory1.mem2[34][2] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\top1.memory1.mem2[3][2] ),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\top1.memory2.mem1[182][1] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\top1.memory1.mem2[179][2] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\top1.memory1.mem1[23][2] ),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\top1.memory1.mem2[116][2] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\top1.memory1.mem1[168][0] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\top1.memory2.mem2[115][0] ),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\top1.memory2.mem1[37][0] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\top1.memory1.mem2[94][0] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\top1.memory2.mem2[128][2] ),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\top1.memory1.mem1[57][1] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\top1.memory2.mem2[94][0] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\top1.memory2.mem1[178][2] ),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\top1.memory2.mem1[23][0] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\top1.memory2.mem2[55][1] ),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\top1.memory1.mem1[110][1] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\top1.memory2.mem1[161][0] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\top1.memory2.mem2[197][1] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\top1.memory1.mem1[57][0] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\top1.memory2.mem2[101][1] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\top1.memory2.mem1[63][2] ),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\top1.memory2.mem2[92][0] ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\top1.memory1.mem2[87][0] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\top1.memory2.mem1[30][2] ),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\top1.memory2.mem1[36][2] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\top1.memory1.mem2[148][0] ),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\top1.memory2.mem1[153][0] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\top1.memory1.mem1[192][0] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\top1.memory1.mem1[166][0] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\top1.memory1.mem1[177][1] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\top1.memory2.mem2[61][2] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\top1.memory2.mem1[106][0] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\top1.memory1.mem1[187][0] ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\top1.memory1.mem2[38][2] ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\top1.memory1.mem2[196][2] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\top1.memory2.mem1[158][0] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\top1.memory1.mem2[181][0] ),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\top1.memory1.mem1[177][0] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\top1.memory1.mem1[107][0] ),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\top1.memory2.mem1[72][2] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\top1.memory1.mem2[185][0] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\top1.memory1.mem2[18][1] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\top1.memory1.mem1[103][1] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\top1.memory1.mem2[196][0] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\top1.memory2.mem2[1][2] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\top1.memory1.mem2[170][1] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\top1.memory1.mem1[189][0] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\top1.memory1.mem1[107][1] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\top1.memory1.mem1[92][1] ),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\top1.memory1.mem2[166][2] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\top1.memory1.mem2[11][2] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\top1.memory2.mem1[38][1] ),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\top1.memory1.mem1[42][1] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\top1.memory2.mem2[80][1] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\top1.memory2.mem1[58][1] ),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\top1.memory2.mem1[66][0] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\top1.memory1.mem2[185][2] ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\top1.memory2.mem1[136][0] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\top1.memory2.mem1[46][0] ),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\top1.memory1.mem1[156][1] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\top1.memory2.mem2[190][1] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\top1.memory1.mem1[28][2] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\top1.memory2.mem1[38][2] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\top1.memory1.mem2[115][1] ),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\top1.memory1.mem1[109][2] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\top1.memory1.mem2[102][2] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\top1.memory2.mem1[54][2] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\top1.memory2.mem1[106][2] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\top1.memory1.mem1[60][0] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\top1.memory2.mem1[172][1] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\top1.memory1.mem2[55][0] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\top1.memory2.mem2[178][2] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\top1.memory2.mem1[49][0] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\top1.memory1.mem1[9][2] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\top1.memory1.mem1[128][2] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\top1.memory1.mem2[117][0] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\top1.memory2.mem1[151][0] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\top1.memory1.mem2[191][2] ),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\top1.memory1.mem2[57][1] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\top1.memory2.mem1[108][1] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\top1.memory2.mem2[155][1] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\top1.memory1.mem2[45][0] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\top1.memory2.mem2[122][2] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\top1.memory1.mem1[29][0] ),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\top1.memory1.mem2[87][1] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\top1.memory1.mem1[114][2] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\top1.memory2.mem2[196][0] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\top1.memory2.mem2[175][1] ),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\top1.memory1.mem1[26][0] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\top1.memory2.mem2[25][1] ),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\top1.memory2.mem1[42][2] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\top1.memory1.mem1[158][2] ),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\top1.memory2.mem1[109][1] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\top1.memory2.mem1[52][1] ),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\top1.memory1.mem2[46][2] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\top1.memory2.mem1[185][0] ),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\top1.memory2.mem2[20][2] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\top1.memory2.mem1[153][1] ),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\top1.memory2.mem1[141][1] ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\top1.memory2.mem2[12][0] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\top1.memory1.mem1[30][2] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\top1.memory2.mem2[57][2] ),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\top1.memory2.mem2[42][2] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\top1.memory2.mem2[78][1] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\top1.memory2.mem2[196][2] ),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\top1.memory2.mem1[22][1] ),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\top1.memory2.mem1[163][2] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\top1.memory1.mem2[123][0] ),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\top1.memory1.mem2[33][0] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\top1.memory1.mem1[151][0] ),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\top1.memory1.mem2[24][0] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\top1.memory2.mem1[188][2] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\top1.memory2.mem2[167][1] ),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\top1.memory1.mem2[178][2] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\top1.memory1.mem1[52][2] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\top1.memory1.mem1[142][0] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\top1.memory2.mem2[117][0] ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\top1.memory2.mem2[148][1] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\top1.memory2.mem1[190][0] ),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\top1.memory1.mem1[53][2] ),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\top1.memory2.mem1[31][0] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\top1.memory1.mem2[14][0] ),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\top1.memory1.mem1[88][0] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\top1.memory2.mem1[16][0] ),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\top1.memory2.mem2[121][1] ),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\top1.memory1.mem2[86][0] ),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\top1.memory2.mem2[68][1] ),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\top1.memory1.mem1[126][2] ),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\top1.memory2.mem1[15][0] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\top1.memory2.mem2[125][0] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\top1.memory1.mem2[92][0] ),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\top1.memory1.mem1[166][2] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\top1.memory1.mem2[42][1] ),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\top1.memory1.mem2[165][2] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\top1.memory2.mem2[62][0] ),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\top1.memory1.mem1[195][0] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\top1.memory1.mem2[10][2] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\top1.memory2.mem2[47][1] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\top1.memory2.mem2[84][2] ),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\top1.memory1.mem2[113][1] ),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\top1.memory1.mem2[18][0] ),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\top1.memory1.mem1[13][1] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\top1.memory2.mem1[85][1] ),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\top1.memory1.mem1[89][1] ),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\top1.memory1.mem2[185][1] ),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\top1.memory1.mem2[162][1] ),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\top1.memory2.mem2[49][1] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\top1.memory2.mem1[118][0] ),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\top1.memory2.mem2[178][1] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\top1.memory2.mem1[157][0] ),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\top1.memory1.mem1[123][0] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\top1.memory1.mem2[32][1] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\top1.memory2.mem2[145][1] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\top1.memory1.mem2[25][1] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\top1.memory1.mem2[109][1] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\top1.memory2.mem1[71][0] ),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\top1.memory1.mem2[177][1] ),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\top1.memory2.mem2[96][1] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\top1.memory1.mem2[47][1] ),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\top1.memory1.mem1[12][1] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\top1.memory2.mem1[75][1] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\top1.memory2.mem1[121][2] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\top1.memory2.mem2[170][1] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\top1.memory1.mem2[146][1] ),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\top1.memory1.mem2[41][0] ),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\top1.memory1.mem2[24][1] ),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\top1.memory2.mem1[29][2] ),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\top1.memory2.mem2[123][1] ),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\top1.memory1.mem2[89][1] ),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\top1.memory2.mem1[116][0] ),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\top1.memory1.mem2[147][1] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\top1.memory1.mem1[10][2] ),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\top1.memory2.mem2[110][0] ),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\top1.memory1.mem1[19][1] ),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\top1.memory2.mem1[152][1] ),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\top1.memory2.mem1[39][2] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\top1.memory1.mem2[124][0] ),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\top1.memory1.mem1[102][1] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\top1.memory2.mem1[189][1] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\top1.memory2.mem1[37][2] ),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\top1.memory1.mem1[25][1] ),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\top1.memory2.mem2[52][2] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\top1.memory1.mem1[34][2] ),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\top1.memory2.mem1[96][1] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\top1.memory1.mem1[39][2] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\top1.memory2.mem1[51][0] ),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\top1.memory1.mem2[174][2] ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\top1.memory1.mem2[149][0] ),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\top1.memory1.mem1[178][2] ),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\top1.memory1.mem1[94][1] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\top1.memory1.mem2[106][2] ),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\top1.memory2.mem2[59][1] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\top1.memory1.mem1[119][2] ),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\top1.memory1.mem1[139][2] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\top1.memory1.mem1[116][1] ),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\top1.memory1.mem2[39][2] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\top1.memory2.mem1[64][2] ),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\top1.memory1.mem2[166][0] ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\top1.memory2.mem2[4][1] ),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\top1.memory1.mem2[182][0] ),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\top1.memory2.mem2[63][1] ),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\top1.memory1.mem1[131][2] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\top1.memory1.mem1[77][2] ),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\top1.memory2.mem1[31][2] ),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\top1.memory2.mem1[14][1] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\top1.memory1.mem1[118][2] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\top1.memory1.mem2[136][1] ),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\top1.memory1.mem2[128][1] ),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\top1.memory1.mem2[67][0] ),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\top1.memory2.mem1[192][0] ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\top1.memory2.mem1[123][2] ),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\top1.memory2.mem1[40][0] ),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\top1.memory1.mem2[119][2] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\top1.memory1.mem2[63][2] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\top1.memory1.mem2[74][1] ),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\top1.memory1.mem1[34][1] ),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\top1.memory1.mem2[78][2] ),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\top1.memory1.mem1[107][2] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\top1.memory2.mem2[67][2] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\top1.memory2.mem1[105][0] ),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\top1.memory1.mem1[16][0] ),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\top1.memory1.mem2[102][1] ),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\top1.memory2.mem2[81][2] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\top1.memory2.mem2[179][0] ),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\top1.memory2.mem1[117][0] ),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\top1.memory2.mem1[72][0] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\top1.memory1.mem2[171][2] ),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\top1.memory1.mem1[69][0] ),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\top1.memory1.mem1[144][2] ),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\top1.memory2.mem2[121][0] ),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\top1.memory2.mem2[186][0] ),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\top1.memory2.mem2[85][0] ),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\top1.memory2.mem2[154][2] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\top1.memory2.mem2[140][1] ),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\top1.memory1.mem2[22][1] ),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\top1.memory1.mem1[175][2] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\top1.memory1.mem2[136][0] ),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\top1.memory2.mem1[9][1] ),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\top1.memory1.mem2[109][0] ),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\top1.memory1.mem2[190][2] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\top1.memory2.mem1[127][1] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\top1.memory1.mem2[91][1] ),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\top1.memory1.mem2[19][1] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\top1.memory2.mem1[60][1] ),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\top1.memory1.mem2[133][0] ),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\top1.memory1.mem1[150][2] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\top1.memory1.mem2[77][0] ),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\top1.memory2.mem2[136][1] ),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\top1.memory1.mem2[197][1] ),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\top1.memory1.mem2[133][1] ),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\top1.memory1.mem2[20][2] ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\top1.memory1.mem2[188][2] ),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\top1.memory2.mem2[17][1] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\top1.memory1.mem1[196][2] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\top1.memory2.mem2[102][1] ),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\top1.memory2.mem2[42][0] ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\top1.memory2.mem1[50][1] ),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\top1.memory1.mem2[75][0] ),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\top1.memory2.mem1[104][0] ),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\top1.memory1.mem1[138][1] ),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\top1.memory1.mem1[4][2] ),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\top1.memory1.mem1[133][2] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\top1.memory1.mem1[13][2] ),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\top1.memory2.mem1[138][0] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\top1.memory1.mem1[100][1] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\top1.memory1.mem1[40][0] ),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\top1.memory1.mem1[122][1] ),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\top1.memory2.mem1[50][0] ),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\top1.memory2.mem2[37][0] ),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\top1.memory2.mem1[133][1] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\top1.memory2.mem2[172][2] ),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\top1.memory1.mem1[137][0] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\top1.memory2.mem2[102][2] ),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\top1.memory1.mem2[178][1] ),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\top1.memory1.mem1[37][2] ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\top1.memory1.mem2[190][1] ),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\top1.memory2.mem1[33][1] ),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\top1.memory1.mem2[25][0] ),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\top1.memory2.mem2[8][2] ),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\top1.memory2.mem2[134][0] ),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\top1.memory1.mem1[81][1] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\top1.memory2.mem1[122][2] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\top1.memory2.mem2[18][2] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\top1.memory1.mem1[115][2] ),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\top1.memory1.mem1[70][2] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\top1.memory2.mem1[166][1] ),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\top1.memory2.mem1[107][1] ),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\top1.memory1.mem1[69][2] ),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\top1.memory2.mem1[124][1] ),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\top1.memory2.mem2[39][0] ),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\top1.memory2.mem1[30][1] ),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\top1.memory2.mem2[142][0] ),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\top1.memory2.mem2[140][0] ),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\top1.memory2.mem2[23][0] ),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\top1.memory1.mem1[55][1] ),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\top1.memory2.mem2[75][1] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\top1.memory1.mem2[33][2] ),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\top1.memory2.mem1[54][1] ),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\top1.memory1.mem2[123][2] ),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\top1.memory1.mem2[27][1] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\top1.memory1.mem1[81][0] ),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\top1.memory2.mem1[174][2] ),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\top1.memory1.mem2[1][2] ),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\top1.memory2.mem1[125][0] ),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\top1.memory2.mem2[33][0] ),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\top1.memory2.mem2[119][2] ),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\top1.memory2.mem1[194][1] ),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\top1.memory2.mem1[189][2] ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\top1.memory1.mem2[26][2] ),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\top1.memory2.mem1[184][1] ),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\top1.memory2.mem1[117][2] ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\top1.memory1.mem1[3][2] ),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\top1.memory1.mem2[49][1] ),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\top1.memory2.mem2[105][2] ),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\top1.memory2.mem1[3][0] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\top1.memory2.mem1[93][0] ),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\top1.memory2.mem1[21][0] ),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\top1.memory2.mem2[150][1] ),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\top1.memory1.mem1[198][2] ),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\top1.memory2.mem1[113][1] ),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\top1.memory2.mem1[88][2] ),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\top1.memory2.mem2[114][1] ),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\top1.memory1.mem1[53][1] ),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\top1.memory1.mem2[129][1] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\top1.memory2.mem2[10][2] ),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\top1.memory1.mem2[12][1] ),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\top1.memory2.mem2[167][2] ),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\top1.memory2.mem1[131][2] ),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\top1.memory1.mem2[19][2] ),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\top1.memory1.mem1[51][0] ),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\top1.memory2.mem1[173][2] ),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\top1.memory1.mem1[140][0] ),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\top1.memory1.mem2[68][1] ),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\top1.memory2.mem2[133][1] ),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\top1.memory1.mem1[54][0] ),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\top1.memory2.mem1[87][1] ),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\top1.memory2.mem1[123][0] ),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\top1.memory2.mem2[118][0] ),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\top1.memory2.mem1[189][0] ),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\top1.memory2.mem1[126][2] ),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\top1.memory1.mem1[37][1] ),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\top1.memory2.mem2[115][1] ),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\top1.memory2.mem2[46][0] ),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\top1.memory1.mem1[131][0] ),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\top1.memory1.mem2[83][1] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\top1.memory2.mem1[5][0] ),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\top1.memory2.mem1[51][1] ),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\top1.memory2.mem1[137][2] ),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\top1.memory1.mem1[65][2] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\top1.memory1.mem2[104][1] ),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\top1.memory2.mem2[123][0] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\top1.memory2.mem1[157][1] ),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\top1.memory2.mem2[106][1] ),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\top1.memory2.mem2[6][0] ),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\top1.memory1.mem2[48][1] ),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\top1.memory2.mem2[153][1] ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\top1.memory2.mem2[26][0] ),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\top1.memory2.mem1[121][0] ),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\top1.memory1.mem1[135][1] ),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\top1.memory2.mem1[105][2] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\top1.memory1.mem1[84][1] ),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\top1.memory2.mem1[23][2] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\top1.memory1.mem1[97][0] ),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\top1.memory2.mem2[83][1] ),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\top1.memory1.mem1[65][0] ),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\top1.memory2.mem1[173][0] ),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\top1.memory1.mem2[9][2] ),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\top1.memory1.mem1[61][1] ),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\top1.memory1.mem2[135][2] ),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\top1.memory1.mem1[169][2] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\top1.memory1.mem2[18][2] ),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\top1.memory2.mem2[128][1] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\top1.memory1.mem2[75][2] ),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\top1.memory1.mem2[15][1] ),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\top1.memory2.mem1[186][2] ),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\top1.memory1.mem1[4][1] ),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\top1.memory1.mem2[40][1] ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\top1.memory2.mem2[0][0] ),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\top1.memory1.mem2[152][2] ),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\top1.memory1.mem2[153][0] ),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold1599 (.A(\top1.memory2.mem2[12][1] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\top1.memory1.mem2[131][0] ),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\top1.memory2.mem1[160][1] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\top1.memory2.mem1[132][1] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\top1.memory1.mem2[119][0] ),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\top1.memory1.mem2[21][2] ),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\top1.memory1.mem1[153][2] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\top1.memory2.mem2[54][0] ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\top1.memory2.mem1[186][1] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\top1.memory1.mem1[102][0] ),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\top1.memory1.mem2[126][1] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\top1.memory1.mem2[90][0] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold1611 (.A(\top1.memory2.mem2[133][0] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\top1.memory1.mem2[37][1] ),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\top1.memory2.mem2[132][2] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\top1.memory1.mem2[189][1] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\top1.memory2.mem1[68][1] ),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\top1.memory1.mem2[51][0] ),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\top1.memory2.mem1[166][0] ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\top1.memory2.mem1[183][1] ),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\top1.memory2.mem1[167][1] ),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\top1.memory1.mem1[187][2] ),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\top1.memory1.mem2[79][1] ),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\top1.memory2.mem1[80][2] ),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\top1.memory1.mem1[72][0] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\top1.memory2.mem2[103][1] ),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\top1.memory1.mem2[142][2] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\top1.memory1.mem1[160][1] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\top1.memory1.mem1[70][0] ),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\top1.memory1.mem1[53][0] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\top1.memory2.mem1[184][0] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\top1.memory2.mem1[178][1] ),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\top1.memory1.mem2[112][2] ),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\top1.memory1.mem1[43][0] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\top1.memory2.mem2[90][2] ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\top1.memory2.mem1[97][2] ),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\top1.memory1.mem1[127][2] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\top1.memory1.mem1[174][2] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\top1.memory1.mem1[159][2] ),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\top1.memory1.mem2[11][0] ),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\top1.memory1.mem1[171][2] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\top1.memory2.mem1[190][2] ),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\top1.memory2.mem2[162][1] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\top1.memory1.mem1[143][1] ),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\top1.memory2.mem2[139][1] ),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\top1.memory2.mem2[52][0] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\top1.memory2.mem1[24][1] ),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\top1.memory2.mem2[1][0] ),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\top1.memory1.mem1[143][2] ),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\top1.memory1.mem1[133][0] ),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\top1.memory2.mem2[5][0] ),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\top1.memory2.mem2[33][1] ),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\top1.memory2.mem2[9][1] ),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\top1.memory1.mem2[64][0] ),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\top1.memory2.mem2[20][0] ),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\top1.memory1.mem2[133][2] ),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\top1.memory1.mem1[29][1] ),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\top1.memory1.mem2[130][0] ),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\top1.memory1.mem2[49][0] ),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\top1.memory2.mem1[62][0] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\top1.memory2.mem2[119][0] ),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\top1.memory2.mem1[144][2] ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\top1.memory2.mem2[170][0] ),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\top1.memory1.mem1[73][2] ),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\top1.memory1.mem2[107][2] ),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\top1.memory1.mem2[52][2] ),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\top1.memory1.mem1[96][2] ),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\top1.memory1.mem2[114][1] ),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\top1.memory1.mem1[42][0] ),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\top1.memory2.mem2[77][1] ),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\top1.memory1.mem2[98][2] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\top1.memory2.mem2[38][0] ),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\top1.memory1.mem1[188][1] ),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\top1.memory2.mem1[2][0] ),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\top1.memory1.mem1[195][1] ),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\top1.memory2.mem1[141][0] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\top1.memory1.mem2[135][1] ),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\top1.memory1.mem2[162][2] ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\top1.memory1.mem2[148][1] ),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\top1.memory1.mem1[75][0] ),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\top1.memory1.mem2[128][0] ),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\top1.memory2.mem2[69][0] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\top1.memory1.mem1[42][2] ),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\top1.memory1.mem2[161][2] ),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\top1.memory2.mem1[9][2] ),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\top1.memory1.mem1[140][2] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\top1.memory2.mem1[167][0] ),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\top1.memory2.mem2[65][0] ),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\top1.memory2.mem2[133][2] ),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\top1.memory1.mem2[43][1] ),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\top1.memory1.mem2[134][1] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\top1.memory1.mem1[46][0] ),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\top1.memory2.mem1[102][2] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\top1.memory2.mem1[83][1] ),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\top1.memory2.mem1[141][2] ),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\top1.memory2.mem1[193][2] ),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\top1.memory2.mem2[2][0] ),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\top1.memory1.mem1[181][1] ),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\top1.memory2.mem1[135][2] ),
    .X(net4135));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\top1.memory1.mem1[24][1] ),
    .X(net4136));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\top1.memory1.mem2[37][0] ),
    .X(net4137));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\top1.memory2.mem2[135][1] ),
    .X(net4138));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\top1.memory2.mem2[139][0] ),
    .X(net4139));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\top1.memory2.mem1[156][1] ),
    .X(net4140));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\top1.memory1.mem1[7][2] ),
    .X(net4141));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\top1.memory2.mem2[135][2] ),
    .X(net4142));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\top1.memory1.mem2[69][1] ),
    .X(net4143));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\top1.memory1.mem2[153][2] ),
    .X(net4144));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\top1.memory2.mem1[140][2] ),
    .X(net4145));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\top1.memory1.mem2[141][1] ),
    .X(net4146));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\top1.memory1.mem1[5][2] ),
    .X(net4147));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\top1.memory1.mem1[43][1] ),
    .X(net4148));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\top1.memory2.mem2[139][2] ),
    .X(net4149));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\top1.memory2.mem1[154][2] ),
    .X(net4150));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\top1.memory2.mem1[174][1] ),
    .X(net4151));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\top1.memory2.mem1[12][2] ),
    .X(net4152));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\top1.memory2.mem1[109][2] ),
    .X(net4153));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\top1.memory2.mem1[98][2] ),
    .X(net4154));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\top1.memory1.mem1[72][1] ),
    .X(net4155));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\top1.memory1.mem2[2][2] ),
    .X(net4156));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\top1.memory1.mem2[3][1] ),
    .X(net4157));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\top1.memory2.mem1[100][0] ),
    .X(net4158));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\top1.memory1.mem1[172][0] ),
    .X(net4159));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\top1.memory1.mem2[151][1] ),
    .X(net4160));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\top1.memory2.mem1[63][0] ),
    .X(net4161));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\top1.memory2.mem2[4][0] ),
    .X(net4162));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\top1.memory1.mem2[74][0] ),
    .X(net4163));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\top1.memory2.mem2[9][2] ),
    .X(net4164));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\top1.memory2.mem2[100][1] ),
    .X(net4165));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\top1.memory2.mem1[137][1] ),
    .X(net4166));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\top1.memory1.mem2[70][2] ),
    .X(net4167));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\top1.memory2.mem2[0][2] ),
    .X(net4168));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\top1.memory1.mem1[132][1] ),
    .X(net4169));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\top1.memory2.mem2[53][1] ),
    .X(net4170));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\top1.memory2.mem2[142][1] ),
    .X(net4171));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\top1.memory1.mem2[175][0] ),
    .X(net4172));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\top1.memory2.mem2[81][1] ),
    .X(net4173));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\top1.memory2.mem1[67][2] ),
    .X(net4174));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\top1.memory1.mem1[0][0] ),
    .X(net4175));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\top1.memory2.mem2[160][2] ),
    .X(net4176));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\top1.memory2.mem2[8][0] ),
    .X(net4177));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\top1.memory1.mem2[70][0] ),
    .X(net4178));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\top1.memory1.mem2[115][2] ),
    .X(net4179));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\top1.memory2.mem1[127][2] ),
    .X(net4180));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\top1.memory2.mem1[142][1] ),
    .X(net4181));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\top1.memory1.mem2[59][0] ),
    .X(net4182));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\top1.memory1.mem1[68][2] ),
    .X(net4183));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\top1.memory2.mem2[60][2] ),
    .X(net4184));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\top1.memory1.mem2[35][2] ),
    .X(net4185));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\top1.memory1.mem1[22][0] ),
    .X(net4186));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\top1.memory1.mem1[67][0] ),
    .X(net4187));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\top1.memory2.mem2[198][1] ),
    .X(net4188));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\top1.memory1.mem2[4][2] ),
    .X(net4189));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\top1.memory2.mem2[144][0] ),
    .X(net4190));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\top1.memory2.mem1[160][2] ),
    .X(net4191));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\top1.memory1.mem2[129][0] ),
    .X(net4192));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\top1.memory1.mem1[161][1] ),
    .X(net4193));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\top1.memory2.mem1[12][0] ),
    .X(net4194));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\top1.memory1.mem2[125][0] ),
    .X(net4195));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\top1.memory2.mem1[133][2] ),
    .X(net4196));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\top1.memory2.mem1[136][1] ),
    .X(net4197));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\top1.memory1.mem1[139][1] ),
    .X(net4198));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\top1.memory1.mem1[63][1] ),
    .X(net4199));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\top1.memory1.mem1[6][2] ),
    .X(net4200));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\top1.memory1.mem1[100][0] ),
    .X(net4201));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\top1.memory2.mem2[170][2] ),
    .X(net4202));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\top1.memory1.mem2[161][0] ),
    .X(net4203));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\top1.memory1.mem2[68][2] ),
    .X(net4204));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\top1.memory2.mem2[143][1] ),
    .X(net4205));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\top1.memory2.mem2[14][0] ),
    .X(net4206));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\top1.memory1.mem1[15][1] ),
    .X(net4207));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\top1.memory2.mem2[69][1] ),
    .X(net4208));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\top1.memory1.mem1[170][2] ),
    .X(net4209));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\top1.memory2.mem1[132][2] ),
    .X(net4210));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\top1.memory1.mem1[163][1] ),
    .X(net4211));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\top1.memory2.mem1[15][2] ),
    .X(net4212));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\top1.memory1.mem1[69][1] ),
    .X(net4213));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\top1.memory1.mem1[129][2] ),
    .X(net4214));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\top1.memory1.mem1[160][0] ),
    .X(net4215));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\top1.memory2.mem1[96][2] ),
    .X(net4216));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\top1.memory1.mem1[79][1] ),
    .X(net4217));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\top1.memory2.mem2[72][2] ),
    .X(net4218));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\top1.memory2.mem1[64][0] ),
    .X(net4219));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\top1.memory1.mem1[96][0] ),
    .X(net4220));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\top1.memory1.mem1[26][2] ),
    .X(net4221));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\top1.memory2.mem2[146][2] ),
    .X(net4222));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\top1.memory2.mem1[5][1] ),
    .X(net4223));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\top1.memory1.mem1[197][1] ),
    .X(net4224));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\top1.memory2.mem2[66][0] ),
    .X(net4225));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\top1.memory1.mem1[160][2] ),
    .X(net4226));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\top1.memory2.mem1[85][2] ),
    .X(net4227));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\top1.memory2.mem2[7][1] ),
    .X(net4228));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\top1.memory2.mem2[88][2] ),
    .X(net4229));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\top1.memory2.mem2[10][0] ),
    .X(net4230));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\top1.memory2.mem2[28][1] ),
    .X(net4231));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\top1.memory2.mem1[13][1] ),
    .X(net4232));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\top1.memory2.mem1[100][2] ),
    .X(net4233));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\top1.memory1.mem2[111][2] ),
    .X(net4234));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\top1.memory2.mem2[137][1] ),
    .X(net4235));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\top1.memory1.mem1[127][0] ),
    .X(net4236));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\top1.memory1.mem1[0][1] ),
    .X(net4237));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\top1.memory1.mem2[143][0] ),
    .X(net4238));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\top1.memory2.mem1[43][0] ),
    .X(net4239));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\top1.memory2.mem1[131][0] ),
    .X(net4240));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\top1.memory1.mem1[171][0] ),
    .X(net4241));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\top1.memory1.mem2[9][0] ),
    .X(net4242));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\top1.memory2.mem2[126][0] ),
    .X(net4243));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\top1.memory1.mem2[99][2] ),
    .X(net4244));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\top1.memory1.mem1[77][1] ),
    .X(net4245));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\top1.memory1.mem1[73][0] ),
    .X(net4246));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\top1.memory2.mem2[122][0] ),
    .X(net4247));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\top1.memory2.mem2[110][1] ),
    .X(net4248));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\top1.memory1.mem2[138][1] ),
    .X(net4249));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\top1.memory1.mem1[73][1] ),
    .X(net4250));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\top1.memory1.mem1[182][1] ),
    .X(net4251));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\top1.memory1.mem1[197][0] ),
    .X(net4252));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\top1.memory1.mem1[2][2] ),
    .X(net4253));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\top1.memory2.mem1[8][2] ),
    .X(net4254));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\top1.memory2.mem2[6][1] ),
    .X(net4255));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\top1.memory1.mem1[135][0] ),
    .X(net4256));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\top1.memory2.mem2[53][0] ),
    .X(net4257));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\top1.memory2.mem1[179][1] ),
    .X(net4258));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\top1.memory2.mem1[12][1] ),
    .X(net4259));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\top1.memory2.mem2[141][1] ),
    .X(net4260));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\top1.memory1.mem1[65][1] ),
    .X(net4261));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\top1.memory1.mem1[56][1] ),
    .X(net4262));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\top1.memory2.mem2[5][1] ),
    .X(net4263));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\top1.memory1.mem1[98][2] ),
    .X(net4264));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\top1.memory2.mem2[99][1] ),
    .X(net4265));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\top1.memory2.mem2[78][2] ),
    .X(net4266));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\top1.memory1.mem1[102][2] ),
    .X(net4267));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\top1.memory2.mem2[109][2] ),
    .X(net4268));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\top1.memory1.mem2[59][1] ),
    .X(net4269));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\top1.memory1.mem1[78][2] ),
    .X(net4270));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\top1.memory1.mem1[27][2] ),
    .X(net4271));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\top1.memory1.mem1[141][0] ),
    .X(net4272));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\top1.memory1.mem1[133][1] ),
    .X(net4273));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\top1.memory2.mem1[128][1] ),
    .X(net4274));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\top1.memory1.mem1[199][1] ),
    .X(net4275));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\top1.memory1.mem2[22][2] ),
    .X(net4276));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\top1.memory1.mem2[128][2] ),
    .X(net4277));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\top1.memory2.mem1[9][0] ),
    .X(net4278));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\top1.memory2.mem2[131][2] ),
    .X(net4279));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\top1.memory1.mem1[98][0] ),
    .X(net4280));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\top1.memory2.mem1[164][1] ),
    .X(net4281));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\top1.memory2.mem1[199][2] ),
    .X(net4282));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\top1.memory1.mem1[99][1] ),
    .X(net4283));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\top1.memory1.mem1[76][1] ),
    .X(net4284));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\top1.memory1.mem2[80][0] ),
    .X(net4285));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\top1.memory1.mem2[138][0] ),
    .X(net4286));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\top1.memory1.mem2[152][0] ),
    .X(net4287));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\top1.memory1.mem1[135][2] ),
    .X(net4288));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\top1.memory1.mem1[128][1] ),
    .X(net4289));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\top1.memory2.mem2[35][1] ),
    .X(net4290));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\top1.memory2.mem1[183][2] ),
    .X(net4291));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\top1.memory1.mem1[118][1] ),
    .X(net4292));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\top1.memory1.mem1[162][0] ),
    .X(net4293));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\top1.memory2.mem2[27][1] ),
    .X(net4294));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\top1.memory2.mem2[131][0] ),
    .X(net4295));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\top1.memory2.mem2[135][0] ),
    .X(net4296));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\top1.memory1.mem1[123][2] ),
    .X(net4297));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\top1.memory1.mem1[1][2] ),
    .X(net4298));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\top1.memory2.mem1[39][1] ),
    .X(net4299));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\top1.memory2.mem1[17][2] ),
    .X(net4300));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\top1.memory2.mem1[139][1] ),
    .X(net4301));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\top1.memory1.mem2[58][1] ),
    .X(net4302));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\top1.fsm.idx_final[7] ),
    .X(net4303));
 sg13g2_dlygate4sd3_1 hold1866 (.A(_01318_),
    .X(net4304));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\top1.memory1.mem2[145][2] ),
    .X(net4305));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\top1.memory1.mem1[112][2] ),
    .X(net4306));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\top1.memory1.mem2[161][1] ),
    .X(net4307));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\top1.memory1.mem1[41][0] ),
    .X(net4308));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\top1.memory1.mem1[50][2] ),
    .X(net4309));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\top1.memory2.mem2[99][2] ),
    .X(net4310));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\top1.memory1.mem2[144][1] ),
    .X(net4311));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\top1.memory2.mem1[100][1] ),
    .X(net4312));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\top1.memory2.mem1[84][1] ),
    .X(net4313));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\top1.memory1.mem2[76][0] ),
    .X(net4314));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\top1.memory1.mem1[5][0] ),
    .X(net4315));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\top1.memory2.mem2[2][1] ),
    .X(net4316));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\top1.memory2.mem2[24][2] ),
    .X(net4317));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\top1.memory1.mem1[177][2] ),
    .X(net4318));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\top1.memory2.mem2[72][1] ),
    .X(net4319));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\top1.memory1.mem1[134][0] ),
    .X(net4320));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\top1.memory1.mem1[80][2] ),
    .X(net4321));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\top1.memory1.mem2[125][1] ),
    .X(net4322));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\top1.memory2.mem1[25][2] ),
    .X(net4323));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\top1.memory1.mem1[74][2] ),
    .X(net4324));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\top1.memory1.mem2[88][2] ),
    .X(net4325));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\top1.memory2.mem1[114][1] ),
    .X(net4326));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\top1.memory1.mem2[100][2] ),
    .X(net4327));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\top1.memory1.mem2[144][2] ),
    .X(net4328));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\top1.memory1.mem2[160][1] ),
    .X(net4329));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\top1.memory2.mem2[3][0] ),
    .X(net4330));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\top1.memory2.mem1[78][2] ),
    .X(net4331));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\top1.memory1.mem2[192][2] ),
    .X(net4332));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\top1.memory2.mem2[129][0] ),
    .X(net4333));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\top1.memory2.mem1[191][2] ),
    .X(net4334));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\top1.memory2.mem1[66][2] ),
    .X(net4335));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\top1.memory2.mem2[8][1] ),
    .X(net4336));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\top1.memory2.mem1[82][2] ),
    .X(net4337));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\top1.memory1.mem1[189][1] ),
    .X(net4338));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\top1.memory2.mem1[4][1] ),
    .X(net4339));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\top1.memory1.mem1[119][1] ),
    .X(net4340));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\top1.memory1.mem2[66][1] ),
    .X(net4341));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\top1.memory1.mem2[72][1] ),
    .X(net4342));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\top1.memory2.mem1[81][0] ),
    .X(net4343));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\top1.memory2.mem2[97][1] ),
    .X(net4344));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\top1.memory2.mem1[184][2] ),
    .X(net4345));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\top1.memory1.mem2[134][2] ),
    .X(net4346));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\top1.memory2.mem1[166][2] ),
    .X(net4347));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\top1.memory1.mem1[2][0] ),
    .X(net4348));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\top1.memory1.mem1[109][0] ),
    .X(net4349));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\top1.memory1.mem2[88][0] ),
    .X(net4350));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\top1.memory2.mem1[103][1] ),
    .X(net4351));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\top1.memory2.mem2[97][0] ),
    .X(net4352));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\top1.memory2.mem1[134][0] ),
    .X(net4353));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\top1.memory1.mem1[156][0] ),
    .X(net4354));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\top1.memory1.mem2[199][1] ),
    .X(net4355));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\top1.memory1.mem2[99][0] ),
    .X(net4356));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\top1.memory1.mem1[131][1] ),
    .X(net4357));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\top1.memory1.mem1[137][2] ),
    .X(net4358));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\top1.memory2.mem1[99][2] ),
    .X(net4359));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\top1.memory2.mem1[55][2] ),
    .X(net4360));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\top1.memory1.mem1[2][1] ),
    .X(net4361));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\top1.memory1.mem2[97][0] ),
    .X(net4362));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\top1.memory1.mem2[5][1] ),
    .X(net4363));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\top1.memory1.mem2[98][0] ),
    .X(net4364));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\top1.memory2.mem2[68][0] ),
    .X(net4365));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\top1.memory2.mem2[156][0] ),
    .X(net4366));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\top1.memory1.mem1[140][1] ),
    .X(net4367));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\top1.memory2.mem1[43][2] ),
    .X(net4368));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\top1.memory2.mem1[65][2] ),
    .X(net4369));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\top1.memory2.mem2[58][0] ),
    .X(net4370));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\top1.memory2.mem2[134][2] ),
    .X(net4371));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\top1.memory1.mem2[145][1] ),
    .X(net4372));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\top1.memory2.mem2[125][1] ),
    .X(net4373));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\top1.memory1.mem1[15][0] ),
    .X(net4374));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\top1.memory2.mem1[82][1] ),
    .X(net4375));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\top1.memory2.mem2[100][0] ),
    .X(net4376));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\top1.memory1.mem2[75][1] ),
    .X(net4377));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\top1.memory1.mem2[80][1] ),
    .X(net4378));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\top1.memory2.mem2[101][0] ),
    .X(net4379));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\top1.memory1.mem1[66][0] ),
    .X(net4380));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\top1.memory2.mem1[81][1] ),
    .X(net4381));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\top1.memory1.mem1[161][0] ),
    .X(net4382));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\top1.memory1.mem2[67][1] ),
    .X(net4383));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\top1.memory2.mem2[46][1] ),
    .X(net4384));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\top1.memory1.mem2[140][2] ),
    .X(net4385));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\top1.memory1.mem1[76][2] ),
    .X(net4386));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\top1.memory2.mem1[75][2] ),
    .X(net4387));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\top1.memory2.mem2[9][0] ),
    .X(net4388));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\top1.memory1.mem2[50][0] ),
    .X(net4389));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\top1.memory1.mem2[73][2] ),
    .X(net4390));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\top1.memory1.mem1[144][0] ),
    .X(net4391));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\top1.memory2.mem1[69][0] ),
    .X(net4392));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\top1.memory1.mem2[139][1] ),
    .X(net4393));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\top1.memory1.mem1[132][0] ),
    .X(net4394));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\top1.memory1.mem2[82][1] ),
    .X(net4395));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\top1.memory1.mem1[154][2] ),
    .X(net4396));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\top1.memory2.mem1[140][1] ),
    .X(net4397));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\top1.memory1.mem1[79][0] ),
    .X(net4398));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\top1.memory2.mem1[101][1] ),
    .X(net4399));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\top1.memory2.mem2[162][2] ),
    .X(net4400));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\top1.memory2.mem2[83][2] ),
    .X(net4401));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\top1.memory2.mem2[199][0] ),
    .X(net4402));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\top1.memory1.mem1[190][1] ),
    .X(net4403));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\top1.memory1.mem2[66][0] ),
    .X(net4404));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\top1.memory2.mem1[96][0] ),
    .X(net4405));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\top1.memory1.mem2[72][2] ),
    .X(net4406));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\top1.memory2.mem1[69][2] ),
    .X(net4407));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\top1.memory2.mem1[68][2] ),
    .X(net4408));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\top1.memory1.mem1[83][1] ),
    .X(net4409));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\top1.memory1.mem2[129][2] ),
    .X(net4410));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\top1.memory2.mem1[138][2] ),
    .X(net4411));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\top1.memory2.mem2[138][0] ),
    .X(net4412));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\top1.memory2.mem1[133][0] ),
    .X(net4413));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\top1.memory1.mem1[145][0] ),
    .X(net4414));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\top1.memory2.mem1[74][0] ),
    .X(net4415));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\top1.memory2.mem1[67][0] ),
    .X(net4416));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\top1.memory1.mem2[70][1] ),
    .X(net4417));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\top1.memory2.mem2[118][1] ),
    .X(net4418));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\top1.memory2.mem2[50][1] ),
    .X(net4419));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\top1.memory2.mem1[77][2] ),
    .X(net4420));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\top1.memory1.mem2[10][1] ),
    .X(net4421));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\top1.memory1.mem2[65][2] ),
    .X(net4422));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\top1.memory2.mem2[5][2] ),
    .X(net4423));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\top1.memory1.mem1[9][0] ),
    .X(net4424));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\top1.memory1.mem2[29][0] ),
    .X(net4425));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\top1.memory2.mem1[127][0] ),
    .X(net4426));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\top1.memory1.mem1[146][2] ),
    .X(net4427));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\top1.memory2.mem2[104][1] ),
    .X(net4428));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\top1.memory2.mem1[129][0] ),
    .X(net4429));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\top1.memory2.mem1[110][2] ),
    .X(net4430));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\top1.memory1.mem1[68][0] ),
    .X(net4431));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\top1.memory1.mem1[20][2] ),
    .X(net4432));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\top1.memory2.mem2[6][2] ),
    .X(net4433));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\top1.memory1.mem2[74][2] ),
    .X(net4434));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\top1.memory2.mem1[135][0] ),
    .X(net4435));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\top1.memory2.mem2[184][2] ),
    .X(net4436));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\top1.memory2.mem2[132][1] ),
    .X(net4437));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\top1.memory1.mem1[139][0] ),
    .X(net4438));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\top1.memory2.mem1[6][1] ),
    .X(net4439));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\top1.memory1.mem1[85][0] ),
    .X(net4440));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\top1.memory1.mem2[73][0] ),
    .X(net4441));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\top1.memory1.mem2[136][2] ),
    .X(net4442));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\top1.memory2.mem1[0][0] ),
    .X(net4443));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\top1.memory2.mem1[76][2] ),
    .X(net4444));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\top1.memory2.mem1[139][2] ),
    .X(net4445));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\top1.memory1.mem1[8][0] ),
    .X(net4446));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\top1.memory1.mem1[67][1] ),
    .X(net4447));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\top1.memory2.mem1[162][1] ),
    .X(net4448));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\top1.memory2.mem1[97][0] ),
    .X(net4449));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\top1.memory2.mem1[78][1] ),
    .X(net4450));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\top1.memory1.mem2[145][0] ),
    .X(net4451));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\top1.memory2.mem1[162][0] ),
    .X(net4452));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\top1.memory2.mem2[137][2] ),
    .X(net4453));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\top1.memory2.mem2[83][0] ),
    .X(net4454));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\top1.memory2.mem2[3][1] ),
    .X(net4455));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\top1.memory1.mem2[137][2] ),
    .X(net4456));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\top1.memory2.mem1[1][2] ),
    .X(net4457));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\top1.memory1.mem2[0][1] ),
    .X(net4458));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\top1.memory2.mem2[144][2] ),
    .X(net4459));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\top1.memory2.mem2[99][0] ),
    .X(net4460));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\top1.memory2.mem2[93][0] ),
    .X(net4461));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\top1.memory1.mem1[191][1] ),
    .X(net4462));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\top1.memory2.mem1[134][2] ),
    .X(net4463));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\top1.memory2.mem2[104][0] ),
    .X(net4464));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\top1.memory2.mem2[145][0] ),
    .X(net4465));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\top1.memory1.mem2[2][1] ),
    .X(net4466));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\top1.memory1.mem2[127][2] ),
    .X(net4467));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\top1.memory2.mem2[96][0] ),
    .X(net4468));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\top1.memory1.mem2[134][0] ),
    .X(net4469));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\top1.memory1.mem2[54][2] ),
    .X(net4470));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\top1.memory2.mem1[81][2] ),
    .X(net4471));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\top1.memory2.mem1[143][0] ),
    .X(net4472));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\top1.memory1.mem2[15][2] ),
    .X(net4473));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\top1.memory2.mem1[145][0] ),
    .X(net4474));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\top1.memory2.mem1[83][2] ),
    .X(net4475));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\top1.memory1.mem2[139][2] ),
    .X(net4476));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\top1.memory1.mem1[66][1] ),
    .X(net4477));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\top1.memory2.mem1[138][1] ),
    .X(net4478));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\top1.memory2.mem1[130][1] ),
    .X(net4479));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\top1.memory1.mem2[132][1] ),
    .X(net4480));
 sg13g2_dlygate4sd3_1 hold2043 (.A(\top1.memory2.mem2[72][0] ),
    .X(net4481));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\top1.fsm.idx_final[0] ),
    .X(net4482));
 sg13g2_dlygate4sd3_1 hold2045 (.A(_01311_),
    .X(net4483));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\top1.memory1.mem2[137][0] ),
    .X(net4484));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\top1.memory2.mem1[98][1] ),
    .X(net4485));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\top1.memory1.mem2[143][1] ),
    .X(net4486));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\top1.memory2.mem2[88][1] ),
    .X(net4487));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\top1.memory1.mem2[100][1] ),
    .X(net4488));
 sg13g2_dlygate4sd3_1 hold2051 (.A(\top1.memory2.mem1[59][0] ),
    .X(net4489));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\top1.memory2.mem1[97][1] ),
    .X(net4490));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\top1.memory2.mem1[145][2] ),
    .X(net4491));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\top1.memory1.mem2[189][2] ),
    .X(net4492));
 sg13g2_dlygate4sd3_1 hold2055 (.A(\top1.memory2.mem1[73][2] ),
    .X(net4493));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\top1.memory1.mem2[24][2] ),
    .X(net4494));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\top1.memory1.mem2[83][2] ),
    .X(net4495));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\top1.memory1.mem1[36][1] ),
    .X(net4496));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\top1.memory1.mem1[83][2] ),
    .X(net4497));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\top1.memory2.mem1[161][2] ),
    .X(net4498));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\top1.memory2.mem2[193][1] ),
    .X(net4499));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\top1.memory1.mem1[64][1] ),
    .X(net4500));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\top1.memory1.mem1[75][2] ),
    .X(net4501));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\top1.memory2.mem1[161][1] ),
    .X(net4502));
 sg13g2_dlygate4sd3_1 hold2065 (.A(\top1.memory2.mem1[65][1] ),
    .X(net4503));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\top1.memory1.mem1[143][0] ),
    .X(net4504));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\top1.memory2.mem1[143][1] ),
    .X(net4505));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\top1.memory2.mem1[0][2] ),
    .X(net4506));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\top1.memory1.mem1[141][2] ),
    .X(net4507));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\top1.memory2.mem1[51][2] ),
    .X(net4508));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\top1.memory2.mem1[70][2] ),
    .X(net4509));
 sg13g2_dlygate4sd3_1 hold2072 (.A(\top1.memory2.mem2[67][1] ),
    .X(net4510));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\top1.memory1.mem2[100][0] ),
    .X(net4511));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\top1.memory1.mem2[67][2] ),
    .X(net4512));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\top1.memory2.mem2[79][1] ),
    .X(net4513));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\top1.memory1.mem2[96][1] ),
    .X(net4514));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\top1.memory1.mem2[29][1] ),
    .X(net4515));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\top1.memory2.mem1[67][1] ),
    .X(net4516));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\top1.memory2.mem1[8][0] ),
    .X(net4517));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\top1.memory1.mem1[82][2] ),
    .X(net4518));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\top1.memory1.mem2[142][1] ),
    .X(net4519));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\top1.memory1.mem2[9][1] ),
    .X(net4520));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\top1.memory1.mem2[4][1] ),
    .X(net4521));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\top1.memory1.mem2[8][2] ),
    .X(net4522));
 sg13g2_dlygate4sd3_1 hold2085 (.A(\top1.memory1.mem2[4][0] ),
    .X(net4523));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\top1.memory2.mem2[141][2] ),
    .X(net4524));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\top1.memory2.mem2[80][0] ),
    .X(net4525));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\top1.memory1.mem1[136][2] ),
    .X(net4526));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\top1.memory2.mem1[79][2] ),
    .X(net4527));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\top1.memory2.mem2[84][1] ),
    .X(net4528));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\top1.memory2.mem2[81][0] ),
    .X(net4529));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\top1.memory1.mem1[84][0] ),
    .X(net4530));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\top1.memory1.mem1[162][2] ),
    .X(net4531));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\top1.memory2.mem2[97][2] ),
    .X(net4532));
 sg13g2_dlygate4sd3_1 hold2095 (.A(\top1.memory1.mem2[97][2] ),
    .X(net4533));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\top1.memory1.mem2[84][1] ),
    .X(net4534));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\top1.memory2.mem1[72][1] ),
    .X(net4535));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\top1.memory1.mem1[146][1] ),
    .X(net4536));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\top1.memory1.mem1[138][0] ),
    .X(net4537));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\top1.memory2.mem2[130][0] ),
    .X(net4538));
 sg13g2_dlygate4sd3_1 hold2101 (.A(\top1.memory1.mem1[127][1] ),
    .X(net4539));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\top1.memory2.mem1[69][1] ),
    .X(net4540));
 sg13g2_dlygate4sd3_1 hold2103 (.A(\top1.memory2.mem1[129][2] ),
    .X(net4541));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\top1.memory1.mem1[132][2] ),
    .X(net4542));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\top1.memory2.mem1[70][1] ),
    .X(net4543));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\top1.memory2.mem1[82][0] ),
    .X(net4544));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\top1.memory2.mem2[59][2] ),
    .X(net4545));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\top1.memory1.mem1[161][2] ),
    .X(net4546));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\top1.memory2.mem1[73][1] ),
    .X(net4547));
 sg13g2_dlygate4sd3_1 hold2110 (.A(\top1.memory1.mem1[130][2] ),
    .X(net4548));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\top1.memory1.mem1[1][1] ),
    .X(net4549));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\top1.memory1.mem2[76][2] ),
    .X(net4550));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\top1.memory1.mem2[127][0] ),
    .X(net4551));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\top1.memory1.mem1[99][0] ),
    .X(net4552));
 sg13g2_dlygate4sd3_1 hold2115 (.A(\top1.memory2.mem1[83][0] ),
    .X(net4553));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\top1.memory1.mem2[135][0] ),
    .X(net4554));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\top1.memory2.mem2[143][0] ),
    .X(net4555));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\top1.memory1.mem2[146][2] ),
    .X(net4556));
 sg13g2_dlygate4sd3_1 hold2119 (.A(\top1.memory2.mem1[68][0] ),
    .X(net4557));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\top1.memory1.mem1[5][1] ),
    .X(net4558));
 sg13g2_dlygate4sd3_1 hold2121 (.A(\top1.memory1.mem2[130][2] ),
    .X(net4559));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\top1.memory1.mem2[132][2] ),
    .X(net4560));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\top1.memory2.mem2[132][0] ),
    .X(net4561));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\top1.memory2.mem1[131][1] ),
    .X(net4562));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\top1.memory1.mem1[84][2] ),
    .X(net4563));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\top1.memory2.mem1[142][0] ),
    .X(net4564));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\top1.memory1.mem2[41][1] ),
    .X(net4565));
 sg13g2_dlygate4sd3_1 hold2128 (.A(\top1.memory2.mem1[88][1] ),
    .X(net4566));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\top1.memory2.mem1[137][0] ),
    .X(net4567));
 sg13g2_dlygate4sd3_1 hold2130 (.A(\top1.memory2.mem2[12][2] ),
    .X(net4568));
 sg13g2_dlygate4sd3_1 hold2131 (.A(\top1.memory2.mem2[146][0] ),
    .X(net4569));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\top1.memory1.mem1[130][1] ),
    .X(net4570));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\top1.memory2.mem1[74][2] ),
    .X(net4571));
 sg13g2_dlygate4sd3_1 hold2134 (.A(\top1.memory1.mem2[1][0] ),
    .X(net4572));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\top1.memory1.mem1[88][2] ),
    .X(net4573));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\top1.memory1.mem1[104][2] ),
    .X(net4574));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\top1.memory2.mem1[146][0] ),
    .X(net4575));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\top1.memory2.mem1[2][2] ),
    .X(net4576));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\top1.memory1.mem2[131][1] ),
    .X(net4577));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\top1.memory2.mem2[73][2] ),
    .X(net4578));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\top1.memory2.mem2[123][2] ),
    .X(net4579));
 sg13g2_dlygate4sd3_1 hold2142 (.A(\top1.memory2.mem1[122][1] ),
    .X(net4580));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\top1.memory2.mem1[135][1] ),
    .X(net4581));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\top1.memory1.mem2[130][1] ),
    .X(net4582));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\top1.memory2.mem2[138][2] ),
    .X(net4583));
 sg13g2_dlygate4sd3_1 hold2146 (.A(\top1.memory2.mem1[77][0] ),
    .X(net4584));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\top1.fsm.idx_final[1] ),
    .X(net4585));
 sg13g2_dlygate4sd3_1 hold2148 (.A(_01312_),
    .X(net4586));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\top1.memory1.mem1[97][1] ),
    .X(net4587));
 sg13g2_dlygate4sd3_1 hold2150 (.A(\top1.memory1.mem1[70][1] ),
    .X(net4588));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\top1.fsm.idx_final[3] ),
    .X(net4589));
 sg13g2_dlygate4sd3_1 hold2152 (.A(_01314_),
    .X(net4590));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\top1.memory1.mem2[81][2] ),
    .X(net4591));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\top1.memory1.mem1[10][1] ),
    .X(net4592));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\top1.memory1.mem1[83][0] ),
    .X(net4593));
 sg13g2_dlygate4sd3_1 hold2156 (.A(\top1.memory1.mem1[74][0] ),
    .X(net4594));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\top1.memory1.mem2[3][0] ),
    .X(net4595));
 sg13g2_dlygate4sd3_1 hold2158 (.A(\top1.memory2.mem2[127][2] ),
    .X(net4596));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\top1.memory2.mem1[146][2] ),
    .X(net4597));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\top1.memory1.mem2[160][2] ),
    .X(net4598));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\top1.memory2.mem1[5][2] ),
    .X(net4599));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\top1.memory1.mem1[8][2] ),
    .X(net4600));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\top1.memory1.mem2[104][2] ),
    .X(net4601));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\top1.memory2.mem1[4][2] ),
    .X(net4602));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\top1.memory2.mem2[105][0] ),
    .X(net4603));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\top1.memory1.mem2[5][2] ),
    .X(net4604));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\top1.memory2.mem1[65][0] ),
    .X(net4605));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\top1.memory1.mem2[142][0] ),
    .X(net4606));
 sg13g2_dlygate4sd3_1 hold2169 (.A(\top1.memory1.mem2[5][0] ),
    .X(net4607));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\top1.memory1.mem2[23][0] ),
    .X(net4608));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\top1.memory1.mem1[145][2] ),
    .X(net4609));
 sg13g2_dlygate4sd3_1 hold2172 (.A(\top1.memory1.mem2[81][1] ),
    .X(net4610));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\top1.memory2.mem2[199][1] ),
    .X(net4611));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\top1.memory2.mem2[74][0] ),
    .X(net4612));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\top1.memory2.mem2[161][0] ),
    .X(net4613));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\top1.memory2.mem2[130][2] ),
    .X(net4614));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\top1.memory1.mem1[130][0] ),
    .X(net4615));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\top1.memory1.mem2[137][1] ),
    .X(net4616));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\top1.memory1.mem2[6][0] ),
    .X(net4617));
 sg13g2_dlygate4sd3_1 hold2180 (.A(\top1.memory1.mem2[84][2] ),
    .X(net4618));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\top1.memory1.mem1[75][1] ),
    .X(net4619));
 sg13g2_dlygate4sd3_1 hold2182 (.A(\top1.memory2.mem1[142][2] ),
    .X(net4620));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\top1.memory1.mem2[199][0] ),
    .X(net4621));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\top1.memory2.mem2[70][1] ),
    .X(net4622));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\top1.memory2.mem1[1][1] ),
    .X(net4623));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\top1.memory2.mem1[84][0] ),
    .X(net4624));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\top1.mem_ctl.state_reg[0] ),
    .X(net4625));
 sg13g2_dlygate4sd3_1 hold2188 (.A(_07202_),
    .X(net4626));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\top1.memory1.mem1[100][2] ),
    .X(net4627));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\top1.memory2.mem2[173][0] ),
    .X(net4628));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\top1.memory2.mem2[64][1] ),
    .X(net4629));
 sg13g2_dlygate4sd3_1 hold2192 (.A(\top1.memory1.mem1[74][1] ),
    .X(net4630));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\top1.memory2.mem2[15][0] ),
    .X(net4631));
 sg13g2_dlygate4sd3_1 hold2194 (.A(\top1.memory1.mem1[142][1] ),
    .X(net4632));
 sg13g2_dlygate4sd3_1 hold2195 (.A(\top1.memory1.mem1[199][2] ),
    .X(net4633));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\top1.memory2.mem2[160][1] ),
    .X(net4634));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\top1.memory2.mem1[79][1] ),
    .X(net4635));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\top1.memory2.mem1[88][0] ),
    .X(net4636));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\top1.memory1.mem2[78][0] ),
    .X(net4637));
 sg13g2_dlygate4sd3_1 hold2200 (.A(\top1.memory1.mem2[127][1] ),
    .X(net4638));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\top1.memory2.mem2[88][0] ),
    .X(net4639));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\top1.memory1.mem2[110][1] ),
    .X(net4640));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\top1.memory1.mem1[104][0] ),
    .X(net4641));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\top1.memory1.mem2[12][2] ),
    .X(net4642));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\top1.memory2.mem2[66][2] ),
    .X(net4643));
 sg13g2_dlygate4sd3_1 hold2206 (.A(\top1.memory2.mem2[65][2] ),
    .X(net4644));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\top1.memory2.mem2[69][2] ),
    .X(net4645));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\top1.memory1.mem2[144][0] ),
    .X(net4646));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\top1.memory2.mem1[146][1] ),
    .X(net4647));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\top1.memory1.mem2[138][2] ),
    .X(net4648));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\top1.memory1.mem1[6][1] ),
    .X(net4649));
 sg13g2_dlygate4sd3_1 hold2212 (.A(\top1.memory2.mem1[74][1] ),
    .X(net4650));
 sg13g2_dlygate4sd3_1 hold2213 (.A(\top1.memory1.mem1[186][2] ),
    .X(net4651));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\top1.memory2.mem1[132][0] ),
    .X(net4652));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\top1.memory2.mem2[70][0] ),
    .X(net4653));
 sg13g2_dlygate4sd3_1 hold2216 (.A(\top1.memory1.mem2[72][0] ),
    .X(net4654));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\top1.memory2.mem1[77][1] ),
    .X(net4655));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\top1.memory2.mem2[76][2] ),
    .X(net4656));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\top1.memory2.mem1[199][0] ),
    .X(net4657));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\top1.memory1.mem1[78][0] ),
    .X(net4658));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\top1.memory2.mem2[129][1] ),
    .X(net4659));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\top1.memory1.mem1[68][1] ),
    .X(net4660));
 sg13g2_dlygate4sd3_1 hold2223 (.A(\top1.memory1.mem1[82][0] ),
    .X(net4661));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\top1.memory2.mem1[10][2] ),
    .X(net4662));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\top1.memory1.mem1[138][2] ),
    .X(net4663));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\top1.memory1.mem2[99][1] ),
    .X(net4664));
 sg13g2_dlygate4sd3_1 hold2227 (.A(\top1.memory1.mem2[64][2] ),
    .X(net4665));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\top1.memory1.mem2[69][2] ),
    .X(net4666));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\top1.memory1.mem2[6][2] ),
    .X(net4667));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\top1.memory2.mem1[99][1] ),
    .X(net4668));
 sg13g2_dlygate4sd3_1 hold2231 (.A(\top1.memory1.mem2[88][1] ),
    .X(net4669));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\top1.memory2.mem1[70][0] ),
    .X(net4670));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\top1.memory1.mem1[12][0] ),
    .X(net4671));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\top1.memory2.mem2[77][0] ),
    .X(net4672));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\top1.memory1.mem1[76][0] ),
    .X(net4673));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\top1.memory1.mem1[104][1] ),
    .X(net4674));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\top1.fsm.idx_final[2] ),
    .X(net4675));
 sg13g2_dlygate4sd3_1 hold2238 (.A(_01313_),
    .X(net4676));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\top1.memory2.mem2[145][2] ),
    .X(net4677));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\top1.memory2.mem1[104][2] ),
    .X(net4678));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\top1.memory2.mem1[1][0] ),
    .X(net4679));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\top1.memory2.mem2[76][1] ),
    .X(net4680));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\top1.memory2.mem2[64][0] ),
    .X(net4681));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\top1.memory1.mem1[67][2] ),
    .X(net4682));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\top1.memory1.mem1[80][1] ),
    .X(net4683));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\top1.memory2.mem1[8][1] ),
    .X(net4684));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\top1.memory1.mem1[137][1] ),
    .X(net4685));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\top1.memory2.mem2[15][1] ),
    .X(net4686));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\top1.memory1.mem1[79][2] ),
    .X(net4687));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\top1.memory2.mem2[68][2] ),
    .X(net4688));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\top1.memory1.mem1[99][2] ),
    .X(net4689));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\top1.memory1.mem1[1][0] ),
    .X(net4690));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\top1.memory2.mem1[2][1] ),
    .X(net4691));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\top1.memory2.mem1[4][0] ),
    .X(net4692));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\top1.memory1.mem1[199][0] ),
    .X(net4693));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\top1.memory2.mem1[199][1] ),
    .X(net4694));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\top1.memory1.mem2[140][0] ),
    .X(net4695));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\top1.memory2.mem2[137][0] ),
    .X(net4696));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\top1.memory1.mem1[3][0] ),
    .X(net4697));
 sg13g2_dlygate4sd3_1 hold2260 (.A(\top1.memory1.mem1[6][0] ),
    .X(net4698));
 sg13g2_dlygate4sd3_1 hold2261 (.A(\top1.memory1.mem1[10][0] ),
    .X(net4699));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\top1.memory1.mem1[97][2] ),
    .X(net4700));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\top1.memory2.mem1[78][0] ),
    .X(net4701));
 sg13g2_dlygate4sd3_1 hold2264 (.A(\top1.memory2.mem2[142][2] ),
    .X(net4702));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\top1.memory1.mem2[65][0] ),
    .X(net4703));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\top1.memory2.mem2[82][2] ),
    .X(net4704));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\top1.fsm.idx_final[6] ),
    .X(net4705));
 sg13g2_dlygate4sd3_1 hold2268 (.A(_01317_),
    .X(net4706));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\top1.memory2.mem2[3][2] ),
    .X(net4707));
 sg13g2_dlygate4sd3_1 hold2270 (.A(\top1.memory2.mem2[138][1] ),
    .X(net4708));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\top1.memory1.mem2[146][0] ),
    .X(net4709));
 sg13g2_dlygate4sd3_1 hold2272 (.A(\top1.memory1.mem1[66][2] ),
    .X(net4710));
 sg13g2_dlygate4sd3_1 hold2273 (.A(\top1.memory2.mem2[10][1] ),
    .X(net4711));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\top1.memory1.mem2[0][0] ),
    .X(net4712));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\top1.fsm.idx_final[5] ),
    .X(net4713));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\top1.memory2.mem2[161][1] ),
    .X(net4714));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\top1.memory2.mem1[80][0] ),
    .X(net4715));
 sg13g2_dlygate4sd3_1 hold2278 (.A(\top1.memory2.mem1[73][0] ),
    .X(net4716));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\top1.memory2.mem2[162][0] ),
    .X(net4717));
 sg13g2_dlygate4sd3_1 hold2280 (.A(\top1.memory2.mem1[6][0] ),
    .X(net4718));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\top1.memory1.mem2[132][0] ),
    .X(net4719));
 sg13g2_dlygate4sd3_1 hold2282 (.A(\top1.memory1.mem2[68][0] ),
    .X(net4720));
 sg13g2_dlygate4sd3_1 hold2283 (.A(\top1.memory1.mem1[12][2] ),
    .X(net4721));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\top1.memory2.mem1[139][0] ),
    .X(net4722));
 sg13g2_dlygate4sd3_1 hold2285 (.A(\top1.memory2.mem2[65][1] ),
    .X(net4723));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\top1.memory1.mem2[82][0] ),
    .X(net4724));
 sg13g2_dlygate4sd3_1 hold2287 (.A(\top1.memory2.mem2[74][2] ),
    .X(net4725));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\top1.memory2.mem2[0][1] ),
    .X(net4726));
 sg13g2_dlygate4sd3_1 hold2289 (.A(\top1.memory2.mem2[82][0] ),
    .X(net4727));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\top1.memory1.mem2[162][0] ),
    .X(net4728));
 sg13g2_dlygate4sd3_1 hold2291 (.A(\top1.memory2.mem2[140][2] ),
    .X(net4729));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\top1.memory1.mem2[98][1] ),
    .X(net4730));
 sg13g2_dlygate4sd3_1 hold2293 (.A(\top1.memory2.mem1[79][0] ),
    .X(net4731));
 sg13g2_dlygate4sd3_1 hold2294 (.A(\top1.memory1.mem1[134][2] ),
    .X(net4732));
 sg13g2_dlygate4sd3_1 hold2295 (.A(\top1.memory2.mem1[80][1] ),
    .X(net4733));
 sg13g2_dlygate4sd3_1 hold2296 (.A(\top1.memory2.mem1[84][2] ),
    .X(net4734));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\top1.memory1.mem1[129][0] ),
    .X(net4735));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\top1.memory2.mem1[10][1] ),
    .X(net4736));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\top1.memory2.mem2[199][2] ),
    .X(net4737));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\top1.memory1.mem2[73][1] ),
    .X(net4738));
 sg13g2_dlygate4sd3_1 hold2301 (.A(\top1.fsm.idx_final[4] ),
    .X(net4739));
 sg13g2_dlygate4sd3_1 hold2302 (.A(_01315_),
    .X(net4740));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\top1.memory1.mem2[84][0] ),
    .X(net4741));
 sg13g2_dlygate4sd3_1 hold2304 (.A(\top1.memory1.mem2[2][0] ),
    .X(net4742));
 sg13g2_dlygate4sd3_1 hold2305 (.A(\top1.memory2.mem2[4][2] ),
    .X(net4743));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\top1.memory1.mem2[131][2] ),
    .X(net4744));
 sg13g2_dlygate4sd3_1 hold2307 (.A(\top1.memory1.mem1[72][2] ),
    .X(net4745));
 sg13g2_dlygate4sd3_1 hold2308 (.A(\top1.memory2.mem1[0][1] ),
    .X(net4746));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\top1.memory1.mem1[142][2] ),
    .X(net4747));
 sg13g2_dlygate4sd3_1 hold2310 (.A(\top1.memory2.mem1[6][2] ),
    .X(net4748));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\top1.memory1.mem1[146][0] ),
    .X(net4749));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\top1.memory2.mem2[130][1] ),
    .X(net4750));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\top1.memory2.mem2[79][2] ),
    .X(net4751));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\top1.memory2.mem2[98][2] ),
    .X(net4752));
 sg13g2_dlygate4sd3_1 hold2315 (.A(\top1.memory2.mem2[2][2] ),
    .X(net4753));
 sg13g2_dlygate4sd3_1 hold2316 (.A(\top1.memory2.mem1[3][1] ),
    .X(net4754));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\top1.memory2.mem2[127][1] ),
    .X(net4755));
 sg13g2_dlygate4sd3_1 hold2318 (.A(\top1.memory1.mem2[1][1] ),
    .X(net4756));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\top1.memory1.mem2[79][0] ),
    .X(net4757));
 sg13g2_dlygate4sd3_1 hold2320 (.A(\top1.memory1.mem1[4][0] ),
    .X(net4758));
 sg13g2_dlygate4sd3_1 hold2321 (.A(\top1.memory2.mem2[127][0] ),
    .X(net4759));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\top1.memory1.mem1[80][0] ),
    .X(net4760));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\top1.memory2.mem2[134][1] ),
    .X(net4761));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\top1.memory2.mem2[64][2] ),
    .X(net4762));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\top1.memory2.mem2[136][2] ),
    .X(net4763));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\top1.memory2.mem2[73][1] ),
    .X(net4764));
 sg13g2_dlygate4sd3_1 hold2327 (.A(\top1.memory2.mem1[129][1] ),
    .X(net4765));
 sg13g2_dlygate4sd3_1 hold2328 (.A(\top1.memory1.mem2[10][0] ),
    .X(net4766));
 sg13g2_dlygate4sd3_1 hold2329 (.A(\top1.memory2.mem1[162][2] ),
    .X(net4767));
 sg13g2_dlygate4sd3_1 hold2330 (.A(\top1.memory1.mem2[64][1] ),
    .X(net4768));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\top1.memory2.mem2[75][2] ),
    .X(net4769));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\top1.memory1.mem2[65][1] ),
    .X(net4770));
 sg13g2_dlygate4sd3_1 hold2333 (.A(\top1.memory1.mem1[144][1] ),
    .X(net4771));
 sg13g2_dlygate4sd3_1 hold2334 (.A(\top1.memory2.mem1[130][2] ),
    .X(net4772));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\top1.memory2.mem1[98][0] ),
    .X(net4773));
 sg13g2_dlygate4sd3_1 hold2336 (.A(\top1.memory2.mem1[66][1] ),
    .X(net4774));
 sg13g2_dlygate4sd3_1 hold2337 (.A(\top1.memory2.mem1[130][0] ),
    .X(net4775));
 sg13g2_dlygate4sd3_1 hold2338 (.A(\top1.memory1.mem1[8][1] ),
    .X(net4776));
 sg13g2_dlygate4sd3_1 hold2339 (.A(\top1.memory2.mem2[143][2] ),
    .X(net4777));
 sg13g2_dlygate4sd3_1 hold2340 (.A(\top1.memory1.mem2[78][1] ),
    .X(net4778));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\top1.memory2.mem2[77][2] ),
    .X(net4779));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\top1.memory2.mem2[100][2] ),
    .X(net4780));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\top1.memory2.mem1[144][0] ),
    .X(net4781));
 sg13g2_dlygate4sd3_1 hold2344 (.A(\top1.memory2.mem1[104][1] ),
    .X(net4782));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\top1.memory2.mem1[160][0] ),
    .X(net4783));
 sg13g2_dlygate4sd3_1 hold2346 (.A(\top1.memory1.mem2[141][2] ),
    .X(net4784));
 sg13g2_dlygate4sd3_1 hold2347 (.A(\top1.memory2.mem1[76][1] ),
    .X(net4785));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\top1.memory1.mem1[64][2] ),
    .X(net4786));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\top1.memory1.mem2[58][0] ),
    .X(net4787));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\top1.memory2.mem2[84][0] ),
    .X(net4788));
 sg13g2_dlygate4sd3_1 hold2351 (.A(\top1.memory2.mem1[134][1] ),
    .X(net4789));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\top1.memory2.mem2[67][0] ),
    .X(net4790));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\top1.memory2.mem2[80][2] ),
    .X(net4791));
 sg13g2_dlygate4sd3_1 hold2354 (.A(\top1.memory1.mem2[8][0] ),
    .X(net4792));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\top1.memory2.mem2[141][0] ),
    .X(net4793));
 sg13g2_dlygate4sd3_1 hold2356 (.A(\top1.memory2.mem2[136][0] ),
    .X(net4794));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\top1.memory1.mem2[77][1] ),
    .X(net4795));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\top1.memory2.mem2[160][0] ),
    .X(net4796));
 sg13g2_dlygate4sd3_1 hold2359 (.A(\top1.memory1.mem2[82][2] ),
    .X(net4797));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\top1.memory1.mem2[6][1] ),
    .X(net4798));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\top1.memory1.mem1[77][0] ),
    .X(net4799));
 sg13g2_dlygate4sd3_1 hold2362 (.A(\top1.memory2.mem2[128][0] ),
    .X(net4800));
 sg13g2_dlygate4sd3_1 hold2363 (.A(\top1.memory2.mem2[98][0] ),
    .X(net4801));
 sg13g2_dlygate4sd3_1 hold2364 (.A(\top1.memory1.mem1[3][1] ),
    .X(net4802));
 sg13g2_dlygate4sd3_1 hold2365 (.A(\top1.memory1.mem2[12][0] ),
    .X(net4803));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\top1.memory2.mem2[96][2] ),
    .X(net4804));
 sg13g2_dlygate4sd3_1 hold2367 (.A(\top1.memory1.mem2[141][0] ),
    .X(net4805));
 sg13g2_dlygate4sd3_1 hold2368 (.A(\top1.memory2.mem2[129][2] ),
    .X(net4806));
 sg13g2_dlygate4sd3_1 hold2369 (.A(\top1.memory2.mem2[73][0] ),
    .X(net4807));
 sg13g2_dlygate4sd3_1 hold2370 (.A(\top1.memory2.mem2[161][2] ),
    .X(net4808));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\top1.memory1.mem2[97][1] ),
    .X(net4809));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\top1.memory2.mem2[78][0] ),
    .X(net4810));
 sg13g2_dlygate4sd3_1 hold2373 (.A(\top1.memory1.mem1[134][1] ),
    .X(net4811));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\top1.memory2.mem2[66][1] ),
    .X(net4812));
 sg13g2_dlygate4sd3_1 hold2375 (.A(\top1.memory1.mem1[96][1] ),
    .X(net4813));
 sg13g2_dlygate4sd3_1 hold2376 (.A(\top1.memory1.mem2[76][1] ),
    .X(net4814));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\top1.memory2.mem1[99][0] ),
    .X(net4815));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\top1.memory1.mem1[82][1] ),
    .X(net4816));
 sg13g2_dlygate4sd3_1 hold2379 (.A(\top1.memory1.mem2[66][2] ),
    .X(net4817));
 sg13g2_dlygate4sd3_1 hold2380 (.A(\top1.memory2.mem2[74][1] ),
    .X(net4818));
 sg13g2_dlygate4sd3_1 hold2381 (.A(\top1.memory2.mem1[64][1] ),
    .X(net4819));
 sg13g2_dlygate4sd3_1 hold2382 (.A(\top1.memory1.mem2[96][2] ),
    .X(net4820));
 sg13g2_dlygate4sd3_1 hold2383 (.A(\top1.memory1.mem1[162][1] ),
    .X(net4821));
 sg13g2_dlygate4sd3_1 hold2384 (.A(\top1.memory1.mem2[81][0] ),
    .X(net4822));
 sg13g2_dlygate4sd3_1 hold2385 (.A(\top1.memory1.mem1[145][1] ),
    .X(net4823));
 sg13g2_dlygate4sd3_1 hold2386 (.A(\top1.memory2.mem1[15][1] ),
    .X(net4824));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\top1.memory2.mem2[1][1] ),
    .X(net4825));
 sg13g2_dlygate4sd3_1 hold2388 (.A(\top1.memory2.mem1[128][2] ),
    .X(net4826));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\top1.memory2.mem1[144][1] ),
    .X(net4827));
 sg13g2_dlygate4sd3_1 hold2390 (.A(\top1.memory2.mem2[98][1] ),
    .X(net4828));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\top1.memory1.mem1[141][1] ),
    .X(net4829));
 sg13g2_dlygate4sd3_1 hold2392 (.A(\top1.memory2.mem2[146][1] ),
    .X(net4830));
 sg13g2_dlygate4sd3_1 hold2393 (.A(\top1.memory2.mem2[79][0] ),
    .X(net4831));
 sg13g2_dlygate4sd3_1 hold2394 (.A(\top1.memory2.mem2[76][0] ),
    .X(net4832));
 sg13g2_dlygate4sd3_1 hold2395 (.A(\top1.memory1.mem2[15][0] ),
    .X(net4833));
 sg13g2_dlygate4sd3_1 hold2396 (.A(\top1.memory1.mem1[0][2] ),
    .X(net4834));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\top1.memory1.mem2[80][2] ),
    .X(net4835));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\top1.memory1.mem1[9][1] ),
    .X(net4836));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\top1.memory2.mem2[70][2] ),
    .X(net4837));
 sg13g2_dlygate4sd3_1 hold2400 (.A(\top1.memory1.mem1[98][1] ),
    .X(net4838));
 sg13g2_dlygate4sd3_1 hold2401 (.A(\top1.memory2.mem1[3][2] ),
    .X(net4839));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\top1.memory1.mem1[128][0] ),
    .X(net4840));
 sg13g2_dlygate4sd3_1 hold2403 (.A(\top1.memory2.mem1[145][1] ),
    .X(net4841));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\top1.memory1.mem2[199][2] ),
    .X(net4842));
 sg13g2_dlygate4sd3_1 hold2405 (.A(\top1.memory2.mem2[104][2] ),
    .X(net4843));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\top1.memory2.mem2[75][0] ),
    .X(net4844));
 sg13g2_dlygate4sd3_1 hold2407 (.A(\top1.memory1.mem2[83][0] ),
    .X(net4845));
 sg13g2_dlygate4sd3_1 hold2408 (.A(\top1.memory2.mem2[82][1] ),
    .X(net4846));
 sg13g2_dlygate4sd3_1 hold2409 (.A(\top1.memory1.mem1[15][2] ),
    .X(net4847));
 sg13g2_dlygate4sd3_1 hold2410 (.A(\top1.memory1.mem2[96][0] ),
    .X(net4848));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\top1.memory1.mem1[81][2] ),
    .X(net4849));
 sg13g2_dlygate4sd3_1 hold2412 (.A(\top1.memory1.mem2[8][1] ),
    .X(net4850));
 sg13g2_dlygate4sd3_1 hold2413 (.A(_00000_),
    .X(net4851));
 sg13g2_dlygate4sd3_1 hold2414 (.A(_01308_),
    .X(net4852));
 sg13g2_dlygate4sd3_1 hold2415 (.A(\top1.memory1.mem1[136][0] ),
    .X(net4853));
 sg13g2_dlygate4sd3_1 hold2416 (.A(\top1.memory1.mem2[79][2] ),
    .X(net4854));
 sg13g2_dlygate4sd3_1 hold2417 (.A(\top1.memory2.mem1[10][0] ),
    .X(net4855));
 sg13g2_dlygate4sd3_1 hold2418 (.A(\top1.memory1.mem2[77][2] ),
    .X(net4856));
 sg13g2_dlygate4sd3_1 hold2419 (.A(\top1.memory1.mem1[78][1] ),
    .X(net4857));
 sg13g2_dlygate4sd3_1 hold2420 (.A(\top1.bank0_full ),
    .X(net4858));
 sg13g2_dlygate4sd3_1 hold2421 (.A(_01310_),
    .X(net4859));
 sg13g2_dlygate4sd3_1 hold2422 (.A(\top1.bank1_full ),
    .X(net4860));
 sg13g2_dlygate4sd3_1 hold2423 (.A(_02616_),
    .X(net4861));
 sg13g2_dlygate4sd3_1 hold2424 (.A(_01319_),
    .X(net4862));
 sg13g2_dlygate4sd3_1 hold2425 (.A(\top1.addr_in[0] ),
    .X(net4863));
 sg13g2_dlygate4sd3_1 hold2426 (.A(\top1.addr_in[2] ),
    .X(net4864));
 sg13g2_dlygate4sd3_1 hold2427 (.A(_04046_),
    .X(net4865));
 sg13g2_dlygate4sd3_1 hold2428 (.A(\top1.addr_in[4] ),
    .X(net4866));
 sg13g2_dlygate4sd3_1 hold2429 (.A(_03846_),
    .X(net4867));
 sg13g2_dlygate4sd3_1 hold2430 (.A(\top1.addr_in[5] ),
    .X(net4868));
 sg13g2_dlygate4sd3_1 hold2431 (.A(\top1.addr_in[7] ),
    .X(net4869));
 sg13g2_dlygate4sd3_1 hold2432 (.A(\top1.mem_ctl.state_reg[1] ),
    .X(net4870));
 sg13g2_antennanp ANTENNA_1 (.A(_00049_));
 sg13g2_antennanp ANTENNA_2 (.A(_04109_));
 sg13g2_antennanp ANTENNA_3 (.A(_04159_));
 sg13g2_antennanp ANTENNA_4 (.A(_04716_));
 sg13g2_antennanp ANTENNA_5 (.A(_04716_));
 sg13g2_antennanp ANTENNA_6 (.A(_04716_));
 sg13g2_antennanp ANTENNA_7 (.A(_05511_));
 sg13g2_antennanp ANTENNA_8 (.A(_05567_));
 sg13g2_antennanp ANTENNA_9 (.A(_05939_));
 sg13g2_antennanp ANTENNA_10 (.A(_06074_));
 sg13g2_antennanp ANTENNA_11 (.A(_06181_));
 sg13g2_antennanp ANTENNA_12 (.A(_06224_));
 sg13g2_antennanp ANTENNA_13 (.A(_06259_));
 sg13g2_antennanp ANTENNA_14 (.A(_06393_));
 sg13g2_antennanp ANTENNA_15 (.A(_06488_));
 sg13g2_antennanp ANTENNA_16 (.A(_06680_));
 sg13g2_antennanp ANTENNA_17 (.A(_06681_));
 sg13g2_antennanp ANTENNA_18 (.A(_06818_));
 sg13g2_antennanp ANTENNA_19 (.A(_06820_));
 sg13g2_antennanp ANTENNA_20 (.A(_06906_));
 sg13g2_antennanp ANTENNA_21 (.A(_07106_));
 sg13g2_antennanp ANTENNA_22 (.A(_07279_));
 sg13g2_antennanp ANTENNA_23 (.A(clk));
 sg13g2_antennanp ANTENNA_24 (.A(clk));
 sg13g2_antennanp ANTENNA_25 (.A(rst_n));
 sg13g2_antennanp ANTENNA_26 (.A(rst_n));
 sg13g2_antennanp ANTENNA_27 (.A(\top1.acquisition_clk ));
 sg13g2_antennanp ANTENNA_28 (.A(net5871));
 sg13g2_antennanp ANTENNA_29 (.A(net5871));
 sg13g2_antennanp ANTENNA_30 (.A(net5871));
 sg13g2_antennanp ANTENNA_31 (.A(net5871));
 sg13g2_antennanp ANTENNA_32 (.A(net5871));
 sg13g2_antennanp ANTENNA_33 (.A(net5871));
 sg13g2_antennanp ANTENNA_34 (.A(net5871));
 sg13g2_antennanp ANTENNA_35 (.A(net5871));
 sg13g2_antennanp ANTENNA_36 (.A(net5871));
 sg13g2_antennanp ANTENNA_37 (.A(net5871));
 sg13g2_antennanp ANTENNA_38 (.A(net5871));
 sg13g2_antennanp ANTENNA_39 (.A(net5871));
 sg13g2_antennanp ANTENNA_40 (.A(net5871));
 sg13g2_antennanp ANTENNA_41 (.A(net5871));
 sg13g2_antennanp ANTENNA_42 (.A(net5871));
 sg13g2_antennanp ANTENNA_43 (.A(net5871));
 sg13g2_antennanp ANTENNA_44 (.A(net5871));
 sg13g2_antennanp ANTENNA_45 (.A(net5871));
 sg13g2_antennanp ANTENNA_46 (.A(net5980));
 sg13g2_antennanp ANTENNA_47 (.A(net5980));
 sg13g2_antennanp ANTENNA_48 (.A(net5980));
 sg13g2_antennanp ANTENNA_49 (.A(net5980));
 sg13g2_antennanp ANTENNA_50 (.A(net5980));
 sg13g2_antennanp ANTENNA_51 (.A(net5980));
 sg13g2_antennanp ANTENNA_52 (.A(net5980));
 sg13g2_antennanp ANTENNA_53 (.A(net5980));
 sg13g2_antennanp ANTENNA_54 (.A(net6107));
 sg13g2_antennanp ANTENNA_55 (.A(net6107));
 sg13g2_antennanp ANTENNA_56 (.A(net6107));
 sg13g2_antennanp ANTENNA_57 (.A(net6107));
 sg13g2_antennanp ANTENNA_58 (.A(net6107));
 sg13g2_antennanp ANTENNA_59 (.A(net6107));
 sg13g2_antennanp ANTENNA_60 (.A(net6107));
 sg13g2_antennanp ANTENNA_61 (.A(net6107));
 sg13g2_antennanp ANTENNA_62 (.A(net6107));
 sg13g2_antennanp ANTENNA_63 (.A(net6107));
 sg13g2_antennanp ANTENNA_64 (.A(net6107));
 sg13g2_antennanp ANTENNA_65 (.A(net6107));
 sg13g2_antennanp ANTENNA_66 (.A(net6107));
 sg13g2_antennanp ANTENNA_67 (.A(net6107));
 sg13g2_antennanp ANTENNA_68 (.A(net6107));
 sg13g2_antennanp ANTENNA_69 (.A(net7065));
 sg13g2_antennanp ANTENNA_70 (.A(net7065));
 sg13g2_antennanp ANTENNA_71 (.A(net7065));
 sg13g2_antennanp ANTENNA_72 (.A(net7065));
 sg13g2_antennanp ANTENNA_73 (.A(net7065));
 sg13g2_antennanp ANTENNA_74 (.A(net7065));
 sg13g2_antennanp ANTENNA_75 (.A(net7065));
 sg13g2_antennanp ANTENNA_76 (.A(net7065));
 sg13g2_antennanp ANTENNA_77 (.A(net7065));
 sg13g2_antennanp ANTENNA_78 (.A(net7065));
 sg13g2_antennanp ANTENNA_79 (.A(net7065));
 sg13g2_antennanp ANTENNA_80 (.A(net7065));
 sg13g2_antennanp ANTENNA_81 (.A(net7065));
 sg13g2_antennanp ANTENNA_82 (.A(net7065));
 sg13g2_antennanp ANTENNA_83 (.A(net7065));
 sg13g2_antennanp ANTENNA_84 (.A(net7065));
 sg13g2_antennanp ANTENNA_85 (.A(net7065));
 sg13g2_antennanp ANTENNA_86 (.A(net7065));
 sg13g2_antennanp ANTENNA_87 (.A(net7065));
 sg13g2_antennanp ANTENNA_88 (.A(net7065));
 sg13g2_antennanp ANTENNA_89 (.A(net7247));
 sg13g2_antennanp ANTENNA_90 (.A(net7247));
 sg13g2_antennanp ANTENNA_91 (.A(net7247));
 sg13g2_antennanp ANTENNA_92 (.A(net7247));
 sg13g2_antennanp ANTENNA_93 (.A(net7247));
 sg13g2_antennanp ANTENNA_94 (.A(net7247));
 sg13g2_antennanp ANTENNA_95 (.A(net7247));
 sg13g2_antennanp ANTENNA_96 (.A(net7247));
 sg13g2_antennanp ANTENNA_97 (.A(net7277));
 sg13g2_antennanp ANTENNA_98 (.A(net7277));
 sg13g2_antennanp ANTENNA_99 (.A(net7277));
 sg13g2_antennanp ANTENNA_100 (.A(net7277));
 sg13g2_antennanp ANTENNA_101 (.A(net7277));
 sg13g2_antennanp ANTENNA_102 (.A(net7277));
 sg13g2_antennanp ANTENNA_103 (.A(net7277));
 sg13g2_antennanp ANTENNA_104 (.A(net7277));
 sg13g2_antennanp ANTENNA_105 (.A(net7277));
 sg13g2_antennanp ANTENNA_106 (.A(net7277));
 sg13g2_antennanp ANTENNA_107 (.A(net7277));
 sg13g2_antennanp ANTENNA_108 (.A(net7277));
 sg13g2_antennanp ANTENNA_109 (.A(net7277));
 sg13g2_antennanp ANTENNA_110 (.A(net7277));
 sg13g2_antennanp ANTENNA_111 (.A(net7277));
 sg13g2_antennanp ANTENNA_112 (.A(net7277));
 sg13g2_antennanp ANTENNA_113 (.A(net7280));
 sg13g2_antennanp ANTENNA_114 (.A(net7280));
 sg13g2_antennanp ANTENNA_115 (.A(net7280));
 sg13g2_antennanp ANTENNA_116 (.A(net7280));
 sg13g2_antennanp ANTENNA_117 (.A(net7280));
 sg13g2_antennanp ANTENNA_118 (.A(net7280));
 sg13g2_antennanp ANTENNA_119 (.A(net7280));
 sg13g2_antennanp ANTENNA_120 (.A(net7280));
 sg13g2_antennanp ANTENNA_121 (.A(net7280));
 sg13g2_antennanp ANTENNA_122 (.A(net7280));
 sg13g2_antennanp ANTENNA_123 (.A(net7280));
 sg13g2_antennanp ANTENNA_124 (.A(net7280));
 sg13g2_antennanp ANTENNA_125 (.A(net7280));
 sg13g2_antennanp ANTENNA_126 (.A(net7280));
 sg13g2_antennanp ANTENNA_127 (.A(net7280));
 sg13g2_antennanp ANTENNA_128 (.A(net7280));
 sg13g2_antennanp ANTENNA_129 (.A(net7280));
 sg13g2_antennanp ANTENNA_130 (.A(net7280));
 sg13g2_antennanp ANTENNA_131 (.A(net7280));
 sg13g2_antennanp ANTENNA_132 (.A(net7284));
 sg13g2_antennanp ANTENNA_133 (.A(net7284));
 sg13g2_antennanp ANTENNA_134 (.A(net7284));
 sg13g2_antennanp ANTENNA_135 (.A(net7284));
 sg13g2_antennanp ANTENNA_136 (.A(net7284));
 sg13g2_antennanp ANTENNA_137 (.A(net7284));
 sg13g2_antennanp ANTENNA_138 (.A(net7284));
 sg13g2_antennanp ANTENNA_139 (.A(net7284));
 sg13g2_antennanp ANTENNA_140 (.A(net7284));
 sg13g2_antennanp ANTENNA_141 (.A(net7284));
 sg13g2_antennanp ANTENNA_142 (.A(net7284));
 sg13g2_antennanp ANTENNA_143 (.A(net7284));
 sg13g2_antennanp ANTENNA_144 (.A(net7284));
 sg13g2_antennanp ANTENNA_145 (.A(net7284));
 sg13g2_antennanp ANTENNA_146 (.A(net7284));
 sg13g2_antennanp ANTENNA_147 (.A(net7284));
 sg13g2_antennanp ANTENNA_148 (.A(net7284));
 sg13g2_antennanp ANTENNA_149 (.A(net7284));
 sg13g2_antennanp ANTENNA_150 (.A(net7361));
 sg13g2_antennanp ANTENNA_151 (.A(net7361));
 sg13g2_antennanp ANTENNA_152 (.A(net7361));
 sg13g2_antennanp ANTENNA_153 (.A(net7361));
 sg13g2_antennanp ANTENNA_154 (.A(net7361));
 sg13g2_antennanp ANTENNA_155 (.A(net7361));
 sg13g2_antennanp ANTENNA_156 (.A(net7361));
 sg13g2_antennanp ANTENNA_157 (.A(net7361));
 sg13g2_antennanp ANTENNA_158 (.A(net7361));
 sg13g2_antennanp ANTENNA_159 (.A(net7361));
 sg13g2_antennanp ANTENNA_160 (.A(net7361));
 sg13g2_antennanp ANTENNA_161 (.A(net7361));
 sg13g2_antennanp ANTENNA_162 (.A(net7361));
 sg13g2_antennanp ANTENNA_163 (.A(net7361));
 sg13g2_antennanp ANTENNA_164 (.A(net7361));
 sg13g2_antennanp ANTENNA_165 (.A(net7361));
 sg13g2_antennanp ANTENNA_166 (.A(net7361));
 sg13g2_antennanp ANTENNA_167 (.A(net7361));
 sg13g2_antennanp ANTENNA_168 (.A(net7361));
 sg13g2_antennanp ANTENNA_169 (.A(net7361));
 sg13g2_antennanp ANTENNA_170 (.A(net7361));
 sg13g2_antennanp ANTENNA_171 (.A(net7361));
 sg13g2_antennanp ANTENNA_172 (.A(net7404));
 sg13g2_antennanp ANTENNA_173 (.A(net7404));
 sg13g2_antennanp ANTENNA_174 (.A(net7404));
 sg13g2_antennanp ANTENNA_175 (.A(net7404));
 sg13g2_antennanp ANTENNA_176 (.A(net7404));
 sg13g2_antennanp ANTENNA_177 (.A(net7404));
 sg13g2_antennanp ANTENNA_178 (.A(net7404));
 sg13g2_antennanp ANTENNA_179 (.A(net7404));
 sg13g2_antennanp ANTENNA_180 (.A(net7404));
 sg13g2_antennanp ANTENNA_181 (.A(net7404));
 sg13g2_antennanp ANTENNA_182 (.A(net7404));
 sg13g2_antennanp ANTENNA_183 (.A(net7404));
 sg13g2_antennanp ANTENNA_184 (.A(net7404));
 sg13g2_antennanp ANTENNA_185 (.A(net7404));
 sg13g2_antennanp ANTENNA_186 (.A(net7404));
 sg13g2_antennanp ANTENNA_187 (.A(net7404));
 sg13g2_antennanp ANTENNA_188 (.A(net7404));
 sg13g2_antennanp ANTENNA_189 (.A(net7404));
 sg13g2_antennanp ANTENNA_190 (.A(net7522));
 sg13g2_antennanp ANTENNA_191 (.A(net7522));
 sg13g2_antennanp ANTENNA_192 (.A(net7522));
 sg13g2_antennanp ANTENNA_193 (.A(net7522));
 sg13g2_antennanp ANTENNA_194 (.A(net7522));
 sg13g2_antennanp ANTENNA_195 (.A(net7522));
 sg13g2_antennanp ANTENNA_196 (.A(net7522));
 sg13g2_antennanp ANTENNA_197 (.A(net7522));
 sg13g2_antennanp ANTENNA_198 (.A(net7522));
 sg13g2_antennanp ANTENNA_199 (.A(net7607));
 sg13g2_antennanp ANTENNA_200 (.A(net7607));
 sg13g2_antennanp ANTENNA_201 (.A(net7607));
 sg13g2_antennanp ANTENNA_202 (.A(net7607));
 sg13g2_antennanp ANTENNA_203 (.A(net7607));
 sg13g2_antennanp ANTENNA_204 (.A(net7607));
 sg13g2_antennanp ANTENNA_205 (.A(net7607));
 sg13g2_antennanp ANTENNA_206 (.A(net7607));
 sg13g2_antennanp ANTENNA_207 (.A(net7607));
 sg13g2_antennanp ANTENNA_208 (.A(net7607));
 sg13g2_antennanp ANTENNA_209 (.A(net7607));
 sg13g2_antennanp ANTENNA_210 (.A(net1));
 sg13g2_antennanp ANTENNA_211 (.A(net1));
 sg13g2_antennanp ANTENNA_212 (.A(net1));
 sg13g2_antennanp ANTENNA_213 (.A(net1));
 sg13g2_antennanp ANTENNA_214 (.A(net2));
 sg13g2_antennanp ANTENNA_215 (.A(net2));
 sg13g2_antennanp ANTENNA_216 (.A(net2));
 sg13g2_antennanp ANTENNA_217 (.A(net2));
 sg13g2_antennanp ANTENNA_218 (.A(net9));
 sg13g2_antennanp ANTENNA_219 (.A(net9));
 sg13g2_antennanp ANTENNA_220 (.A(net9));
 sg13g2_antennanp ANTENNA_221 (.A(net9));
 sg13g2_antennanp ANTENNA_222 (.A(net10));
 sg13g2_antennanp ANTENNA_223 (.A(net10));
 sg13g2_antennanp ANTENNA_224 (.A(net10));
 sg13g2_antennanp ANTENNA_225 (.A(net10));
 sg13g2_antennanp ANTENNA_226 (.A(net11));
 sg13g2_antennanp ANTENNA_227 (.A(net11));
 sg13g2_antennanp ANTENNA_228 (.A(net11));
 sg13g2_antennanp ANTENNA_229 (.A(net11));
 sg13g2_antennanp ANTENNA_230 (.A(net16));
 sg13g2_antennanp ANTENNA_231 (.A(_00049_));
 sg13g2_antennanp ANTENNA_232 (.A(_04109_));
 sg13g2_antennanp ANTENNA_233 (.A(_04159_));
 sg13g2_antennanp ANTENNA_234 (.A(_04716_));
 sg13g2_antennanp ANTENNA_235 (.A(_04716_));
 sg13g2_antennanp ANTENNA_236 (.A(_04716_));
 sg13g2_antennanp ANTENNA_237 (.A(_04716_));
 sg13g2_antennanp ANTENNA_238 (.A(_05511_));
 sg13g2_antennanp ANTENNA_239 (.A(_05567_));
 sg13g2_antennanp ANTENNA_240 (.A(_05595_));
 sg13g2_antennanp ANTENNA_241 (.A(_05620_));
 sg13g2_antennanp ANTENNA_242 (.A(_05939_));
 sg13g2_antennanp ANTENNA_243 (.A(_06181_));
 sg13g2_antennanp ANTENNA_244 (.A(_06224_));
 sg13g2_antennanp ANTENNA_245 (.A(_06259_));
 sg13g2_antennanp ANTENNA_246 (.A(_06393_));
 sg13g2_antennanp ANTENNA_247 (.A(_06680_));
 sg13g2_antennanp ANTENNA_248 (.A(_06681_));
 sg13g2_antennanp ANTENNA_249 (.A(_06730_));
 sg13g2_antennanp ANTENNA_250 (.A(_06818_));
 sg13g2_antennanp ANTENNA_251 (.A(_06906_));
 sg13g2_antennanp ANTENNA_252 (.A(_07106_));
 sg13g2_antennanp ANTENNA_253 (.A(_07279_));
 sg13g2_antennanp ANTENNA_254 (.A(clk));
 sg13g2_antennanp ANTENNA_255 (.A(clk));
 sg13g2_antennanp ANTENNA_256 (.A(rst_n));
 sg13g2_antennanp ANTENNA_257 (.A(rst_n));
 sg13g2_antennanp ANTENNA_258 (.A(net5980));
 sg13g2_antennanp ANTENNA_259 (.A(net5980));
 sg13g2_antennanp ANTENNA_260 (.A(net5980));
 sg13g2_antennanp ANTENNA_261 (.A(net5980));
 sg13g2_antennanp ANTENNA_262 (.A(net5980));
 sg13g2_antennanp ANTENNA_263 (.A(net7065));
 sg13g2_antennanp ANTENNA_264 (.A(net7065));
 sg13g2_antennanp ANTENNA_265 (.A(net7065));
 sg13g2_antennanp ANTENNA_266 (.A(net7065));
 sg13g2_antennanp ANTENNA_267 (.A(net7065));
 sg13g2_antennanp ANTENNA_268 (.A(net7065));
 sg13g2_antennanp ANTENNA_269 (.A(net7065));
 sg13g2_antennanp ANTENNA_270 (.A(net7065));
 sg13g2_antennanp ANTENNA_271 (.A(net7065));
 sg13g2_antennanp ANTENNA_272 (.A(net7065));
 sg13g2_antennanp ANTENNA_273 (.A(net7065));
 sg13g2_antennanp ANTENNA_274 (.A(net7065));
 sg13g2_antennanp ANTENNA_275 (.A(net7065));
 sg13g2_antennanp ANTENNA_276 (.A(net7065));
 sg13g2_antennanp ANTENNA_277 (.A(net7065));
 sg13g2_antennanp ANTENNA_278 (.A(net7065));
 sg13g2_antennanp ANTENNA_279 (.A(net7065));
 sg13g2_antennanp ANTENNA_280 (.A(net7065));
 sg13g2_antennanp ANTENNA_281 (.A(net7065));
 sg13g2_antennanp ANTENNA_282 (.A(net7065));
 sg13g2_antennanp ANTENNA_283 (.A(net7273));
 sg13g2_antennanp ANTENNA_284 (.A(net7273));
 sg13g2_antennanp ANTENNA_285 (.A(net7273));
 sg13g2_antennanp ANTENNA_286 (.A(net7273));
 sg13g2_antennanp ANTENNA_287 (.A(net7273));
 sg13g2_antennanp ANTENNA_288 (.A(net7273));
 sg13g2_antennanp ANTENNA_289 (.A(net7273));
 sg13g2_antennanp ANTENNA_290 (.A(net7273));
 sg13g2_antennanp ANTENNA_291 (.A(net7273));
 sg13g2_antennanp ANTENNA_292 (.A(net7273));
 sg13g2_antennanp ANTENNA_293 (.A(net7273));
 sg13g2_antennanp ANTENNA_294 (.A(net7273));
 sg13g2_antennanp ANTENNA_295 (.A(net7273));
 sg13g2_antennanp ANTENNA_296 (.A(net7273));
 sg13g2_antennanp ANTENNA_297 (.A(net7273));
 sg13g2_antennanp ANTENNA_298 (.A(net7273));
 sg13g2_antennanp ANTENNA_299 (.A(net7273));
 sg13g2_antennanp ANTENNA_300 (.A(net7275));
 sg13g2_antennanp ANTENNA_301 (.A(net7275));
 sg13g2_antennanp ANTENNA_302 (.A(net7275));
 sg13g2_antennanp ANTENNA_303 (.A(net7275));
 sg13g2_antennanp ANTENNA_304 (.A(net7275));
 sg13g2_antennanp ANTENNA_305 (.A(net7275));
 sg13g2_antennanp ANTENNA_306 (.A(net7275));
 sg13g2_antennanp ANTENNA_307 (.A(net7275));
 sg13g2_antennanp ANTENNA_308 (.A(net7275));
 sg13g2_antennanp ANTENNA_309 (.A(net7275));
 sg13g2_antennanp ANTENNA_310 (.A(net7275));
 sg13g2_antennanp ANTENNA_311 (.A(net7275));
 sg13g2_antennanp ANTENNA_312 (.A(net7275));
 sg13g2_antennanp ANTENNA_313 (.A(net7275));
 sg13g2_antennanp ANTENNA_314 (.A(net7275));
 sg13g2_antennanp ANTENNA_315 (.A(net7275));
 sg13g2_antennanp ANTENNA_316 (.A(net7275));
 sg13g2_antennanp ANTENNA_317 (.A(net7275));
 sg13g2_antennanp ANTENNA_318 (.A(net7277));
 sg13g2_antennanp ANTENNA_319 (.A(net7277));
 sg13g2_antennanp ANTENNA_320 (.A(net7277));
 sg13g2_antennanp ANTENNA_321 (.A(net7277));
 sg13g2_antennanp ANTENNA_322 (.A(net7277));
 sg13g2_antennanp ANTENNA_323 (.A(net7277));
 sg13g2_antennanp ANTENNA_324 (.A(net7277));
 sg13g2_antennanp ANTENNA_325 (.A(net7277));
 sg13g2_antennanp ANTENNA_326 (.A(net7277));
 sg13g2_antennanp ANTENNA_327 (.A(net7277));
 sg13g2_antennanp ANTENNA_328 (.A(net7277));
 sg13g2_antennanp ANTENNA_329 (.A(net7277));
 sg13g2_antennanp ANTENNA_330 (.A(net7277));
 sg13g2_antennanp ANTENNA_331 (.A(net7277));
 sg13g2_antennanp ANTENNA_332 (.A(net7277));
 sg13g2_antennanp ANTENNA_333 (.A(net7277));
 sg13g2_antennanp ANTENNA_334 (.A(net7284));
 sg13g2_antennanp ANTENNA_335 (.A(net7284));
 sg13g2_antennanp ANTENNA_336 (.A(net7284));
 sg13g2_antennanp ANTENNA_337 (.A(net7284));
 sg13g2_antennanp ANTENNA_338 (.A(net7284));
 sg13g2_antennanp ANTENNA_339 (.A(net7284));
 sg13g2_antennanp ANTENNA_340 (.A(net7284));
 sg13g2_antennanp ANTENNA_341 (.A(net7284));
 sg13g2_antennanp ANTENNA_342 (.A(net7361));
 sg13g2_antennanp ANTENNA_343 (.A(net7361));
 sg13g2_antennanp ANTENNA_344 (.A(net7361));
 sg13g2_antennanp ANTENNA_345 (.A(net7361));
 sg13g2_antennanp ANTENNA_346 (.A(net7361));
 sg13g2_antennanp ANTENNA_347 (.A(net7361));
 sg13g2_antennanp ANTENNA_348 (.A(net7361));
 sg13g2_antennanp ANTENNA_349 (.A(net7361));
 sg13g2_antennanp ANTENNA_350 (.A(net7522));
 sg13g2_antennanp ANTENNA_351 (.A(net7522));
 sg13g2_antennanp ANTENNA_352 (.A(net7522));
 sg13g2_antennanp ANTENNA_353 (.A(net7522));
 sg13g2_antennanp ANTENNA_354 (.A(net7522));
 sg13g2_antennanp ANTENNA_355 (.A(net7522));
 sg13g2_antennanp ANTENNA_356 (.A(net7522));
 sg13g2_antennanp ANTENNA_357 (.A(net7522));
 sg13g2_antennanp ANTENNA_358 (.A(net7522));
 sg13g2_antennanp ANTENNA_359 (.A(net7522));
 sg13g2_antennanp ANTENNA_360 (.A(net7522));
 sg13g2_antennanp ANTENNA_361 (.A(net7607));
 sg13g2_antennanp ANTENNA_362 (.A(net7607));
 sg13g2_antennanp ANTENNA_363 (.A(net7607));
 sg13g2_antennanp ANTENNA_364 (.A(net7607));
 sg13g2_antennanp ANTENNA_365 (.A(net7607));
 sg13g2_antennanp ANTENNA_366 (.A(net7607));
 sg13g2_antennanp ANTENNA_367 (.A(net7607));
 sg13g2_antennanp ANTENNA_368 (.A(net7607));
 sg13g2_antennanp ANTENNA_369 (.A(net7607));
 sg13g2_antennanp ANTENNA_370 (.A(net7607));
 sg13g2_antennanp ANTENNA_371 (.A(net7607));
 sg13g2_antennanp ANTENNA_372 (.A(net1));
 sg13g2_antennanp ANTENNA_373 (.A(net1));
 sg13g2_antennanp ANTENNA_374 (.A(net1));
 sg13g2_antennanp ANTENNA_375 (.A(net1));
 sg13g2_antennanp ANTENNA_376 (.A(net2));
 sg13g2_antennanp ANTENNA_377 (.A(net2));
 sg13g2_antennanp ANTENNA_378 (.A(net2));
 sg13g2_antennanp ANTENNA_379 (.A(net2));
 sg13g2_antennanp ANTENNA_380 (.A(net9));
 sg13g2_antennanp ANTENNA_381 (.A(net9));
 sg13g2_antennanp ANTENNA_382 (.A(net9));
 sg13g2_antennanp ANTENNA_383 (.A(net9));
 sg13g2_antennanp ANTENNA_384 (.A(net10));
 sg13g2_antennanp ANTENNA_385 (.A(net10));
 sg13g2_antennanp ANTENNA_386 (.A(net10));
 sg13g2_antennanp ANTENNA_387 (.A(net10));
 sg13g2_antennanp ANTENNA_388 (.A(net11));
 sg13g2_antennanp ANTENNA_389 (.A(net11));
 sg13g2_antennanp ANTENNA_390 (.A(net11));
 sg13g2_antennanp ANTENNA_391 (.A(net11));
 sg13g2_antennanp ANTENNA_392 (.A(_00049_));
 sg13g2_antennanp ANTENNA_393 (.A(_04109_));
 sg13g2_antennanp ANTENNA_394 (.A(_04159_));
 sg13g2_antennanp ANTENNA_395 (.A(_04716_));
 sg13g2_antennanp ANTENNA_396 (.A(_04716_));
 sg13g2_antennanp ANTENNA_397 (.A(_04716_));
 sg13g2_antennanp ANTENNA_398 (.A(_04716_));
 sg13g2_antennanp ANTENNA_399 (.A(_05511_));
 sg13g2_antennanp ANTENNA_400 (.A(_05567_));
 sg13g2_antennanp ANTENNA_401 (.A(_05595_));
 sg13g2_antennanp ANTENNA_402 (.A(_05939_));
 sg13g2_antennanp ANTENNA_403 (.A(_06224_));
 sg13g2_antennanp ANTENNA_404 (.A(_06259_));
 sg13g2_antennanp ANTENNA_405 (.A(_06680_));
 sg13g2_antennanp ANTENNA_406 (.A(_06730_));
 sg13g2_antennanp ANTENNA_407 (.A(_06818_));
 sg13g2_antennanp ANTENNA_408 (.A(_06906_));
 sg13g2_antennanp ANTENNA_409 (.A(_07279_));
 sg13g2_antennanp ANTENNA_410 (.A(clk));
 sg13g2_antennanp ANTENNA_411 (.A(clk));
 sg13g2_antennanp ANTENNA_412 (.A(rst_n));
 sg13g2_antennanp ANTENNA_413 (.A(rst_n));
 sg13g2_antennanp ANTENNA_414 (.A(net7065));
 sg13g2_antennanp ANTENNA_415 (.A(net7065));
 sg13g2_antennanp ANTENNA_416 (.A(net7065));
 sg13g2_antennanp ANTENNA_417 (.A(net7065));
 sg13g2_antennanp ANTENNA_418 (.A(net7065));
 sg13g2_antennanp ANTENNA_419 (.A(net7065));
 sg13g2_antennanp ANTENNA_420 (.A(net7065));
 sg13g2_antennanp ANTENNA_421 (.A(net7065));
 sg13g2_antennanp ANTENNA_422 (.A(net7065));
 sg13g2_antennanp ANTENNA_423 (.A(net7065));
 sg13g2_antennanp ANTENNA_424 (.A(net7065));
 sg13g2_antennanp ANTENNA_425 (.A(net7065));
 sg13g2_antennanp ANTENNA_426 (.A(net7065));
 sg13g2_antennanp ANTENNA_427 (.A(net7065));
 sg13g2_antennanp ANTENNA_428 (.A(net7065));
 sg13g2_antennanp ANTENNA_429 (.A(net7065));
 sg13g2_antennanp ANTENNA_430 (.A(net7065));
 sg13g2_antennanp ANTENNA_431 (.A(net7065));
 sg13g2_antennanp ANTENNA_432 (.A(net7065));
 sg13g2_antennanp ANTENNA_433 (.A(net7065));
 sg13g2_antennanp ANTENNA_434 (.A(net7273));
 sg13g2_antennanp ANTENNA_435 (.A(net7273));
 sg13g2_antennanp ANTENNA_436 (.A(net7273));
 sg13g2_antennanp ANTENNA_437 (.A(net7273));
 sg13g2_antennanp ANTENNA_438 (.A(net7273));
 sg13g2_antennanp ANTENNA_439 (.A(net7273));
 sg13g2_antennanp ANTENNA_440 (.A(net7273));
 sg13g2_antennanp ANTENNA_441 (.A(net7273));
 sg13g2_antennanp ANTENNA_442 (.A(net7273));
 sg13g2_antennanp ANTENNA_443 (.A(net7273));
 sg13g2_antennanp ANTENNA_444 (.A(net7273));
 sg13g2_antennanp ANTENNA_445 (.A(net7273));
 sg13g2_antennanp ANTENNA_446 (.A(net7277));
 sg13g2_antennanp ANTENNA_447 (.A(net7277));
 sg13g2_antennanp ANTENNA_448 (.A(net7277));
 sg13g2_antennanp ANTENNA_449 (.A(net7277));
 sg13g2_antennanp ANTENNA_450 (.A(net7277));
 sg13g2_antennanp ANTENNA_451 (.A(net7277));
 sg13g2_antennanp ANTENNA_452 (.A(net7277));
 sg13g2_antennanp ANTENNA_453 (.A(net7277));
 sg13g2_antennanp ANTENNA_454 (.A(net7277));
 sg13g2_antennanp ANTENNA_455 (.A(net7277));
 sg13g2_antennanp ANTENNA_456 (.A(net7277));
 sg13g2_antennanp ANTENNA_457 (.A(net7277));
 sg13g2_antennanp ANTENNA_458 (.A(net7277));
 sg13g2_antennanp ANTENNA_459 (.A(net7277));
 sg13g2_antennanp ANTENNA_460 (.A(net7277));
 sg13g2_antennanp ANTENNA_461 (.A(net7277));
 sg13g2_antennanp ANTENNA_462 (.A(net7522));
 sg13g2_antennanp ANTENNA_463 (.A(net7522));
 sg13g2_antennanp ANTENNA_464 (.A(net7522));
 sg13g2_antennanp ANTENNA_465 (.A(net7522));
 sg13g2_antennanp ANTENNA_466 (.A(net7522));
 sg13g2_antennanp ANTENNA_467 (.A(net7522));
 sg13g2_antennanp ANTENNA_468 (.A(net7522));
 sg13g2_antennanp ANTENNA_469 (.A(net7522));
 sg13g2_antennanp ANTENNA_470 (.A(net7522));
 sg13g2_antennanp ANTENNA_471 (.A(net7522));
 sg13g2_antennanp ANTENNA_472 (.A(net7522));
 sg13g2_antennanp ANTENNA_473 (.A(net7522));
 sg13g2_antennanp ANTENNA_474 (.A(net7522));
 sg13g2_antennanp ANTENNA_475 (.A(net2));
 sg13g2_antennanp ANTENNA_476 (.A(net2));
 sg13g2_antennanp ANTENNA_477 (.A(net2));
 sg13g2_antennanp ANTENNA_478 (.A(net2));
 sg13g2_antennanp ANTENNA_479 (.A(net9));
 sg13g2_antennanp ANTENNA_480 (.A(net9));
 sg13g2_antennanp ANTENNA_481 (.A(net9));
 sg13g2_antennanp ANTENNA_482 (.A(net9));
 sg13g2_antennanp ANTENNA_483 (.A(net10));
 sg13g2_antennanp ANTENNA_484 (.A(net10));
 sg13g2_antennanp ANTENNA_485 (.A(net10));
 sg13g2_antennanp ANTENNA_486 (.A(net10));
 sg13g2_antennanp ANTENNA_487 (.A(net11));
 sg13g2_antennanp ANTENNA_488 (.A(net11));
 sg13g2_antennanp ANTENNA_489 (.A(net11));
 sg13g2_antennanp ANTENNA_490 (.A(net11));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_fill_1 FILLER_0_567 ();
 sg13g2_fill_1 FILLER_0_594 ();
 sg13g2_fill_1 FILLER_0_603 ();
 sg13g2_fill_1 FILLER_0_608 ();
 sg13g2_fill_1 FILLER_0_613 ();
 sg13g2_decap_4 FILLER_0_640 ();
 sg13g2_fill_2 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_654 ();
 sg13g2_decap_4 FILLER_0_661 ();
 sg13g2_fill_1 FILLER_0_665 ();
 sg13g2_fill_2 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_676 ();
 sg13g2_decap_4 FILLER_0_683 ();
 sg13g2_fill_1 FILLER_0_687 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_fill_1 FILLER_0_704 ();
 sg13g2_decap_8 FILLER_0_709 ();
 sg13g2_decap_8 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_730 ();
 sg13g2_decap_4 FILLER_0_737 ();
 sg13g2_fill_2 FILLER_0_741 ();
 sg13g2_fill_2 FILLER_0_776 ();
 sg13g2_fill_1 FILLER_0_778 ();
 sg13g2_fill_2 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_fill_1 FILLER_0_840 ();
 sg13g2_decap_4 FILLER_0_892 ();
 sg13g2_fill_1 FILLER_0_896 ();
 sg13g2_fill_1 FILLER_0_914 ();
 sg13g2_fill_2 FILLER_0_978 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_8 FILLER_0_1025 ();
 sg13g2_fill_2 FILLER_0_1032 ();
 sg13g2_fill_1 FILLER_0_1034 ();
 sg13g2_fill_2 FILLER_0_1065 ();
 sg13g2_fill_1 FILLER_0_1067 ();
 sg13g2_fill_2 FILLER_0_1119 ();
 sg13g2_decap_8 FILLER_0_1169 ();
 sg13g2_decap_8 FILLER_0_1176 ();
 sg13g2_decap_8 FILLER_0_1183 ();
 sg13g2_fill_2 FILLER_0_1190 ();
 sg13g2_fill_1 FILLER_0_1192 ();
 sg13g2_decap_8 FILLER_0_1197 ();
 sg13g2_decap_4 FILLER_0_1204 ();
 sg13g2_fill_1 FILLER_0_1208 ();
 sg13g2_decap_4 FILLER_0_1247 ();
 sg13g2_decap_4 FILLER_0_1277 ();
 sg13g2_fill_1 FILLER_0_1281 ();
 sg13g2_fill_1 FILLER_0_1334 ();
 sg13g2_decap_8 FILLER_0_1344 ();
 sg13g2_decap_4 FILLER_0_1351 ();
 sg13g2_fill_2 FILLER_0_1355 ();
 sg13g2_fill_2 FILLER_0_1361 ();
 sg13g2_decap_4 FILLER_0_1367 ();
 sg13g2_fill_2 FILLER_0_1371 ();
 sg13g2_fill_2 FILLER_0_1377 ();
 sg13g2_fill_2 FILLER_0_1387 ();
 sg13g2_fill_1 FILLER_0_1398 ();
 sg13g2_fill_2 FILLER_0_1403 ();
 sg13g2_fill_2 FILLER_0_1424 ();
 sg13g2_fill_2 FILLER_0_1434 ();
 sg13g2_fill_1 FILLER_0_1436 ();
 sg13g2_fill_1 FILLER_0_1454 ();
 sg13g2_fill_2 FILLER_0_1463 ();
 sg13g2_fill_1 FILLER_0_1465 ();
 sg13g2_decap_8 FILLER_0_1474 ();
 sg13g2_decap_8 FILLER_0_1481 ();
 sg13g2_decap_8 FILLER_0_1509 ();
 sg13g2_decap_4 FILLER_0_1516 ();
 sg13g2_fill_1 FILLER_0_1520 ();
 sg13g2_fill_2 FILLER_0_1526 ();
 sg13g2_fill_2 FILLER_0_1537 ();
 sg13g2_decap_4 FILLER_0_1556 ();
 sg13g2_fill_1 FILLER_0_1560 ();
 sg13g2_fill_1 FILLER_0_1583 ();
 sg13g2_fill_2 FILLER_0_1605 ();
 sg13g2_decap_4 FILLER_0_1678 ();
 sg13g2_fill_1 FILLER_0_1682 ();
 sg13g2_fill_2 FILLER_0_1688 ();
 sg13g2_fill_1 FILLER_0_1690 ();
 sg13g2_fill_2 FILLER_0_1700 ();
 sg13g2_fill_1 FILLER_0_1702 ();
 sg13g2_decap_8 FILLER_0_1707 ();
 sg13g2_decap_8 FILLER_0_1714 ();
 sg13g2_fill_2 FILLER_0_1721 ();
 sg13g2_fill_1 FILLER_0_1723 ();
 sg13g2_decap_8 FILLER_0_1728 ();
 sg13g2_decap_8 FILLER_0_1735 ();
 sg13g2_decap_8 FILLER_0_1742 ();
 sg13g2_decap_8 FILLER_0_1749 ();
 sg13g2_decap_8 FILLER_0_1756 ();
 sg13g2_decap_8 FILLER_0_1763 ();
 sg13g2_decap_4 FILLER_0_1770 ();
 sg13g2_fill_1 FILLER_0_1774 ();
 sg13g2_decap_4 FILLER_0_1784 ();
 sg13g2_fill_1 FILLER_0_1788 ();
 sg13g2_fill_2 FILLER_0_1810 ();
 sg13g2_fill_1 FILLER_0_1812 ();
 sg13g2_fill_1 FILLER_0_1818 ();
 sg13g2_fill_2 FILLER_0_1831 ();
 sg13g2_fill_1 FILLER_0_1833 ();
 sg13g2_fill_2 FILLER_0_1847 ();
 sg13g2_fill_1 FILLER_0_1849 ();
 sg13g2_decap_8 FILLER_0_1884 ();
 sg13g2_decap_8 FILLER_0_1891 ();
 sg13g2_decap_8 FILLER_0_1898 ();
 sg13g2_decap_8 FILLER_0_1905 ();
 sg13g2_decap_8 FILLER_0_1912 ();
 sg13g2_decap_8 FILLER_0_1919 ();
 sg13g2_decap_4 FILLER_0_1926 ();
 sg13g2_decap_8 FILLER_0_1947 ();
 sg13g2_decap_4 FILLER_0_1954 ();
 sg13g2_fill_2 FILLER_0_1958 ();
 sg13g2_fill_2 FILLER_0_1965 ();
 sg13g2_fill_1 FILLER_0_1967 ();
 sg13g2_decap_8 FILLER_0_1985 ();
 sg13g2_fill_2 FILLER_0_1992 ();
 sg13g2_fill_1 FILLER_0_1994 ();
 sg13g2_fill_1 FILLER_0_2003 ();
 sg13g2_fill_1 FILLER_0_2008 ();
 sg13g2_fill_2 FILLER_0_2027 ();
 sg13g2_decap_8 FILLER_0_2046 ();
 sg13g2_fill_2 FILLER_0_2057 ();
 sg13g2_fill_1 FILLER_0_2059 ();
 sg13g2_decap_4 FILLER_0_2064 ();
 sg13g2_decap_8 FILLER_0_2085 ();
 sg13g2_decap_8 FILLER_0_2092 ();
 sg13g2_fill_2 FILLER_0_2099 ();
 sg13g2_decap_4 FILLER_0_2166 ();
 sg13g2_fill_1 FILLER_0_2170 ();
 sg13g2_fill_2 FILLER_0_2249 ();
 sg13g2_fill_1 FILLER_0_2251 ();
 sg13g2_fill_2 FILLER_0_2283 ();
 sg13g2_fill_2 FILLER_0_2307 ();
 sg13g2_fill_1 FILLER_0_2309 ();
 sg13g2_fill_1 FILLER_0_2323 ();
 sg13g2_fill_1 FILLER_0_2350 ();
 sg13g2_fill_2 FILLER_0_2373 ();
 sg13g2_fill_1 FILLER_0_2375 ();
 sg13g2_fill_2 FILLER_0_2397 ();
 sg13g2_decap_8 FILLER_0_2416 ();
 sg13g2_decap_8 FILLER_0_2423 ();
 sg13g2_decap_8 FILLER_0_2430 ();
 sg13g2_decap_8 FILLER_0_2437 ();
 sg13g2_decap_8 FILLER_0_2444 ();
 sg13g2_decap_8 FILLER_0_2451 ();
 sg13g2_decap_8 FILLER_0_2458 ();
 sg13g2_decap_8 FILLER_0_2465 ();
 sg13g2_decap_8 FILLER_0_2472 ();
 sg13g2_decap_8 FILLER_0_2479 ();
 sg13g2_decap_8 FILLER_0_2486 ();
 sg13g2_decap_8 FILLER_0_2493 ();
 sg13g2_decap_8 FILLER_0_2500 ();
 sg13g2_decap_8 FILLER_0_2507 ();
 sg13g2_decap_8 FILLER_0_2514 ();
 sg13g2_decap_8 FILLER_0_2521 ();
 sg13g2_decap_8 FILLER_0_2528 ();
 sg13g2_decap_8 FILLER_0_2535 ();
 sg13g2_decap_8 FILLER_0_2542 ();
 sg13g2_decap_8 FILLER_0_2549 ();
 sg13g2_decap_8 FILLER_0_2556 ();
 sg13g2_decap_8 FILLER_0_2563 ();
 sg13g2_decap_8 FILLER_0_2570 ();
 sg13g2_decap_8 FILLER_0_2577 ();
 sg13g2_decap_8 FILLER_0_2584 ();
 sg13g2_decap_8 FILLER_0_2591 ();
 sg13g2_decap_8 FILLER_0_2598 ();
 sg13g2_decap_8 FILLER_0_2605 ();
 sg13g2_decap_8 FILLER_0_2612 ();
 sg13g2_decap_8 FILLER_0_2619 ();
 sg13g2_decap_8 FILLER_0_2626 ();
 sg13g2_decap_8 FILLER_0_2633 ();
 sg13g2_decap_8 FILLER_0_2640 ();
 sg13g2_decap_8 FILLER_0_2647 ();
 sg13g2_decap_8 FILLER_0_2654 ();
 sg13g2_decap_8 FILLER_0_2661 ();
 sg13g2_decap_4 FILLER_0_2668 ();
 sg13g2_fill_2 FILLER_0_2672 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_fill_1 FILLER_1_567 ();
 sg13g2_fill_2 FILLER_1_594 ();
 sg13g2_fill_1 FILLER_1_596 ();
 sg13g2_fill_1 FILLER_1_649 ();
 sg13g2_fill_1 FILLER_1_693 ();
 sg13g2_decap_4 FILLER_1_729 ();
 sg13g2_fill_2 FILLER_1_733 ();
 sg13g2_fill_2 FILLER_1_761 ();
 sg13g2_fill_2 FILLER_1_772 ();
 sg13g2_decap_8 FILLER_1_818 ();
 sg13g2_decap_4 FILLER_1_825 ();
 sg13g2_fill_1 FILLER_1_855 ();
 sg13g2_fill_1 FILLER_1_887 ();
 sg13g2_decap_8 FILLER_1_897 ();
 sg13g2_fill_1 FILLER_1_943 ();
 sg13g2_fill_1 FILLER_1_983 ();
 sg13g2_fill_1 FILLER_1_1019 ();
 sg13g2_fill_2 FILLER_1_1028 ();
 sg13g2_fill_1 FILLER_1_1030 ();
 sg13g2_fill_2 FILLER_1_1061 ();
 sg13g2_fill_1 FILLER_1_1063 ();
 sg13g2_fill_1 FILLER_1_1103 ();
 sg13g2_fill_2 FILLER_1_1135 ();
 sg13g2_decap_8 FILLER_1_1172 ();
 sg13g2_decap_8 FILLER_1_1278 ();
 sg13g2_decap_4 FILLER_1_1285 ();
 sg13g2_fill_2 FILLER_1_1289 ();
 sg13g2_fill_2 FILLER_1_1382 ();
 sg13g2_fill_1 FILLER_1_1384 ();
 sg13g2_fill_1 FILLER_1_1459 ();
 sg13g2_fill_2 FILLER_1_1552 ();
 sg13g2_fill_1 FILLER_1_1554 ();
 sg13g2_fill_1 FILLER_1_1563 ();
 sg13g2_fill_1 FILLER_1_1671 ();
 sg13g2_fill_1 FILLER_1_1676 ();
 sg13g2_fill_1 FILLER_1_1712 ();
 sg13g2_decap_8 FILLER_1_1753 ();
 sg13g2_fill_2 FILLER_1_1760 ();
 sg13g2_fill_1 FILLER_1_1762 ();
 sg13g2_fill_2 FILLER_1_1789 ();
 sg13g2_fill_1 FILLER_1_1791 ();
 sg13g2_decap_8 FILLER_1_1892 ();
 sg13g2_decap_8 FILLER_1_1899 ();
 sg13g2_decap_8 FILLER_1_1906 ();
 sg13g2_decap_8 FILLER_1_1913 ();
 sg13g2_fill_2 FILLER_1_1920 ();
 sg13g2_fill_1 FILLER_1_1922 ();
 sg13g2_decap_4 FILLER_1_1953 ();
 sg13g2_fill_1 FILLER_1_1987 ();
 sg13g2_fill_2 FILLER_1_2048 ();
 sg13g2_fill_2 FILLER_1_2055 ();
 sg13g2_fill_2 FILLER_1_2127 ();
 sg13g2_fill_2 FILLER_1_2203 ();
 sg13g2_fill_2 FILLER_1_2235 ();
 sg13g2_fill_1 FILLER_1_2237 ();
 sg13g2_fill_2 FILLER_1_2264 ();
 sg13g2_fill_1 FILLER_1_2266 ();
 sg13g2_fill_2 FILLER_1_2349 ();
 sg13g2_fill_1 FILLER_1_2351 ();
 sg13g2_fill_2 FILLER_1_2378 ();
 sg13g2_fill_1 FILLER_1_2380 ();
 sg13g2_fill_2 FILLER_1_2394 ();
 sg13g2_decap_8 FILLER_1_2435 ();
 sg13g2_decap_8 FILLER_1_2442 ();
 sg13g2_decap_8 FILLER_1_2449 ();
 sg13g2_decap_8 FILLER_1_2456 ();
 sg13g2_decap_8 FILLER_1_2463 ();
 sg13g2_decap_8 FILLER_1_2470 ();
 sg13g2_decap_8 FILLER_1_2477 ();
 sg13g2_decap_8 FILLER_1_2484 ();
 sg13g2_decap_8 FILLER_1_2491 ();
 sg13g2_decap_8 FILLER_1_2498 ();
 sg13g2_decap_8 FILLER_1_2505 ();
 sg13g2_decap_8 FILLER_1_2512 ();
 sg13g2_decap_8 FILLER_1_2519 ();
 sg13g2_decap_8 FILLER_1_2526 ();
 sg13g2_decap_8 FILLER_1_2533 ();
 sg13g2_decap_8 FILLER_1_2540 ();
 sg13g2_decap_8 FILLER_1_2547 ();
 sg13g2_decap_8 FILLER_1_2554 ();
 sg13g2_decap_8 FILLER_1_2561 ();
 sg13g2_decap_8 FILLER_1_2568 ();
 sg13g2_decap_8 FILLER_1_2575 ();
 sg13g2_decap_8 FILLER_1_2582 ();
 sg13g2_decap_8 FILLER_1_2589 ();
 sg13g2_decap_8 FILLER_1_2596 ();
 sg13g2_decap_8 FILLER_1_2603 ();
 sg13g2_decap_8 FILLER_1_2610 ();
 sg13g2_decap_8 FILLER_1_2617 ();
 sg13g2_decap_8 FILLER_1_2624 ();
 sg13g2_decap_8 FILLER_1_2631 ();
 sg13g2_decap_8 FILLER_1_2638 ();
 sg13g2_decap_8 FILLER_1_2645 ();
 sg13g2_decap_8 FILLER_1_2652 ();
 sg13g2_decap_8 FILLER_1_2659 ();
 sg13g2_decap_8 FILLER_1_2666 ();
 sg13g2_fill_1 FILLER_1_2673 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_fill_2 FILLER_2_644 ();
 sg13g2_fill_2 FILLER_2_663 ();
 sg13g2_fill_1 FILLER_2_665 ();
 sg13g2_fill_1 FILLER_2_696 ();
 sg13g2_fill_1 FILLER_2_702 ();
 sg13g2_fill_2 FILLER_2_764 ();
 sg13g2_fill_2 FILLER_2_826 ();
 sg13g2_fill_1 FILLER_2_828 ();
 sg13g2_fill_1 FILLER_2_982 ();
 sg13g2_fill_2 FILLER_2_993 ();
 sg13g2_fill_1 FILLER_2_1034 ();
 sg13g2_fill_1 FILLER_2_1065 ();
 sg13g2_fill_2 FILLER_2_1106 ();
 sg13g2_fill_2 FILLER_2_1138 ();
 sg13g2_fill_1 FILLER_2_1140 ();
 sg13g2_fill_2 FILLER_2_1176 ();
 sg13g2_fill_2 FILLER_2_1223 ();
 sg13g2_fill_2 FILLER_2_1282 ();
 sg13g2_fill_1 FILLER_2_1471 ();
 sg13g2_fill_2 FILLER_2_1503 ();
 sg13g2_fill_1 FILLER_2_1505 ();
 sg13g2_fill_2 FILLER_2_1589 ();
 sg13g2_fill_2 FILLER_2_1751 ();
 sg13g2_fill_1 FILLER_2_1753 ();
 sg13g2_fill_1 FILLER_2_1846 ();
 sg13g2_fill_2 FILLER_2_1873 ();
 sg13g2_fill_1 FILLER_2_1875 ();
 sg13g2_fill_2 FILLER_2_1889 ();
 sg13g2_fill_1 FILLER_2_1891 ();
 sg13g2_decap_8 FILLER_2_1900 ();
 sg13g2_decap_4 FILLER_2_1907 ();
 sg13g2_fill_1 FILLER_2_1951 ();
 sg13g2_fill_1 FILLER_2_1983 ();
 sg13g2_fill_2 FILLER_2_2019 ();
 sg13g2_fill_1 FILLER_2_2021 ();
 sg13g2_fill_2 FILLER_2_2100 ();
 sg13g2_fill_1 FILLER_2_2102 ();
 sg13g2_fill_1 FILLER_2_2107 ();
 sg13g2_fill_1 FILLER_2_2210 ();
 sg13g2_fill_2 FILLER_2_2226 ();
 sg13g2_fill_1 FILLER_2_2228 ();
 sg13g2_fill_1 FILLER_2_2242 ();
 sg13g2_fill_2 FILLER_2_2253 ();
 sg13g2_fill_1 FILLER_2_2278 ();
 sg13g2_decap_8 FILLER_2_2444 ();
 sg13g2_decap_8 FILLER_2_2451 ();
 sg13g2_decap_8 FILLER_2_2458 ();
 sg13g2_decap_8 FILLER_2_2465 ();
 sg13g2_decap_8 FILLER_2_2472 ();
 sg13g2_decap_8 FILLER_2_2479 ();
 sg13g2_decap_8 FILLER_2_2486 ();
 sg13g2_decap_8 FILLER_2_2493 ();
 sg13g2_decap_8 FILLER_2_2500 ();
 sg13g2_decap_8 FILLER_2_2507 ();
 sg13g2_decap_8 FILLER_2_2514 ();
 sg13g2_decap_8 FILLER_2_2521 ();
 sg13g2_decap_8 FILLER_2_2528 ();
 sg13g2_decap_8 FILLER_2_2535 ();
 sg13g2_decap_8 FILLER_2_2542 ();
 sg13g2_decap_8 FILLER_2_2549 ();
 sg13g2_decap_8 FILLER_2_2556 ();
 sg13g2_decap_8 FILLER_2_2563 ();
 sg13g2_decap_8 FILLER_2_2570 ();
 sg13g2_decap_8 FILLER_2_2577 ();
 sg13g2_decap_8 FILLER_2_2584 ();
 sg13g2_decap_8 FILLER_2_2591 ();
 sg13g2_decap_8 FILLER_2_2598 ();
 sg13g2_decap_8 FILLER_2_2605 ();
 sg13g2_decap_8 FILLER_2_2612 ();
 sg13g2_decap_8 FILLER_2_2619 ();
 sg13g2_decap_8 FILLER_2_2626 ();
 sg13g2_decap_8 FILLER_2_2633 ();
 sg13g2_decap_8 FILLER_2_2640 ();
 sg13g2_decap_8 FILLER_2_2647 ();
 sg13g2_decap_8 FILLER_2_2654 ();
 sg13g2_decap_8 FILLER_2_2661 ();
 sg13g2_decap_4 FILLER_2_2668 ();
 sg13g2_fill_2 FILLER_2_2672 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_fill_2 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_524 ();
 sg13g2_decap_8 FILLER_3_531 ();
 sg13g2_decap_8 FILLER_3_538 ();
 sg13g2_decap_8 FILLER_3_545 ();
 sg13g2_decap_4 FILLER_3_552 ();
 sg13g2_fill_1 FILLER_3_556 ();
 sg13g2_fill_1 FILLER_3_578 ();
 sg13g2_fill_1 FILLER_3_619 ();
 sg13g2_fill_2 FILLER_3_655 ();
 sg13g2_fill_2 FILLER_3_687 ();
 sg13g2_fill_2 FILLER_3_732 ();
 sg13g2_fill_2 FILLER_3_829 ();
 sg13g2_fill_1 FILLER_3_888 ();
 sg13g2_fill_2 FILLER_3_938 ();
 sg13g2_fill_1 FILLER_3_1019 ();
 sg13g2_fill_1 FILLER_3_1068 ();
 sg13g2_fill_2 FILLER_3_1099 ();
 sg13g2_fill_2 FILLER_3_1132 ();
 sg13g2_fill_1 FILLER_3_1134 ();
 sg13g2_fill_2 FILLER_3_1240 ();
 sg13g2_fill_2 FILLER_3_1265 ();
 sg13g2_fill_2 FILLER_3_1280 ();
 sg13g2_fill_2 FILLER_3_1324 ();
 sg13g2_fill_1 FILLER_3_1394 ();
 sg13g2_fill_2 FILLER_3_1421 ();
 sg13g2_fill_1 FILLER_3_1423 ();
 sg13g2_fill_1 FILLER_3_1590 ();
 sg13g2_fill_1 FILLER_3_1609 ();
 sg13g2_fill_2 FILLER_3_1673 ();
 sg13g2_fill_1 FILLER_3_1675 ();
 sg13g2_fill_1 FILLER_3_1763 ();
 sg13g2_fill_1 FILLER_3_1848 ();
 sg13g2_fill_1 FILLER_3_1884 ();
 sg13g2_fill_2 FILLER_3_1924 ();
 sg13g2_fill_1 FILLER_3_1926 ();
 sg13g2_fill_1 FILLER_3_1953 ();
 sg13g2_fill_2 FILLER_3_1959 ();
 sg13g2_fill_1 FILLER_3_1961 ();
 sg13g2_fill_1 FILLER_3_2015 ();
 sg13g2_fill_2 FILLER_3_2054 ();
 sg13g2_fill_1 FILLER_3_2056 ();
 sg13g2_decap_8 FILLER_3_2165 ();
 sg13g2_fill_1 FILLER_3_2172 ();
 sg13g2_fill_2 FILLER_3_2203 ();
 sg13g2_fill_1 FILLER_3_2205 ();
 sg13g2_fill_2 FILLER_3_2245 ();
 sg13g2_fill_1 FILLER_3_2247 ();
 sg13g2_fill_2 FILLER_3_2274 ();
 sg13g2_fill_1 FILLER_3_2276 ();
 sg13g2_fill_2 FILLER_3_2311 ();
 sg13g2_fill_1 FILLER_3_2357 ();
 sg13g2_fill_2 FILLER_3_2384 ();
 sg13g2_fill_1 FILLER_3_2386 ();
 sg13g2_decap_8 FILLER_3_2448 ();
 sg13g2_decap_8 FILLER_3_2455 ();
 sg13g2_decap_8 FILLER_3_2462 ();
 sg13g2_decap_8 FILLER_3_2469 ();
 sg13g2_decap_8 FILLER_3_2476 ();
 sg13g2_decap_8 FILLER_3_2483 ();
 sg13g2_decap_8 FILLER_3_2490 ();
 sg13g2_decap_8 FILLER_3_2497 ();
 sg13g2_decap_8 FILLER_3_2504 ();
 sg13g2_decap_8 FILLER_3_2511 ();
 sg13g2_decap_8 FILLER_3_2518 ();
 sg13g2_decap_8 FILLER_3_2525 ();
 sg13g2_decap_8 FILLER_3_2532 ();
 sg13g2_decap_8 FILLER_3_2539 ();
 sg13g2_decap_8 FILLER_3_2546 ();
 sg13g2_decap_8 FILLER_3_2553 ();
 sg13g2_decap_8 FILLER_3_2560 ();
 sg13g2_decap_8 FILLER_3_2567 ();
 sg13g2_decap_8 FILLER_3_2574 ();
 sg13g2_decap_8 FILLER_3_2581 ();
 sg13g2_decap_8 FILLER_3_2588 ();
 sg13g2_decap_8 FILLER_3_2595 ();
 sg13g2_decap_8 FILLER_3_2602 ();
 sg13g2_decap_8 FILLER_3_2609 ();
 sg13g2_decap_8 FILLER_3_2616 ();
 sg13g2_decap_8 FILLER_3_2623 ();
 sg13g2_decap_8 FILLER_3_2630 ();
 sg13g2_decap_8 FILLER_3_2637 ();
 sg13g2_decap_8 FILLER_3_2644 ();
 sg13g2_decap_8 FILLER_3_2651 ();
 sg13g2_decap_8 FILLER_3_2658 ();
 sg13g2_decap_8 FILLER_3_2665 ();
 sg13g2_fill_2 FILLER_3_2672 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_4 FILLER_4_534 ();
 sg13g2_fill_1 FILLER_4_538 ();
 sg13g2_decap_4 FILLER_4_548 ();
 sg13g2_fill_1 FILLER_4_557 ();
 sg13g2_fill_2 FILLER_4_611 ();
 sg13g2_fill_1 FILLER_4_613 ();
 sg13g2_fill_1 FILLER_4_645 ();
 sg13g2_fill_2 FILLER_4_660 ();
 sg13g2_fill_1 FILLER_4_662 ();
 sg13g2_fill_2 FILLER_4_672 ();
 sg13g2_fill_2 FILLER_4_688 ();
 sg13g2_fill_1 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_fill_2 FILLER_4_720 ();
 sg13g2_fill_2 FILLER_4_744 ();
 sg13g2_decap_4 FILLER_4_769 ();
 sg13g2_fill_2 FILLER_4_773 ();
 sg13g2_fill_2 FILLER_4_805 ();
 sg13g2_fill_1 FILLER_4_807 ();
 sg13g2_fill_2 FILLER_4_817 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_4 FILLER_4_830 ();
 sg13g2_decap_4 FILLER_4_838 ();
 sg13g2_fill_2 FILLER_4_842 ();
 sg13g2_decap_4 FILLER_4_883 ();
 sg13g2_fill_1 FILLER_4_887 ();
 sg13g2_fill_2 FILLER_4_892 ();
 sg13g2_fill_1 FILLER_4_894 ();
 sg13g2_fill_2 FILLER_4_933 ();
 sg13g2_fill_1 FILLER_4_935 ();
 sg13g2_fill_2 FILLER_4_946 ();
 sg13g2_fill_1 FILLER_4_948 ();
 sg13g2_fill_2 FILLER_4_1028 ();
 sg13g2_fill_1 FILLER_4_1030 ();
 sg13g2_fill_2 FILLER_4_1131 ();
 sg13g2_fill_2 FILLER_4_1173 ();
 sg13g2_fill_2 FILLER_4_1188 ();
 sg13g2_fill_1 FILLER_4_1190 ();
 sg13g2_fill_1 FILLER_4_1204 ();
 sg13g2_fill_1 FILLER_4_1210 ();
 sg13g2_fill_1 FILLER_4_1254 ();
 sg13g2_fill_2 FILLER_4_1281 ();
 sg13g2_fill_1 FILLER_4_1283 ();
 sg13g2_decap_8 FILLER_4_1349 ();
 sg13g2_fill_1 FILLER_4_1356 ();
 sg13g2_fill_2 FILLER_4_1400 ();
 sg13g2_fill_2 FILLER_4_1407 ();
 sg13g2_fill_2 FILLER_4_1444 ();
 sg13g2_fill_1 FILLER_4_1446 ();
 sg13g2_fill_1 FILLER_4_1478 ();
 sg13g2_fill_2 FILLER_4_1528 ();
 sg13g2_fill_1 FILLER_4_1559 ();
 sg13g2_fill_1 FILLER_4_1635 ();
 sg13g2_fill_2 FILLER_4_1709 ();
 sg13g2_fill_2 FILLER_4_1764 ();
 sg13g2_fill_1 FILLER_4_1766 ();
 sg13g2_fill_2 FILLER_4_1777 ();
 sg13g2_fill_2 FILLER_4_1784 ();
 sg13g2_fill_1 FILLER_4_1786 ();
 sg13g2_fill_2 FILLER_4_1842 ();
 sg13g2_fill_2 FILLER_4_1854 ();
 sg13g2_decap_8 FILLER_4_1885 ();
 sg13g2_decap_8 FILLER_4_1892 ();
 sg13g2_decap_4 FILLER_4_1899 ();
 sg13g2_fill_2 FILLER_4_1903 ();
 sg13g2_fill_2 FILLER_4_1913 ();
 sg13g2_fill_1 FILLER_4_1920 ();
 sg13g2_fill_2 FILLER_4_1994 ();
 sg13g2_fill_1 FILLER_4_2032 ();
 sg13g2_fill_2 FILLER_4_2057 ();
 sg13g2_fill_1 FILLER_4_2059 ();
 sg13g2_fill_1 FILLER_4_2117 ();
 sg13g2_fill_1 FILLER_4_2132 ();
 sg13g2_decap_8 FILLER_4_2159 ();
 sg13g2_decap_4 FILLER_4_2166 ();
 sg13g2_fill_1 FILLER_4_2240 ();
 sg13g2_fill_2 FILLER_4_2300 ();
 sg13g2_fill_1 FILLER_4_2302 ();
 sg13g2_fill_2 FILLER_4_2321 ();
 sg13g2_fill_1 FILLER_4_2323 ();
 sg13g2_fill_2 FILLER_4_2345 ();
 sg13g2_fill_1 FILLER_4_2347 ();
 sg13g2_decap_4 FILLER_4_2447 ();
 sg13g2_fill_2 FILLER_4_2451 ();
 sg13g2_decap_4 FILLER_4_2470 ();
 sg13g2_fill_1 FILLER_4_2482 ();
 sg13g2_decap_8 FILLER_4_2487 ();
 sg13g2_decap_8 FILLER_4_2494 ();
 sg13g2_decap_8 FILLER_4_2501 ();
 sg13g2_decap_8 FILLER_4_2508 ();
 sg13g2_decap_8 FILLER_4_2515 ();
 sg13g2_decap_8 FILLER_4_2522 ();
 sg13g2_decap_8 FILLER_4_2529 ();
 sg13g2_decap_8 FILLER_4_2536 ();
 sg13g2_decap_8 FILLER_4_2543 ();
 sg13g2_decap_8 FILLER_4_2550 ();
 sg13g2_decap_8 FILLER_4_2557 ();
 sg13g2_decap_8 FILLER_4_2564 ();
 sg13g2_decap_8 FILLER_4_2571 ();
 sg13g2_decap_8 FILLER_4_2578 ();
 sg13g2_decap_8 FILLER_4_2585 ();
 sg13g2_decap_8 FILLER_4_2592 ();
 sg13g2_decap_8 FILLER_4_2599 ();
 sg13g2_decap_8 FILLER_4_2606 ();
 sg13g2_decap_8 FILLER_4_2613 ();
 sg13g2_decap_8 FILLER_4_2620 ();
 sg13g2_decap_8 FILLER_4_2627 ();
 sg13g2_decap_8 FILLER_4_2634 ();
 sg13g2_decap_8 FILLER_4_2641 ();
 sg13g2_decap_8 FILLER_4_2648 ();
 sg13g2_decap_8 FILLER_4_2655 ();
 sg13g2_decap_8 FILLER_4_2662 ();
 sg13g2_decap_4 FILLER_4_2669 ();
 sg13g2_fill_1 FILLER_4_2673 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_fill_2 FILLER_5_497 ();
 sg13g2_fill_1 FILLER_5_499 ();
 sg13g2_fill_2 FILLER_5_564 ();
 sg13g2_fill_1 FILLER_5_583 ();
 sg13g2_fill_2 FILLER_5_597 ();
 sg13g2_fill_2 FILLER_5_637 ();
 sg13g2_fill_1 FILLER_5_639 ();
 sg13g2_fill_2 FILLER_5_692 ();
 sg13g2_fill_1 FILLER_5_694 ();
 sg13g2_fill_1 FILLER_5_747 ();
 sg13g2_fill_2 FILLER_5_766 ();
 sg13g2_fill_2 FILLER_5_820 ();
 sg13g2_fill_1 FILLER_5_939 ();
 sg13g2_fill_1 FILLER_5_945 ();
 sg13g2_fill_1 FILLER_5_963 ();
 sg13g2_fill_1 FILLER_5_968 ();
 sg13g2_fill_1 FILLER_5_982 ();
 sg13g2_fill_1 FILLER_5_995 ();
 sg13g2_fill_2 FILLER_5_1041 ();
 sg13g2_fill_1 FILLER_5_1043 ();
 sg13g2_fill_2 FILLER_5_1062 ();
 sg13g2_fill_1 FILLER_5_1142 ();
 sg13g2_fill_2 FILLER_5_1194 ();
 sg13g2_fill_2 FILLER_5_1201 ();
 sg13g2_fill_1 FILLER_5_1256 ();
 sg13g2_decap_4 FILLER_5_1283 ();
 sg13g2_decap_8 FILLER_5_1342 ();
 sg13g2_decap_8 FILLER_5_1349 ();
 sg13g2_decap_4 FILLER_5_1356 ();
 sg13g2_fill_1 FILLER_5_1360 ();
 sg13g2_decap_8 FILLER_5_1390 ();
 sg13g2_fill_1 FILLER_5_1397 ();
 sg13g2_fill_1 FILLER_5_1406 ();
 sg13g2_fill_1 FILLER_5_1415 ();
 sg13g2_decap_8 FILLER_5_1469 ();
 sg13g2_decap_8 FILLER_5_1476 ();
 sg13g2_fill_1 FILLER_5_1483 ();
 sg13g2_fill_1 FILLER_5_1514 ();
 sg13g2_fill_2 FILLER_5_1525 ();
 sg13g2_decap_4 FILLER_5_1548 ();
 sg13g2_fill_1 FILLER_5_1552 ();
 sg13g2_fill_1 FILLER_5_1557 ();
 sg13g2_fill_2 FILLER_5_1658 ();
 sg13g2_fill_1 FILLER_5_1660 ();
 sg13g2_fill_1 FILLER_5_1700 ();
 sg13g2_fill_2 FILLER_5_1710 ();
 sg13g2_fill_2 FILLER_5_1725 ();
 sg13g2_fill_1 FILLER_5_1727 ();
 sg13g2_decap_8 FILLER_5_1753 ();
 sg13g2_fill_1 FILLER_5_1764 ();
 sg13g2_fill_2 FILLER_5_1813 ();
 sg13g2_fill_2 FILLER_5_1893 ();
 sg13g2_fill_2 FILLER_5_1921 ();
 sg13g2_fill_1 FILLER_5_1923 ();
 sg13g2_fill_2 FILLER_5_1969 ();
 sg13g2_fill_1 FILLER_5_1971 ();
 sg13g2_fill_2 FILLER_5_1981 ();
 sg13g2_fill_1 FILLER_5_1996 ();
 sg13g2_fill_2 FILLER_5_2064 ();
 sg13g2_fill_1 FILLER_5_2066 ();
 sg13g2_fill_2 FILLER_5_2089 ();
 sg13g2_fill_1 FILLER_5_2091 ();
 sg13g2_decap_8 FILLER_5_2167 ();
 sg13g2_fill_2 FILLER_5_2174 ();
 sg13g2_fill_2 FILLER_5_2212 ();
 sg13g2_fill_1 FILLER_5_2235 ();
 sg13g2_fill_1 FILLER_5_2245 ();
 sg13g2_fill_2 FILLER_5_2276 ();
 sg13g2_fill_1 FILLER_5_2343 ();
 sg13g2_fill_2 FILLER_5_2353 ();
 sg13g2_fill_1 FILLER_5_2355 ();
 sg13g2_fill_2 FILLER_5_2366 ();
 sg13g2_fill_1 FILLER_5_2368 ();
 sg13g2_fill_2 FILLER_5_2390 ();
 sg13g2_fill_2 FILLER_5_2411 ();
 sg13g2_fill_2 FILLER_5_2443 ();
 sg13g2_decap_8 FILLER_5_2493 ();
 sg13g2_fill_2 FILLER_5_2505 ();
 sg13g2_fill_1 FILLER_5_2507 ();
 sg13g2_decap_8 FILLER_5_2538 ();
 sg13g2_decap_8 FILLER_5_2545 ();
 sg13g2_decap_8 FILLER_5_2552 ();
 sg13g2_decap_8 FILLER_5_2559 ();
 sg13g2_decap_8 FILLER_5_2566 ();
 sg13g2_decap_8 FILLER_5_2573 ();
 sg13g2_decap_8 FILLER_5_2580 ();
 sg13g2_decap_8 FILLER_5_2587 ();
 sg13g2_decap_8 FILLER_5_2594 ();
 sg13g2_decap_8 FILLER_5_2601 ();
 sg13g2_decap_8 FILLER_5_2608 ();
 sg13g2_decap_8 FILLER_5_2615 ();
 sg13g2_decap_8 FILLER_5_2622 ();
 sg13g2_decap_8 FILLER_5_2629 ();
 sg13g2_decap_8 FILLER_5_2636 ();
 sg13g2_decap_8 FILLER_5_2643 ();
 sg13g2_decap_8 FILLER_5_2650 ();
 sg13g2_decap_8 FILLER_5_2657 ();
 sg13g2_decap_8 FILLER_5_2664 ();
 sg13g2_fill_2 FILLER_5_2671 ();
 sg13g2_fill_1 FILLER_5_2673 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_4 FILLER_6_483 ();
 sg13g2_fill_1 FILLER_6_487 ();
 sg13g2_fill_2 FILLER_6_519 ();
 sg13g2_fill_2 FILLER_6_573 ();
 sg13g2_fill_2 FILLER_6_605 ();
 sg13g2_fill_1 FILLER_6_607 ();
 sg13g2_fill_2 FILLER_6_617 ();
 sg13g2_fill_1 FILLER_6_704 ();
 sg13g2_fill_2 FILLER_6_766 ();
 sg13g2_fill_1 FILLER_6_834 ();
 sg13g2_fill_2 FILLER_6_980 ();
 sg13g2_fill_1 FILLER_6_986 ();
 sg13g2_fill_1 FILLER_6_997 ();
 sg13g2_fill_2 FILLER_6_1024 ();
 sg13g2_fill_2 FILLER_6_1040 ();
 sg13g2_fill_1 FILLER_6_1042 ();
 sg13g2_fill_1 FILLER_6_1064 ();
 sg13g2_fill_1 FILLER_6_1093 ();
 sg13g2_fill_1 FILLER_6_1108 ();
 sg13g2_fill_2 FILLER_6_1136 ();
 sg13g2_fill_1 FILLER_6_1178 ();
 sg13g2_fill_1 FILLER_6_1215 ();
 sg13g2_fill_2 FILLER_6_1225 ();
 sg13g2_fill_1 FILLER_6_1227 ();
 sg13g2_fill_1 FILLER_6_1258 ();
 sg13g2_fill_1 FILLER_6_1282 ();
 sg13g2_decap_8 FILLER_6_1331 ();
 sg13g2_fill_2 FILLER_6_1338 ();
 sg13g2_fill_2 FILLER_6_1344 ();
 sg13g2_fill_1 FILLER_6_1367 ();
 sg13g2_fill_1 FILLER_6_1399 ();
 sg13g2_fill_1 FILLER_6_1419 ();
 sg13g2_decap_8 FILLER_6_1471 ();
 sg13g2_decap_8 FILLER_6_1478 ();
 sg13g2_decap_8 FILLER_6_1485 ();
 sg13g2_decap_8 FILLER_6_1496 ();
 sg13g2_fill_2 FILLER_6_1508 ();
 sg13g2_fill_2 FILLER_6_1514 ();
 sg13g2_fill_1 FILLER_6_1516 ();
 sg13g2_fill_1 FILLER_6_1556 ();
 sg13g2_fill_1 FILLER_6_1592 ();
 sg13g2_fill_1 FILLER_6_1619 ();
 sg13g2_fill_2 FILLER_6_1667 ();
 sg13g2_fill_1 FILLER_6_1669 ();
 sg13g2_decap_8 FILLER_6_1696 ();
 sg13g2_decap_8 FILLER_6_1703 ();
 sg13g2_fill_2 FILLER_6_1710 ();
 sg13g2_fill_2 FILLER_6_1751 ();
 sg13g2_fill_1 FILLER_6_1779 ();
 sg13g2_fill_2 FILLER_6_1785 ();
 sg13g2_fill_1 FILLER_6_1787 ();
 sg13g2_fill_1 FILLER_6_1823 ();
 sg13g2_fill_2 FILLER_6_1847 ();
 sg13g2_fill_1 FILLER_6_1858 ();
 sg13g2_fill_2 FILLER_6_1863 ();
 sg13g2_fill_1 FILLER_6_1865 ();
 sg13g2_fill_1 FILLER_6_1913 ();
 sg13g2_fill_2 FILLER_6_1923 ();
 sg13g2_fill_1 FILLER_6_1939 ();
 sg13g2_fill_2 FILLER_6_2001 ();
 sg13g2_fill_1 FILLER_6_2003 ();
 sg13g2_fill_2 FILLER_6_2014 ();
 sg13g2_fill_1 FILLER_6_2016 ();
 sg13g2_fill_1 FILLER_6_2064 ();
 sg13g2_fill_1 FILLER_6_2085 ();
 sg13g2_fill_2 FILLER_6_2116 ();
 sg13g2_fill_1 FILLER_6_2118 ();
 sg13g2_decap_8 FILLER_6_2183 ();
 sg13g2_decap_4 FILLER_6_2190 ();
 sg13g2_fill_1 FILLER_6_2194 ();
 sg13g2_decap_4 FILLER_6_2203 ();
 sg13g2_fill_1 FILLER_6_2207 ();
 sg13g2_fill_2 FILLER_6_2214 ();
 sg13g2_fill_1 FILLER_6_2220 ();
 sg13g2_fill_1 FILLER_6_2227 ();
 sg13g2_fill_1 FILLER_6_2241 ();
 sg13g2_fill_1 FILLER_6_2246 ();
 sg13g2_fill_1 FILLER_6_2297 ();
 sg13g2_fill_2 FILLER_6_2379 ();
 sg13g2_fill_1 FILLER_6_2381 ();
 sg13g2_fill_2 FILLER_6_2414 ();
 sg13g2_fill_1 FILLER_6_2438 ();
 sg13g2_fill_2 FILLER_6_2470 ();
 sg13g2_decap_8 FILLER_6_2550 ();
 sg13g2_decap_8 FILLER_6_2557 ();
 sg13g2_decap_8 FILLER_6_2564 ();
 sg13g2_decap_8 FILLER_6_2571 ();
 sg13g2_decap_8 FILLER_6_2578 ();
 sg13g2_decap_8 FILLER_6_2585 ();
 sg13g2_decap_8 FILLER_6_2592 ();
 sg13g2_decap_8 FILLER_6_2599 ();
 sg13g2_decap_8 FILLER_6_2606 ();
 sg13g2_decap_8 FILLER_6_2613 ();
 sg13g2_decap_8 FILLER_6_2620 ();
 sg13g2_decap_8 FILLER_6_2627 ();
 sg13g2_decap_8 FILLER_6_2634 ();
 sg13g2_decap_8 FILLER_6_2641 ();
 sg13g2_decap_8 FILLER_6_2648 ();
 sg13g2_decap_8 FILLER_6_2655 ();
 sg13g2_decap_8 FILLER_6_2662 ();
 sg13g2_decap_4 FILLER_6_2669 ();
 sg13g2_fill_1 FILLER_6_2673 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_4 FILLER_7_483 ();
 sg13g2_fill_2 FILLER_7_570 ();
 sg13g2_fill_2 FILLER_7_577 ();
 sg13g2_fill_2 FILLER_7_610 ();
 sg13g2_fill_1 FILLER_7_612 ();
 sg13g2_fill_2 FILLER_7_622 ();
 sg13g2_fill_2 FILLER_7_650 ();
 sg13g2_fill_2 FILLER_7_709 ();
 sg13g2_fill_1 FILLER_7_711 ();
 sg13g2_fill_1 FILLER_7_760 ();
 sg13g2_fill_1 FILLER_7_839 ();
 sg13g2_fill_2 FILLER_7_849 ();
 sg13g2_fill_1 FILLER_7_885 ();
 sg13g2_fill_1 FILLER_7_938 ();
 sg13g2_fill_2 FILLER_7_965 ();
 sg13g2_fill_2 FILLER_7_1037 ();
 sg13g2_fill_1 FILLER_7_1065 ();
 sg13g2_fill_1 FILLER_7_1092 ();
 sg13g2_fill_2 FILLER_7_1117 ();
 sg13g2_fill_1 FILLER_7_1119 ();
 sg13g2_fill_2 FILLER_7_1158 ();
 sg13g2_fill_2 FILLER_7_1165 ();
 sg13g2_fill_1 FILLER_7_1232 ();
 sg13g2_fill_1 FILLER_7_1271 ();
 sg13g2_decap_4 FILLER_7_1284 ();
 sg13g2_fill_2 FILLER_7_1288 ();
 sg13g2_fill_1 FILLER_7_1299 ();
 sg13g2_fill_2 FILLER_7_1309 ();
 sg13g2_fill_1 FILLER_7_1311 ();
 sg13g2_decap_4 FILLER_7_1320 ();
 sg13g2_fill_1 FILLER_7_1324 ();
 sg13g2_fill_1 FILLER_7_1333 ();
 sg13g2_fill_2 FILLER_7_1369 ();
 sg13g2_fill_1 FILLER_7_1371 ();
 sg13g2_fill_2 FILLER_7_1407 ();
 sg13g2_decap_8 FILLER_7_1482 ();
 sg13g2_decap_4 FILLER_7_1489 ();
 sg13g2_fill_1 FILLER_7_1545 ();
 sg13g2_fill_2 FILLER_7_1559 ();
 sg13g2_fill_1 FILLER_7_1561 ();
 sg13g2_fill_2 FILLER_7_1618 ();
 sg13g2_fill_1 FILLER_7_1620 ();
 sg13g2_fill_1 FILLER_7_1630 ();
 sg13g2_fill_1 FILLER_7_1636 ();
 sg13g2_fill_1 FILLER_7_1664 ();
 sg13g2_fill_2 FILLER_7_1734 ();
 sg13g2_fill_1 FILLER_7_1736 ();
 sg13g2_fill_2 FILLER_7_1763 ();
 sg13g2_fill_1 FILLER_7_1765 ();
 sg13g2_fill_1 FILLER_7_1828 ();
 sg13g2_fill_2 FILLER_7_1883 ();
 sg13g2_fill_1 FILLER_7_1885 ();
 sg13g2_fill_1 FILLER_7_1944 ();
 sg13g2_fill_2 FILLER_7_1994 ();
 sg13g2_fill_2 FILLER_7_2009 ();
 sg13g2_fill_2 FILLER_7_2021 ();
 sg13g2_fill_1 FILLER_7_2023 ();
 sg13g2_fill_1 FILLER_7_2055 ();
 sg13g2_decap_8 FILLER_7_2090 ();
 sg13g2_fill_2 FILLER_7_2105 ();
 sg13g2_fill_1 FILLER_7_2116 ();
 sg13g2_fill_2 FILLER_7_2174 ();
 sg13g2_fill_1 FILLER_7_2176 ();
 sg13g2_fill_2 FILLER_7_2186 ();
 sg13g2_decap_4 FILLER_7_2209 ();
 sg13g2_fill_1 FILLER_7_2213 ();
 sg13g2_fill_2 FILLER_7_2223 ();
 sg13g2_fill_2 FILLER_7_2246 ();
 sg13g2_fill_1 FILLER_7_2248 ();
 sg13g2_fill_1 FILLER_7_2257 ();
 sg13g2_fill_2 FILLER_7_2266 ();
 sg13g2_fill_1 FILLER_7_2268 ();
 sg13g2_decap_4 FILLER_7_2277 ();
 sg13g2_fill_1 FILLER_7_2281 ();
 sg13g2_fill_2 FILLER_7_2399 ();
 sg13g2_fill_2 FILLER_7_2440 ();
 sg13g2_fill_1 FILLER_7_2442 ();
 sg13g2_fill_2 FILLER_7_2483 ();
 sg13g2_fill_1 FILLER_7_2485 ();
 sg13g2_decap_8 FILLER_7_2560 ();
 sg13g2_decap_8 FILLER_7_2567 ();
 sg13g2_decap_8 FILLER_7_2574 ();
 sg13g2_decap_8 FILLER_7_2581 ();
 sg13g2_decap_8 FILLER_7_2588 ();
 sg13g2_decap_8 FILLER_7_2595 ();
 sg13g2_decap_8 FILLER_7_2602 ();
 sg13g2_decap_8 FILLER_7_2609 ();
 sg13g2_decap_8 FILLER_7_2616 ();
 sg13g2_decap_8 FILLER_7_2623 ();
 sg13g2_decap_8 FILLER_7_2630 ();
 sg13g2_decap_8 FILLER_7_2637 ();
 sg13g2_decap_8 FILLER_7_2644 ();
 sg13g2_decap_8 FILLER_7_2651 ();
 sg13g2_decap_8 FILLER_7_2658 ();
 sg13g2_decap_8 FILLER_7_2665 ();
 sg13g2_fill_2 FILLER_7_2672 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_fill_1 FILLER_8_483 ();
 sg13g2_fill_1 FILLER_8_540 ();
 sg13g2_fill_2 FILLER_8_576 ();
 sg13g2_fill_1 FILLER_8_578 ();
 sg13g2_fill_1 FILLER_8_631 ();
 sg13g2_fill_1 FILLER_8_663 ();
 sg13g2_decap_4 FILLER_8_720 ();
 sg13g2_fill_2 FILLER_8_749 ();
 sg13g2_fill_1 FILLER_8_751 ();
 sg13g2_fill_1 FILLER_8_799 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_fill_2 FILLER_8_847 ();
 sg13g2_fill_1 FILLER_8_849 ();
 sg13g2_decap_8 FILLER_8_858 ();
 sg13g2_fill_1 FILLER_8_865 ();
 sg13g2_decap_4 FILLER_8_875 ();
 sg13g2_fill_2 FILLER_8_905 ();
 sg13g2_decap_8 FILLER_8_963 ();
 sg13g2_decap_8 FILLER_8_970 ();
 sg13g2_fill_1 FILLER_8_977 ();
 sg13g2_fill_1 FILLER_8_1025 ();
 sg13g2_decap_8 FILLER_8_1065 ();
 sg13g2_fill_1 FILLER_8_1072 ();
 sg13g2_decap_4 FILLER_8_1076 ();
 sg13g2_fill_1 FILLER_8_1080 ();
 sg13g2_fill_1 FILLER_8_1133 ();
 sg13g2_fill_2 FILLER_8_1169 ();
 sg13g2_fill_2 FILLER_8_1248 ();
 sg13g2_fill_1 FILLER_8_1250 ();
 sg13g2_decap_8 FILLER_8_1287 ();
 sg13g2_decap_8 FILLER_8_1294 ();
 sg13g2_fill_2 FILLER_8_1301 ();
 sg13g2_fill_2 FILLER_8_1312 ();
 sg13g2_fill_1 FILLER_8_1314 ();
 sg13g2_fill_2 FILLER_8_1325 ();
 sg13g2_fill_1 FILLER_8_1327 ();
 sg13g2_fill_1 FILLER_8_1439 ();
 sg13g2_fill_1 FILLER_8_1454 ();
 sg13g2_fill_2 FILLER_8_1498 ();
 sg13g2_fill_1 FILLER_8_1500 ();
 sg13g2_fill_2 FILLER_8_1510 ();
 sg13g2_fill_1 FILLER_8_1512 ();
 sg13g2_fill_1 FILLER_8_1548 ();
 sg13g2_decap_8 FILLER_8_1553 ();
 sg13g2_decap_8 FILLER_8_1560 ();
 sg13g2_fill_2 FILLER_8_1567 ();
 sg13g2_fill_1 FILLER_8_1569 ();
 sg13g2_fill_2 FILLER_8_1603 ();
 sg13g2_decap_8 FILLER_8_1620 ();
 sg13g2_decap_8 FILLER_8_1627 ();
 sg13g2_fill_2 FILLER_8_1634 ();
 sg13g2_decap_4 FILLER_8_1640 ();
 sg13g2_decap_4 FILLER_8_1648 ();
 sg13g2_fill_2 FILLER_8_1688 ();
 sg13g2_fill_1 FILLER_8_1696 ();
 sg13g2_fill_2 FILLER_8_1746 ();
 sg13g2_fill_2 FILLER_8_1854 ();
 sg13g2_fill_1 FILLER_8_1856 ();
 sg13g2_fill_2 FILLER_8_1876 ();
 sg13g2_fill_1 FILLER_8_1878 ();
 sg13g2_fill_2 FILLER_8_1893 ();
 sg13g2_fill_2 FILLER_8_1944 ();
 sg13g2_fill_2 FILLER_8_1977 ();
 sg13g2_fill_1 FILLER_8_1984 ();
 sg13g2_fill_2 FILLER_8_2082 ();
 sg13g2_fill_1 FILLER_8_2097 ();
 sg13g2_decap_4 FILLER_8_2102 ();
 sg13g2_fill_1 FILLER_8_2106 ();
 sg13g2_fill_1 FILLER_8_2209 ();
 sg13g2_fill_2 FILLER_8_2285 ();
 sg13g2_fill_2 FILLER_8_2291 ();
 sg13g2_fill_1 FILLER_8_2293 ();
 sg13g2_fill_1 FILLER_8_2299 ();
 sg13g2_fill_2 FILLER_8_2353 ();
 sg13g2_fill_2 FILLER_8_2461 ();
 sg13g2_fill_1 FILLER_8_2463 ();
 sg13g2_fill_2 FILLER_8_2485 ();
 sg13g2_fill_1 FILLER_8_2487 ();
 sg13g2_fill_2 FILLER_8_2512 ();
 sg13g2_fill_1 FILLER_8_2514 ();
 sg13g2_decap_8 FILLER_8_2549 ();
 sg13g2_decap_8 FILLER_8_2556 ();
 sg13g2_decap_8 FILLER_8_2563 ();
 sg13g2_decap_8 FILLER_8_2570 ();
 sg13g2_decap_8 FILLER_8_2577 ();
 sg13g2_decap_8 FILLER_8_2584 ();
 sg13g2_decap_8 FILLER_8_2591 ();
 sg13g2_decap_8 FILLER_8_2598 ();
 sg13g2_decap_8 FILLER_8_2605 ();
 sg13g2_decap_8 FILLER_8_2612 ();
 sg13g2_decap_8 FILLER_8_2619 ();
 sg13g2_decap_8 FILLER_8_2626 ();
 sg13g2_decap_8 FILLER_8_2633 ();
 sg13g2_decap_8 FILLER_8_2640 ();
 sg13g2_decap_8 FILLER_8_2647 ();
 sg13g2_decap_8 FILLER_8_2654 ();
 sg13g2_decap_8 FILLER_8_2661 ();
 sg13g2_decap_4 FILLER_8_2668 ();
 sg13g2_fill_2 FILLER_8_2672 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_4 FILLER_9_490 ();
 sg13g2_fill_1 FILLER_9_542 ();
 sg13g2_fill_2 FILLER_9_572 ();
 sg13g2_fill_2 FILLER_9_682 ();
 sg13g2_fill_1 FILLER_9_688 ();
 sg13g2_decap_8 FILLER_9_718 ();
 sg13g2_fill_2 FILLER_9_725 ();
 sg13g2_decap_8 FILLER_9_850 ();
 sg13g2_fill_1 FILLER_9_857 ();
 sg13g2_fill_2 FILLER_9_863 ();
 sg13g2_fill_1 FILLER_9_873 ();
 sg13g2_fill_1 FILLER_9_945 ();
 sg13g2_fill_1 FILLER_9_985 ();
 sg13g2_fill_1 FILLER_9_991 ();
 sg13g2_fill_1 FILLER_9_1015 ();
 sg13g2_fill_2 FILLER_9_1063 ();
 sg13g2_fill_2 FILLER_9_1083 ();
 sg13g2_fill_1 FILLER_9_1085 ();
 sg13g2_fill_2 FILLER_9_1125 ();
 sg13g2_fill_1 FILLER_9_1127 ();
 sg13g2_fill_2 FILLER_9_1158 ();
 sg13g2_fill_1 FILLER_9_1178 ();
 sg13g2_fill_1 FILLER_9_1188 ();
 sg13g2_fill_2 FILLER_9_1214 ();
 sg13g2_fill_1 FILLER_9_1216 ();
 sg13g2_decap_4 FILLER_9_1288 ();
 sg13g2_fill_1 FILLER_9_1292 ();
 sg13g2_fill_1 FILLER_9_1328 ();
 sg13g2_fill_2 FILLER_9_1402 ();
 sg13g2_fill_2 FILLER_9_1418 ();
 sg13g2_fill_1 FILLER_9_1420 ();
 sg13g2_fill_1 FILLER_9_1455 ();
 sg13g2_fill_1 FILLER_9_1461 ();
 sg13g2_decap_4 FILLER_9_1500 ();
 sg13g2_fill_1 FILLER_9_1504 ();
 sg13g2_fill_2 FILLER_9_1514 ();
 sg13g2_fill_1 FILLER_9_1516 ();
 sg13g2_fill_2 FILLER_9_1535 ();
 sg13g2_fill_2 FILLER_9_1584 ();
 sg13g2_fill_1 FILLER_9_1586 ();
 sg13g2_fill_1 FILLER_9_1606 ();
 sg13g2_fill_2 FILLER_9_1628 ();
 sg13g2_fill_1 FILLER_9_1630 ();
 sg13g2_decap_8 FILLER_9_1635 ();
 sg13g2_decap_4 FILLER_9_1642 ();
 sg13g2_fill_1 FILLER_9_1646 ();
 sg13g2_fill_2 FILLER_9_1669 ();
 sg13g2_fill_1 FILLER_9_1702 ();
 sg13g2_fill_2 FILLER_9_1756 ();
 sg13g2_fill_1 FILLER_9_1762 ();
 sg13g2_fill_2 FILLER_9_1768 ();
 sg13g2_fill_1 FILLER_9_1770 ();
 sg13g2_fill_2 FILLER_9_1793 ();
 sg13g2_fill_2 FILLER_9_1825 ();
 sg13g2_fill_2 FILLER_9_1835 ();
 sg13g2_fill_1 FILLER_9_1837 ();
 sg13g2_fill_1 FILLER_9_1853 ();
 sg13g2_fill_1 FILLER_9_1859 ();
 sg13g2_fill_2 FILLER_9_1904 ();
 sg13g2_fill_1 FILLER_9_1906 ();
 sg13g2_fill_1 FILLER_9_1985 ();
 sg13g2_fill_2 FILLER_9_2012 ();
 sg13g2_fill_2 FILLER_9_2044 ();
 sg13g2_fill_1 FILLER_9_2102 ();
 sg13g2_fill_2 FILLER_9_2156 ();
 sg13g2_fill_1 FILLER_9_2162 ();
 sg13g2_fill_2 FILLER_9_2246 ();
 sg13g2_fill_2 FILLER_9_2262 ();
 sg13g2_fill_2 FILLER_9_2308 ();
 sg13g2_decap_8 FILLER_9_2335 ();
 sg13g2_decap_8 FILLER_9_2342 ();
 sg13g2_fill_1 FILLER_9_2349 ();
 sg13g2_fill_1 FILLER_9_2393 ();
 sg13g2_decap_8 FILLER_9_2441 ();
 sg13g2_fill_1 FILLER_9_2448 ();
 sg13g2_decap_8 FILLER_9_2534 ();
 sg13g2_decap_8 FILLER_9_2541 ();
 sg13g2_decap_8 FILLER_9_2548 ();
 sg13g2_decap_8 FILLER_9_2555 ();
 sg13g2_decap_8 FILLER_9_2562 ();
 sg13g2_decap_8 FILLER_9_2569 ();
 sg13g2_decap_8 FILLER_9_2576 ();
 sg13g2_decap_8 FILLER_9_2583 ();
 sg13g2_decap_8 FILLER_9_2590 ();
 sg13g2_decap_8 FILLER_9_2597 ();
 sg13g2_decap_8 FILLER_9_2604 ();
 sg13g2_decap_8 FILLER_9_2611 ();
 sg13g2_decap_8 FILLER_9_2618 ();
 sg13g2_decap_8 FILLER_9_2625 ();
 sg13g2_decap_8 FILLER_9_2632 ();
 sg13g2_decap_8 FILLER_9_2639 ();
 sg13g2_decap_8 FILLER_9_2646 ();
 sg13g2_decap_8 FILLER_9_2653 ();
 sg13g2_decap_8 FILLER_9_2660 ();
 sg13g2_decap_8 FILLER_9_2667 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_fill_2 FILLER_10_483 ();
 sg13g2_fill_1 FILLER_10_521 ();
 sg13g2_fill_2 FILLER_10_601 ();
 sg13g2_fill_1 FILLER_10_603 ();
 sg13g2_fill_2 FILLER_10_613 ();
 sg13g2_fill_1 FILLER_10_629 ();
 sg13g2_fill_2 FILLER_10_639 ();
 sg13g2_fill_2 FILLER_10_653 ();
 sg13g2_fill_1 FILLER_10_672 ();
 sg13g2_fill_2 FILLER_10_689 ();
 sg13g2_fill_1 FILLER_10_691 ();
 sg13g2_decap_8 FILLER_10_709 ();
 sg13g2_decap_8 FILLER_10_716 ();
 sg13g2_fill_2 FILLER_10_723 ();
 sg13g2_fill_2 FILLER_10_751 ();
 sg13g2_fill_1 FILLER_10_753 ();
 sg13g2_fill_1 FILLER_10_805 ();
 sg13g2_fill_2 FILLER_10_815 ();
 sg13g2_fill_2 FILLER_10_851 ();
 sg13g2_decap_4 FILLER_10_858 ();
 sg13g2_fill_1 FILLER_10_862 ();
 sg13g2_fill_1 FILLER_10_987 ();
 sg13g2_fill_1 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1031 ();
 sg13g2_fill_1 FILLER_10_1061 ();
 sg13g2_decap_8 FILLER_10_1088 ();
 sg13g2_fill_1 FILLER_10_1095 ();
 sg13g2_decap_8 FILLER_10_1102 ();
 sg13g2_fill_2 FILLER_10_1125 ();
 sg13g2_fill_1 FILLER_10_1127 ();
 sg13g2_fill_1 FILLER_10_1133 ();
 sg13g2_fill_2 FILLER_10_1148 ();
 sg13g2_fill_1 FILLER_10_1150 ();
 sg13g2_decap_8 FILLER_10_1208 ();
 sg13g2_fill_2 FILLER_10_1215 ();
 sg13g2_fill_2 FILLER_10_1230 ();
 sg13g2_fill_1 FILLER_10_1232 ();
 sg13g2_fill_2 FILLER_10_1289 ();
 sg13g2_fill_1 FILLER_10_1291 ();
 sg13g2_decap_4 FILLER_10_1376 ();
 sg13g2_fill_2 FILLER_10_1445 ();
 sg13g2_fill_2 FILLER_10_1556 ();
 sg13g2_fill_2 FILLER_10_1610 ();
 sg13g2_fill_1 FILLER_10_1612 ();
 sg13g2_fill_2 FILLER_10_1707 ();
 sg13g2_fill_1 FILLER_10_1709 ();
 sg13g2_fill_2 FILLER_10_1744 ();
 sg13g2_fill_1 FILLER_10_1781 ();
 sg13g2_fill_2 FILLER_10_1817 ();
 sg13g2_fill_2 FILLER_10_1854 ();
 sg13g2_fill_1 FILLER_10_1856 ();
 sg13g2_fill_2 FILLER_10_1870 ();
 sg13g2_fill_1 FILLER_10_1910 ();
 sg13g2_fill_1 FILLER_10_1945 ();
 sg13g2_fill_2 FILLER_10_1960 ();
 sg13g2_fill_2 FILLER_10_2006 ();
 sg13g2_fill_1 FILLER_10_2008 ();
 sg13g2_fill_1 FILLER_10_2051 ();
 sg13g2_fill_1 FILLER_10_2090 ();
 sg13g2_fill_2 FILLER_10_2122 ();
 sg13g2_fill_1 FILLER_10_2133 ();
 sg13g2_fill_2 FILLER_10_2252 ();
 sg13g2_fill_2 FILLER_10_2259 ();
 sg13g2_fill_1 FILLER_10_2287 ();
 sg13g2_decap_8 FILLER_10_2340 ();
 sg13g2_decap_8 FILLER_10_2347 ();
 sg13g2_decap_4 FILLER_10_2354 ();
 sg13g2_fill_1 FILLER_10_2358 ();
 sg13g2_fill_2 FILLER_10_2369 ();
 sg13g2_fill_2 FILLER_10_2383 ();
 sg13g2_fill_1 FILLER_10_2385 ();
 sg13g2_fill_2 FILLER_10_2406 ();
 sg13g2_decap_4 FILLER_10_2429 ();
 sg13g2_fill_2 FILLER_10_2433 ();
 sg13g2_fill_2 FILLER_10_2461 ();
 sg13g2_fill_1 FILLER_10_2498 ();
 sg13g2_fill_1 FILLER_10_2543 ();
 sg13g2_fill_1 FILLER_10_2549 ();
 sg13g2_decap_8 FILLER_10_2571 ();
 sg13g2_decap_8 FILLER_10_2578 ();
 sg13g2_decap_8 FILLER_10_2585 ();
 sg13g2_decap_8 FILLER_10_2592 ();
 sg13g2_decap_8 FILLER_10_2599 ();
 sg13g2_decap_8 FILLER_10_2606 ();
 sg13g2_decap_8 FILLER_10_2613 ();
 sg13g2_decap_8 FILLER_10_2620 ();
 sg13g2_decap_8 FILLER_10_2627 ();
 sg13g2_decap_8 FILLER_10_2634 ();
 sg13g2_decap_8 FILLER_10_2641 ();
 sg13g2_decap_8 FILLER_10_2648 ();
 sg13g2_decap_8 FILLER_10_2655 ();
 sg13g2_decap_8 FILLER_10_2662 ();
 sg13g2_decap_4 FILLER_10_2669 ();
 sg13g2_fill_1 FILLER_10_2673 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_4 FILLER_11_476 ();
 sg13g2_fill_1 FILLER_11_480 ();
 sg13g2_fill_1 FILLER_11_542 ();
 sg13g2_fill_2 FILLER_11_583 ();
 sg13g2_fill_1 FILLER_11_620 ();
 sg13g2_fill_2 FILLER_11_636 ();
 sg13g2_fill_2 FILLER_11_666 ();
 sg13g2_fill_1 FILLER_11_668 ();
 sg13g2_fill_1 FILLER_11_711 ();
 sg13g2_fill_2 FILLER_11_720 ();
 sg13g2_fill_1 FILLER_11_757 ();
 sg13g2_fill_2 FILLER_11_778 ();
 sg13g2_fill_2 FILLER_11_842 ();
 sg13g2_fill_2 FILLER_11_857 ();
 sg13g2_decap_8 FILLER_11_867 ();
 sg13g2_fill_1 FILLER_11_874 ();
 sg13g2_fill_1 FILLER_11_901 ();
 sg13g2_decap_8 FILLER_11_936 ();
 sg13g2_fill_2 FILLER_11_943 ();
 sg13g2_fill_1 FILLER_11_988 ();
 sg13g2_fill_2 FILLER_11_1002 ();
 sg13g2_fill_1 FILLER_11_1004 ();
 sg13g2_fill_1 FILLER_11_1014 ();
 sg13g2_fill_2 FILLER_11_1109 ();
 sg13g2_fill_1 FILLER_11_1111 ();
 sg13g2_fill_1 FILLER_11_1121 ();
 sg13g2_fill_2 FILLER_11_1143 ();
 sg13g2_fill_2 FILLER_11_1184 ();
 sg13g2_decap_8 FILLER_11_1219 ();
 sg13g2_decap_8 FILLER_11_1280 ();
 sg13g2_decap_4 FILLER_11_1287 ();
 sg13g2_fill_1 FILLER_11_1326 ();
 sg13g2_decap_4 FILLER_11_1333 ();
 sg13g2_fill_1 FILLER_11_1341 ();
 sg13g2_fill_1 FILLER_11_1351 ();
 sg13g2_decap_8 FILLER_11_1406 ();
 sg13g2_fill_2 FILLER_11_1413 ();
 sg13g2_fill_1 FILLER_11_1415 ();
 sg13g2_decap_4 FILLER_11_1424 ();
 sg13g2_fill_2 FILLER_11_1428 ();
 sg13g2_fill_1 FILLER_11_1456 ();
 sg13g2_fill_2 FILLER_11_1488 ();
 sg13g2_fill_1 FILLER_11_1490 ();
 sg13g2_fill_1 FILLER_11_1504 ();
 sg13g2_fill_2 FILLER_11_1552 ();
 sg13g2_decap_4 FILLER_11_1558 ();
 sg13g2_fill_2 FILLER_11_1588 ();
 sg13g2_fill_1 FILLER_11_1616 ();
 sg13g2_fill_1 FILLER_11_1682 ();
 sg13g2_fill_1 FILLER_11_1710 ();
 sg13g2_fill_2 FILLER_11_1715 ();
 sg13g2_fill_1 FILLER_11_1717 ();
 sg13g2_fill_2 FILLER_11_1728 ();
 sg13g2_fill_2 FILLER_11_1782 ();
 sg13g2_fill_2 FILLER_11_1815 ();
 sg13g2_fill_1 FILLER_11_1817 ();
 sg13g2_fill_2 FILLER_11_1857 ();
 sg13g2_fill_1 FILLER_11_1944 ();
 sg13g2_decap_4 FILLER_11_1988 ();
 sg13g2_decap_8 FILLER_11_1996 ();
 sg13g2_fill_1 FILLER_11_2037 ();
 sg13g2_fill_2 FILLER_11_2074 ();
 sg13g2_fill_1 FILLER_11_2089 ();
 sg13g2_fill_2 FILLER_11_2095 ();
 sg13g2_fill_1 FILLER_11_2097 ();
 sg13g2_fill_2 FILLER_11_2107 ();
 sg13g2_fill_1 FILLER_11_2109 ();
 sg13g2_fill_1 FILLER_11_2173 ();
 sg13g2_fill_2 FILLER_11_2192 ();
 sg13g2_fill_2 FILLER_11_2207 ();
 sg13g2_fill_1 FILLER_11_2209 ();
 sg13g2_fill_1 FILLER_11_2233 ();
 sg13g2_fill_2 FILLER_11_2259 ();
 sg13g2_fill_1 FILLER_11_2261 ();
 sg13g2_fill_1 FILLER_11_2303 ();
 sg13g2_fill_2 FILLER_11_2343 ();
 sg13g2_fill_1 FILLER_11_2345 ();
 sg13g2_fill_2 FILLER_11_2385 ();
 sg13g2_fill_1 FILLER_11_2387 ();
 sg13g2_fill_2 FILLER_11_2396 ();
 sg13g2_fill_1 FILLER_11_2408 ();
 sg13g2_decap_8 FILLER_11_2426 ();
 sg13g2_fill_2 FILLER_11_2441 ();
 sg13g2_fill_1 FILLER_11_2443 ();
 sg13g2_fill_2 FILLER_11_2449 ();
 sg13g2_fill_1 FILLER_11_2451 ();
 sg13g2_decap_8 FILLER_11_2579 ();
 sg13g2_decap_8 FILLER_11_2586 ();
 sg13g2_decap_8 FILLER_11_2593 ();
 sg13g2_decap_8 FILLER_11_2600 ();
 sg13g2_decap_8 FILLER_11_2607 ();
 sg13g2_decap_8 FILLER_11_2614 ();
 sg13g2_decap_8 FILLER_11_2621 ();
 sg13g2_decap_8 FILLER_11_2628 ();
 sg13g2_decap_8 FILLER_11_2635 ();
 sg13g2_decap_8 FILLER_11_2642 ();
 sg13g2_decap_8 FILLER_11_2649 ();
 sg13g2_decap_8 FILLER_11_2656 ();
 sg13g2_decap_8 FILLER_11_2663 ();
 sg13g2_decap_4 FILLER_11_2670 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_fill_2 FILLER_12_476 ();
 sg13g2_fill_2 FILLER_12_534 ();
 sg13g2_fill_1 FILLER_12_536 ();
 sg13g2_fill_1 FILLER_12_542 ();
 sg13g2_fill_1 FILLER_12_578 ();
 sg13g2_fill_2 FILLER_12_623 ();
 sg13g2_fill_1 FILLER_12_625 ();
 sg13g2_fill_2 FILLER_12_635 ();
 sg13g2_fill_1 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_fill_2 FILLER_12_762 ();
 sg13g2_fill_1 FILLER_12_790 ();
 sg13g2_fill_2 FILLER_12_799 ();
 sg13g2_fill_2 FILLER_12_820 ();
 sg13g2_fill_1 FILLER_12_831 ();
 sg13g2_fill_2 FILLER_12_878 ();
 sg13g2_fill_2 FILLER_12_925 ();
 sg13g2_decap_8 FILLER_12_942 ();
 sg13g2_fill_1 FILLER_12_949 ();
 sg13g2_fill_2 FILLER_12_959 ();
 sg13g2_fill_1 FILLER_12_961 ();
 sg13g2_fill_1 FILLER_12_968 ();
 sg13g2_fill_2 FILLER_12_1025 ();
 sg13g2_fill_1 FILLER_12_1051 ();
 sg13g2_fill_2 FILLER_12_1112 ();
 sg13g2_fill_1 FILLER_12_1114 ();
 sg13g2_fill_2 FILLER_12_1141 ();
 sg13g2_fill_1 FILLER_12_1143 ();
 sg13g2_fill_1 FILLER_12_1174 ();
 sg13g2_fill_2 FILLER_12_1188 ();
 sg13g2_fill_2 FILLER_12_1195 ();
 sg13g2_fill_1 FILLER_12_1202 ();
 sg13g2_fill_2 FILLER_12_1251 ();
 sg13g2_fill_1 FILLER_12_1262 ();
 sg13g2_decap_8 FILLER_12_1289 ();
 sg13g2_fill_1 FILLER_12_1296 ();
 sg13g2_fill_1 FILLER_12_1332 ();
 sg13g2_decap_4 FILLER_12_1341 ();
 sg13g2_fill_1 FILLER_12_1345 ();
 sg13g2_fill_2 FILLER_12_1382 ();
 sg13g2_fill_1 FILLER_12_1384 ();
 sg13g2_fill_2 FILLER_12_1394 ();
 sg13g2_fill_1 FILLER_12_1396 ();
 sg13g2_fill_2 FILLER_12_1416 ();
 sg13g2_decap_4 FILLER_12_1499 ();
 sg13g2_fill_2 FILLER_12_1503 ();
 sg13g2_fill_1 FILLER_12_1518 ();
 sg13g2_fill_2 FILLER_12_1558 ();
 sg13g2_fill_1 FILLER_12_1560 ();
 sg13g2_fill_1 FILLER_12_1565 ();
 sg13g2_fill_2 FILLER_12_1606 ();
 sg13g2_fill_1 FILLER_12_1622 ();
 sg13g2_fill_2 FILLER_12_1649 ();
 sg13g2_fill_1 FILLER_12_1651 ();
 sg13g2_fill_2 FILLER_12_1670 ();
 sg13g2_fill_1 FILLER_12_1686 ();
 sg13g2_fill_2 FILLER_12_1717 ();
 sg13g2_fill_1 FILLER_12_1719 ();
 sg13g2_fill_2 FILLER_12_1725 ();
 sg13g2_fill_2 FILLER_12_1757 ();
 sg13g2_fill_1 FILLER_12_1785 ();
 sg13g2_fill_2 FILLER_12_1846 ();
 sg13g2_fill_2 FILLER_12_1870 ();
 sg13g2_fill_1 FILLER_12_1872 ();
 sg13g2_decap_8 FILLER_12_1908 ();
 sg13g2_fill_2 FILLER_12_1988 ();
 sg13g2_fill_1 FILLER_12_1990 ();
 sg13g2_fill_2 FILLER_12_2050 ();
 sg13g2_fill_2 FILLER_12_2057 ();
 sg13g2_fill_2 FILLER_12_2088 ();
 sg13g2_fill_1 FILLER_12_2090 ();
 sg13g2_fill_1 FILLER_12_2121 ();
 sg13g2_fill_1 FILLER_12_2127 ();
 sg13g2_fill_2 FILLER_12_2171 ();
 sg13g2_fill_2 FILLER_12_2221 ();
 sg13g2_fill_2 FILLER_12_2250 ();
 sg13g2_fill_2 FILLER_12_2261 ();
 sg13g2_fill_2 FILLER_12_2289 ();
 sg13g2_fill_1 FILLER_12_2291 ();
 sg13g2_fill_2 FILLER_12_2396 ();
 sg13g2_fill_2 FILLER_12_2454 ();
 sg13g2_fill_1 FILLER_12_2456 ();
 sg13g2_fill_2 FILLER_12_2501 ();
 sg13g2_decap_8 FILLER_12_2599 ();
 sg13g2_decap_8 FILLER_12_2606 ();
 sg13g2_decap_8 FILLER_12_2613 ();
 sg13g2_decap_8 FILLER_12_2620 ();
 sg13g2_decap_8 FILLER_12_2627 ();
 sg13g2_decap_8 FILLER_12_2634 ();
 sg13g2_decap_8 FILLER_12_2641 ();
 sg13g2_decap_8 FILLER_12_2648 ();
 sg13g2_decap_8 FILLER_12_2655 ();
 sg13g2_decap_8 FILLER_12_2662 ();
 sg13g2_decap_4 FILLER_12_2669 ();
 sg13g2_fill_1 FILLER_12_2673 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_4 FILLER_13_469 ();
 sg13g2_fill_2 FILLER_13_473 ();
 sg13g2_fill_1 FILLER_13_509 ();
 sg13g2_fill_2 FILLER_13_575 ();
 sg13g2_fill_1 FILLER_13_577 ();
 sg13g2_fill_1 FILLER_13_584 ();
 sg13g2_fill_1 FILLER_13_675 ();
 sg13g2_fill_1 FILLER_13_702 ();
 sg13g2_fill_1 FILLER_13_729 ();
 sg13g2_fill_2 FILLER_13_770 ();
 sg13g2_fill_1 FILLER_13_790 ();
 sg13g2_fill_2 FILLER_13_831 ();
 sg13g2_fill_2 FILLER_13_988 ();
 sg13g2_fill_1 FILLER_13_1010 ();
 sg13g2_fill_1 FILLER_13_1101 ();
 sg13g2_fill_1 FILLER_13_1116 ();
 sg13g2_fill_1 FILLER_13_1215 ();
 sg13g2_fill_2 FILLER_13_1256 ();
 sg13g2_decap_8 FILLER_13_1289 ();
 sg13g2_fill_2 FILLER_13_1378 ();
 sg13g2_fill_2 FILLER_13_1397 ();
 sg13g2_fill_2 FILLER_13_1407 ();
 sg13g2_fill_2 FILLER_13_1424 ();
 sg13g2_fill_1 FILLER_13_1426 ();
 sg13g2_fill_2 FILLER_13_1431 ();
 sg13g2_fill_2 FILLER_13_1459 ();
 sg13g2_fill_1 FILLER_13_1497 ();
 sg13g2_fill_1 FILLER_13_1553 ();
 sg13g2_fill_2 FILLER_13_1562 ();
 sg13g2_fill_1 FILLER_13_1564 ();
 sg13g2_fill_1 FILLER_13_1578 ();
 sg13g2_fill_2 FILLER_13_1584 ();
 sg13g2_fill_2 FILLER_13_1607 ();
 sg13g2_fill_1 FILLER_13_1609 ();
 sg13g2_fill_1 FILLER_13_1645 ();
 sg13g2_fill_1 FILLER_13_1711 ();
 sg13g2_fill_1 FILLER_13_1752 ();
 sg13g2_fill_2 FILLER_13_1770 ();
 sg13g2_fill_1 FILLER_13_1772 ();
 sg13g2_fill_2 FILLER_13_1792 ();
 sg13g2_fill_1 FILLER_13_1820 ();
 sg13g2_fill_1 FILLER_13_1825 ();
 sg13g2_fill_2 FILLER_13_1835 ();
 sg13g2_fill_1 FILLER_13_1837 ();
 sg13g2_fill_2 FILLER_13_1851 ();
 sg13g2_fill_1 FILLER_13_1858 ();
 sg13g2_fill_1 FILLER_13_1876 ();
 sg13g2_fill_1 FILLER_13_1882 ();
 sg13g2_fill_2 FILLER_13_1896 ();
 sg13g2_decap_8 FILLER_13_1907 ();
 sg13g2_fill_1 FILLER_13_1927 ();
 sg13g2_fill_2 FILLER_13_1933 ();
 sg13g2_fill_2 FILLER_13_1950 ();
 sg13g2_fill_2 FILLER_13_1978 ();
 sg13g2_fill_1 FILLER_13_1980 ();
 sg13g2_fill_1 FILLER_13_2033 ();
 sg13g2_fill_1 FILLER_13_2043 ();
 sg13g2_fill_2 FILLER_13_2074 ();
 sg13g2_fill_2 FILLER_13_2085 ();
 sg13g2_fill_2 FILLER_13_2128 ();
 sg13g2_fill_1 FILLER_13_2130 ();
 sg13g2_decap_8 FILLER_13_2158 ();
 sg13g2_fill_1 FILLER_13_2179 ();
 sg13g2_fill_2 FILLER_13_2206 ();
 sg13g2_fill_2 FILLER_13_2217 ();
 sg13g2_fill_1 FILLER_13_2219 ();
 sg13g2_fill_1 FILLER_13_2251 ();
 sg13g2_fill_2 FILLER_13_2265 ();
 sg13g2_fill_2 FILLER_13_2297 ();
 sg13g2_fill_1 FILLER_13_2299 ();
 sg13g2_fill_1 FILLER_13_2345 ();
 sg13g2_fill_2 FILLER_13_2387 ();
 sg13g2_fill_1 FILLER_13_2389 ();
 sg13g2_fill_1 FILLER_13_2395 ();
 sg13g2_fill_1 FILLER_13_2440 ();
 sg13g2_fill_1 FILLER_13_2461 ();
 sg13g2_fill_2 FILLER_13_2493 ();
 sg13g2_fill_1 FILLER_13_2495 ();
 sg13g2_fill_2 FILLER_13_2500 ();
 sg13g2_fill_1 FILLER_13_2502 ();
 sg13g2_decap_8 FILLER_13_2591 ();
 sg13g2_decap_8 FILLER_13_2598 ();
 sg13g2_decap_8 FILLER_13_2605 ();
 sg13g2_decap_8 FILLER_13_2612 ();
 sg13g2_decap_8 FILLER_13_2619 ();
 sg13g2_decap_8 FILLER_13_2626 ();
 sg13g2_decap_8 FILLER_13_2633 ();
 sg13g2_decap_8 FILLER_13_2640 ();
 sg13g2_decap_8 FILLER_13_2647 ();
 sg13g2_decap_8 FILLER_13_2654 ();
 sg13g2_decap_8 FILLER_13_2661 ();
 sg13g2_decap_4 FILLER_13_2668 ();
 sg13g2_fill_2 FILLER_13_2672 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_fill_1 FILLER_14_483 ();
 sg13g2_fill_1 FILLER_14_501 ();
 sg13g2_fill_1 FILLER_14_511 ();
 sg13g2_fill_2 FILLER_14_543 ();
 sg13g2_fill_2 FILLER_14_625 ();
 sg13g2_fill_1 FILLER_14_627 ();
 sg13g2_fill_1 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_737 ();
 sg13g2_fill_2 FILLER_14_744 ();
 sg13g2_fill_2 FILLER_14_750 ();
 sg13g2_fill_2 FILLER_14_940 ();
 sg13g2_fill_2 FILLER_14_1232 ();
 sg13g2_fill_2 FILLER_14_1254 ();
 sg13g2_decap_4 FILLER_14_1292 ();
 sg13g2_fill_2 FILLER_14_1296 ();
 sg13g2_fill_2 FILLER_14_1315 ();
 sg13g2_fill_1 FILLER_14_1317 ();
 sg13g2_fill_2 FILLER_14_1327 ();
 sg13g2_fill_1 FILLER_14_1329 ();
 sg13g2_fill_1 FILLER_14_1374 ();
 sg13g2_fill_2 FILLER_14_1396 ();
 sg13g2_fill_2 FILLER_14_1439 ();
 sg13g2_fill_1 FILLER_14_1441 ();
 sg13g2_fill_2 FILLER_14_1542 ();
 sg13g2_fill_1 FILLER_14_1583 ();
 sg13g2_fill_1 FILLER_14_1616 ();
 sg13g2_fill_2 FILLER_14_1634 ();
 sg13g2_fill_1 FILLER_14_1649 ();
 sg13g2_fill_2 FILLER_14_1654 ();
 sg13g2_fill_1 FILLER_14_1661 ();
 sg13g2_fill_2 FILLER_14_1722 ();
 sg13g2_fill_2 FILLER_14_1734 ();
 sg13g2_fill_2 FILLER_14_1766 ();
 sg13g2_fill_1 FILLER_14_1768 ();
 sg13g2_decap_4 FILLER_14_1829 ();
 sg13g2_decap_8 FILLER_14_1902 ();
 sg13g2_fill_1 FILLER_14_1935 ();
 sg13g2_fill_2 FILLER_14_1954 ();
 sg13g2_fill_1 FILLER_14_1956 ();
 sg13g2_fill_2 FILLER_14_2071 ();
 sg13g2_fill_2 FILLER_14_2104 ();
 sg13g2_fill_2 FILLER_14_2146 ();
 sg13g2_decap_4 FILLER_14_2152 ();
 sg13g2_fill_2 FILLER_14_2156 ();
 sg13g2_fill_2 FILLER_14_2210 ();
 sg13g2_decap_4 FILLER_14_2272 ();
 sg13g2_fill_2 FILLER_14_2276 ();
 sg13g2_fill_2 FILLER_14_2291 ();
 sg13g2_fill_1 FILLER_14_2307 ();
 sg13g2_fill_2 FILLER_14_2316 ();
 sg13g2_fill_2 FILLER_14_2347 ();
 sg13g2_fill_1 FILLER_14_2349 ();
 sg13g2_fill_2 FILLER_14_2354 ();
 sg13g2_fill_1 FILLER_14_2356 ();
 sg13g2_fill_2 FILLER_14_2436 ();
 sg13g2_fill_1 FILLER_14_2443 ();
 sg13g2_fill_2 FILLER_14_2458 ();
 sg13g2_fill_1 FILLER_14_2460 ();
 sg13g2_fill_2 FILLER_14_2471 ();
 sg13g2_fill_1 FILLER_14_2512 ();
 sg13g2_fill_2 FILLER_14_2521 ();
 sg13g2_fill_1 FILLER_14_2527 ();
 sg13g2_fill_2 FILLER_14_2544 ();
 sg13g2_fill_1 FILLER_14_2546 ();
 sg13g2_fill_1 FILLER_14_2570 ();
 sg13g2_decap_8 FILLER_14_2588 ();
 sg13g2_decap_8 FILLER_14_2595 ();
 sg13g2_decap_8 FILLER_14_2602 ();
 sg13g2_decap_8 FILLER_14_2609 ();
 sg13g2_decap_8 FILLER_14_2616 ();
 sg13g2_decap_8 FILLER_14_2623 ();
 sg13g2_decap_8 FILLER_14_2630 ();
 sg13g2_decap_8 FILLER_14_2637 ();
 sg13g2_decap_8 FILLER_14_2644 ();
 sg13g2_decap_8 FILLER_14_2651 ();
 sg13g2_decap_8 FILLER_14_2658 ();
 sg13g2_decap_8 FILLER_14_2665 ();
 sg13g2_fill_2 FILLER_14_2672 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_fill_1 FILLER_15_483 ();
 sg13g2_fill_2 FILLER_15_514 ();
 sg13g2_fill_1 FILLER_15_516 ();
 sg13g2_fill_2 FILLER_15_557 ();
 sg13g2_decap_8 FILLER_15_573 ();
 sg13g2_decap_4 FILLER_15_580 ();
 sg13g2_fill_2 FILLER_15_584 ();
 sg13g2_fill_2 FILLER_15_678 ();
 sg13g2_fill_2 FILLER_15_703 ();
 sg13g2_fill_1 FILLER_15_705 ();
 sg13g2_fill_1 FILLER_15_710 ();
 sg13g2_fill_2 FILLER_15_720 ();
 sg13g2_fill_1 FILLER_15_722 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_decap_4 FILLER_15_751 ();
 sg13g2_fill_2 FILLER_15_755 ();
 sg13g2_fill_2 FILLER_15_786 ();
 sg13g2_fill_1 FILLER_15_817 ();
 sg13g2_fill_2 FILLER_15_844 ();
 sg13g2_fill_2 FILLER_15_863 ();
 sg13g2_fill_1 FILLER_15_865 ();
 sg13g2_fill_1 FILLER_15_896 ();
 sg13g2_decap_4 FILLER_15_906 ();
 sg13g2_fill_1 FILLER_15_910 ();
 sg13g2_fill_2 FILLER_15_926 ();
 sg13g2_fill_1 FILLER_15_984 ();
 sg13g2_fill_2 FILLER_15_993 ();
 sg13g2_fill_1 FILLER_15_995 ();
 sg13g2_fill_2 FILLER_15_1004 ();
 sg13g2_fill_1 FILLER_15_1006 ();
 sg13g2_fill_1 FILLER_15_1017 ();
 sg13g2_fill_2 FILLER_15_1057 ();
 sg13g2_fill_1 FILLER_15_1181 ();
 sg13g2_fill_2 FILLER_15_1227 ();
 sg13g2_fill_1 FILLER_15_1239 ();
 sg13g2_decap_8 FILLER_15_1285 ();
 sg13g2_fill_2 FILLER_15_1292 ();
 sg13g2_fill_1 FILLER_15_1395 ();
 sg13g2_fill_2 FILLER_15_1414 ();
 sg13g2_decap_8 FILLER_15_1443 ();
 sg13g2_fill_1 FILLER_15_1474 ();
 sg13g2_fill_2 FILLER_15_1506 ();
 sg13g2_fill_2 FILLER_15_1542 ();
 sg13g2_fill_2 FILLER_15_1634 ();
 sg13g2_fill_1 FILLER_15_1636 ();
 sg13g2_fill_2 FILLER_15_1658 ();
 sg13g2_fill_1 FILLER_15_1701 ();
 sg13g2_fill_2 FILLER_15_1731 ();
 sg13g2_fill_2 FILLER_15_1794 ();
 sg13g2_fill_1 FILLER_15_1796 ();
 sg13g2_fill_1 FILLER_15_1806 ();
 sg13g2_fill_1 FILLER_15_1813 ();
 sg13g2_decap_8 FILLER_15_1892 ();
 sg13g2_fill_1 FILLER_15_1899 ();
 sg13g2_fill_1 FILLER_15_1951 ();
 sg13g2_fill_1 FILLER_15_1991 ();
 sg13g2_fill_1 FILLER_15_1997 ();
 sg13g2_decap_8 FILLER_15_2024 ();
 sg13g2_decap_8 FILLER_15_2035 ();
 sg13g2_fill_2 FILLER_15_2042 ();
 sg13g2_fill_2 FILLER_15_2146 ();
 sg13g2_fill_1 FILLER_15_2148 ();
 sg13g2_fill_2 FILLER_15_2165 ();
 sg13g2_decap_8 FILLER_15_2279 ();
 sg13g2_fill_2 FILLER_15_2286 ();
 sg13g2_decap_4 FILLER_15_2293 ();
 sg13g2_fill_1 FILLER_15_2297 ();
 sg13g2_fill_2 FILLER_15_2308 ();
 sg13g2_fill_1 FILLER_15_2310 ();
 sg13g2_decap_8 FILLER_15_2328 ();
 sg13g2_decap_8 FILLER_15_2335 ();
 sg13g2_decap_8 FILLER_15_2342 ();
 sg13g2_decap_8 FILLER_15_2349 ();
 sg13g2_fill_1 FILLER_15_2396 ();
 sg13g2_fill_2 FILLER_15_2402 ();
 sg13g2_fill_1 FILLER_15_2404 ();
 sg13g2_fill_1 FILLER_15_2430 ();
 sg13g2_fill_2 FILLER_15_2488 ();
 sg13g2_fill_1 FILLER_15_2503 ();
 sg13g2_fill_2 FILLER_15_2521 ();
 sg13g2_fill_1 FILLER_15_2523 ();
 sg13g2_fill_2 FILLER_15_2529 ();
 sg13g2_fill_1 FILLER_15_2531 ();
 sg13g2_fill_1 FILLER_15_2537 ();
 sg13g2_decap_8 FILLER_15_2581 ();
 sg13g2_decap_8 FILLER_15_2588 ();
 sg13g2_decap_8 FILLER_15_2595 ();
 sg13g2_decap_8 FILLER_15_2602 ();
 sg13g2_decap_8 FILLER_15_2609 ();
 sg13g2_decap_8 FILLER_15_2616 ();
 sg13g2_decap_8 FILLER_15_2623 ();
 sg13g2_decap_8 FILLER_15_2630 ();
 sg13g2_decap_8 FILLER_15_2637 ();
 sg13g2_decap_8 FILLER_15_2644 ();
 sg13g2_decap_8 FILLER_15_2651 ();
 sg13g2_decap_8 FILLER_15_2658 ();
 sg13g2_decap_8 FILLER_15_2665 ();
 sg13g2_fill_2 FILLER_15_2672 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_4 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_579 ();
 sg13g2_fill_2 FILLER_16_586 ();
 sg13g2_fill_1 FILLER_16_588 ();
 sg13g2_fill_2 FILLER_16_598 ();
 sg13g2_fill_1 FILLER_16_609 ();
 sg13g2_fill_2 FILLER_16_648 ();
 sg13g2_fill_1 FILLER_16_655 ();
 sg13g2_fill_1 FILLER_16_673 ();
 sg13g2_decap_8 FILLER_16_729 ();
 sg13g2_fill_2 FILLER_16_736 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_decap_4 FILLER_16_760 ();
 sg13g2_fill_1 FILLER_16_764 ();
 sg13g2_fill_2 FILLER_16_811 ();
 sg13g2_fill_2 FILLER_16_821 ();
 sg13g2_fill_2 FILLER_16_827 ();
 sg13g2_fill_2 FILLER_16_833 ();
 sg13g2_fill_2 FILLER_16_886 ();
 sg13g2_fill_1 FILLER_16_888 ();
 sg13g2_fill_2 FILLER_16_903 ();
 sg13g2_fill_1 FILLER_16_915 ();
 sg13g2_decap_8 FILLER_16_926 ();
 sg13g2_fill_2 FILLER_16_933 ();
 sg13g2_fill_1 FILLER_16_935 ();
 sg13g2_decap_4 FILLER_16_941 ();
 sg13g2_fill_1 FILLER_16_945 ();
 sg13g2_fill_2 FILLER_16_986 ();
 sg13g2_fill_2 FILLER_16_1031 ();
 sg13g2_fill_1 FILLER_16_1033 ();
 sg13g2_decap_8 FILLER_16_1049 ();
 sg13g2_decap_4 FILLER_16_1056 ();
 sg13g2_fill_2 FILLER_16_1060 ();
 sg13g2_decap_8 FILLER_16_1066 ();
 sg13g2_decap_4 FILLER_16_1090 ();
 sg13g2_fill_2 FILLER_16_1094 ();
 sg13g2_fill_1 FILLER_16_1100 ();
 sg13g2_fill_1 FILLER_16_1149 ();
 sg13g2_fill_2 FILLER_16_1158 ();
 sg13g2_fill_2 FILLER_16_1185 ();
 sg13g2_decap_4 FILLER_16_1195 ();
 sg13g2_decap_4 FILLER_16_1207 ();
 sg13g2_fill_1 FILLER_16_1211 ();
 sg13g2_fill_2 FILLER_16_1221 ();
 sg13g2_fill_1 FILLER_16_1223 ();
 sg13g2_decap_8 FILLER_16_1285 ();
 sg13g2_decap_4 FILLER_16_1292 ();
 sg13g2_fill_1 FILLER_16_1296 ();
 sg13g2_fill_2 FILLER_16_1323 ();
 sg13g2_fill_1 FILLER_16_1325 ();
 sg13g2_fill_2 FILLER_16_1352 ();
 sg13g2_fill_2 FILLER_16_1504 ();
 sg13g2_fill_2 FILLER_16_1532 ();
 sg13g2_fill_1 FILLER_16_1534 ();
 sg13g2_fill_2 FILLER_16_1556 ();
 sg13g2_fill_2 FILLER_16_1571 ();
 sg13g2_fill_2 FILLER_16_1682 ();
 sg13g2_fill_1 FILLER_16_1684 ();
 sg13g2_fill_2 FILLER_16_1703 ();
 sg13g2_fill_2 FILLER_16_1735 ();
 sg13g2_fill_1 FILLER_16_1737 ();
 sg13g2_fill_2 FILLER_16_1772 ();
 sg13g2_decap_8 FILLER_16_1824 ();
 sg13g2_fill_2 FILLER_16_1831 ();
 sg13g2_fill_1 FILLER_16_1833 ();
 sg13g2_fill_2 FILLER_16_1842 ();
 sg13g2_fill_1 FILLER_16_1844 ();
 sg13g2_fill_2 FILLER_16_1871 ();
 sg13g2_fill_2 FILLER_16_1878 ();
 sg13g2_fill_1 FILLER_16_1880 ();
 sg13g2_decap_4 FILLER_16_1903 ();
 sg13g2_fill_2 FILLER_16_1981 ();
 sg13g2_fill_2 FILLER_16_2032 ();
 sg13g2_fill_2 FILLER_16_2045 ();
 sg13g2_fill_1 FILLER_16_2052 ();
 sg13g2_fill_2 FILLER_16_2069 ();
 sg13g2_fill_1 FILLER_16_2084 ();
 sg13g2_fill_2 FILLER_16_2098 ();
 sg13g2_fill_2 FILLER_16_2209 ();
 sg13g2_fill_1 FILLER_16_2211 ();
 sg13g2_fill_2 FILLER_16_2237 ();
 sg13g2_decap_8 FILLER_16_2272 ();
 sg13g2_decap_8 FILLER_16_2279 ();
 sg13g2_decap_4 FILLER_16_2286 ();
 sg13g2_fill_2 FILLER_16_2330 ();
 sg13g2_fill_2 FILLER_16_2378 ();
 sg13g2_fill_2 FILLER_16_2499 ();
 sg13g2_fill_1 FILLER_16_2536 ();
 sg13g2_decap_8 FILLER_16_2581 ();
 sg13g2_decap_8 FILLER_16_2588 ();
 sg13g2_decap_8 FILLER_16_2595 ();
 sg13g2_decap_8 FILLER_16_2602 ();
 sg13g2_decap_8 FILLER_16_2609 ();
 sg13g2_decap_8 FILLER_16_2616 ();
 sg13g2_decap_8 FILLER_16_2623 ();
 sg13g2_decap_8 FILLER_16_2630 ();
 sg13g2_decap_8 FILLER_16_2637 ();
 sg13g2_decap_8 FILLER_16_2644 ();
 sg13g2_decap_8 FILLER_16_2651 ();
 sg13g2_decap_8 FILLER_16_2658 ();
 sg13g2_decap_8 FILLER_16_2665 ();
 sg13g2_fill_2 FILLER_16_2672 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_fill_2 FILLER_17_483 ();
 sg13g2_fill_1 FILLER_17_485 ();
 sg13g2_fill_2 FILLER_17_564 ();
 sg13g2_fill_2 FILLER_17_571 ();
 sg13g2_fill_1 FILLER_17_613 ();
 sg13g2_decap_8 FILLER_17_745 ();
 sg13g2_decap_8 FILLER_17_752 ();
 sg13g2_fill_1 FILLER_17_759 ();
 sg13g2_fill_1 FILLER_17_786 ();
 sg13g2_fill_2 FILLER_17_796 ();
 sg13g2_fill_1 FILLER_17_798 ();
 sg13g2_fill_1 FILLER_17_839 ();
 sg13g2_decap_8 FILLER_17_869 ();
 sg13g2_fill_2 FILLER_17_876 ();
 sg13g2_fill_2 FILLER_17_886 ();
 sg13g2_fill_1 FILLER_17_888 ();
 sg13g2_fill_1 FILLER_17_911 ();
 sg13g2_decap_8 FILLER_17_918 ();
 sg13g2_fill_2 FILLER_17_925 ();
 sg13g2_fill_2 FILLER_17_939 ();
 sg13g2_decap_8 FILLER_17_1029 ();
 sg13g2_fill_2 FILLER_17_1044 ();
 sg13g2_fill_2 FILLER_17_1055 ();
 sg13g2_fill_1 FILLER_17_1057 ();
 sg13g2_decap_8 FILLER_17_1063 ();
 sg13g2_decap_4 FILLER_17_1074 ();
 sg13g2_fill_2 FILLER_17_1078 ();
 sg13g2_decap_8 FILLER_17_1084 ();
 sg13g2_decap_8 FILLER_17_1091 ();
 sg13g2_fill_2 FILLER_17_1102 ();
 sg13g2_fill_2 FILLER_17_1125 ();
 sg13g2_fill_2 FILLER_17_1136 ();
 sg13g2_fill_1 FILLER_17_1163 ();
 sg13g2_fill_2 FILLER_17_1216 ();
 sg13g2_fill_2 FILLER_17_1248 ();
 sg13g2_decap_8 FILLER_17_1285 ();
 sg13g2_decap_4 FILLER_17_1292 ();
 sg13g2_fill_1 FILLER_17_1296 ();
 sg13g2_decap_4 FILLER_17_1329 ();
 sg13g2_fill_2 FILLER_17_1347 ();
 sg13g2_fill_1 FILLER_17_1349 ();
 sg13g2_fill_2 FILLER_17_1355 ();
 sg13g2_fill_1 FILLER_17_1357 ();
 sg13g2_fill_1 FILLER_17_1362 ();
 sg13g2_fill_2 FILLER_17_1389 ();
 sg13g2_fill_2 FILLER_17_1427 ();
 sg13g2_fill_2 FILLER_17_1459 ();
 sg13g2_fill_2 FILLER_17_1531 ();
 sg13g2_fill_1 FILLER_17_1533 ();
 sg13g2_fill_2 FILLER_17_1569 ();
 sg13g2_fill_2 FILLER_17_1595 ();
 sg13g2_fill_1 FILLER_17_1597 ();
 sg13g2_fill_1 FILLER_17_1607 ();
 sg13g2_fill_2 FILLER_17_1617 ();
 sg13g2_fill_2 FILLER_17_1654 ();
 sg13g2_fill_1 FILLER_17_1656 ();
 sg13g2_fill_2 FILLER_17_1725 ();
 sg13g2_fill_1 FILLER_17_1727 ();
 sg13g2_fill_1 FILLER_17_1749 ();
 sg13g2_fill_2 FILLER_17_1772 ();
 sg13g2_fill_1 FILLER_17_1821 ();
 sg13g2_fill_2 FILLER_17_1835 ();
 sg13g2_fill_1 FILLER_17_1837 ();
 sg13g2_fill_2 FILLER_17_1846 ();
 sg13g2_fill_2 FILLER_17_1875 ();
 sg13g2_fill_2 FILLER_17_1907 ();
 sg13g2_fill_2 FILLER_17_1921 ();
 sg13g2_fill_2 FILLER_17_1936 ();
 sg13g2_fill_1 FILLER_17_1938 ();
 sg13g2_fill_2 FILLER_17_1980 ();
 sg13g2_fill_2 FILLER_17_2102 ();
 sg13g2_fill_1 FILLER_17_2135 ();
 sg13g2_fill_2 FILLER_17_2158 ();
 sg13g2_fill_1 FILLER_17_2160 ();
 sg13g2_fill_1 FILLER_17_2200 ();
 sg13g2_decap_8 FILLER_17_2205 ();
 sg13g2_decap_8 FILLER_17_2212 ();
 sg13g2_fill_2 FILLER_17_2219 ();
 sg13g2_fill_1 FILLER_17_2221 ();
 sg13g2_decap_8 FILLER_17_2226 ();
 sg13g2_fill_2 FILLER_17_2254 ();
 sg13g2_fill_1 FILLER_17_2256 ();
 sg13g2_fill_2 FILLER_17_2283 ();
 sg13g2_fill_1 FILLER_17_2285 ();
 sg13g2_fill_2 FILLER_17_2312 ();
 sg13g2_fill_1 FILLER_17_2314 ();
 sg13g2_fill_1 FILLER_17_2371 ();
 sg13g2_fill_2 FILLER_17_2389 ();
 sg13g2_decap_4 FILLER_17_2399 ();
 sg13g2_decap_4 FILLER_17_2456 ();
 sg13g2_fill_2 FILLER_17_2464 ();
 sg13g2_fill_1 FILLER_17_2466 ();
 sg13g2_fill_2 FILLER_17_2524 ();
 sg13g2_fill_2 FILLER_17_2530 ();
 sg13g2_fill_1 FILLER_17_2532 ();
 sg13g2_decap_8 FILLER_17_2598 ();
 sg13g2_decap_8 FILLER_17_2605 ();
 sg13g2_decap_8 FILLER_17_2612 ();
 sg13g2_decap_8 FILLER_17_2619 ();
 sg13g2_decap_8 FILLER_17_2626 ();
 sg13g2_decap_8 FILLER_17_2633 ();
 sg13g2_decap_8 FILLER_17_2640 ();
 sg13g2_decap_8 FILLER_17_2647 ();
 sg13g2_decap_8 FILLER_17_2654 ();
 sg13g2_decap_8 FILLER_17_2661 ();
 sg13g2_decap_4 FILLER_17_2668 ();
 sg13g2_fill_2 FILLER_17_2672 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_4 FILLER_18_483 ();
 sg13g2_fill_1 FILLER_18_487 ();
 sg13g2_fill_2 FILLER_18_533 ();
 sg13g2_fill_2 FILLER_18_548 ();
 sg13g2_fill_2 FILLER_18_568 ();
 sg13g2_fill_2 FILLER_18_605 ();
 sg13g2_fill_2 FILLER_18_652 ();
 sg13g2_fill_1 FILLER_18_654 ();
 sg13g2_fill_1 FILLER_18_660 ();
 sg13g2_fill_2 FILLER_18_710 ();
 sg13g2_fill_1 FILLER_18_809 ();
 sg13g2_fill_2 FILLER_18_869 ();
 sg13g2_fill_2 FILLER_18_885 ();
 sg13g2_fill_1 FILLER_18_929 ();
 sg13g2_decap_8 FILLER_18_1043 ();
 sg13g2_decap_4 FILLER_18_1050 ();
 sg13g2_fill_1 FILLER_18_1073 ();
 sg13g2_fill_2 FILLER_18_1079 ();
 sg13g2_fill_1 FILLER_18_1081 ();
 sg13g2_fill_1 FILLER_18_1247 ();
 sg13g2_decap_4 FILLER_18_1291 ();
 sg13g2_fill_1 FILLER_18_1295 ();
 sg13g2_decap_8 FILLER_18_1335 ();
 sg13g2_fill_1 FILLER_18_1373 ();
 sg13g2_fill_2 FILLER_18_1425 ();
 sg13g2_fill_1 FILLER_18_1489 ();
 sg13g2_fill_1 FILLER_18_1507 ();
 sg13g2_fill_2 FILLER_18_1513 ();
 sg13g2_fill_1 FILLER_18_1515 ();
 sg13g2_fill_2 FILLER_18_1521 ();
 sg13g2_fill_2 FILLER_18_1529 ();
 sg13g2_fill_2 FILLER_18_1621 ();
 sg13g2_fill_2 FILLER_18_1657 ();
 sg13g2_fill_1 FILLER_18_1659 ();
 sg13g2_fill_2 FILLER_18_1712 ();
 sg13g2_fill_1 FILLER_18_1714 ();
 sg13g2_fill_2 FILLER_18_1741 ();
 sg13g2_fill_2 FILLER_18_1768 ();
 sg13g2_fill_1 FILLER_18_1770 ();
 sg13g2_fill_2 FILLER_18_1797 ();
 sg13g2_fill_1 FILLER_18_1799 ();
 sg13g2_decap_4 FILLER_18_1806 ();
 sg13g2_fill_1 FILLER_18_1810 ();
 sg13g2_fill_2 FILLER_18_1867 ();
 sg13g2_fill_2 FILLER_18_1953 ();
 sg13g2_fill_1 FILLER_18_1955 ();
 sg13g2_fill_1 FILLER_18_1974 ();
 sg13g2_fill_2 FILLER_18_2001 ();
 sg13g2_fill_1 FILLER_18_2003 ();
 sg13g2_fill_2 FILLER_18_2013 ();
 sg13g2_fill_1 FILLER_18_2111 ();
 sg13g2_fill_2 FILLER_18_2150 ();
 sg13g2_fill_1 FILLER_18_2152 ();
 sg13g2_fill_2 FILLER_18_2200 ();
 sg13g2_fill_2 FILLER_18_2224 ();
 sg13g2_fill_1 FILLER_18_2294 ();
 sg13g2_fill_2 FILLER_18_2331 ();
 sg13g2_fill_1 FILLER_18_2333 ();
 sg13g2_decap_4 FILLER_18_2386 ();
 sg13g2_decap_8 FILLER_18_2396 ();
 sg13g2_decap_4 FILLER_18_2403 ();
 sg13g2_fill_2 FILLER_18_2452 ();
 sg13g2_fill_1 FILLER_18_2454 ();
 sg13g2_decap_4 FILLER_18_2472 ();
 sg13g2_fill_1 FILLER_18_2545 ();
 sg13g2_fill_2 FILLER_18_2584 ();
 sg13g2_decap_8 FILLER_18_2595 ();
 sg13g2_decap_8 FILLER_18_2602 ();
 sg13g2_decap_8 FILLER_18_2609 ();
 sg13g2_decap_8 FILLER_18_2616 ();
 sg13g2_decap_8 FILLER_18_2623 ();
 sg13g2_decap_8 FILLER_18_2630 ();
 sg13g2_decap_8 FILLER_18_2637 ();
 sg13g2_decap_8 FILLER_18_2644 ();
 sg13g2_decap_8 FILLER_18_2651 ();
 sg13g2_decap_8 FILLER_18_2658 ();
 sg13g2_decap_8 FILLER_18_2665 ();
 sg13g2_fill_2 FILLER_18_2672 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_fill_2 FILLER_19_533 ();
 sg13g2_fill_1 FILLER_19_535 ();
 sg13g2_decap_4 FILLER_19_540 ();
 sg13g2_fill_1 FILLER_19_544 ();
 sg13g2_fill_2 FILLER_19_549 ();
 sg13g2_fill_1 FILLER_19_551 ();
 sg13g2_fill_1 FILLER_19_569 ();
 sg13g2_decap_4 FILLER_19_612 ();
 sg13g2_fill_1 FILLER_19_616 ();
 sg13g2_fill_1 FILLER_19_622 ();
 sg13g2_fill_1 FILLER_19_632 ();
 sg13g2_fill_2 FILLER_19_651 ();
 sg13g2_fill_1 FILLER_19_764 ();
 sg13g2_fill_1 FILLER_19_788 ();
 sg13g2_fill_1 FILLER_19_875 ();
 sg13g2_fill_2 FILLER_19_928 ();
 sg13g2_fill_2 FILLER_19_956 ();
 sg13g2_fill_1 FILLER_19_958 ();
 sg13g2_fill_1 FILLER_19_1011 ();
 sg13g2_fill_2 FILLER_19_1046 ();
 sg13g2_fill_2 FILLER_19_1078 ();
 sg13g2_fill_1 FILLER_19_1080 ();
 sg13g2_fill_2 FILLER_19_1142 ();
 sg13g2_fill_1 FILLER_19_1144 ();
 sg13g2_fill_1 FILLER_19_1150 ();
 sg13g2_fill_1 FILLER_19_1174 ();
 sg13g2_fill_2 FILLER_19_1242 ();
 sg13g2_fill_1 FILLER_19_1287 ();
 sg13g2_decap_8 FILLER_19_1333 ();
 sg13g2_decap_8 FILLER_19_1340 ();
 sg13g2_decap_4 FILLER_19_1347 ();
 sg13g2_fill_2 FILLER_19_1351 ();
 sg13g2_fill_2 FILLER_19_1362 ();
 sg13g2_decap_4 FILLER_19_1398 ();
 sg13g2_fill_1 FILLER_19_1402 ();
 sg13g2_fill_2 FILLER_19_1441 ();
 sg13g2_fill_1 FILLER_19_1504 ();
 sg13g2_fill_1 FILLER_19_1510 ();
 sg13g2_fill_2 FILLER_19_1516 ();
 sg13g2_fill_1 FILLER_19_1518 ();
 sg13g2_fill_1 FILLER_19_1534 ();
 sg13g2_fill_2 FILLER_19_1545 ();
 sg13g2_fill_1 FILLER_19_1547 ();
 sg13g2_fill_2 FILLER_19_1578 ();
 sg13g2_fill_1 FILLER_19_1580 ();
 sg13g2_fill_2 FILLER_19_1621 ();
 sg13g2_fill_1 FILLER_19_1662 ();
 sg13g2_fill_2 FILLER_19_1671 ();
 sg13g2_fill_2 FILLER_19_1698 ();
 sg13g2_fill_1 FILLER_19_1757 ();
 sg13g2_fill_1 FILLER_19_1796 ();
 sg13g2_decap_8 FILLER_19_1912 ();
 sg13g2_decap_4 FILLER_19_1919 ();
 sg13g2_decap_4 FILLER_19_1926 ();
 sg13g2_fill_2 FILLER_19_1930 ();
 sg13g2_fill_2 FILLER_19_1984 ();
 sg13g2_decap_4 FILLER_19_2020 ();
 sg13g2_fill_2 FILLER_19_2024 ();
 sg13g2_decap_4 FILLER_19_2031 ();
 sg13g2_fill_2 FILLER_19_2039 ();
 sg13g2_fill_1 FILLER_19_2041 ();
 sg13g2_fill_1 FILLER_19_2081 ();
 sg13g2_fill_1 FILLER_19_2173 ();
 sg13g2_decap_4 FILLER_19_2200 ();
 sg13g2_decap_4 FILLER_19_2214 ();
 sg13g2_fill_1 FILLER_19_2218 ();
 sg13g2_fill_1 FILLER_19_2275 ();
 sg13g2_fill_1 FILLER_19_2305 ();
 sg13g2_decap_4 FILLER_19_2332 ();
 sg13g2_fill_2 FILLER_19_2372 ();
 sg13g2_fill_1 FILLER_19_2374 ();
 sg13g2_fill_2 FILLER_19_2384 ();
 sg13g2_fill_1 FILLER_19_2402 ();
 sg13g2_fill_2 FILLER_19_2443 ();
 sg13g2_fill_1 FILLER_19_2445 ();
 sg13g2_fill_2 FILLER_19_2530 ();
 sg13g2_fill_1 FILLER_19_2548 ();
 sg13g2_decap_8 FILLER_19_2579 ();
 sg13g2_decap_8 FILLER_19_2586 ();
 sg13g2_decap_8 FILLER_19_2593 ();
 sg13g2_decap_8 FILLER_19_2600 ();
 sg13g2_decap_8 FILLER_19_2607 ();
 sg13g2_decap_8 FILLER_19_2614 ();
 sg13g2_decap_8 FILLER_19_2621 ();
 sg13g2_decap_8 FILLER_19_2628 ();
 sg13g2_decap_8 FILLER_19_2635 ();
 sg13g2_decap_8 FILLER_19_2642 ();
 sg13g2_decap_8 FILLER_19_2649 ();
 sg13g2_decap_8 FILLER_19_2656 ();
 sg13g2_decap_8 FILLER_19_2663 ();
 sg13g2_decap_4 FILLER_19_2670 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_fill_2 FILLER_20_490 ();
 sg13g2_fill_2 FILLER_20_519 ();
 sg13g2_decap_8 FILLER_20_556 ();
 sg13g2_fill_1 FILLER_20_563 ();
 sg13g2_fill_2 FILLER_20_590 ();
 sg13g2_fill_1 FILLER_20_592 ();
 sg13g2_fill_2 FILLER_20_642 ();
 sg13g2_decap_8 FILLER_20_660 ();
 sg13g2_fill_1 FILLER_20_667 ();
 sg13g2_fill_2 FILLER_20_676 ();
 sg13g2_fill_2 FILLER_20_704 ();
 sg13g2_fill_1 FILLER_20_777 ();
 sg13g2_fill_1 FILLER_20_787 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_decap_4 FILLER_20_799 ();
 sg13g2_decap_8 FILLER_20_807 ();
 sg13g2_decap_8 FILLER_20_814 ();
 sg13g2_fill_2 FILLER_20_821 ();
 sg13g2_fill_2 FILLER_20_841 ();
 sg13g2_fill_2 FILLER_20_857 ();
 sg13g2_fill_1 FILLER_20_864 ();
 sg13g2_fill_1 FILLER_20_927 ();
 sg13g2_fill_1 FILLER_20_969 ();
 sg13g2_fill_2 FILLER_20_1000 ();
 sg13g2_fill_2 FILLER_20_1109 ();
 sg13g2_fill_1 FILLER_20_1116 ();
 sg13g2_fill_2 FILLER_20_1155 ();
 sg13g2_fill_2 FILLER_20_1292 ();
 sg13g2_fill_1 FILLER_20_1294 ();
 sg13g2_decap_8 FILLER_20_1340 ();
 sg13g2_fill_2 FILLER_20_1347 ();
 sg13g2_fill_1 FILLER_20_1349 ();
 sg13g2_fill_1 FILLER_20_1376 ();
 sg13g2_fill_1 FILLER_20_1395 ();
 sg13g2_fill_2 FILLER_20_1496 ();
 sg13g2_fill_1 FILLER_20_1524 ();
 sg13g2_fill_2 FILLER_20_1560 ();
 sg13g2_fill_2 FILLER_20_1578 ();
 sg13g2_fill_1 FILLER_20_1594 ();
 sg13g2_decap_4 FILLER_20_1598 ();
 sg13g2_fill_1 FILLER_20_1636 ();
 sg13g2_fill_1 FILLER_20_1693 ();
 sg13g2_fill_2 FILLER_20_1708 ();
 sg13g2_fill_2 FILLER_20_1740 ();
 sg13g2_fill_1 FILLER_20_1742 ();
 sg13g2_fill_2 FILLER_20_1778 ();
 sg13g2_fill_1 FILLER_20_1780 ();
 sg13g2_fill_2 FILLER_20_1790 ();
 sg13g2_fill_1 FILLER_20_1792 ();
 sg13g2_decap_8 FILLER_20_1850 ();
 sg13g2_fill_1 FILLER_20_1857 ();
 sg13g2_decap_8 FILLER_20_1927 ();
 sg13g2_fill_1 FILLER_20_1934 ();
 sg13g2_fill_2 FILLER_20_1940 ();
 sg13g2_fill_1 FILLER_20_1942 ();
 sg13g2_fill_2 FILLER_20_1982 ();
 sg13g2_decap_4 FILLER_20_2033 ();
 sg13g2_fill_1 FILLER_20_2037 ();
 sg13g2_fill_2 FILLER_20_2043 ();
 sg13g2_fill_1 FILLER_20_2045 ();
 sg13g2_fill_1 FILLER_20_2064 ();
 sg13g2_fill_2 FILLER_20_2073 ();
 sg13g2_fill_1 FILLER_20_2075 ();
 sg13g2_fill_2 FILLER_20_2086 ();
 sg13g2_fill_1 FILLER_20_2114 ();
 sg13g2_fill_2 FILLER_20_2193 ();
 sg13g2_fill_1 FILLER_20_2195 ();
 sg13g2_fill_2 FILLER_20_2240 ();
 sg13g2_fill_1 FILLER_20_2242 ();
 sg13g2_fill_2 FILLER_20_2285 ();
 sg13g2_fill_1 FILLER_20_2304 ();
 sg13g2_fill_1 FILLER_20_2314 ();
 sg13g2_fill_2 FILLER_20_2332 ();
 sg13g2_fill_1 FILLER_20_2334 ();
 sg13g2_fill_2 FILLER_20_2343 ();
 sg13g2_fill_2 FILLER_20_2353 ();
 sg13g2_fill_1 FILLER_20_2369 ();
 sg13g2_fill_2 FILLER_20_2379 ();
 sg13g2_fill_1 FILLER_20_2386 ();
 sg13g2_fill_2 FILLER_20_2401 ();
 sg13g2_fill_1 FILLER_20_2427 ();
 sg13g2_fill_2 FILLER_20_2492 ();
 sg13g2_fill_1 FILLER_20_2494 ();
 sg13g2_fill_1 FILLER_20_2500 ();
 sg13g2_fill_1 FILLER_20_2531 ();
 sg13g2_fill_1 FILLER_20_2558 ();
 sg13g2_decap_8 FILLER_20_2589 ();
 sg13g2_decap_8 FILLER_20_2596 ();
 sg13g2_decap_8 FILLER_20_2603 ();
 sg13g2_decap_8 FILLER_20_2610 ();
 sg13g2_decap_8 FILLER_20_2617 ();
 sg13g2_decap_8 FILLER_20_2624 ();
 sg13g2_decap_8 FILLER_20_2631 ();
 sg13g2_decap_8 FILLER_20_2638 ();
 sg13g2_decap_8 FILLER_20_2645 ();
 sg13g2_decap_8 FILLER_20_2652 ();
 sg13g2_decap_8 FILLER_20_2659 ();
 sg13g2_decap_8 FILLER_20_2666 ();
 sg13g2_fill_1 FILLER_20_2673 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_fill_2 FILLER_21_483 ();
 sg13g2_fill_1 FILLER_21_572 ();
 sg13g2_fill_1 FILLER_21_603 ();
 sg13g2_fill_1 FILLER_21_644 ();
 sg13g2_fill_2 FILLER_21_650 ();
 sg13g2_decap_8 FILLER_21_660 ();
 sg13g2_decap_4 FILLER_21_667 ();
 sg13g2_fill_2 FILLER_21_671 ();
 sg13g2_fill_2 FILLER_21_729 ();
 sg13g2_fill_2 FILLER_21_774 ();
 sg13g2_fill_1 FILLER_21_776 ();
 sg13g2_fill_1 FILLER_21_791 ();
 sg13g2_fill_2 FILLER_21_800 ();
 sg13g2_fill_1 FILLER_21_812 ();
 sg13g2_decap_4 FILLER_21_822 ();
 sg13g2_fill_2 FILLER_21_826 ();
 sg13g2_decap_4 FILLER_21_832 ();
 sg13g2_fill_1 FILLER_21_836 ();
 sg13g2_fill_2 FILLER_21_846 ();
 sg13g2_decap_4 FILLER_21_865 ();
 sg13g2_fill_2 FILLER_21_873 ();
 sg13g2_fill_1 FILLER_21_896 ();
 sg13g2_fill_2 FILLER_21_919 ();
 sg13g2_fill_1 FILLER_21_926 ();
 sg13g2_fill_1 FILLER_21_970 ();
 sg13g2_decap_4 FILLER_21_1041 ();
 sg13g2_fill_2 FILLER_21_1045 ();
 sg13g2_fill_2 FILLER_21_1073 ();
 sg13g2_fill_1 FILLER_21_1084 ();
 sg13g2_fill_2 FILLER_21_1090 ();
 sg13g2_fill_1 FILLER_21_1149 ();
 sg13g2_fill_1 FILLER_21_1185 ();
 sg13g2_fill_2 FILLER_21_1218 ();
 sg13g2_fill_2 FILLER_21_1232 ();
 sg13g2_decap_8 FILLER_21_1282 ();
 sg13g2_fill_2 FILLER_21_1289 ();
 sg13g2_fill_1 FILLER_21_1291 ();
 sg13g2_fill_1 FILLER_21_1334 ();
 sg13g2_fill_2 FILLER_21_1343 ();
 sg13g2_fill_1 FILLER_21_1345 ();
 sg13g2_fill_1 FILLER_21_1377 ();
 sg13g2_fill_1 FILLER_21_1388 ();
 sg13g2_fill_1 FILLER_21_1424 ();
 sg13g2_fill_2 FILLER_21_1447 ();
 sg13g2_fill_2 FILLER_21_1457 ();
 sg13g2_fill_1 FILLER_21_1499 ();
 sg13g2_fill_1 FILLER_21_1566 ();
 sg13g2_fill_1 FILLER_21_1577 ();
 sg13g2_fill_2 FILLER_21_1600 ();
 sg13g2_fill_2 FILLER_21_1690 ();
 sg13g2_fill_1 FILLER_21_1692 ();
 sg13g2_fill_2 FILLER_21_1707 ();
 sg13g2_fill_1 FILLER_21_1709 ();
 sg13g2_fill_1 FILLER_21_1736 ();
 sg13g2_decap_8 FILLER_21_1794 ();
 sg13g2_fill_2 FILLER_21_1801 ();
 sg13g2_fill_1 FILLER_21_1803 ();
 sg13g2_fill_1 FILLER_21_1812 ();
 sg13g2_fill_2 FILLER_21_1828 ();
 sg13g2_fill_1 FILLER_21_1865 ();
 sg13g2_fill_2 FILLER_21_1871 ();
 sg13g2_fill_2 FILLER_21_1881 ();
 sg13g2_fill_2 FILLER_21_1892 ();
 sg13g2_fill_1 FILLER_21_1894 ();
 sg13g2_fill_2 FILLER_21_1939 ();
 sg13g2_fill_1 FILLER_21_1941 ();
 sg13g2_decap_4 FILLER_21_2035 ();
 sg13g2_fill_1 FILLER_21_2098 ();
 sg13g2_fill_2 FILLER_21_2107 ();
 sg13g2_fill_1 FILLER_21_2131 ();
 sg13g2_decap_8 FILLER_21_2141 ();
 sg13g2_decap_8 FILLER_21_2148 ();
 sg13g2_fill_2 FILLER_21_2155 ();
 sg13g2_fill_1 FILLER_21_2157 ();
 sg13g2_fill_1 FILLER_21_2163 ();
 sg13g2_fill_1 FILLER_21_2181 ();
 sg13g2_decap_4 FILLER_21_2191 ();
 sg13g2_fill_2 FILLER_21_2204 ();
 sg13g2_fill_1 FILLER_21_2206 ();
 sg13g2_fill_1 FILLER_21_2220 ();
 sg13g2_fill_2 FILLER_21_2234 ();
 sg13g2_fill_2 FILLER_21_2240 ();
 sg13g2_fill_1 FILLER_21_2242 ();
 sg13g2_fill_1 FILLER_21_2257 ();
 sg13g2_fill_2 FILLER_21_2271 ();
 sg13g2_fill_2 FILLER_21_2299 ();
 sg13g2_fill_1 FILLER_21_2301 ();
 sg13g2_fill_1 FILLER_21_2306 ();
 sg13g2_fill_1 FILLER_21_2329 ();
 sg13g2_fill_2 FILLER_21_2396 ();
 sg13g2_fill_1 FILLER_21_2398 ();
 sg13g2_fill_1 FILLER_21_2443 ();
 sg13g2_fill_1 FILLER_21_2449 ();
 sg13g2_fill_2 FILLER_21_2490 ();
 sg13g2_fill_1 FILLER_21_2492 ();
 sg13g2_fill_1 FILLER_21_2522 ();
 sg13g2_fill_2 FILLER_21_2527 ();
 sg13g2_fill_1 FILLER_21_2555 ();
 sg13g2_decap_8 FILLER_21_2599 ();
 sg13g2_decap_8 FILLER_21_2606 ();
 sg13g2_decap_8 FILLER_21_2613 ();
 sg13g2_decap_8 FILLER_21_2620 ();
 sg13g2_decap_8 FILLER_21_2627 ();
 sg13g2_decap_8 FILLER_21_2634 ();
 sg13g2_decap_8 FILLER_21_2641 ();
 sg13g2_decap_8 FILLER_21_2648 ();
 sg13g2_decap_8 FILLER_21_2655 ();
 sg13g2_decap_8 FILLER_21_2662 ();
 sg13g2_decap_4 FILLER_21_2669 ();
 sg13g2_fill_1 FILLER_21_2673 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_4 FILLER_22_476 ();
 sg13g2_fill_2 FILLER_22_480 ();
 sg13g2_fill_2 FILLER_22_521 ();
 sg13g2_fill_2 FILLER_22_554 ();
 sg13g2_fill_1 FILLER_22_570 ();
 sg13g2_fill_2 FILLER_22_593 ();
 sg13g2_fill_2 FILLER_22_608 ();
 sg13g2_fill_1 FILLER_22_610 ();
 sg13g2_fill_2 FILLER_22_620 ();
 sg13g2_fill_1 FILLER_22_622 ();
 sg13g2_fill_1 FILLER_22_637 ();
 sg13g2_fill_2 FILLER_22_695 ();
 sg13g2_fill_1 FILLER_22_697 ();
 sg13g2_fill_2 FILLER_22_724 ();
 sg13g2_fill_1 FILLER_22_734 ();
 sg13g2_fill_2 FILLER_22_784 ();
 sg13g2_fill_1 FILLER_22_811 ();
 sg13g2_fill_2 FILLER_22_817 ();
 sg13g2_fill_2 FILLER_22_878 ();
 sg13g2_fill_2 FILLER_22_889 ();
 sg13g2_decap_4 FILLER_22_1032 ();
 sg13g2_fill_2 FILLER_22_1036 ();
 sg13g2_fill_1 FILLER_22_1079 ();
 sg13g2_fill_2 FILLER_22_1085 ();
 sg13g2_fill_1 FILLER_22_1087 ();
 sg13g2_fill_2 FILLER_22_1131 ();
 sg13g2_fill_1 FILLER_22_1133 ();
 sg13g2_fill_2 FILLER_22_1144 ();
 sg13g2_fill_2 FILLER_22_1206 ();
 sg13g2_fill_1 FILLER_22_1239 ();
 sg13g2_fill_2 FILLER_22_1254 ();
 sg13g2_decap_4 FILLER_22_1288 ();
 sg13g2_fill_1 FILLER_22_1330 ();
 sg13g2_fill_2 FILLER_22_1345 ();
 sg13g2_fill_2 FILLER_22_1353 ();
 sg13g2_fill_1 FILLER_22_1355 ();
 sg13g2_fill_1 FILLER_22_1404 ();
 sg13g2_fill_1 FILLER_22_1413 ();
 sg13g2_fill_2 FILLER_22_1502 ();
 sg13g2_fill_1 FILLER_22_1504 ();
 sg13g2_fill_2 FILLER_22_1510 ();
 sg13g2_decap_8 FILLER_22_1547 ();
 sg13g2_decap_8 FILLER_22_1554 ();
 sg13g2_fill_1 FILLER_22_1561 ();
 sg13g2_fill_1 FILLER_22_1567 ();
 sg13g2_fill_1 FILLER_22_1636 ();
 sg13g2_fill_1 FILLER_22_1671 ();
 sg13g2_fill_1 FILLER_22_1744 ();
 sg13g2_fill_2 FILLER_22_1758 ();
 sg13g2_fill_2 FILLER_22_1770 ();
 sg13g2_fill_1 FILLER_22_1782 ();
 sg13g2_decap_8 FILLER_22_1796 ();
 sg13g2_fill_1 FILLER_22_1803 ();
 sg13g2_fill_1 FILLER_22_1821 ();
 sg13g2_fill_1 FILLER_22_1878 ();
 sg13g2_fill_1 FILLER_22_1894 ();
 sg13g2_decap_8 FILLER_22_1935 ();
 sg13g2_decap_4 FILLER_22_1942 ();
 sg13g2_fill_2 FILLER_22_1972 ();
 sg13g2_fill_1 FILLER_22_1974 ();
 sg13g2_fill_1 FILLER_22_2066 ();
 sg13g2_decap_4 FILLER_22_2098 ();
 sg13g2_fill_1 FILLER_22_2102 ();
 sg13g2_fill_2 FILLER_22_2111 ();
 sg13g2_fill_1 FILLER_22_2113 ();
 sg13g2_fill_2 FILLER_22_2128 ();
 sg13g2_fill_1 FILLER_22_2134 ();
 sg13g2_decap_8 FILLER_22_2139 ();
 sg13g2_decap_4 FILLER_22_2146 ();
 sg13g2_decap_4 FILLER_22_2180 ();
 sg13g2_fill_1 FILLER_22_2184 ();
 sg13g2_decap_4 FILLER_22_2202 ();
 sg13g2_decap_8 FILLER_22_2223 ();
 sg13g2_decap_8 FILLER_22_2230 ();
 sg13g2_fill_2 FILLER_22_2237 ();
 sg13g2_fill_1 FILLER_22_2239 ();
 sg13g2_fill_2 FILLER_22_2245 ();
 sg13g2_fill_1 FILLER_22_2247 ();
 sg13g2_fill_1 FILLER_22_2258 ();
 sg13g2_fill_2 FILLER_22_2306 ();
 sg13g2_fill_1 FILLER_22_2308 ();
 sg13g2_fill_2 FILLER_22_2343 ();
 sg13g2_fill_2 FILLER_22_2371 ();
 sg13g2_fill_2 FILLER_22_2439 ();
 sg13g2_fill_1 FILLER_22_2441 ();
 sg13g2_fill_1 FILLER_22_2491 ();
 sg13g2_fill_2 FILLER_22_2500 ();
 sg13g2_fill_2 FILLER_22_2507 ();
 sg13g2_fill_1 FILLER_22_2509 ();
 sg13g2_fill_2 FILLER_22_2519 ();
 sg13g2_fill_1 FILLER_22_2521 ();
 sg13g2_fill_2 FILLER_22_2558 ();
 sg13g2_decap_8 FILLER_22_2604 ();
 sg13g2_decap_8 FILLER_22_2611 ();
 sg13g2_decap_8 FILLER_22_2618 ();
 sg13g2_decap_8 FILLER_22_2625 ();
 sg13g2_decap_8 FILLER_22_2632 ();
 sg13g2_decap_8 FILLER_22_2639 ();
 sg13g2_decap_8 FILLER_22_2646 ();
 sg13g2_decap_8 FILLER_22_2653 ();
 sg13g2_decap_8 FILLER_22_2660 ();
 sg13g2_decap_8 FILLER_22_2667 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_4 FILLER_23_476 ();
 sg13g2_fill_2 FILLER_23_480 ();
 sg13g2_fill_1 FILLER_23_543 ();
 sg13g2_fill_2 FILLER_23_598 ();
 sg13g2_fill_1 FILLER_23_600 ();
 sg13g2_fill_2 FILLER_23_617 ();
 sg13g2_fill_1 FILLER_23_619 ();
 sg13g2_fill_2 FILLER_23_625 ();
 sg13g2_fill_2 FILLER_23_641 ();
 sg13g2_fill_2 FILLER_23_684 ();
 sg13g2_fill_1 FILLER_23_686 ();
 sg13g2_fill_1 FILLER_23_702 ();
 sg13g2_fill_2 FILLER_23_738 ();
 sg13g2_decap_8 FILLER_23_766 ();
 sg13g2_fill_1 FILLER_23_773 ();
 sg13g2_fill_2 FILLER_23_810 ();
 sg13g2_fill_1 FILLER_23_856 ();
 sg13g2_fill_1 FILLER_23_883 ();
 sg13g2_fill_2 FILLER_23_916 ();
 sg13g2_fill_1 FILLER_23_924 ();
 sg13g2_fill_1 FILLER_23_954 ();
 sg13g2_fill_1 FILLER_23_964 ();
 sg13g2_fill_2 FILLER_23_989 ();
 sg13g2_decap_8 FILLER_23_1028 ();
 sg13g2_decap_4 FILLER_23_1035 ();
 sg13g2_fill_2 FILLER_23_1039 ();
 sg13g2_fill_1 FILLER_23_1049 ();
 sg13g2_fill_2 FILLER_23_1063 ();
 sg13g2_fill_1 FILLER_23_1065 ();
 sg13g2_fill_2 FILLER_23_1071 ();
 sg13g2_fill_1 FILLER_23_1078 ();
 sg13g2_fill_2 FILLER_23_1096 ();
 sg13g2_fill_2 FILLER_23_1128 ();
 sg13g2_fill_1 FILLER_23_1130 ();
 sg13g2_fill_2 FILLER_23_1145 ();
 sg13g2_fill_1 FILLER_23_1147 ();
 sg13g2_fill_1 FILLER_23_1156 ();
 sg13g2_fill_2 FILLER_23_1180 ();
 sg13g2_fill_2 FILLER_23_1196 ();
 sg13g2_fill_1 FILLER_23_1240 ();
 sg13g2_fill_1 FILLER_23_1274 ();
 sg13g2_decap_4 FILLER_23_1284 ();
 sg13g2_fill_1 FILLER_23_1294 ();
 sg13g2_fill_2 FILLER_23_1298 ();
 sg13g2_fill_1 FILLER_23_1300 ();
 sg13g2_fill_1 FILLER_23_1331 ();
 sg13g2_fill_1 FILLER_23_1341 ();
 sg13g2_fill_2 FILLER_23_1373 ();
 sg13g2_fill_1 FILLER_23_1385 ();
 sg13g2_fill_1 FILLER_23_1407 ();
 sg13g2_fill_1 FILLER_23_1416 ();
 sg13g2_decap_8 FILLER_23_1430 ();
 sg13g2_fill_2 FILLER_23_1462 ();
 sg13g2_fill_2 FILLER_23_1468 ();
 sg13g2_fill_1 FILLER_23_1474 ();
 sg13g2_decap_8 FILLER_23_1488 ();
 sg13g2_decap_4 FILLER_23_1495 ();
 sg13g2_fill_2 FILLER_23_1516 ();
 sg13g2_fill_1 FILLER_23_1518 ();
 sg13g2_fill_2 FILLER_23_1544 ();
 sg13g2_fill_1 FILLER_23_1546 ();
 sg13g2_decap_4 FILLER_23_1599 ();
 sg13g2_fill_2 FILLER_23_1608 ();
 sg13g2_fill_1 FILLER_23_1620 ();
 sg13g2_fill_1 FILLER_23_1642 ();
 sg13g2_fill_2 FILLER_23_1657 ();
 sg13g2_fill_2 FILLER_23_1688 ();
 sg13g2_fill_1 FILLER_23_1690 ();
 sg13g2_fill_2 FILLER_23_1749 ();
 sg13g2_fill_1 FILLER_23_1751 ();
 sg13g2_fill_2 FILLER_23_1760 ();
 sg13g2_fill_2 FILLER_23_1771 ();
 sg13g2_fill_1 FILLER_23_1773 ();
 sg13g2_decap_8 FILLER_23_1791 ();
 sg13g2_decap_8 FILLER_23_1798 ();
 sg13g2_decap_8 FILLER_23_1805 ();
 sg13g2_fill_2 FILLER_23_1817 ();
 sg13g2_fill_2 FILLER_23_1824 ();
 sg13g2_fill_1 FILLER_23_1826 ();
 sg13g2_decap_8 FILLER_23_1836 ();
 sg13g2_decap_8 FILLER_23_1843 ();
 sg13g2_decap_4 FILLER_23_1850 ();
 sg13g2_fill_2 FILLER_23_1854 ();
 sg13g2_fill_2 FILLER_23_1861 ();
 sg13g2_fill_1 FILLER_23_1863 ();
 sg13g2_fill_2 FILLER_23_1873 ();
 sg13g2_fill_1 FILLER_23_1875 ();
 sg13g2_fill_2 FILLER_23_1902 ();
 sg13g2_fill_1 FILLER_23_1904 ();
 sg13g2_decap_4 FILLER_23_1985 ();
 sg13g2_fill_1 FILLER_23_1989 ();
 sg13g2_fill_2 FILLER_23_2004 ();
 sg13g2_fill_1 FILLER_23_2006 ();
 sg13g2_fill_2 FILLER_23_2015 ();
 sg13g2_fill_1 FILLER_23_2029 ();
 sg13g2_fill_2 FILLER_23_2056 ();
 sg13g2_fill_1 FILLER_23_2058 ();
 sg13g2_fill_1 FILLER_23_2080 ();
 sg13g2_fill_2 FILLER_23_2091 ();
 sg13g2_fill_2 FILLER_23_2102 ();
 sg13g2_fill_2 FILLER_23_2141 ();
 sg13g2_fill_2 FILLER_23_2191 ();
 sg13g2_fill_1 FILLER_23_2232 ();
 sg13g2_fill_2 FILLER_23_2362 ();
 sg13g2_decap_8 FILLER_23_2490 ();
 sg13g2_decap_8 FILLER_23_2497 ();
 sg13g2_fill_1 FILLER_23_2504 ();
 sg13g2_fill_2 FILLER_23_2547 ();
 sg13g2_fill_2 FILLER_23_2563 ();
 sg13g2_decap_8 FILLER_23_2595 ();
 sg13g2_decap_8 FILLER_23_2602 ();
 sg13g2_decap_8 FILLER_23_2609 ();
 sg13g2_decap_8 FILLER_23_2616 ();
 sg13g2_decap_8 FILLER_23_2623 ();
 sg13g2_decap_8 FILLER_23_2630 ();
 sg13g2_decap_8 FILLER_23_2637 ();
 sg13g2_decap_8 FILLER_23_2644 ();
 sg13g2_decap_8 FILLER_23_2651 ();
 sg13g2_decap_8 FILLER_23_2658 ();
 sg13g2_decap_8 FILLER_23_2665 ();
 sg13g2_fill_2 FILLER_23_2672 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_fill_1 FILLER_24_490 ();
 sg13g2_fill_2 FILLER_24_522 ();
 sg13g2_fill_2 FILLER_24_599 ();
 sg13g2_fill_2 FILLER_24_679 ();
 sg13g2_fill_1 FILLER_24_690 ();
 sg13g2_fill_2 FILLER_24_704 ();
 sg13g2_fill_1 FILLER_24_725 ();
 sg13g2_decap_8 FILLER_24_768 ();
 sg13g2_decap_8 FILLER_24_775 ();
 sg13g2_fill_1 FILLER_24_804 ();
 sg13g2_fill_2 FILLER_24_847 ();
 sg13g2_fill_2 FILLER_24_889 ();
 sg13g2_fill_1 FILLER_24_922 ();
 sg13g2_fill_2 FILLER_24_982 ();
 sg13g2_fill_2 FILLER_24_1031 ();
 sg13g2_fill_2 FILLER_24_1150 ();
 sg13g2_fill_1 FILLER_24_1152 ();
 sg13g2_fill_2 FILLER_24_1157 ();
 sg13g2_fill_1 FILLER_24_1174 ();
 sg13g2_fill_1 FILLER_24_1180 ();
 sg13g2_fill_1 FILLER_24_1194 ();
 sg13g2_fill_2 FILLER_24_1204 ();
 sg13g2_fill_2 FILLER_24_1249 ();
 sg13g2_decap_4 FILLER_24_1310 ();
 sg13g2_fill_2 FILLER_24_1314 ();
 sg13g2_decap_8 FILLER_24_1381 ();
 sg13g2_fill_2 FILLER_24_1388 ();
 sg13g2_fill_1 FILLER_24_1390 ();
 sg13g2_fill_2 FILLER_24_1426 ();
 sg13g2_fill_2 FILLER_24_1433 ();
 sg13g2_fill_1 FILLER_24_1435 ();
 sg13g2_decap_4 FILLER_24_1444 ();
 sg13g2_fill_1 FILLER_24_1448 ();
 sg13g2_decap_8 FILLER_24_1458 ();
 sg13g2_fill_1 FILLER_24_1465 ();
 sg13g2_decap_4 FILLER_24_1476 ();
 sg13g2_decap_8 FILLER_24_1498 ();
 sg13g2_decap_8 FILLER_24_1505 ();
 sg13g2_fill_1 FILLER_24_1512 ();
 sg13g2_decap_4 FILLER_24_1567 ();
 sg13g2_fill_2 FILLER_24_1571 ();
 sg13g2_decap_4 FILLER_24_1577 ();
 sg13g2_fill_2 FILLER_24_1581 ();
 sg13g2_decap_8 FILLER_24_1589 ();
 sg13g2_fill_2 FILLER_24_1596 ();
 sg13g2_fill_1 FILLER_24_1598 ();
 sg13g2_fill_2 FILLER_24_1607 ();
 sg13g2_fill_1 FILLER_24_1683 ();
 sg13g2_fill_2 FILLER_24_1688 ();
 sg13g2_fill_2 FILLER_24_1726 ();
 sg13g2_fill_1 FILLER_24_1728 ();
 sg13g2_fill_1 FILLER_24_1738 ();
 sg13g2_fill_2 FILLER_24_1744 ();
 sg13g2_fill_1 FILLER_24_1746 ();
 sg13g2_fill_2 FILLER_24_1760 ();
 sg13g2_decap_4 FILLER_24_1793 ();
 sg13g2_fill_1 FILLER_24_1933 ();
 sg13g2_decap_8 FILLER_24_1948 ();
 sg13g2_decap_4 FILLER_24_1976 ();
 sg13g2_fill_1 FILLER_24_1980 ();
 sg13g2_decap_8 FILLER_24_2020 ();
 sg13g2_fill_2 FILLER_24_2027 ();
 sg13g2_fill_1 FILLER_24_2029 ();
 sg13g2_fill_1 FILLER_24_2040 ();
 sg13g2_fill_1 FILLER_24_2072 ();
 sg13g2_fill_2 FILLER_24_2104 ();
 sg13g2_fill_1 FILLER_24_2106 ();
 sg13g2_fill_1 FILLER_24_2133 ();
 sg13g2_fill_2 FILLER_24_2140 ();
 sg13g2_fill_1 FILLER_24_2142 ();
 sg13g2_fill_2 FILLER_24_2169 ();
 sg13g2_fill_1 FILLER_24_2360 ();
 sg13g2_decap_8 FILLER_24_2419 ();
 sg13g2_fill_1 FILLER_24_2426 ();
 sg13g2_fill_1 FILLER_24_2458 ();
 sg13g2_fill_2 FILLER_24_2485 ();
 sg13g2_decap_8 FILLER_24_2491 ();
 sg13g2_fill_1 FILLER_24_2498 ();
 sg13g2_fill_1 FILLER_24_2543 ();
 sg13g2_fill_2 FILLER_24_2549 ();
 sg13g2_fill_1 FILLER_24_2551 ();
 sg13g2_decap_8 FILLER_24_2595 ();
 sg13g2_decap_8 FILLER_24_2602 ();
 sg13g2_decap_8 FILLER_24_2609 ();
 sg13g2_decap_8 FILLER_24_2616 ();
 sg13g2_decap_8 FILLER_24_2623 ();
 sg13g2_decap_8 FILLER_24_2630 ();
 sg13g2_decap_8 FILLER_24_2637 ();
 sg13g2_decap_8 FILLER_24_2644 ();
 sg13g2_decap_8 FILLER_24_2651 ();
 sg13g2_decap_8 FILLER_24_2658 ();
 sg13g2_decap_8 FILLER_24_2665 ();
 sg13g2_fill_2 FILLER_24_2672 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_4 FILLER_25_483 ();
 sg13g2_fill_2 FILLER_25_517 ();
 sg13g2_fill_1 FILLER_25_568 ();
 sg13g2_fill_1 FILLER_25_584 ();
 sg13g2_fill_2 FILLER_25_595 ();
 sg13g2_fill_1 FILLER_25_597 ();
 sg13g2_fill_2 FILLER_25_614 ();
 sg13g2_fill_2 FILLER_25_624 ();
 sg13g2_fill_1 FILLER_25_626 ();
 sg13g2_fill_2 FILLER_25_636 ();
 sg13g2_fill_2 FILLER_25_657 ();
 sg13g2_fill_2 FILLER_25_677 ();
 sg13g2_fill_1 FILLER_25_685 ();
 sg13g2_fill_2 FILLER_25_707 ();
 sg13g2_fill_1 FILLER_25_738 ();
 sg13g2_fill_1 FILLER_25_755 ();
 sg13g2_decap_8 FILLER_25_775 ();
 sg13g2_fill_2 FILLER_25_793 ();
 sg13g2_fill_2 FILLER_25_799 ();
 sg13g2_fill_2 FILLER_25_813 ();
 sg13g2_fill_1 FILLER_25_828 ();
 sg13g2_fill_2 FILLER_25_834 ();
 sg13g2_fill_2 FILLER_25_884 ();
 sg13g2_fill_1 FILLER_25_886 ();
 sg13g2_fill_2 FILLER_25_936 ();
 sg13g2_fill_2 FILLER_25_946 ();
 sg13g2_fill_2 FILLER_25_992 ();
 sg13g2_fill_2 FILLER_25_1016 ();
 sg13g2_fill_2 FILLER_25_1110 ();
 sg13g2_fill_1 FILLER_25_1112 ();
 sg13g2_fill_1 FILLER_25_1118 ();
 sg13g2_fill_2 FILLER_25_1129 ();
 sg13g2_fill_1 FILLER_25_1136 ();
 sg13g2_fill_2 FILLER_25_1153 ();
 sg13g2_fill_1 FILLER_25_1155 ();
 sg13g2_fill_2 FILLER_25_1216 ();
 sg13g2_fill_2 FILLER_25_1248 ();
 sg13g2_fill_1 FILLER_25_1250 ();
 sg13g2_fill_2 FILLER_25_1256 ();
 sg13g2_fill_1 FILLER_25_1258 ();
 sg13g2_fill_1 FILLER_25_1294 ();
 sg13g2_decap_4 FILLER_25_1381 ();
 sg13g2_fill_2 FILLER_25_1385 ();
 sg13g2_fill_2 FILLER_25_1422 ();
 sg13g2_fill_1 FILLER_25_1424 ();
 sg13g2_decap_8 FILLER_25_1442 ();
 sg13g2_decap_8 FILLER_25_1449 ();
 sg13g2_fill_2 FILLER_25_1456 ();
 sg13g2_fill_1 FILLER_25_1458 ();
 sg13g2_fill_1 FILLER_25_1501 ();
 sg13g2_decap_4 FILLER_25_1528 ();
 sg13g2_decap_4 FILLER_25_1545 ();
 sg13g2_fill_2 FILLER_25_1549 ();
 sg13g2_fill_1 FILLER_25_1568 ();
 sg13g2_fill_2 FILLER_25_1601 ();
 sg13g2_fill_1 FILLER_25_1660 ();
 sg13g2_decap_8 FILLER_25_1691 ();
 sg13g2_fill_2 FILLER_25_1698 ();
 sg13g2_fill_1 FILLER_25_1734 ();
 sg13g2_fill_1 FILLER_25_1761 ();
 sg13g2_fill_1 FILLER_25_1921 ();
 sg13g2_decap_8 FILLER_25_1957 ();
 sg13g2_decap_4 FILLER_25_1964 ();
 sg13g2_fill_1 FILLER_25_1968 ();
 sg13g2_fill_2 FILLER_25_2030 ();
 sg13g2_decap_8 FILLER_25_2045 ();
 sg13g2_fill_2 FILLER_25_2052 ();
 sg13g2_fill_1 FILLER_25_2084 ();
 sg13g2_fill_2 FILLER_25_2089 ();
 sg13g2_fill_1 FILLER_25_2091 ();
 sg13g2_fill_2 FILLER_25_2101 ();
 sg13g2_fill_1 FILLER_25_2103 ();
 sg13g2_decap_4 FILLER_25_2134 ();
 sg13g2_fill_2 FILLER_25_2138 ();
 sg13g2_decap_4 FILLER_25_2237 ();
 sg13g2_fill_2 FILLER_25_2272 ();
 sg13g2_fill_2 FILLER_25_2293 ();
 sg13g2_fill_2 FILLER_25_2318 ();
 sg13g2_fill_1 FILLER_25_2320 ();
 sg13g2_fill_1 FILLER_25_2338 ();
 sg13g2_fill_2 FILLER_25_2344 ();
 sg13g2_fill_2 FILLER_25_2351 ();
 sg13g2_fill_2 FILLER_25_2377 ();
 sg13g2_fill_1 FILLER_25_2379 ();
 sg13g2_fill_1 FILLER_25_2397 ();
 sg13g2_decap_4 FILLER_25_2406 ();
 sg13g2_fill_2 FILLER_25_2493 ();
 sg13g2_fill_1 FILLER_25_2539 ();
 sg13g2_decap_8 FILLER_25_2591 ();
 sg13g2_decap_8 FILLER_25_2598 ();
 sg13g2_decap_8 FILLER_25_2605 ();
 sg13g2_decap_8 FILLER_25_2612 ();
 sg13g2_decap_8 FILLER_25_2619 ();
 sg13g2_decap_8 FILLER_25_2626 ();
 sg13g2_decap_8 FILLER_25_2633 ();
 sg13g2_decap_8 FILLER_25_2640 ();
 sg13g2_decap_8 FILLER_25_2647 ();
 sg13g2_decap_8 FILLER_25_2654 ();
 sg13g2_decap_8 FILLER_25_2661 ();
 sg13g2_decap_4 FILLER_25_2668 ();
 sg13g2_fill_2 FILLER_25_2672 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_fill_1 FILLER_26_497 ();
 sg13g2_fill_1 FILLER_26_515 ();
 sg13g2_fill_1 FILLER_26_618 ();
 sg13g2_fill_2 FILLER_26_647 ();
 sg13g2_fill_1 FILLER_26_685 ();
 sg13g2_fill_2 FILLER_26_769 ();
 sg13g2_fill_1 FILLER_26_771 ();
 sg13g2_fill_2 FILLER_26_785 ();
 sg13g2_fill_1 FILLER_26_787 ();
 sg13g2_decap_4 FILLER_26_791 ();
 sg13g2_fill_2 FILLER_26_795 ();
 sg13g2_fill_1 FILLER_26_845 ();
 sg13g2_fill_1 FILLER_26_875 ();
 sg13g2_fill_2 FILLER_26_891 ();
 sg13g2_fill_1 FILLER_26_893 ();
 sg13g2_decap_4 FILLER_26_919 ();
 sg13g2_fill_2 FILLER_26_988 ();
 sg13g2_fill_2 FILLER_26_1016 ();
 sg13g2_fill_1 FILLER_26_1095 ();
 sg13g2_fill_2 FILLER_26_1152 ();
 sg13g2_fill_1 FILLER_26_1154 ();
 sg13g2_fill_2 FILLER_26_1181 ();
 sg13g2_fill_1 FILLER_26_1183 ();
 sg13g2_fill_2 FILLER_26_1201 ();
 sg13g2_fill_1 FILLER_26_1203 ();
 sg13g2_fill_2 FILLER_26_1232 ();
 sg13g2_fill_2 FILLER_26_1248 ();
 sg13g2_fill_1 FILLER_26_1250 ();
 sg13g2_fill_2 FILLER_26_1296 ();
 sg13g2_fill_1 FILLER_26_1358 ();
 sg13g2_fill_2 FILLER_26_1378 ();
 sg13g2_fill_2 FILLER_26_1394 ();
 sg13g2_fill_2 FILLER_26_1406 ();
 sg13g2_decap_4 FILLER_26_1448 ();
 sg13g2_fill_1 FILLER_26_1452 ();
 sg13g2_fill_1 FILLER_26_1456 ();
 sg13g2_fill_2 FILLER_26_1550 ();
 sg13g2_fill_1 FILLER_26_1552 ();
 sg13g2_fill_2 FILLER_26_1566 ();
 sg13g2_fill_2 FILLER_26_1578 ();
 sg13g2_decap_4 FILLER_26_1588 ();
 sg13g2_fill_2 FILLER_26_1592 ();
 sg13g2_fill_1 FILLER_26_1598 ();
 sg13g2_decap_4 FILLER_26_1698 ();
 sg13g2_fill_2 FILLER_26_1710 ();
 sg13g2_fill_1 FILLER_26_1712 ();
 sg13g2_decap_4 FILLER_26_1721 ();
 sg13g2_fill_1 FILLER_26_1725 ();
 sg13g2_fill_1 FILLER_26_1730 ();
 sg13g2_fill_2 FILLER_26_1807 ();
 sg13g2_fill_1 FILLER_26_1809 ();
 sg13g2_fill_2 FILLER_26_1867 ();
 sg13g2_fill_1 FILLER_26_1869 ();
 sg13g2_fill_1 FILLER_26_1965 ();
 sg13g2_fill_1 FILLER_26_1987 ();
 sg13g2_fill_2 FILLER_26_1997 ();
 sg13g2_decap_8 FILLER_26_2051 ();
 sg13g2_decap_8 FILLER_26_2058 ();
 sg13g2_decap_4 FILLER_26_2065 ();
 sg13g2_fill_2 FILLER_26_2077 ();
 sg13g2_decap_8 FILLER_26_2092 ();
 sg13g2_decap_8 FILLER_26_2099 ();
 sg13g2_decap_4 FILLER_26_2106 ();
 sg13g2_fill_1 FILLER_26_2110 ();
 sg13g2_fill_1 FILLER_26_2120 ();
 sg13g2_decap_8 FILLER_26_2130 ();
 sg13g2_decap_4 FILLER_26_2137 ();
 sg13g2_fill_2 FILLER_26_2141 ();
 sg13g2_fill_2 FILLER_26_2148 ();
 sg13g2_fill_1 FILLER_26_2150 ();
 sg13g2_fill_2 FILLER_26_2170 ();
 sg13g2_fill_1 FILLER_26_2181 ();
 sg13g2_fill_2 FILLER_26_2196 ();
 sg13g2_fill_1 FILLER_26_2215 ();
 sg13g2_decap_8 FILLER_26_2225 ();
 sg13g2_fill_2 FILLER_26_2232 ();
 sg13g2_decap_4 FILLER_26_2240 ();
 sg13g2_fill_1 FILLER_26_2244 ();
 sg13g2_fill_2 FILLER_26_2250 ();
 sg13g2_fill_1 FILLER_26_2252 ();
 sg13g2_fill_2 FILLER_26_2309 ();
 sg13g2_fill_1 FILLER_26_2311 ();
 sg13g2_fill_2 FILLER_26_2328 ();
 sg13g2_fill_1 FILLER_26_2330 ();
 sg13g2_fill_2 FILLER_26_2342 ();
 sg13g2_fill_1 FILLER_26_2382 ();
 sg13g2_fill_1 FILLER_26_2438 ();
 sg13g2_fill_1 FILLER_26_2448 ();
 sg13g2_decap_8 FILLER_26_2581 ();
 sg13g2_decap_8 FILLER_26_2588 ();
 sg13g2_decap_8 FILLER_26_2595 ();
 sg13g2_decap_8 FILLER_26_2602 ();
 sg13g2_decap_8 FILLER_26_2609 ();
 sg13g2_decap_8 FILLER_26_2616 ();
 sg13g2_decap_8 FILLER_26_2623 ();
 sg13g2_decap_8 FILLER_26_2630 ();
 sg13g2_decap_8 FILLER_26_2637 ();
 sg13g2_decap_8 FILLER_26_2644 ();
 sg13g2_decap_8 FILLER_26_2651 ();
 sg13g2_decap_8 FILLER_26_2658 ();
 sg13g2_decap_8 FILLER_26_2665 ();
 sg13g2_fill_2 FILLER_26_2672 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_fill_2 FILLER_27_523 ();
 sg13g2_fill_2 FILLER_27_534 ();
 sg13g2_fill_1 FILLER_27_541 ();
 sg13g2_fill_1 FILLER_27_560 ();
 sg13g2_fill_2 FILLER_27_585 ();
 sg13g2_fill_1 FILLER_27_657 ();
 sg13g2_fill_2 FILLER_27_684 ();
 sg13g2_fill_1 FILLER_27_712 ();
 sg13g2_decap_4 FILLER_27_727 ();
 sg13g2_fill_1 FILLER_27_731 ();
 sg13g2_fill_1 FILLER_27_785 ();
 sg13g2_fill_1 FILLER_27_812 ();
 sg13g2_fill_2 FILLER_27_862 ();
 sg13g2_fill_2 FILLER_27_873 ();
 sg13g2_fill_1 FILLER_27_875 ();
 sg13g2_fill_1 FILLER_27_911 ();
 sg13g2_fill_2 FILLER_27_917 ();
 sg13g2_fill_2 FILLER_27_931 ();
 sg13g2_fill_2 FILLER_27_986 ();
 sg13g2_fill_1 FILLER_27_988 ();
 sg13g2_fill_2 FILLER_27_1014 ();
 sg13g2_fill_1 FILLER_27_1025 ();
 sg13g2_fill_2 FILLER_27_1039 ();
 sg13g2_fill_2 FILLER_27_1062 ();
 sg13g2_fill_1 FILLER_27_1064 ();
 sg13g2_fill_2 FILLER_27_1082 ();
 sg13g2_fill_2 FILLER_27_1152 ();
 sg13g2_fill_2 FILLER_27_1193 ();
 sg13g2_fill_2 FILLER_27_1221 ();
 sg13g2_fill_1 FILLER_27_1223 ();
 sg13g2_fill_1 FILLER_27_1236 ();
 sg13g2_fill_1 FILLER_27_1242 ();
 sg13g2_fill_2 FILLER_27_1265 ();
 sg13g2_fill_1 FILLER_27_1267 ();
 sg13g2_fill_1 FILLER_27_1297 ();
 sg13g2_fill_1 FILLER_27_1309 ();
 sg13g2_fill_2 FILLER_27_1417 ();
 sg13g2_fill_1 FILLER_27_1465 ();
 sg13g2_fill_2 FILLER_27_1489 ();
 sg13g2_fill_1 FILLER_27_1491 ();
 sg13g2_fill_1 FILLER_27_1520 ();
 sg13g2_decap_8 FILLER_27_1547 ();
 sg13g2_decap_8 FILLER_27_1554 ();
 sg13g2_fill_1 FILLER_27_1561 ();
 sg13g2_decap_8 FILLER_27_1588 ();
 sg13g2_fill_2 FILLER_27_1595 ();
 sg13g2_fill_1 FILLER_27_1623 ();
 sg13g2_fill_1 FILLER_27_1710 ();
 sg13g2_decap_4 FILLER_27_1728 ();
 sg13g2_fill_2 FILLER_27_1732 ();
 sg13g2_decap_4 FILLER_27_1766 ();
 sg13g2_fill_2 FILLER_27_1770 ();
 sg13g2_fill_2 FILLER_27_1778 ();
 sg13g2_fill_1 FILLER_27_1780 ();
 sg13g2_fill_1 FILLER_27_1806 ();
 sg13g2_fill_2 FILLER_27_1846 ();
 sg13g2_fill_1 FILLER_27_1857 ();
 sg13g2_fill_1 FILLER_27_1881 ();
 sg13g2_fill_2 FILLER_27_1896 ();
 sg13g2_fill_2 FILLER_27_1963 ();
 sg13g2_fill_2 FILLER_27_1969 ();
 sg13g2_fill_1 FILLER_27_2071 ();
 sg13g2_fill_2 FILLER_27_2117 ();
 sg13g2_fill_1 FILLER_27_2119 ();
 sg13g2_fill_1 FILLER_27_2124 ();
 sg13g2_fill_2 FILLER_27_2131 ();
 sg13g2_fill_2 FILLER_27_2137 ();
 sg13g2_fill_1 FILLER_27_2139 ();
 sg13g2_fill_1 FILLER_27_2182 ();
 sg13g2_fill_2 FILLER_27_2195 ();
 sg13g2_fill_2 FILLER_27_2205 ();
 sg13g2_fill_1 FILLER_27_2207 ();
 sg13g2_decap_8 FILLER_27_2220 ();
 sg13g2_fill_2 FILLER_27_2227 ();
 sg13g2_fill_1 FILLER_27_2229 ();
 sg13g2_fill_1 FILLER_27_2246 ();
 sg13g2_fill_1 FILLER_27_2300 ();
 sg13g2_fill_2 FILLER_27_2314 ();
 sg13g2_fill_1 FILLER_27_2316 ();
 sg13g2_fill_1 FILLER_27_2408 ();
 sg13g2_fill_2 FILLER_27_2414 ();
 sg13g2_fill_1 FILLER_27_2428 ();
 sg13g2_fill_2 FILLER_27_2434 ();
 sg13g2_fill_1 FILLER_27_2477 ();
 sg13g2_fill_1 FILLER_27_2505 ();
 sg13g2_fill_2 FILLER_27_2532 ();
 sg13g2_decap_8 FILLER_27_2590 ();
 sg13g2_decap_8 FILLER_27_2597 ();
 sg13g2_decap_8 FILLER_27_2604 ();
 sg13g2_decap_8 FILLER_27_2611 ();
 sg13g2_decap_8 FILLER_27_2618 ();
 sg13g2_decap_8 FILLER_27_2625 ();
 sg13g2_decap_8 FILLER_27_2632 ();
 sg13g2_decap_8 FILLER_27_2639 ();
 sg13g2_decap_8 FILLER_27_2646 ();
 sg13g2_decap_8 FILLER_27_2653 ();
 sg13g2_decap_8 FILLER_27_2660 ();
 sg13g2_decap_8 FILLER_27_2667 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_decap_8 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_462 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_4 FILLER_28_483 ();
 sg13g2_fill_2 FILLER_28_487 ();
 sg13g2_fill_2 FILLER_28_591 ();
 sg13g2_fill_2 FILLER_28_647 ();
 sg13g2_fill_1 FILLER_28_649 ();
 sg13g2_fill_2 FILLER_28_659 ();
 sg13g2_fill_1 FILLER_28_670 ();
 sg13g2_fill_2 FILLER_28_692 ();
 sg13g2_fill_1 FILLER_28_791 ();
 sg13g2_fill_2 FILLER_28_837 ();
 sg13g2_fill_1 FILLER_28_839 ();
 sg13g2_fill_1 FILLER_28_930 ();
 sg13g2_fill_2 FILLER_28_991 ();
 sg13g2_fill_1 FILLER_28_1011 ();
 sg13g2_fill_1 FILLER_28_1022 ();
 sg13g2_fill_2 FILLER_28_1033 ();
 sg13g2_fill_1 FILLER_28_1044 ();
 sg13g2_fill_1 FILLER_28_1144 ();
 sg13g2_decap_8 FILLER_28_1162 ();
 sg13g2_fill_1 FILLER_28_1169 ();
 sg13g2_fill_2 FILLER_28_1183 ();
 sg13g2_fill_1 FILLER_28_1185 ();
 sg13g2_fill_1 FILLER_28_1204 ();
 sg13g2_fill_2 FILLER_28_1223 ();
 sg13g2_fill_1 FILLER_28_1225 ();
 sg13g2_fill_2 FILLER_28_1252 ();
 sg13g2_fill_2 FILLER_28_1271 ();
 sg13g2_fill_2 FILLER_28_1355 ();
 sg13g2_fill_1 FILLER_28_1357 ();
 sg13g2_fill_2 FILLER_28_1411 ();
 sg13g2_fill_2 FILLER_28_1432 ();
 sg13g2_fill_1 FILLER_28_1434 ();
 sg13g2_fill_1 FILLER_28_1473 ();
 sg13g2_fill_2 FILLER_28_1486 ();
 sg13g2_fill_2 FILLER_28_1494 ();
 sg13g2_fill_1 FILLER_28_1496 ();
 sg13g2_fill_2 FILLER_28_1512 ();
 sg13g2_fill_1 FILLER_28_1514 ();
 sg13g2_decap_4 FILLER_28_1562 ();
 sg13g2_fill_2 FILLER_28_1566 ();
 sg13g2_fill_2 FILLER_28_1602 ();
 sg13g2_fill_1 FILLER_28_1634 ();
 sg13g2_fill_1 FILLER_28_1644 ();
 sg13g2_fill_2 FILLER_28_1659 ();
 sg13g2_fill_1 FILLER_28_1661 ();
 sg13g2_fill_1 FILLER_28_1676 ();
 sg13g2_fill_2 FILLER_28_1686 ();
 sg13g2_fill_1 FILLER_28_1754 ();
 sg13g2_decap_8 FILLER_28_1765 ();
 sg13g2_fill_2 FILLER_28_1772 ();
 sg13g2_decap_4 FILLER_28_1796 ();
 sg13g2_fill_2 FILLER_28_1809 ();
 sg13g2_fill_1 FILLER_28_1811 ();
 sg13g2_fill_1 FILLER_28_1817 ();
 sg13g2_fill_2 FILLER_28_1832 ();
 sg13g2_fill_1 FILLER_28_1834 ();
 sg13g2_fill_2 FILLER_28_1852 ();
 sg13g2_fill_1 FILLER_28_1854 ();
 sg13g2_fill_2 FILLER_28_1863 ();
 sg13g2_fill_2 FILLER_28_1870 ();
 sg13g2_fill_1 FILLER_28_1902 ();
 sg13g2_fill_2 FILLER_28_1935 ();
 sg13g2_fill_2 FILLER_28_1967 ();
 sg13g2_fill_1 FILLER_28_1990 ();
 sg13g2_fill_2 FILLER_28_2070 ();
 sg13g2_fill_1 FILLER_28_2114 ();
 sg13g2_fill_2 FILLER_28_2165 ();
 sg13g2_fill_2 FILLER_28_2189 ();
 sg13g2_fill_2 FILLER_28_2210 ();
 sg13g2_decap_8 FILLER_28_2230 ();
 sg13g2_fill_1 FILLER_28_2287 ();
 sg13g2_fill_2 FILLER_28_2317 ();
 sg13g2_fill_1 FILLER_28_2373 ();
 sg13g2_fill_2 FILLER_28_2387 ();
 sg13g2_fill_2 FILLER_28_2404 ();
 sg13g2_fill_1 FILLER_28_2406 ();
 sg13g2_fill_2 FILLER_28_2416 ();
 sg13g2_fill_2 FILLER_28_2440 ();
 sg13g2_fill_1 FILLER_28_2448 ();
 sg13g2_fill_2 FILLER_28_2485 ();
 sg13g2_fill_1 FILLER_28_2520 ();
 sg13g2_decap_8 FILLER_28_2578 ();
 sg13g2_decap_8 FILLER_28_2585 ();
 sg13g2_decap_8 FILLER_28_2592 ();
 sg13g2_decap_8 FILLER_28_2599 ();
 sg13g2_decap_8 FILLER_28_2606 ();
 sg13g2_decap_8 FILLER_28_2613 ();
 sg13g2_decap_8 FILLER_28_2620 ();
 sg13g2_decap_8 FILLER_28_2627 ();
 sg13g2_decap_8 FILLER_28_2634 ();
 sg13g2_decap_8 FILLER_28_2641 ();
 sg13g2_decap_8 FILLER_28_2648 ();
 sg13g2_decap_8 FILLER_28_2655 ();
 sg13g2_decap_8 FILLER_28_2662 ();
 sg13g2_decap_4 FILLER_28_2669 ();
 sg13g2_fill_1 FILLER_28_2673 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_4 FILLER_29_490 ();
 sg13g2_fill_2 FILLER_29_537 ();
 sg13g2_fill_1 FILLER_29_604 ();
 sg13g2_fill_2 FILLER_29_631 ();
 sg13g2_fill_2 FILLER_29_668 ();
 sg13g2_fill_1 FILLER_29_670 ();
 sg13g2_fill_2 FILLER_29_676 ();
 sg13g2_fill_1 FILLER_29_678 ();
 sg13g2_fill_2 FILLER_29_692 ();
 sg13g2_fill_1 FILLER_29_694 ();
 sg13g2_fill_1 FILLER_29_706 ();
 sg13g2_fill_2 FILLER_29_753 ();
 sg13g2_fill_1 FILLER_29_795 ();
 sg13g2_fill_1 FILLER_29_800 ();
 sg13g2_fill_2 FILLER_29_804 ();
 sg13g2_decap_4 FILLER_29_809 ();
 sg13g2_fill_1 FILLER_29_813 ();
 sg13g2_fill_2 FILLER_29_850 ();
 sg13g2_fill_1 FILLER_29_852 ();
 sg13g2_fill_1 FILLER_29_935 ();
 sg13g2_fill_2 FILLER_29_1024 ();
 sg13g2_fill_1 FILLER_29_1026 ();
 sg13g2_fill_1 FILLER_29_1045 ();
 sg13g2_fill_2 FILLER_29_1055 ();
 sg13g2_fill_1 FILLER_29_1097 ();
 sg13g2_fill_2 FILLER_29_1133 ();
 sg13g2_fill_1 FILLER_29_1143 ();
 sg13g2_decap_8 FILLER_29_1169 ();
 sg13g2_fill_2 FILLER_29_1236 ();
 sg13g2_fill_2 FILLER_29_1271 ();
 sg13g2_fill_1 FILLER_29_1285 ();
 sg13g2_fill_2 FILLER_29_1327 ();
 sg13g2_fill_2 FILLER_29_1384 ();
 sg13g2_fill_1 FILLER_29_1391 ();
 sg13g2_fill_2 FILLER_29_1432 ();
 sg13g2_fill_1 FILLER_29_1434 ();
 sg13g2_fill_1 FILLER_29_1470 ();
 sg13g2_fill_1 FILLER_29_1506 ();
 sg13g2_decap_4 FILLER_29_1576 ();
 sg13g2_fill_1 FILLER_29_1580 ();
 sg13g2_fill_2 FILLER_29_1619 ();
 sg13g2_fill_2 FILLER_29_1681 ();
 sg13g2_fill_2 FILLER_29_1772 ();
 sg13g2_fill_2 FILLER_29_1779 ();
 sg13g2_fill_1 FILLER_29_1781 ();
 sg13g2_fill_2 FILLER_29_1791 ();
 sg13g2_fill_2 FILLER_29_1844 ();
 sg13g2_fill_1 FILLER_29_1846 ();
 sg13g2_fill_2 FILLER_29_1865 ();
 sg13g2_fill_2 FILLER_29_1899 ();
 sg13g2_fill_1 FILLER_29_1909 ();
 sg13g2_fill_2 FILLER_29_1951 ();
 sg13g2_fill_1 FILLER_29_1953 ();
 sg13g2_fill_2 FILLER_29_1990 ();
 sg13g2_fill_1 FILLER_29_1992 ();
 sg13g2_fill_1 FILLER_29_2015 ();
 sg13g2_fill_2 FILLER_29_2061 ();
 sg13g2_fill_1 FILLER_29_2063 ();
 sg13g2_fill_1 FILLER_29_2095 ();
 sg13g2_fill_1 FILLER_29_2126 ();
 sg13g2_fill_2 FILLER_29_2143 ();
 sg13g2_fill_2 FILLER_29_2265 ();
 sg13g2_fill_1 FILLER_29_2271 ();
 sg13g2_fill_1 FILLER_29_2295 ();
 sg13g2_fill_2 FILLER_29_2378 ();
 sg13g2_fill_2 FILLER_29_2418 ();
 sg13g2_fill_1 FILLER_29_2483 ();
 sg13g2_decap_4 FILLER_29_2518 ();
 sg13g2_fill_1 FILLER_29_2522 ();
 sg13g2_decap_8 FILLER_29_2584 ();
 sg13g2_decap_8 FILLER_29_2591 ();
 sg13g2_decap_8 FILLER_29_2598 ();
 sg13g2_decap_8 FILLER_29_2605 ();
 sg13g2_decap_8 FILLER_29_2612 ();
 sg13g2_decap_8 FILLER_29_2619 ();
 sg13g2_decap_8 FILLER_29_2626 ();
 sg13g2_decap_8 FILLER_29_2633 ();
 sg13g2_decap_8 FILLER_29_2640 ();
 sg13g2_decap_8 FILLER_29_2647 ();
 sg13g2_decap_8 FILLER_29_2654 ();
 sg13g2_decap_8 FILLER_29_2661 ();
 sg13g2_decap_4 FILLER_29_2668 ();
 sg13g2_fill_2 FILLER_29_2672 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_fill_2 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_533 ();
 sg13g2_fill_2 FILLER_30_540 ();
 sg13g2_fill_1 FILLER_30_572 ();
 sg13g2_fill_1 FILLER_30_587 ();
 sg13g2_fill_2 FILLER_30_665 ();
 sg13g2_fill_2 FILLER_30_702 ();
 sg13g2_fill_1 FILLER_30_704 ();
 sg13g2_fill_1 FILLER_30_739 ();
 sg13g2_fill_2 FILLER_30_772 ();
 sg13g2_fill_1 FILLER_30_774 ();
 sg13g2_fill_2 FILLER_30_785 ();
 sg13g2_fill_2 FILLER_30_795 ();
 sg13g2_fill_1 FILLER_30_797 ();
 sg13g2_fill_1 FILLER_30_811 ();
 sg13g2_fill_2 FILLER_30_837 ();
 sg13g2_fill_1 FILLER_30_839 ();
 sg13g2_fill_2 FILLER_30_849 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_fill_1 FILLER_30_867 ();
 sg13g2_fill_2 FILLER_30_885 ();
 sg13g2_fill_1 FILLER_30_887 ();
 sg13g2_fill_1 FILLER_30_892 ();
 sg13g2_fill_2 FILLER_30_898 ();
 sg13g2_fill_2 FILLER_30_913 ();
 sg13g2_fill_2 FILLER_30_1006 ();
 sg13g2_fill_1 FILLER_30_1069 ();
 sg13g2_decap_4 FILLER_30_1078 ();
 sg13g2_fill_1 FILLER_30_1082 ();
 sg13g2_decap_4 FILLER_30_1091 ();
 sg13g2_fill_2 FILLER_30_1103 ();
 sg13g2_decap_4 FILLER_30_1122 ();
 sg13g2_fill_2 FILLER_30_1178 ();
 sg13g2_fill_1 FILLER_30_1180 ();
 sg13g2_fill_1 FILLER_30_1186 ();
 sg13g2_fill_2 FILLER_30_1373 ();
 sg13g2_fill_1 FILLER_30_1375 ();
 sg13g2_fill_1 FILLER_30_1402 ();
 sg13g2_fill_1 FILLER_30_1458 ();
 sg13g2_fill_2 FILLER_30_1585 ();
 sg13g2_fill_1 FILLER_30_1587 ();
 sg13g2_decap_4 FILLER_30_1593 ();
 sg13g2_fill_1 FILLER_30_1597 ();
 sg13g2_fill_1 FILLER_30_1637 ();
 sg13g2_fill_2 FILLER_30_1664 ();
 sg13g2_fill_1 FILLER_30_1712 ();
 sg13g2_fill_2 FILLER_30_1718 ();
 sg13g2_fill_1 FILLER_30_1737 ();
 sg13g2_fill_2 FILLER_30_1884 ();
 sg13g2_fill_2 FILLER_30_1921 ();
 sg13g2_fill_1 FILLER_30_1988 ();
 sg13g2_fill_2 FILLER_30_2023 ();
 sg13g2_fill_1 FILLER_30_2025 ();
 sg13g2_fill_1 FILLER_30_2031 ();
 sg13g2_fill_2 FILLER_30_2040 ();
 sg13g2_fill_1 FILLER_30_2061 ();
 sg13g2_fill_2 FILLER_30_2067 ();
 sg13g2_fill_1 FILLER_30_2069 ();
 sg13g2_fill_2 FILLER_30_2097 ();
 sg13g2_fill_1 FILLER_30_2124 ();
 sg13g2_fill_2 FILLER_30_2134 ();
 sg13g2_fill_1 FILLER_30_2136 ();
 sg13g2_fill_2 FILLER_30_2218 ();
 sg13g2_decap_8 FILLER_30_2241 ();
 sg13g2_decap_8 FILLER_30_2248 ();
 sg13g2_decap_4 FILLER_30_2255 ();
 sg13g2_decap_8 FILLER_30_2277 ();
 sg13g2_fill_2 FILLER_30_2318 ();
 sg13g2_fill_1 FILLER_30_2320 ();
 sg13g2_fill_2 FILLER_30_2366 ();
 sg13g2_fill_2 FILLER_30_2419 ();
 sg13g2_fill_1 FILLER_30_2421 ();
 sg13g2_fill_1 FILLER_30_2448 ();
 sg13g2_fill_1 FILLER_30_2460 ();
 sg13g2_fill_1 FILLER_30_2534 ();
 sg13g2_decap_8 FILLER_30_2565 ();
 sg13g2_decap_8 FILLER_30_2572 ();
 sg13g2_decap_8 FILLER_30_2579 ();
 sg13g2_decap_8 FILLER_30_2586 ();
 sg13g2_decap_8 FILLER_30_2593 ();
 sg13g2_decap_8 FILLER_30_2600 ();
 sg13g2_decap_8 FILLER_30_2607 ();
 sg13g2_decap_8 FILLER_30_2614 ();
 sg13g2_decap_8 FILLER_30_2621 ();
 sg13g2_decap_8 FILLER_30_2628 ();
 sg13g2_decap_8 FILLER_30_2635 ();
 sg13g2_decap_8 FILLER_30_2642 ();
 sg13g2_decap_8 FILLER_30_2649 ();
 sg13g2_decap_8 FILLER_30_2656 ();
 sg13g2_decap_8 FILLER_30_2663 ();
 sg13g2_decap_4 FILLER_30_2670 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_4 FILLER_31_511 ();
 sg13g2_fill_1 FILLER_31_515 ();
 sg13g2_fill_2 FILLER_31_534 ();
 sg13g2_fill_1 FILLER_31_536 ();
 sg13g2_fill_2 FILLER_31_583 ();
 sg13g2_fill_2 FILLER_31_624 ();
 sg13g2_fill_1 FILLER_31_626 ();
 sg13g2_fill_2 FILLER_31_655 ();
 sg13g2_fill_2 FILLER_31_731 ();
 sg13g2_fill_1 FILLER_31_771 ();
 sg13g2_fill_2 FILLER_31_807 ();
 sg13g2_fill_2 FILLER_31_835 ();
 sg13g2_fill_1 FILLER_31_857 ();
 sg13g2_decap_4 FILLER_31_862 ();
 sg13g2_fill_2 FILLER_31_866 ();
 sg13g2_fill_2 FILLER_31_933 ();
 sg13g2_fill_1 FILLER_31_935 ();
 sg13g2_fill_2 FILLER_31_945 ();
 sg13g2_fill_1 FILLER_31_978 ();
 sg13g2_fill_1 FILLER_31_993 ();
 sg13g2_fill_1 FILLER_31_1020 ();
 sg13g2_fill_1 FILLER_31_1059 ();
 sg13g2_fill_2 FILLER_31_1086 ();
 sg13g2_fill_1 FILLER_31_1088 ();
 sg13g2_fill_1 FILLER_31_1097 ();
 sg13g2_fill_1 FILLER_31_1106 ();
 sg13g2_fill_1 FILLER_31_1116 ();
 sg13g2_fill_1 FILLER_31_1120 ();
 sg13g2_fill_2 FILLER_31_1184 ();
 sg13g2_fill_1 FILLER_31_1186 ();
 sg13g2_fill_1 FILLER_31_1201 ();
 sg13g2_fill_2 FILLER_31_1272 ();
 sg13g2_fill_2 FILLER_31_1295 ();
 sg13g2_decap_8 FILLER_31_1329 ();
 sg13g2_fill_2 FILLER_31_1336 ();
 sg13g2_fill_1 FILLER_31_1338 ();
 sg13g2_decap_8 FILLER_31_1347 ();
 sg13g2_decap_4 FILLER_31_1354 ();
 sg13g2_decap_8 FILLER_31_1370 ();
 sg13g2_fill_1 FILLER_31_1386 ();
 sg13g2_fill_2 FILLER_31_1391 ();
 sg13g2_fill_1 FILLER_31_1393 ();
 sg13g2_fill_2 FILLER_31_1403 ();
 sg13g2_fill_1 FILLER_31_1405 ();
 sg13g2_fill_1 FILLER_31_1414 ();
 sg13g2_fill_2 FILLER_31_1427 ();
 sg13g2_fill_1 FILLER_31_1438 ();
 sg13g2_fill_2 FILLER_31_1484 ();
 sg13g2_fill_2 FILLER_31_1505 ();
 sg13g2_fill_1 FILLER_31_1507 ();
 sg13g2_fill_2 FILLER_31_1516 ();
 sg13g2_fill_1 FILLER_31_1518 ();
 sg13g2_fill_2 FILLER_31_1528 ();
 sg13g2_fill_2 FILLER_31_1560 ();
 sg13g2_fill_1 FILLER_31_1562 ();
 sg13g2_decap_8 FILLER_31_1589 ();
 sg13g2_decap_4 FILLER_31_1596 ();
 sg13g2_fill_2 FILLER_31_1604 ();
 sg13g2_fill_1 FILLER_31_1633 ();
 sg13g2_fill_1 FILLER_31_1664 ();
 sg13g2_fill_1 FILLER_31_1673 ();
 sg13g2_fill_2 FILLER_31_1744 ();
 sg13g2_decap_8 FILLER_31_1785 ();
 sg13g2_decap_4 FILLER_31_1792 ();
 sg13g2_fill_2 FILLER_31_1879 ();
 sg13g2_fill_1 FILLER_31_1906 ();
 sg13g2_fill_2 FILLER_31_1926 ();
 sg13g2_fill_2 FILLER_31_1985 ();
 sg13g2_fill_2 FILLER_31_2017 ();
 sg13g2_decap_8 FILLER_31_2043 ();
 sg13g2_fill_2 FILLER_31_2050 ();
 sg13g2_decap_4 FILLER_31_2057 ();
 sg13g2_fill_1 FILLER_31_2061 ();
 sg13g2_fill_1 FILLER_31_2066 ();
 sg13g2_fill_2 FILLER_31_2081 ();
 sg13g2_fill_1 FILLER_31_2083 ();
 sg13g2_fill_1 FILLER_31_2107 ();
 sg13g2_fill_1 FILLER_31_2134 ();
 sg13g2_fill_1 FILLER_31_2161 ();
 sg13g2_fill_1 FILLER_31_2185 ();
 sg13g2_fill_2 FILLER_31_2225 ();
 sg13g2_fill_2 FILLER_31_2236 ();
 sg13g2_fill_1 FILLER_31_2238 ();
 sg13g2_fill_1 FILLER_31_2259 ();
 sg13g2_fill_2 FILLER_31_2265 ();
 sg13g2_fill_1 FILLER_31_2267 ();
 sg13g2_fill_1 FILLER_31_2307 ();
 sg13g2_fill_2 FILLER_31_2313 ();
 sg13g2_fill_2 FILLER_31_2355 ();
 sg13g2_fill_2 FILLER_31_2397 ();
 sg13g2_fill_1 FILLER_31_2399 ();
 sg13g2_fill_1 FILLER_31_2457 ();
 sg13g2_fill_2 FILLER_31_2494 ();
 sg13g2_fill_1 FILLER_31_2496 ();
 sg13g2_fill_2 FILLER_31_2532 ();
 sg13g2_fill_1 FILLER_31_2534 ();
 sg13g2_decap_8 FILLER_31_2570 ();
 sg13g2_decap_8 FILLER_31_2577 ();
 sg13g2_decap_8 FILLER_31_2584 ();
 sg13g2_decap_8 FILLER_31_2591 ();
 sg13g2_decap_8 FILLER_31_2598 ();
 sg13g2_decap_8 FILLER_31_2605 ();
 sg13g2_decap_8 FILLER_31_2612 ();
 sg13g2_decap_8 FILLER_31_2619 ();
 sg13g2_decap_8 FILLER_31_2626 ();
 sg13g2_decap_8 FILLER_31_2633 ();
 sg13g2_decap_8 FILLER_31_2640 ();
 sg13g2_decap_8 FILLER_31_2647 ();
 sg13g2_decap_8 FILLER_31_2654 ();
 sg13g2_decap_8 FILLER_31_2661 ();
 sg13g2_decap_4 FILLER_31_2668 ();
 sg13g2_fill_2 FILLER_31_2672 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_8 FILLER_32_434 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_8 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_469 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_fill_1 FILLER_32_511 ();
 sg13g2_fill_2 FILLER_32_547 ();
 sg13g2_fill_1 FILLER_32_557 ();
 sg13g2_fill_1 FILLER_32_577 ();
 sg13g2_fill_2 FILLER_32_618 ();
 sg13g2_fill_2 FILLER_32_632 ();
 sg13g2_fill_1 FILLER_32_634 ();
 sg13g2_fill_2 FILLER_32_644 ();
 sg13g2_fill_1 FILLER_32_699 ();
 sg13g2_fill_1 FILLER_32_712 ();
 sg13g2_fill_2 FILLER_32_734 ();
 sg13g2_fill_1 FILLER_32_736 ();
 sg13g2_fill_2 FILLER_32_741 ();
 sg13g2_fill_1 FILLER_32_747 ();
 sg13g2_fill_1 FILLER_32_756 ();
 sg13g2_decap_4 FILLER_32_771 ();
 sg13g2_fill_2 FILLER_32_775 ();
 sg13g2_fill_1 FILLER_32_782 ();
 sg13g2_fill_1 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_858 ();
 sg13g2_fill_2 FILLER_32_873 ();
 sg13g2_fill_2 FILLER_32_902 ();
 sg13g2_fill_1 FILLER_32_904 ();
 sg13g2_fill_1 FILLER_32_909 ();
 sg13g2_decap_4 FILLER_32_914 ();
 sg13g2_fill_2 FILLER_32_918 ();
 sg13g2_fill_2 FILLER_32_924 ();
 sg13g2_decap_8 FILLER_32_934 ();
 sg13g2_fill_1 FILLER_32_963 ();
 sg13g2_fill_2 FILLER_32_980 ();
 sg13g2_decap_4 FILLER_32_987 ();
 sg13g2_fill_1 FILLER_32_999 ();
 sg13g2_fill_2 FILLER_32_1013 ();
 sg13g2_fill_2 FILLER_32_1029 ();
 sg13g2_fill_1 FILLER_32_1052 ();
 sg13g2_fill_1 FILLER_32_1146 ();
 sg13g2_fill_2 FILLER_32_1190 ();
 sg13g2_fill_2 FILLER_32_1205 ();
 sg13g2_fill_1 FILLER_32_1207 ();
 sg13g2_fill_2 FILLER_32_1264 ();
 sg13g2_fill_2 FILLER_32_1310 ();
 sg13g2_fill_2 FILLER_32_1356 ();
 sg13g2_fill_1 FILLER_32_1358 ();
 sg13g2_fill_1 FILLER_32_1403 ();
 sg13g2_fill_1 FILLER_32_1426 ();
 sg13g2_fill_2 FILLER_32_1436 ();
 sg13g2_fill_2 FILLER_32_1481 ();
 sg13g2_fill_1 FILLER_32_1483 ();
 sg13g2_fill_2 FILLER_32_1586 ();
 sg13g2_fill_1 FILLER_32_1588 ();
 sg13g2_fill_2 FILLER_32_1615 ();
 sg13g2_fill_1 FILLER_32_1617 ();
 sg13g2_fill_2 FILLER_32_1648 ();
 sg13g2_fill_1 FILLER_32_1663 ();
 sg13g2_decap_8 FILLER_32_1787 ();
 sg13g2_fill_2 FILLER_32_1794 ();
 sg13g2_fill_1 FILLER_32_1796 ();
 sg13g2_fill_2 FILLER_32_1818 ();
 sg13g2_fill_2 FILLER_32_1847 ();
 sg13g2_fill_1 FILLER_32_1849 ();
 sg13g2_fill_2 FILLER_32_1870 ();
 sg13g2_fill_2 FILLER_32_1963 ();
 sg13g2_fill_1 FILLER_32_1992 ();
 sg13g2_fill_2 FILLER_32_2055 ();
 sg13g2_fill_1 FILLER_32_2057 ();
 sg13g2_fill_2 FILLER_32_2067 ();
 sg13g2_fill_1 FILLER_32_2069 ();
 sg13g2_fill_2 FILLER_32_2096 ();
 sg13g2_fill_1 FILLER_32_2142 ();
 sg13g2_fill_1 FILLER_32_2165 ();
 sg13g2_fill_1 FILLER_32_2179 ();
 sg13g2_fill_1 FILLER_32_2189 ();
 sg13g2_fill_1 FILLER_32_2210 ();
 sg13g2_fill_1 FILLER_32_2312 ();
 sg13g2_decap_4 FILLER_32_2364 ();
 sg13g2_fill_2 FILLER_32_2372 ();
 sg13g2_fill_2 FILLER_32_2502 ();
 sg13g2_fill_1 FILLER_32_2525 ();
 sg13g2_decap_8 FILLER_32_2565 ();
 sg13g2_decap_8 FILLER_32_2572 ();
 sg13g2_decap_8 FILLER_32_2579 ();
 sg13g2_decap_8 FILLER_32_2586 ();
 sg13g2_decap_8 FILLER_32_2593 ();
 sg13g2_decap_8 FILLER_32_2600 ();
 sg13g2_decap_8 FILLER_32_2607 ();
 sg13g2_decap_8 FILLER_32_2614 ();
 sg13g2_decap_8 FILLER_32_2621 ();
 sg13g2_decap_8 FILLER_32_2628 ();
 sg13g2_decap_8 FILLER_32_2635 ();
 sg13g2_decap_8 FILLER_32_2642 ();
 sg13g2_decap_8 FILLER_32_2649 ();
 sg13g2_decap_8 FILLER_32_2656 ();
 sg13g2_decap_8 FILLER_32_2663 ();
 sg13g2_decap_4 FILLER_32_2670 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_fill_1 FILLER_33_537 ();
 sg13g2_decap_4 FILLER_33_565 ();
 sg13g2_fill_1 FILLER_33_569 ();
 sg13g2_fill_2 FILLER_33_626 ();
 sg13g2_fill_1 FILLER_33_701 ();
 sg13g2_fill_2 FILLER_33_728 ();
 sg13g2_fill_2 FILLER_33_744 ();
 sg13g2_fill_1 FILLER_33_746 ();
 sg13g2_fill_2 FILLER_33_786 ();
 sg13g2_fill_1 FILLER_33_788 ();
 sg13g2_fill_1 FILLER_33_794 ();
 sg13g2_fill_2 FILLER_33_870 ();
 sg13g2_fill_1 FILLER_33_872 ();
 sg13g2_fill_2 FILLER_33_904 ();
 sg13g2_fill_1 FILLER_33_906 ();
 sg13g2_fill_2 FILLER_33_919 ();
 sg13g2_fill_1 FILLER_33_921 ();
 sg13g2_fill_2 FILLER_33_935 ();
 sg13g2_fill_1 FILLER_33_937 ();
 sg13g2_decap_4 FILLER_33_982 ();
 sg13g2_fill_2 FILLER_33_986 ();
 sg13g2_fill_2 FILLER_33_997 ();
 sg13g2_fill_1 FILLER_33_999 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_4 FILLER_33_1020 ();
 sg13g2_fill_2 FILLER_33_1064 ();
 sg13g2_fill_2 FILLER_33_1116 ();
 sg13g2_fill_1 FILLER_33_1158 ();
 sg13g2_fill_1 FILLER_33_1267 ();
 sg13g2_fill_2 FILLER_33_1323 ();
 sg13g2_fill_2 FILLER_33_1392 ();
 sg13g2_fill_1 FILLER_33_1394 ();
 sg13g2_fill_1 FILLER_33_1452 ();
 sg13g2_fill_2 FILLER_33_1490 ();
 sg13g2_fill_1 FILLER_33_1492 ();
 sg13g2_fill_1 FILLER_33_1506 ();
 sg13g2_fill_1 FILLER_33_1550 ();
 sg13g2_fill_2 FILLER_33_1584 ();
 sg13g2_fill_1 FILLER_33_1687 ();
 sg13g2_fill_2 FILLER_33_1714 ();
 sg13g2_fill_1 FILLER_33_1737 ();
 sg13g2_fill_1 FILLER_33_1764 ();
 sg13g2_decap_4 FILLER_33_1794 ();
 sg13g2_fill_1 FILLER_33_1798 ();
 sg13g2_fill_1 FILLER_33_1820 ();
 sg13g2_fill_2 FILLER_33_1834 ();
 sg13g2_fill_1 FILLER_33_1836 ();
 sg13g2_fill_1 FILLER_33_1851 ();
 sg13g2_fill_2 FILLER_33_1868 ();
 sg13g2_decap_4 FILLER_33_1884 ();
 sg13g2_fill_1 FILLER_33_1888 ();
 sg13g2_fill_1 FILLER_33_1893 ();
 sg13g2_fill_2 FILLER_33_1899 ();
 sg13g2_fill_1 FILLER_33_1901 ();
 sg13g2_fill_1 FILLER_33_1951 ();
 sg13g2_decap_8 FILLER_33_1960 ();
 sg13g2_fill_2 FILLER_33_1967 ();
 sg13g2_fill_1 FILLER_33_1969 ();
 sg13g2_fill_1 FILLER_33_2005 ();
 sg13g2_fill_1 FILLER_33_2011 ();
 sg13g2_fill_1 FILLER_33_2028 ();
 sg13g2_decap_4 FILLER_33_2124 ();
 sg13g2_fill_1 FILLER_33_2128 ();
 sg13g2_decap_8 FILLER_33_2134 ();
 sg13g2_fill_1 FILLER_33_2141 ();
 sg13g2_fill_1 FILLER_33_2160 ();
 sg13g2_fill_1 FILLER_33_2174 ();
 sg13g2_fill_2 FILLER_33_2201 ();
 sg13g2_fill_1 FILLER_33_2203 ();
 sg13g2_fill_2 FILLER_33_2230 ();
 sg13g2_fill_2 FILLER_33_2241 ();
 sg13g2_fill_1 FILLER_33_2243 ();
 sg13g2_fill_2 FILLER_33_2249 ();
 sg13g2_fill_2 FILLER_33_2321 ();
 sg13g2_decap_8 FILLER_33_2357 ();
 sg13g2_decap_8 FILLER_33_2369 ();
 sg13g2_fill_2 FILLER_33_2376 ();
 sg13g2_fill_2 FILLER_33_2396 ();
 sg13g2_fill_1 FILLER_33_2398 ();
 sg13g2_decap_4 FILLER_33_2430 ();
 sg13g2_fill_1 FILLER_33_2434 ();
 sg13g2_fill_2 FILLER_33_2439 ();
 sg13g2_fill_2 FILLER_33_2493 ();
 sg13g2_fill_1 FILLER_33_2495 ();
 sg13g2_fill_1 FILLER_33_2510 ();
 sg13g2_fill_2 FILLER_33_2525 ();
 sg13g2_fill_1 FILLER_33_2527 ();
 sg13g2_decap_8 FILLER_33_2561 ();
 sg13g2_decap_8 FILLER_33_2568 ();
 sg13g2_decap_8 FILLER_33_2575 ();
 sg13g2_decap_8 FILLER_33_2582 ();
 sg13g2_decap_8 FILLER_33_2589 ();
 sg13g2_decap_8 FILLER_33_2596 ();
 sg13g2_decap_8 FILLER_33_2603 ();
 sg13g2_decap_8 FILLER_33_2610 ();
 sg13g2_decap_8 FILLER_33_2617 ();
 sg13g2_decap_8 FILLER_33_2624 ();
 sg13g2_decap_8 FILLER_33_2631 ();
 sg13g2_decap_8 FILLER_33_2638 ();
 sg13g2_decap_8 FILLER_33_2645 ();
 sg13g2_decap_8 FILLER_33_2652 ();
 sg13g2_decap_8 FILLER_33_2659 ();
 sg13g2_decap_8 FILLER_33_2666 ();
 sg13g2_fill_1 FILLER_33_2673 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_decap_8 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_8 FILLER_34_483 ();
 sg13g2_decap_8 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_497 ();
 sg13g2_fill_2 FILLER_34_538 ();
 sg13g2_fill_2 FILLER_34_579 ();
 sg13g2_fill_1 FILLER_34_581 ();
 sg13g2_fill_2 FILLER_34_586 ();
 sg13g2_fill_2 FILLER_34_598 ();
 sg13g2_fill_1 FILLER_34_654 ();
 sg13g2_fill_1 FILLER_34_669 ();
 sg13g2_fill_1 FILLER_34_678 ();
 sg13g2_fill_2 FILLER_34_684 ();
 sg13g2_fill_1 FILLER_34_691 ();
 sg13g2_fill_2 FILLER_34_697 ();
 sg13g2_fill_2 FILLER_34_755 ();
 sg13g2_decap_4 FILLER_34_790 ();
 sg13g2_fill_2 FILLER_34_803 ();
 sg13g2_fill_1 FILLER_34_835 ();
 sg13g2_fill_2 FILLER_34_970 ();
 sg13g2_fill_2 FILLER_34_998 ();
 sg13g2_fill_1 FILLER_34_1000 ();
 sg13g2_fill_1 FILLER_34_1007 ();
 sg13g2_fill_1 FILLER_34_1016 ();
 sg13g2_fill_1 FILLER_34_1026 ();
 sg13g2_fill_2 FILLER_34_1074 ();
 sg13g2_fill_1 FILLER_34_1076 ();
 sg13g2_fill_1 FILLER_34_1096 ();
 sg13g2_fill_2 FILLER_34_1140 ();
 sg13g2_fill_2 FILLER_34_1151 ();
 sg13g2_fill_1 FILLER_34_1153 ();
 sg13g2_fill_1 FILLER_34_1176 ();
 sg13g2_fill_2 FILLER_34_1185 ();
 sg13g2_fill_1 FILLER_34_1187 ();
 sg13g2_fill_2 FILLER_34_1289 ();
 sg13g2_fill_1 FILLER_34_1317 ();
 sg13g2_fill_2 FILLER_34_1386 ();
 sg13g2_fill_1 FILLER_34_1388 ();
 sg13g2_fill_1 FILLER_34_1429 ();
 sg13g2_fill_2 FILLER_34_1440 ();
 sg13g2_fill_1 FILLER_34_1451 ();
 sg13g2_fill_2 FILLER_34_1499 ();
 sg13g2_fill_1 FILLER_34_1501 ();
 sg13g2_fill_2 FILLER_34_1508 ();
 sg13g2_fill_1 FILLER_34_1510 ();
 sg13g2_fill_2 FILLER_34_1516 ();
 sg13g2_fill_2 FILLER_34_1528 ();
 sg13g2_fill_2 FILLER_34_1538 ();
 sg13g2_fill_2 FILLER_34_1548 ();
 sg13g2_fill_1 FILLER_34_1550 ();
 sg13g2_decap_4 FILLER_34_1589 ();
 sg13g2_fill_1 FILLER_34_1598 ();
 sg13g2_fill_2 FILLER_34_1604 ();
 sg13g2_fill_1 FILLER_34_1670 ();
 sg13g2_fill_2 FILLER_34_1697 ();
 sg13g2_fill_2 FILLER_34_1738 ();
 sg13g2_fill_1 FILLER_34_1764 ();
 sg13g2_fill_2 FILLER_34_1796 ();
 sg13g2_fill_2 FILLER_34_1886 ();
 sg13g2_decap_8 FILLER_34_1942 ();
 sg13g2_decap_8 FILLER_34_1949 ();
 sg13g2_fill_2 FILLER_34_1982 ();
 sg13g2_fill_1 FILLER_34_1984 ();
 sg13g2_fill_2 FILLER_34_2068 ();
 sg13g2_decap_8 FILLER_34_2119 ();
 sg13g2_decap_4 FILLER_34_2136 ();
 sg13g2_fill_2 FILLER_34_2150 ();
 sg13g2_fill_2 FILLER_34_2157 ();
 sg13g2_fill_2 FILLER_34_2172 ();
 sg13g2_fill_1 FILLER_34_2234 ();
 sg13g2_fill_1 FILLER_34_2253 ();
 sg13g2_fill_2 FILLER_34_2275 ();
 sg13g2_fill_2 FILLER_34_2295 ();
 sg13g2_fill_1 FILLER_34_2297 ();
 sg13g2_fill_1 FILLER_34_2320 ();
 sg13g2_fill_2 FILLER_34_2325 ();
 sg13g2_decap_8 FILLER_34_2344 ();
 sg13g2_fill_2 FILLER_34_2351 ();
 sg13g2_fill_2 FILLER_34_2357 ();
 sg13g2_fill_1 FILLER_34_2359 ();
 sg13g2_fill_1 FILLER_34_2379 ();
 sg13g2_decap_8 FILLER_34_2401 ();
 sg13g2_decap_4 FILLER_34_2408 ();
 sg13g2_fill_2 FILLER_34_2412 ();
 sg13g2_decap_4 FILLER_34_2422 ();
 sg13g2_fill_1 FILLER_34_2426 ();
 sg13g2_fill_1 FILLER_34_2449 ();
 sg13g2_fill_2 FILLER_34_2454 ();
 sg13g2_fill_1 FILLER_34_2456 ();
 sg13g2_fill_1 FILLER_34_2498 ();
 sg13g2_fill_1 FILLER_34_2525 ();
 sg13g2_decap_8 FILLER_34_2568 ();
 sg13g2_decap_8 FILLER_34_2575 ();
 sg13g2_decap_8 FILLER_34_2582 ();
 sg13g2_decap_8 FILLER_34_2589 ();
 sg13g2_decap_8 FILLER_34_2596 ();
 sg13g2_decap_8 FILLER_34_2603 ();
 sg13g2_decap_8 FILLER_34_2610 ();
 sg13g2_decap_8 FILLER_34_2617 ();
 sg13g2_decap_8 FILLER_34_2624 ();
 sg13g2_decap_8 FILLER_34_2631 ();
 sg13g2_decap_8 FILLER_34_2638 ();
 sg13g2_decap_8 FILLER_34_2645 ();
 sg13g2_decap_8 FILLER_34_2652 ();
 sg13g2_decap_8 FILLER_34_2659 ();
 sg13g2_decap_8 FILLER_34_2666 ();
 sg13g2_fill_1 FILLER_34_2673 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_decap_8 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_fill_2 FILLER_35_511 ();
 sg13g2_fill_1 FILLER_35_513 ();
 sg13g2_fill_2 FILLER_35_533 ();
 sg13g2_fill_1 FILLER_35_565 ();
 sg13g2_fill_2 FILLER_35_575 ();
 sg13g2_fill_2 FILLER_35_586 ();
 sg13g2_fill_1 FILLER_35_592 ();
 sg13g2_fill_1 FILLER_35_626 ();
 sg13g2_fill_1 FILLER_35_679 ();
 sg13g2_fill_2 FILLER_35_688 ();
 sg13g2_fill_1 FILLER_35_690 ();
 sg13g2_fill_1 FILLER_35_695 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_fill_2 FILLER_35_747 ();
 sg13g2_decap_8 FILLER_35_807 ();
 sg13g2_fill_2 FILLER_35_814 ();
 sg13g2_decap_4 FILLER_35_820 ();
 sg13g2_fill_1 FILLER_35_824 ();
 sg13g2_fill_1 FILLER_35_833 ();
 sg13g2_fill_2 FILLER_35_872 ();
 sg13g2_fill_2 FILLER_35_879 ();
 sg13g2_fill_1 FILLER_35_881 ();
 sg13g2_fill_1 FILLER_35_891 ();
 sg13g2_fill_1 FILLER_35_906 ();
 sg13g2_fill_1 FILLER_35_926 ();
 sg13g2_fill_1 FILLER_35_956 ();
 sg13g2_fill_1 FILLER_35_967 ();
 sg13g2_fill_2 FILLER_35_989 ();
 sg13g2_fill_1 FILLER_35_991 ();
 sg13g2_fill_2 FILLER_35_1027 ();
 sg13g2_fill_2 FILLER_35_1037 ();
 sg13g2_fill_1 FILLER_35_1039 ();
 sg13g2_fill_1 FILLER_35_1044 ();
 sg13g2_fill_2 FILLER_35_1068 ();
 sg13g2_fill_2 FILLER_35_1100 ();
 sg13g2_fill_1 FILLER_35_1118 ();
 sg13g2_fill_2 FILLER_35_1129 ();
 sg13g2_decap_8 FILLER_35_1183 ();
 sg13g2_decap_4 FILLER_35_1190 ();
 sg13g2_fill_1 FILLER_35_1194 ();
 sg13g2_decap_4 FILLER_35_1251 ();
 sg13g2_fill_1 FILLER_35_1262 ();
 sg13g2_fill_1 FILLER_35_1272 ();
 sg13g2_decap_4 FILLER_35_1333 ();
 sg13g2_fill_2 FILLER_35_1337 ();
 sg13g2_fill_1 FILLER_35_1352 ();
 sg13g2_fill_2 FILLER_35_1410 ();
 sg13g2_fill_1 FILLER_35_1412 ();
 sg13g2_fill_2 FILLER_35_1430 ();
 sg13g2_fill_2 FILLER_35_1458 ();
 sg13g2_fill_2 FILLER_35_1474 ();
 sg13g2_fill_1 FILLER_35_1532 ();
 sg13g2_decap_8 FILLER_35_1592 ();
 sg13g2_fill_2 FILLER_35_1599 ();
 sg13g2_fill_1 FILLER_35_1610 ();
 sg13g2_fill_2 FILLER_35_1628 ();
 sg13g2_fill_2 FILLER_35_1635 ();
 sg13g2_fill_1 FILLER_35_1642 ();
 sg13g2_fill_2 FILLER_35_1690 ();
 sg13g2_fill_1 FILLER_35_1797 ();
 sg13g2_fill_2 FILLER_35_1850 ();
 sg13g2_fill_1 FILLER_35_1852 ();
 sg13g2_decap_8 FILLER_35_1942 ();
 sg13g2_fill_2 FILLER_35_1949 ();
 sg13g2_fill_1 FILLER_35_1951 ();
 sg13g2_fill_2 FILLER_35_2007 ();
 sg13g2_fill_2 FILLER_35_2062 ();
 sg13g2_fill_2 FILLER_35_2068 ();
 sg13g2_fill_1 FILLER_35_2070 ();
 sg13g2_fill_2 FILLER_35_2075 ();
 sg13g2_fill_1 FILLER_35_2077 ();
 sg13g2_fill_2 FILLER_35_2082 ();
 sg13g2_decap_4 FILLER_35_2115 ();
 sg13g2_fill_2 FILLER_35_2141 ();
 sg13g2_fill_2 FILLER_35_2169 ();
 sg13g2_fill_1 FILLER_35_2183 ();
 sg13g2_fill_1 FILLER_35_2197 ();
 sg13g2_fill_2 FILLER_35_2203 ();
 sg13g2_fill_1 FILLER_35_2215 ();
 sg13g2_fill_2 FILLER_35_2235 ();
 sg13g2_fill_1 FILLER_35_2237 ();
 sg13g2_decap_8 FILLER_35_2264 ();
 sg13g2_decap_4 FILLER_35_2271 ();
 sg13g2_decap_8 FILLER_35_2295 ();
 sg13g2_decap_8 FILLER_35_2302 ();
 sg13g2_fill_2 FILLER_35_2309 ();
 sg13g2_fill_1 FILLER_35_2311 ();
 sg13g2_fill_2 FILLER_35_2321 ();
 sg13g2_decap_8 FILLER_35_2332 ();
 sg13g2_decap_4 FILLER_35_2365 ();
 sg13g2_fill_1 FILLER_35_2390 ();
 sg13g2_fill_2 FILLER_35_2417 ();
 sg13g2_fill_1 FILLER_35_2419 ();
 sg13g2_fill_1 FILLER_35_2453 ();
 sg13g2_fill_1 FILLER_35_2544 ();
 sg13g2_decap_8 FILLER_35_2580 ();
 sg13g2_decap_8 FILLER_35_2587 ();
 sg13g2_decap_8 FILLER_35_2594 ();
 sg13g2_decap_8 FILLER_35_2601 ();
 sg13g2_decap_8 FILLER_35_2608 ();
 sg13g2_decap_8 FILLER_35_2615 ();
 sg13g2_decap_8 FILLER_35_2622 ();
 sg13g2_decap_8 FILLER_35_2629 ();
 sg13g2_decap_8 FILLER_35_2636 ();
 sg13g2_decap_8 FILLER_35_2643 ();
 sg13g2_decap_8 FILLER_35_2650 ();
 sg13g2_decap_8 FILLER_35_2657 ();
 sg13g2_decap_8 FILLER_35_2664 ();
 sg13g2_fill_2 FILLER_35_2671 ();
 sg13g2_fill_1 FILLER_35_2673 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_8 FILLER_36_448 ();
 sg13g2_decap_8 FILLER_36_455 ();
 sg13g2_decap_8 FILLER_36_462 ();
 sg13g2_decap_8 FILLER_36_469 ();
 sg13g2_decap_8 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_483 ();
 sg13g2_decap_8 FILLER_36_490 ();
 sg13g2_decap_8 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_decap_4 FILLER_36_511 ();
 sg13g2_fill_2 FILLER_36_515 ();
 sg13g2_fill_1 FILLER_36_539 ();
 sg13g2_fill_2 FILLER_36_549 ();
 sg13g2_fill_2 FILLER_36_607 ();
 sg13g2_fill_1 FILLER_36_622 ();
 sg13g2_fill_2 FILLER_36_627 ();
 sg13g2_fill_1 FILLER_36_629 ();
 sg13g2_fill_1 FILLER_36_661 ();
 sg13g2_fill_1 FILLER_36_668 ();
 sg13g2_decap_8 FILLER_36_699 ();
 sg13g2_decap_4 FILLER_36_706 ();
 sg13g2_fill_2 FILLER_36_710 ();
 sg13g2_fill_2 FILLER_36_742 ();
 sg13g2_fill_1 FILLER_36_744 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_fill_1 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_816 ();
 sg13g2_fill_1 FILLER_36_857 ();
 sg13g2_fill_1 FILLER_36_867 ();
 sg13g2_fill_2 FILLER_36_908 ();
 sg13g2_fill_1 FILLER_36_910 ();
 sg13g2_fill_2 FILLER_36_929 ();
 sg13g2_fill_1 FILLER_36_953 ();
 sg13g2_fill_2 FILLER_36_964 ();
 sg13g2_fill_2 FILLER_36_1001 ();
 sg13g2_fill_1 FILLER_36_1003 ();
 sg13g2_fill_1 FILLER_36_1043 ();
 sg13g2_fill_2 FILLER_36_1070 ();
 sg13g2_fill_1 FILLER_36_1077 ();
 sg13g2_fill_2 FILLER_36_1102 ();
 sg13g2_decap_4 FILLER_36_1189 ();
 sg13g2_fill_2 FILLER_36_1193 ();
 sg13g2_fill_1 FILLER_36_1205 ();
 sg13g2_fill_1 FILLER_36_1232 ();
 sg13g2_fill_2 FILLER_36_1242 ();
 sg13g2_fill_1 FILLER_36_1244 ();
 sg13g2_fill_2 FILLER_36_1251 ();
 sg13g2_fill_1 FILLER_36_1253 ();
 sg13g2_decap_8 FILLER_36_1262 ();
 sg13g2_decap_8 FILLER_36_1273 ();
 sg13g2_fill_1 FILLER_36_1307 ();
 sg13g2_fill_1 FILLER_36_1317 ();
 sg13g2_decap_8 FILLER_36_1326 ();
 sg13g2_decap_8 FILLER_36_1333 ();
 sg13g2_decap_4 FILLER_36_1340 ();
 sg13g2_fill_2 FILLER_36_1344 ();
 sg13g2_fill_2 FILLER_36_1354 ();
 sg13g2_fill_1 FILLER_36_1356 ();
 sg13g2_fill_2 FILLER_36_1366 ();
 sg13g2_fill_1 FILLER_36_1368 ();
 sg13g2_decap_4 FILLER_36_1373 ();
 sg13g2_fill_2 FILLER_36_1381 ();
 sg13g2_decap_8 FILLER_36_1419 ();
 sg13g2_decap_4 FILLER_36_1426 ();
 sg13g2_decap_8 FILLER_36_1434 ();
 sg13g2_fill_1 FILLER_36_1479 ();
 sg13g2_fill_1 FILLER_36_1515 ();
 sg13g2_fill_2 FILLER_36_1524 ();
 sg13g2_fill_1 FILLER_36_1526 ();
 sg13g2_fill_2 FILLER_36_1582 ();
 sg13g2_fill_1 FILLER_36_1584 ();
 sg13g2_fill_2 FILLER_36_1598 ();
 sg13g2_fill_1 FILLER_36_1600 ();
 sg13g2_fill_2 FILLER_36_1620 ();
 sg13g2_fill_1 FILLER_36_1622 ();
 sg13g2_fill_2 FILLER_36_1628 ();
 sg13g2_fill_2 FILLER_36_1635 ();
 sg13g2_fill_2 FILLER_36_1642 ();
 sg13g2_fill_1 FILLER_36_1644 ();
 sg13g2_fill_2 FILLER_36_1686 ();
 sg13g2_fill_1 FILLER_36_1721 ();
 sg13g2_fill_2 FILLER_36_1757 ();
 sg13g2_decap_8 FILLER_36_1793 ();
 sg13g2_fill_2 FILLER_36_1800 ();
 sg13g2_fill_1 FILLER_36_1802 ();
 sg13g2_fill_2 FILLER_36_1817 ();
 sg13g2_fill_2 FILLER_36_1838 ();
 sg13g2_fill_1 FILLER_36_1840 ();
 sg13g2_fill_1 FILLER_36_1850 ();
 sg13g2_fill_2 FILLER_36_1908 ();
 sg13g2_fill_1 FILLER_36_1910 ();
 sg13g2_fill_1 FILLER_36_1960 ();
 sg13g2_fill_2 FILLER_36_1992 ();
 sg13g2_fill_1 FILLER_36_1994 ();
 sg13g2_fill_2 FILLER_36_2020 ();
 sg13g2_fill_2 FILLER_36_2056 ();
 sg13g2_fill_1 FILLER_36_2058 ();
 sg13g2_decap_4 FILLER_36_2068 ();
 sg13g2_fill_2 FILLER_36_2072 ();
 sg13g2_fill_2 FILLER_36_2084 ();
 sg13g2_fill_1 FILLER_36_2086 ();
 sg13g2_fill_1 FILLER_36_2133 ();
 sg13g2_fill_1 FILLER_36_2173 ();
 sg13g2_fill_2 FILLER_36_2203 ();
 sg13g2_fill_2 FILLER_36_2242 ();
 sg13g2_fill_1 FILLER_36_2244 ();
 sg13g2_fill_2 FILLER_36_2275 ();
 sg13g2_decap_8 FILLER_36_2282 ();
 sg13g2_decap_8 FILLER_36_2289 ();
 sg13g2_fill_2 FILLER_36_2296 ();
 sg13g2_fill_1 FILLER_36_2298 ();
 sg13g2_fill_1 FILLER_36_2351 ();
 sg13g2_fill_1 FILLER_36_2404 ();
 sg13g2_fill_1 FILLER_36_2440 ();
 sg13g2_fill_1 FILLER_36_2495 ();
 sg13g2_fill_2 FILLER_36_2531 ();
 sg13g2_fill_1 FILLER_36_2533 ();
 sg13g2_fill_2 FILLER_36_2544 ();
 sg13g2_decap_8 FILLER_36_2582 ();
 sg13g2_decap_8 FILLER_36_2589 ();
 sg13g2_decap_8 FILLER_36_2596 ();
 sg13g2_decap_8 FILLER_36_2603 ();
 sg13g2_decap_8 FILLER_36_2610 ();
 sg13g2_decap_8 FILLER_36_2617 ();
 sg13g2_decap_8 FILLER_36_2624 ();
 sg13g2_decap_8 FILLER_36_2631 ();
 sg13g2_decap_8 FILLER_36_2638 ();
 sg13g2_decap_8 FILLER_36_2645 ();
 sg13g2_decap_8 FILLER_36_2652 ();
 sg13g2_decap_8 FILLER_36_2659 ();
 sg13g2_decap_8 FILLER_36_2666 ();
 sg13g2_fill_1 FILLER_36_2673 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_fill_2 FILLER_37_511 ();
 sg13g2_fill_1 FILLER_37_513 ();
 sg13g2_fill_2 FILLER_37_540 ();
 sg13g2_fill_2 FILLER_37_560 ();
 sg13g2_fill_2 FILLER_37_623 ();
 sg13g2_decap_4 FILLER_37_639 ();
 sg13g2_fill_1 FILLER_37_643 ();
 sg13g2_fill_2 FILLER_37_655 ();
 sg13g2_fill_1 FILLER_37_673 ();
 sg13g2_decap_8 FILLER_37_713 ();
 sg13g2_fill_2 FILLER_37_720 ();
 sg13g2_fill_1 FILLER_37_722 ();
 sg13g2_fill_2 FILLER_37_735 ();
 sg13g2_fill_2 FILLER_37_746 ();
 sg13g2_decap_4 FILLER_37_773 ();
 sg13g2_fill_2 FILLER_37_781 ();
 sg13g2_fill_1 FILLER_37_783 ();
 sg13g2_fill_1 FILLER_37_819 ();
 sg13g2_fill_2 FILLER_37_864 ();
 sg13g2_fill_1 FILLER_37_866 ();
 sg13g2_fill_2 FILLER_37_931 ();
 sg13g2_fill_1 FILLER_37_933 ();
 sg13g2_fill_2 FILLER_37_978 ();
 sg13g2_fill_2 FILLER_37_1000 ();
 sg13g2_fill_1 FILLER_37_1002 ();
 sg13g2_fill_1 FILLER_37_1011 ();
 sg13g2_fill_2 FILLER_37_1036 ();
 sg13g2_fill_1 FILLER_37_1141 ();
 sg13g2_fill_2 FILLER_37_1156 ();
 sg13g2_fill_2 FILLER_37_1163 ();
 sg13g2_fill_1 FILLER_37_1165 ();
 sg13g2_fill_2 FILLER_37_1174 ();
 sg13g2_fill_2 FILLER_37_1185 ();
 sg13g2_decap_4 FILLER_37_1193 ();
 sg13g2_decap_8 FILLER_37_1254 ();
 sg13g2_fill_1 FILLER_37_1261 ();
 sg13g2_decap_8 FILLER_37_1266 ();
 sg13g2_fill_2 FILLER_37_1273 ();
 sg13g2_decap_4 FILLER_37_1285 ();
 sg13g2_decap_8 FILLER_37_1297 ();
 sg13g2_decap_4 FILLER_37_1304 ();
 sg13g2_fill_1 FILLER_37_1311 ();
 sg13g2_decap_8 FILLER_37_1316 ();
 sg13g2_fill_1 FILLER_37_1323 ();
 sg13g2_fill_2 FILLER_37_1329 ();
 sg13g2_fill_1 FILLER_37_1339 ();
 sg13g2_decap_4 FILLER_37_1349 ();
 sg13g2_fill_1 FILLER_37_1353 ();
 sg13g2_decap_8 FILLER_37_1362 ();
 sg13g2_decap_8 FILLER_37_1369 ();
 sg13g2_decap_8 FILLER_37_1376 ();
 sg13g2_decap_4 FILLER_37_1383 ();
 sg13g2_fill_1 FILLER_37_1387 ();
 sg13g2_decap_8 FILLER_37_1400 ();
 sg13g2_decap_8 FILLER_37_1407 ();
 sg13g2_fill_2 FILLER_37_1414 ();
 sg13g2_decap_4 FILLER_37_1429 ();
 sg13g2_fill_1 FILLER_37_1433 ();
 sg13g2_fill_2 FILLER_37_1469 ();
 sg13g2_decap_8 FILLER_37_1476 ();
 sg13g2_fill_2 FILLER_37_1483 ();
 sg13g2_fill_2 FILLER_37_1503 ();
 sg13g2_fill_1 FILLER_37_1505 ();
 sg13g2_decap_4 FILLER_37_1510 ();
 sg13g2_fill_1 FILLER_37_1514 ();
 sg13g2_decap_4 FILLER_37_1521 ();
 sg13g2_fill_1 FILLER_37_1525 ();
 sg13g2_fill_2 FILLER_37_1544 ();
 sg13g2_decap_8 FILLER_37_1580 ();
 sg13g2_fill_2 FILLER_37_1587 ();
 sg13g2_fill_1 FILLER_37_1589 ();
 sg13g2_fill_1 FILLER_37_1681 ();
 sg13g2_fill_1 FILLER_37_1722 ();
 sg13g2_decap_8 FILLER_37_1795 ();
 sg13g2_fill_1 FILLER_37_1802 ();
 sg13g2_decap_8 FILLER_37_1808 ();
 sg13g2_fill_1 FILLER_37_1815 ();
 sg13g2_decap_4 FILLER_37_1825 ();
 sg13g2_fill_2 FILLER_37_1829 ();
 sg13g2_fill_2 FILLER_37_1860 ();
 sg13g2_fill_1 FILLER_37_1894 ();
 sg13g2_fill_1 FILLER_37_1921 ();
 sg13g2_fill_1 FILLER_37_1926 ();
 sg13g2_fill_1 FILLER_37_1985 ();
 sg13g2_fill_2 FILLER_37_2016 ();
 sg13g2_fill_1 FILLER_37_2018 ();
 sg13g2_fill_1 FILLER_37_2123 ();
 sg13g2_fill_1 FILLER_37_2136 ();
 sg13g2_fill_1 FILLER_37_2234 ();
 sg13g2_decap_4 FILLER_37_2274 ();
 sg13g2_fill_1 FILLER_37_2278 ();
 sg13g2_decap_4 FILLER_37_2288 ();
 sg13g2_fill_2 FILLER_37_2318 ();
 sg13g2_fill_2 FILLER_37_2338 ();
 sg13g2_fill_1 FILLER_37_2354 ();
 sg13g2_fill_2 FILLER_37_2386 ();
 sg13g2_fill_2 FILLER_37_2398 ();
 sg13g2_fill_2 FILLER_37_2451 ();
 sg13g2_fill_1 FILLER_37_2468 ();
 sg13g2_fill_1 FILLER_37_2517 ();
 sg13g2_fill_2 FILLER_37_2527 ();
 sg13g2_fill_1 FILLER_37_2542 ();
 sg13g2_fill_2 FILLER_37_2548 ();
 sg13g2_fill_1 FILLER_37_2550 ();
 sg13g2_decap_8 FILLER_37_2590 ();
 sg13g2_decap_8 FILLER_37_2597 ();
 sg13g2_decap_8 FILLER_37_2604 ();
 sg13g2_decap_8 FILLER_37_2611 ();
 sg13g2_decap_8 FILLER_37_2618 ();
 sg13g2_decap_8 FILLER_37_2625 ();
 sg13g2_decap_8 FILLER_37_2632 ();
 sg13g2_decap_8 FILLER_37_2639 ();
 sg13g2_decap_8 FILLER_37_2646 ();
 sg13g2_decap_8 FILLER_37_2653 ();
 sg13g2_decap_8 FILLER_37_2660 ();
 sg13g2_decap_8 FILLER_37_2667 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_441 ();
 sg13g2_decap_8 FILLER_38_448 ();
 sg13g2_decap_8 FILLER_38_455 ();
 sg13g2_decap_8 FILLER_38_462 ();
 sg13g2_decap_8 FILLER_38_469 ();
 sg13g2_decap_8 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_decap_8 FILLER_38_497 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_fill_1 FILLER_38_511 ();
 sg13g2_fill_1 FILLER_38_578 ();
 sg13g2_fill_1 FILLER_38_619 ();
 sg13g2_fill_1 FILLER_38_657 ();
 sg13g2_fill_2 FILLER_38_666 ();
 sg13g2_fill_1 FILLER_38_668 ();
 sg13g2_fill_2 FILLER_38_674 ();
 sg13g2_fill_2 FILLER_38_718 ();
 sg13g2_fill_1 FILLER_38_720 ();
 sg13g2_decap_8 FILLER_38_725 ();
 sg13g2_fill_1 FILLER_38_732 ();
 sg13g2_decap_8 FILLER_38_741 ();
 sg13g2_decap_8 FILLER_38_748 ();
 sg13g2_decap_4 FILLER_38_755 ();
 sg13g2_fill_2 FILLER_38_759 ();
 sg13g2_decap_8 FILLER_38_765 ();
 sg13g2_decap_4 FILLER_38_776 ();
 sg13g2_fill_2 FILLER_38_780 ();
 sg13g2_decap_8 FILLER_38_808 ();
 sg13g2_fill_1 FILLER_38_831 ();
 sg13g2_fill_2 FILLER_38_876 ();
 sg13g2_fill_1 FILLER_38_878 ();
 sg13g2_fill_1 FILLER_38_914 ();
 sg13g2_fill_2 FILLER_38_941 ();
 sg13g2_decap_4 FILLER_38_1012 ();
 sg13g2_fill_1 FILLER_38_1032 ();
 sg13g2_fill_2 FILLER_38_1068 ();
 sg13g2_fill_2 FILLER_38_1092 ();
 sg13g2_fill_1 FILLER_38_1094 ();
 sg13g2_fill_1 FILLER_38_1100 ();
 sg13g2_fill_2 FILLER_38_1104 ();
 sg13g2_fill_1 FILLER_38_1106 ();
 sg13g2_fill_2 FILLER_38_1129 ();
 sg13g2_fill_1 FILLER_38_1131 ();
 sg13g2_decap_8 FILLER_38_1160 ();
 sg13g2_decap_4 FILLER_38_1167 ();
 sg13g2_fill_1 FILLER_38_1171 ();
 sg13g2_fill_2 FILLER_38_1187 ();
 sg13g2_fill_2 FILLER_38_1224 ();
 sg13g2_fill_1 FILLER_38_1226 ();
 sg13g2_fill_2 FILLER_38_1259 ();
 sg13g2_fill_2 FILLER_38_1267 ();
 sg13g2_decap_4 FILLER_38_1291 ();
 sg13g2_fill_2 FILLER_38_1295 ();
 sg13g2_fill_2 FILLER_38_1339 ();
 sg13g2_fill_1 FILLER_38_1341 ();
 sg13g2_decap_4 FILLER_38_1355 ();
 sg13g2_fill_1 FILLER_38_1359 ();
 sg13g2_fill_2 FILLER_38_1378 ();
 sg13g2_decap_8 FILLER_38_1386 ();
 sg13g2_decap_4 FILLER_38_1393 ();
 sg13g2_decap_4 FILLER_38_1423 ();
 sg13g2_fill_1 FILLER_38_1427 ();
 sg13g2_decap_4 FILLER_38_1468 ();
 sg13g2_fill_1 FILLER_38_1472 ();
 sg13g2_decap_4 FILLER_38_1483 ();
 sg13g2_fill_2 FILLER_38_1505 ();
 sg13g2_fill_2 FILLER_38_1533 ();
 sg13g2_fill_1 FILLER_38_1535 ();
 sg13g2_fill_1 FILLER_38_1546 ();
 sg13g2_fill_2 FILLER_38_1557 ();
 sg13g2_fill_1 FILLER_38_1559 ();
 sg13g2_decap_8 FILLER_38_1573 ();
 sg13g2_decap_8 FILLER_38_1580 ();
 sg13g2_fill_1 FILLER_38_1587 ();
 sg13g2_fill_2 FILLER_38_1641 ();
 sg13g2_fill_1 FILLER_38_1643 ();
 sg13g2_fill_2 FILLER_38_1744 ();
 sg13g2_fill_1 FILLER_38_1767 ();
 sg13g2_decap_4 FILLER_38_1786 ();
 sg13g2_fill_2 FILLER_38_1790 ();
 sg13g2_decap_4 FILLER_38_1809 ();
 sg13g2_fill_1 FILLER_38_1813 ();
 sg13g2_fill_2 FILLER_38_1831 ();
 sg13g2_fill_1 FILLER_38_1833 ();
 sg13g2_decap_8 FILLER_38_1899 ();
 sg13g2_decap_4 FILLER_38_1906 ();
 sg13g2_fill_2 FILLER_38_1943 ();
 sg13g2_fill_1 FILLER_38_1945 ();
 sg13g2_fill_2 FILLER_38_1955 ();
 sg13g2_decap_4 FILLER_38_1965 ();
 sg13g2_fill_1 FILLER_38_1969 ();
 sg13g2_fill_2 FILLER_38_2069 ();
 sg13g2_fill_2 FILLER_38_2115 ();
 sg13g2_fill_2 FILLER_38_2134 ();
 sg13g2_fill_1 FILLER_38_2236 ();
 sg13g2_fill_2 FILLER_38_2263 ();
 sg13g2_fill_1 FILLER_38_2265 ();
 sg13g2_fill_2 FILLER_38_2348 ();
 sg13g2_fill_2 FILLER_38_2354 ();
 sg13g2_fill_2 FILLER_38_2382 ();
 sg13g2_fill_1 FILLER_38_2397 ();
 sg13g2_fill_1 FILLER_38_2444 ();
 sg13g2_fill_2 FILLER_38_2461 ();
 sg13g2_fill_1 FILLER_38_2463 ();
 sg13g2_fill_2 FILLER_38_2526 ();
 sg13g2_fill_2 FILLER_38_2546 ();
 sg13g2_decap_8 FILLER_38_2591 ();
 sg13g2_decap_8 FILLER_38_2598 ();
 sg13g2_decap_8 FILLER_38_2605 ();
 sg13g2_decap_8 FILLER_38_2612 ();
 sg13g2_decap_8 FILLER_38_2619 ();
 sg13g2_decap_8 FILLER_38_2626 ();
 sg13g2_decap_8 FILLER_38_2633 ();
 sg13g2_decap_8 FILLER_38_2640 ();
 sg13g2_decap_8 FILLER_38_2647 ();
 sg13g2_decap_8 FILLER_38_2654 ();
 sg13g2_decap_8 FILLER_38_2661 ();
 sg13g2_decap_4 FILLER_38_2668 ();
 sg13g2_fill_2 FILLER_38_2672 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_504 ();
 sg13g2_fill_2 FILLER_39_511 ();
 sg13g2_fill_2 FILLER_39_543 ();
 sg13g2_fill_1 FILLER_39_570 ();
 sg13g2_decap_8 FILLER_39_580 ();
 sg13g2_fill_1 FILLER_39_587 ();
 sg13g2_fill_1 FILLER_39_597 ();
 sg13g2_fill_2 FILLER_39_616 ();
 sg13g2_fill_2 FILLER_39_655 ();
 sg13g2_fill_1 FILLER_39_657 ();
 sg13g2_fill_1 FILLER_39_709 ();
 sg13g2_fill_2 FILLER_39_745 ();
 sg13g2_fill_2 FILLER_39_773 ();
 sg13g2_fill_1 FILLER_39_817 ();
 sg13g2_fill_2 FILLER_39_826 ();
 sg13g2_fill_1 FILLER_39_859 ();
 sg13g2_decap_4 FILLER_39_935 ();
 sg13g2_fill_2 FILLER_39_939 ();
 sg13g2_fill_2 FILLER_39_997 ();
 sg13g2_fill_1 FILLER_39_999 ();
 sg13g2_decap_8 FILLER_39_1009 ();
 sg13g2_fill_1 FILLER_39_1016 ();
 sg13g2_decap_8 FILLER_39_1025 ();
 sg13g2_decap_4 FILLER_39_1032 ();
 sg13g2_fill_2 FILLER_39_1067 ();
 sg13g2_fill_2 FILLER_39_1109 ();
 sg13g2_fill_1 FILLER_39_1133 ();
 sg13g2_fill_2 FILLER_39_1160 ();
 sg13g2_fill_1 FILLER_39_1201 ();
 sg13g2_fill_2 FILLER_39_1208 ();
 sg13g2_fill_2 FILLER_39_1258 ();
 sg13g2_fill_2 FILLER_39_1268 ();
 sg13g2_fill_1 FILLER_39_1270 ();
 sg13g2_fill_2 FILLER_39_1289 ();
 sg13g2_fill_1 FILLER_39_1291 ();
 sg13g2_fill_1 FILLER_39_1299 ();
 sg13g2_decap_8 FILLER_39_1323 ();
 sg13g2_decap_8 FILLER_39_1330 ();
 sg13g2_decap_8 FILLER_39_1337 ();
 sg13g2_decap_8 FILLER_39_1344 ();
 sg13g2_fill_2 FILLER_39_1351 ();
 sg13g2_fill_1 FILLER_39_1353 ();
 sg13g2_fill_2 FILLER_39_1385 ();
 sg13g2_fill_1 FILLER_39_1387 ();
 sg13g2_fill_2 FILLER_39_1395 ();
 sg13g2_fill_2 FILLER_39_1441 ();
 sg13g2_decap_4 FILLER_39_1457 ();
 sg13g2_fill_1 FILLER_39_1461 ();
 sg13g2_fill_1 FILLER_39_1491 ();
 sg13g2_fill_1 FILLER_39_1509 ();
 sg13g2_decap_4 FILLER_39_1514 ();
 sg13g2_fill_2 FILLER_39_1527 ();
 sg13g2_fill_1 FILLER_39_1529 ();
 sg13g2_fill_1 FILLER_39_1547 ();
 sg13g2_fill_2 FILLER_39_1556 ();
 sg13g2_fill_2 FILLER_39_1596 ();
 sg13g2_fill_1 FILLER_39_1598 ();
 sg13g2_fill_2 FILLER_39_1646 ();
 sg13g2_fill_1 FILLER_39_1648 ();
 sg13g2_fill_1 FILLER_39_1690 ();
 sg13g2_fill_2 FILLER_39_1714 ();
 sg13g2_fill_2 FILLER_39_1725 ();
 sg13g2_fill_2 FILLER_39_1763 ();
 sg13g2_decap_8 FILLER_39_1891 ();
 sg13g2_decap_4 FILLER_39_1898 ();
 sg13g2_fill_1 FILLER_39_1902 ();
 sg13g2_fill_1 FILLER_39_1919 ();
 sg13g2_fill_2 FILLER_39_1928 ();
 sg13g2_fill_2 FILLER_39_1939 ();
 sg13g2_fill_1 FILLER_39_1941 ();
 sg13g2_fill_2 FILLER_39_1955 ();
 sg13g2_fill_1 FILLER_39_1957 ();
 sg13g2_fill_2 FILLER_39_1966 ();
 sg13g2_fill_1 FILLER_39_1968 ();
 sg13g2_fill_2 FILLER_39_2009 ();
 sg13g2_fill_1 FILLER_39_2011 ();
 sg13g2_fill_2 FILLER_39_2026 ();
 sg13g2_fill_1 FILLER_39_2028 ();
 sg13g2_fill_2 FILLER_39_2070 ();
 sg13g2_fill_1 FILLER_39_2072 ();
 sg13g2_fill_2 FILLER_39_2103 ();
 sg13g2_decap_4 FILLER_39_2138 ();
 sg13g2_fill_2 FILLER_39_2142 ();
 sg13g2_fill_2 FILLER_39_2157 ();
 sg13g2_fill_1 FILLER_39_2159 ();
 sg13g2_decap_8 FILLER_39_2169 ();
 sg13g2_fill_1 FILLER_39_2176 ();
 sg13g2_decap_4 FILLER_39_2182 ();
 sg13g2_fill_1 FILLER_39_2199 ();
 sg13g2_fill_2 FILLER_39_2204 ();
 sg13g2_fill_1 FILLER_39_2236 ();
 sg13g2_fill_2 FILLER_39_2246 ();
 sg13g2_fill_1 FILLER_39_2252 ();
 sg13g2_decap_4 FILLER_39_2279 ();
 sg13g2_fill_1 FILLER_39_2304 ();
 sg13g2_fill_1 FILLER_39_2319 ();
 sg13g2_decap_4 FILLER_39_2347 ();
 sg13g2_fill_2 FILLER_39_2351 ();
 sg13g2_fill_2 FILLER_39_2375 ();
 sg13g2_fill_2 FILLER_39_2381 ();
 sg13g2_fill_2 FILLER_39_2403 ();
 sg13g2_fill_1 FILLER_39_2405 ();
 sg13g2_fill_2 FILLER_39_2427 ();
 sg13g2_fill_1 FILLER_39_2429 ();
 sg13g2_fill_2 FILLER_39_2456 ();
 sg13g2_fill_1 FILLER_39_2458 ();
 sg13g2_decap_8 FILLER_39_2577 ();
 sg13g2_decap_8 FILLER_39_2584 ();
 sg13g2_decap_8 FILLER_39_2591 ();
 sg13g2_decap_8 FILLER_39_2598 ();
 sg13g2_decap_8 FILLER_39_2605 ();
 sg13g2_decap_8 FILLER_39_2612 ();
 sg13g2_decap_8 FILLER_39_2619 ();
 sg13g2_decap_8 FILLER_39_2626 ();
 sg13g2_decap_8 FILLER_39_2633 ();
 sg13g2_decap_8 FILLER_39_2640 ();
 sg13g2_decap_8 FILLER_39_2647 ();
 sg13g2_decap_8 FILLER_39_2654 ();
 sg13g2_decap_8 FILLER_39_2661 ();
 sg13g2_decap_4 FILLER_39_2668 ();
 sg13g2_fill_2 FILLER_39_2672 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_4 FILLER_40_511 ();
 sg13g2_fill_2 FILLER_40_532 ();
 sg13g2_fill_1 FILLER_40_534 ();
 sg13g2_fill_2 FILLER_40_544 ();
 sg13g2_fill_1 FILLER_40_580 ();
 sg13g2_fill_2 FILLER_40_589 ();
 sg13g2_fill_1 FILLER_40_591 ();
 sg13g2_decap_8 FILLER_40_624 ();
 sg13g2_fill_1 FILLER_40_631 ();
 sg13g2_fill_2 FILLER_40_658 ();
 sg13g2_decap_4 FILLER_40_699 ();
 sg13g2_fill_2 FILLER_40_703 ();
 sg13g2_fill_2 FILLER_40_822 ();
 sg13g2_fill_1 FILLER_40_824 ();
 sg13g2_fill_2 FILLER_40_851 ();
 sg13g2_fill_2 FILLER_40_862 ();
 sg13g2_fill_1 FILLER_40_864 ();
 sg13g2_fill_1 FILLER_40_875 ();
 sg13g2_fill_1 FILLER_40_889 ();
 sg13g2_fill_1 FILLER_40_916 ();
 sg13g2_decap_8 FILLER_40_921 ();
 sg13g2_decap_8 FILLER_40_928 ();
 sg13g2_decap_8 FILLER_40_935 ();
 sg13g2_decap_4 FILLER_40_942 ();
 sg13g2_fill_2 FILLER_40_946 ();
 sg13g2_decap_8 FILLER_40_952 ();
 sg13g2_decap_8 FILLER_40_959 ();
 sg13g2_decap_4 FILLER_40_966 ();
 sg13g2_fill_2 FILLER_40_970 ();
 sg13g2_fill_2 FILLER_40_976 ();
 sg13g2_fill_1 FILLER_40_982 ();
 sg13g2_fill_2 FILLER_40_996 ();
 sg13g2_fill_1 FILLER_40_998 ();
 sg13g2_decap_4 FILLER_40_1029 ();
 sg13g2_fill_1 FILLER_40_1089 ();
 sg13g2_fill_2 FILLER_40_1148 ();
 sg13g2_fill_2 FILLER_40_1202 ();
 sg13g2_fill_2 FILLER_40_1211 ();
 sg13g2_fill_1 FILLER_40_1213 ();
 sg13g2_fill_2 FILLER_40_1236 ();
 sg13g2_fill_1 FILLER_40_1238 ();
 sg13g2_fill_1 FILLER_40_1253 ();
 sg13g2_fill_1 FILLER_40_1263 ();
 sg13g2_fill_2 FILLER_40_1288 ();
 sg13g2_decap_8 FILLER_40_1295 ();
 sg13g2_decap_4 FILLER_40_1302 ();
 sg13g2_fill_2 FILLER_40_1306 ();
 sg13g2_fill_2 FILLER_40_1344 ();
 sg13g2_fill_1 FILLER_40_1346 ();
 sg13g2_decap_4 FILLER_40_1360 ();
 sg13g2_fill_1 FILLER_40_1390 ();
 sg13g2_fill_2 FILLER_40_1408 ();
 sg13g2_decap_4 FILLER_40_1418 ();
 sg13g2_decap_4 FILLER_40_1447 ();
 sg13g2_fill_2 FILLER_40_1451 ();
 sg13g2_fill_2 FILLER_40_1461 ();
 sg13g2_fill_1 FILLER_40_1463 ();
 sg13g2_fill_1 FILLER_40_1493 ();
 sg13g2_decap_8 FILLER_40_1507 ();
 sg13g2_decap_4 FILLER_40_1514 ();
 sg13g2_fill_1 FILLER_40_1518 ();
 sg13g2_decap_8 FILLER_40_1530 ();
 sg13g2_fill_1 FILLER_40_1560 ();
 sg13g2_decap_8 FILLER_40_1587 ();
 sg13g2_fill_2 FILLER_40_1594 ();
 sg13g2_fill_2 FILLER_40_1633 ();
 sg13g2_fill_1 FILLER_40_1635 ();
 sg13g2_fill_2 FILLER_40_1646 ();
 sg13g2_decap_4 FILLER_40_1683 ();
 sg13g2_fill_1 FILLER_40_1687 ();
 sg13g2_fill_2 FILLER_40_1760 ();
 sg13g2_fill_1 FILLER_40_1762 ();
 sg13g2_fill_1 FILLER_40_1873 ();
 sg13g2_fill_1 FILLER_40_1892 ();
 sg13g2_decap_4 FILLER_40_1919 ();
 sg13g2_fill_2 FILLER_40_1950 ();
 sg13g2_fill_1 FILLER_40_1952 ();
 sg13g2_fill_2 FILLER_40_1964 ();
 sg13g2_fill_1 FILLER_40_1966 ();
 sg13g2_fill_2 FILLER_40_2023 ();
 sg13g2_fill_1 FILLER_40_2025 ();
 sg13g2_fill_2 FILLER_40_2039 ();
 sg13g2_fill_2 FILLER_40_2053 ();
 sg13g2_fill_1 FILLER_40_2055 ();
 sg13g2_fill_1 FILLER_40_2060 ();
 sg13g2_fill_1 FILLER_40_2065 ();
 sg13g2_decap_4 FILLER_40_2071 ();
 sg13g2_fill_1 FILLER_40_2075 ();
 sg13g2_decap_8 FILLER_40_2141 ();
 sg13g2_decap_8 FILLER_40_2148 ();
 sg13g2_fill_2 FILLER_40_2155 ();
 sg13g2_decap_8 FILLER_40_2161 ();
 sg13g2_fill_1 FILLER_40_2168 ();
 sg13g2_fill_2 FILLER_40_2177 ();
 sg13g2_decap_8 FILLER_40_2184 ();
 sg13g2_decap_8 FILLER_40_2191 ();
 sg13g2_decap_4 FILLER_40_2198 ();
 sg13g2_fill_2 FILLER_40_2202 ();
 sg13g2_decap_4 FILLER_40_2208 ();
 sg13g2_fill_1 FILLER_40_2212 ();
 sg13g2_fill_1 FILLER_40_2217 ();
 sg13g2_decap_8 FILLER_40_2239 ();
 sg13g2_decap_8 FILLER_40_2246 ();
 sg13g2_fill_2 FILLER_40_2411 ();
 sg13g2_fill_1 FILLER_40_2413 ();
 sg13g2_decap_4 FILLER_40_2466 ();
 sg13g2_fill_1 FILLER_40_2474 ();
 sg13g2_decap_4 FILLER_40_2483 ();
 sg13g2_fill_1 FILLER_40_2487 ();
 sg13g2_fill_2 FILLER_40_2558 ();
 sg13g2_decap_8 FILLER_40_2569 ();
 sg13g2_decap_8 FILLER_40_2576 ();
 sg13g2_decap_8 FILLER_40_2583 ();
 sg13g2_decap_8 FILLER_40_2590 ();
 sg13g2_decap_8 FILLER_40_2597 ();
 sg13g2_decap_8 FILLER_40_2604 ();
 sg13g2_decap_8 FILLER_40_2611 ();
 sg13g2_decap_8 FILLER_40_2618 ();
 sg13g2_decap_8 FILLER_40_2625 ();
 sg13g2_decap_8 FILLER_40_2632 ();
 sg13g2_decap_8 FILLER_40_2639 ();
 sg13g2_decap_8 FILLER_40_2646 ();
 sg13g2_decap_8 FILLER_40_2653 ();
 sg13g2_decap_8 FILLER_40_2660 ();
 sg13g2_decap_8 FILLER_40_2667 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_4 FILLER_41_504 ();
 sg13g2_fill_2 FILLER_41_508 ();
 sg13g2_fill_1 FILLER_41_541 ();
 sg13g2_fill_2 FILLER_41_551 ();
 sg13g2_fill_2 FILLER_41_588 ();
 sg13g2_fill_1 FILLER_41_616 ();
 sg13g2_decap_4 FILLER_41_637 ();
 sg13g2_fill_1 FILLER_41_641 ();
 sg13g2_fill_2 FILLER_41_672 ();
 sg13g2_fill_1 FILLER_41_674 ();
 sg13g2_decap_8 FILLER_41_690 ();
 sg13g2_fill_2 FILLER_41_697 ();
 sg13g2_fill_2 FILLER_41_708 ();
 sg13g2_fill_1 FILLER_41_710 ();
 sg13g2_fill_1 FILLER_41_740 ();
 sg13g2_fill_1 FILLER_41_766 ();
 sg13g2_fill_1 FILLER_41_772 ();
 sg13g2_fill_1 FILLER_41_791 ();
 sg13g2_fill_2 FILLER_41_796 ();
 sg13g2_fill_1 FILLER_41_798 ();
 sg13g2_fill_1 FILLER_41_809 ();
 sg13g2_decap_4 FILLER_41_828 ();
 sg13g2_fill_1 FILLER_41_832 ();
 sg13g2_fill_2 FILLER_41_849 ();
 sg13g2_fill_2 FILLER_41_868 ();
 sg13g2_fill_1 FILLER_41_870 ();
 sg13g2_decap_8 FILLER_41_909 ();
 sg13g2_fill_1 FILLER_41_916 ();
 sg13g2_decap_4 FILLER_41_928 ();
 sg13g2_fill_2 FILLER_41_932 ();
 sg13g2_fill_1 FILLER_41_1017 ();
 sg13g2_decap_8 FILLER_41_1026 ();
 sg13g2_decap_4 FILLER_41_1033 ();
 sg13g2_fill_2 FILLER_41_1037 ();
 sg13g2_fill_1 FILLER_41_1066 ();
 sg13g2_fill_2 FILLER_41_1133 ();
 sg13g2_fill_1 FILLER_41_1135 ();
 sg13g2_fill_1 FILLER_41_1149 ();
 sg13g2_fill_2 FILLER_41_1203 ();
 sg13g2_fill_1 FILLER_41_1205 ();
 sg13g2_fill_2 FILLER_41_1212 ();
 sg13g2_decap_8 FILLER_41_1223 ();
 sg13g2_decap_4 FILLER_41_1230 ();
 sg13g2_fill_2 FILLER_41_1234 ();
 sg13g2_fill_1 FILLER_41_1241 ();
 sg13g2_decap_4 FILLER_41_1248 ();
 sg13g2_fill_1 FILLER_41_1252 ();
 sg13g2_fill_2 FILLER_41_1276 ();
 sg13g2_decap_8 FILLER_41_1283 ();
 sg13g2_fill_1 FILLER_41_1290 ();
 sg13g2_fill_1 FILLER_41_1303 ();
 sg13g2_decap_4 FILLER_41_1339 ();
 sg13g2_fill_2 FILLER_41_1343 ();
 sg13g2_fill_2 FILLER_41_1358 ();
 sg13g2_decap_4 FILLER_41_1374 ();
 sg13g2_fill_2 FILLER_41_1472 ();
 sg13g2_fill_1 FILLER_41_1499 ();
 sg13g2_decap_8 FILLER_41_1525 ();
 sg13g2_fill_1 FILLER_41_1532 ();
 sg13g2_fill_2 FILLER_41_1538 ();
 sg13g2_fill_1 FILLER_41_1540 ();
 sg13g2_decap_8 FILLER_41_1593 ();
 sg13g2_fill_2 FILLER_41_1624 ();
 sg13g2_fill_1 FILLER_41_1626 ();
 sg13g2_fill_2 FILLER_41_1666 ();
 sg13g2_fill_1 FILLER_41_1668 ();
 sg13g2_fill_2 FILLER_41_1674 ();
 sg13g2_fill_1 FILLER_41_1676 ();
 sg13g2_fill_2 FILLER_41_1682 ();
 sg13g2_decap_4 FILLER_41_1752 ();
 sg13g2_fill_1 FILLER_41_1756 ();
 sg13g2_decap_4 FILLER_41_1783 ();
 sg13g2_fill_1 FILLER_41_1891 ();
 sg13g2_decap_8 FILLER_41_1905 ();
 sg13g2_fill_1 FILLER_41_1912 ();
 sg13g2_fill_1 FILLER_41_1916 ();
 sg13g2_fill_2 FILLER_41_1948 ();
 sg13g2_fill_1 FILLER_41_1978 ();
 sg13g2_fill_1 FILLER_41_2025 ();
 sg13g2_decap_4 FILLER_41_2047 ();
 sg13g2_fill_1 FILLER_41_2055 ();
 sg13g2_fill_1 FILLER_41_2061 ();
 sg13g2_fill_2 FILLER_41_2085 ();
 sg13g2_fill_1 FILLER_41_2087 ();
 sg13g2_fill_2 FILLER_41_2100 ();
 sg13g2_decap_4 FILLER_41_2137 ();
 sg13g2_fill_2 FILLER_41_2141 ();
 sg13g2_fill_2 FILLER_41_2206 ();
 sg13g2_fill_1 FILLER_41_2213 ();
 sg13g2_decap_8 FILLER_41_2245 ();
 sg13g2_decap_8 FILLER_41_2252 ();
 sg13g2_decap_4 FILLER_41_2271 ();
 sg13g2_fill_1 FILLER_41_2275 ();
 sg13g2_fill_1 FILLER_41_2292 ();
 sg13g2_fill_2 FILLER_41_2302 ();
 sg13g2_fill_1 FILLER_41_2304 ();
 sg13g2_decap_4 FILLER_41_2343 ();
 sg13g2_fill_1 FILLER_41_2347 ();
 sg13g2_fill_2 FILLER_41_2440 ();
 sg13g2_fill_1 FILLER_41_2442 ();
 sg13g2_decap_8 FILLER_41_2469 ();
 sg13g2_decap_8 FILLER_41_2476 ();
 sg13g2_decap_8 FILLER_41_2483 ();
 sg13g2_decap_4 FILLER_41_2490 ();
 sg13g2_fill_1 FILLER_41_2494 ();
 sg13g2_fill_2 FILLER_41_2554 ();
 sg13g2_fill_2 FILLER_41_2582 ();
 sg13g2_fill_1 FILLER_41_2584 ();
 sg13g2_decap_8 FILLER_41_2606 ();
 sg13g2_decap_8 FILLER_41_2613 ();
 sg13g2_decap_8 FILLER_41_2620 ();
 sg13g2_decap_8 FILLER_41_2627 ();
 sg13g2_decap_8 FILLER_41_2634 ();
 sg13g2_decap_8 FILLER_41_2641 ();
 sg13g2_decap_8 FILLER_41_2648 ();
 sg13g2_decap_8 FILLER_41_2655 ();
 sg13g2_decap_8 FILLER_41_2662 ();
 sg13g2_decap_4 FILLER_41_2669 ();
 sg13g2_fill_1 FILLER_41_2673 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_434 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_fill_2 FILLER_42_511 ();
 sg13g2_fill_2 FILLER_42_544 ();
 sg13g2_fill_2 FILLER_42_637 ();
 sg13g2_fill_1 FILLER_42_639 ();
 sg13g2_decap_8 FILLER_42_645 ();
 sg13g2_decap_8 FILLER_42_652 ();
 sg13g2_fill_1 FILLER_42_659 ();
 sg13g2_fill_2 FILLER_42_674 ();
 sg13g2_decap_4 FILLER_42_681 ();
 sg13g2_fill_1 FILLER_42_685 ();
 sg13g2_fill_1 FILLER_42_712 ();
 sg13g2_fill_1 FILLER_42_755 ();
 sg13g2_fill_1 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_842 ();
 sg13g2_decap_8 FILLER_42_849 ();
 sg13g2_decap_4 FILLER_42_874 ();
 sg13g2_fill_1 FILLER_42_878 ();
 sg13g2_fill_1 FILLER_42_883 ();
 sg13g2_fill_1 FILLER_42_922 ();
 sg13g2_decap_8 FILLER_42_975 ();
 sg13g2_decap_4 FILLER_42_982 ();
 sg13g2_fill_1 FILLER_42_986 ();
 sg13g2_fill_2 FILLER_42_991 ();
 sg13g2_fill_1 FILLER_42_993 ();
 sg13g2_fill_1 FILLER_42_1020 ();
 sg13g2_fill_1 FILLER_42_1029 ();
 sg13g2_fill_1 FILLER_42_1038 ();
 sg13g2_fill_1 FILLER_42_1047 ();
 sg13g2_fill_1 FILLER_42_1074 ();
 sg13g2_fill_1 FILLER_42_1105 ();
 sg13g2_fill_2 FILLER_42_1128 ();
 sg13g2_fill_2 FILLER_42_1139 ();
 sg13g2_fill_2 FILLER_42_1156 ();
 sg13g2_fill_1 FILLER_42_1167 ();
 sg13g2_decap_8 FILLER_42_1204 ();
 sg13g2_fill_2 FILLER_42_1211 ();
 sg13g2_decap_8 FILLER_42_1221 ();
 sg13g2_decap_4 FILLER_42_1228 ();
 sg13g2_fill_2 FILLER_42_1232 ();
 sg13g2_decap_4 FILLER_42_1246 ();
 sg13g2_decap_4 FILLER_42_1254 ();
 sg13g2_fill_2 FILLER_42_1258 ();
 sg13g2_decap_8 FILLER_42_1264 ();
 sg13g2_decap_8 FILLER_42_1271 ();
 sg13g2_fill_2 FILLER_42_1278 ();
 sg13g2_fill_1 FILLER_42_1280 ();
 sg13g2_fill_1 FILLER_42_1311 ();
 sg13g2_fill_2 FILLER_42_1338 ();
 sg13g2_fill_1 FILLER_42_1340 ();
 sg13g2_decap_8 FILLER_42_1346 ();
 sg13g2_fill_1 FILLER_42_1353 ();
 sg13g2_decap_4 FILLER_42_1362 ();
 sg13g2_fill_1 FILLER_42_1366 ();
 sg13g2_decap_4 FILLER_42_1385 ();
 sg13g2_decap_8 FILLER_42_1457 ();
 sg13g2_decap_8 FILLER_42_1464 ();
 sg13g2_decap_8 FILLER_42_1471 ();
 sg13g2_fill_2 FILLER_42_1478 ();
 sg13g2_fill_1 FILLER_42_1480 ();
 sg13g2_fill_2 FILLER_42_1507 ();
 sg13g2_fill_2 FILLER_42_1521 ();
 sg13g2_fill_2 FILLER_42_1553 ();
 sg13g2_fill_1 FILLER_42_1555 ();
 sg13g2_fill_2 FILLER_42_1567 ();
 sg13g2_fill_1 FILLER_42_1569 ();
 sg13g2_decap_8 FILLER_42_1593 ();
 sg13g2_decap_8 FILLER_42_1600 ();
 sg13g2_decap_8 FILLER_42_1607 ();
 sg13g2_decap_8 FILLER_42_1614 ();
 sg13g2_decap_8 FILLER_42_1621 ();
 sg13g2_fill_2 FILLER_42_1628 ();
 sg13g2_fill_2 FILLER_42_1639 ();
 sg13g2_decap_4 FILLER_42_1651 ();
 sg13g2_fill_1 FILLER_42_1655 ();
 sg13g2_fill_1 FILLER_42_1661 ();
 sg13g2_fill_2 FILLER_42_1666 ();
 sg13g2_decap_4 FILLER_42_1691 ();
 sg13g2_decap_8 FILLER_42_1703 ();
 sg13g2_decap_4 FILLER_42_1710 ();
 sg13g2_decap_8 FILLER_42_1751 ();
 sg13g2_decap_4 FILLER_42_1758 ();
 sg13g2_fill_1 FILLER_42_1762 ();
 sg13g2_fill_2 FILLER_42_1777 ();
 sg13g2_fill_1 FILLER_42_1779 ();
 sg13g2_fill_2 FILLER_42_1806 ();
 sg13g2_fill_1 FILLER_42_1808 ();
 sg13g2_decap_4 FILLER_42_1843 ();
 sg13g2_fill_1 FILLER_42_1855 ();
 sg13g2_fill_2 FILLER_42_1911 ();
 sg13g2_fill_1 FILLER_42_1946 ();
 sg13g2_fill_2 FILLER_42_2006 ();
 sg13g2_fill_2 FILLER_42_2038 ();
 sg13g2_fill_1 FILLER_42_2040 ();
 sg13g2_fill_1 FILLER_42_2128 ();
 sg13g2_fill_2 FILLER_42_2159 ();
 sg13g2_fill_1 FILLER_42_2201 ();
 sg13g2_fill_2 FILLER_42_2228 ();
 sg13g2_fill_1 FILLER_42_2230 ();
 sg13g2_fill_2 FILLER_42_2265 ();
 sg13g2_fill_1 FILLER_42_2267 ();
 sg13g2_decap_8 FILLER_42_2294 ();
 sg13g2_decap_8 FILLER_42_2301 ();
 sg13g2_fill_2 FILLER_42_2320 ();
 sg13g2_fill_2 FILLER_42_2343 ();
 sg13g2_fill_1 FILLER_42_2345 ();
 sg13g2_fill_1 FILLER_42_2423 ();
 sg13g2_decap_8 FILLER_42_2464 ();
 sg13g2_fill_2 FILLER_42_2471 ();
 sg13g2_decap_4 FILLER_42_2507 ();
 sg13g2_fill_2 FILLER_42_2511 ();
 sg13g2_fill_2 FILLER_42_2521 ();
 sg13g2_fill_2 FILLER_42_2527 ();
 sg13g2_fill_1 FILLER_42_2529 ();
 sg13g2_decap_4 FILLER_42_2540 ();
 sg13g2_fill_1 FILLER_42_2544 ();
 sg13g2_decap_8 FILLER_42_2615 ();
 sg13g2_decap_8 FILLER_42_2622 ();
 sg13g2_decap_8 FILLER_42_2629 ();
 sg13g2_decap_8 FILLER_42_2636 ();
 sg13g2_decap_8 FILLER_42_2643 ();
 sg13g2_decap_8 FILLER_42_2650 ();
 sg13g2_decap_8 FILLER_42_2657 ();
 sg13g2_decap_8 FILLER_42_2664 ();
 sg13g2_fill_2 FILLER_42_2671 ();
 sg13g2_fill_1 FILLER_42_2673 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_8 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_497 ();
 sg13g2_fill_2 FILLER_43_504 ();
 sg13g2_fill_1 FILLER_43_545 ();
 sg13g2_fill_1 FILLER_43_581 ();
 sg13g2_fill_2 FILLER_43_610 ();
 sg13g2_fill_2 FILLER_43_668 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_fill_1 FILLER_43_686 ();
 sg13g2_fill_1 FILLER_43_700 ();
 sg13g2_fill_1 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_754 ();
 sg13g2_fill_1 FILLER_43_789 ();
 sg13g2_fill_1 FILLER_43_814 ();
 sg13g2_decap_4 FILLER_43_841 ();
 sg13g2_fill_2 FILLER_43_850 ();
 sg13g2_fill_1 FILLER_43_852 ();
 sg13g2_fill_2 FILLER_43_888 ();
 sg13g2_fill_1 FILLER_43_890 ();
 sg13g2_fill_2 FILLER_43_920 ();
 sg13g2_fill_1 FILLER_43_922 ();
 sg13g2_fill_1 FILLER_43_994 ();
 sg13g2_decap_8 FILLER_43_1010 ();
 sg13g2_fill_1 FILLER_43_1017 ();
 sg13g2_decap_4 FILLER_43_1039 ();
 sg13g2_fill_2 FILLER_43_1043 ();
 sg13g2_fill_2 FILLER_43_1097 ();
 sg13g2_fill_2 FILLER_43_1132 ();
 sg13g2_fill_1 FILLER_43_1134 ();
 sg13g2_fill_1 FILLER_43_1164 ();
 sg13g2_fill_1 FILLER_43_1177 ();
 sg13g2_decap_4 FILLER_43_1200 ();
 sg13g2_fill_1 FILLER_43_1204 ();
 sg13g2_fill_2 FILLER_43_1279 ();
 sg13g2_fill_1 FILLER_43_1307 ();
 sg13g2_fill_2 FILLER_43_1342 ();
 sg13g2_fill_1 FILLER_43_1344 ();
 sg13g2_fill_2 FILLER_43_1398 ();
 sg13g2_decap_8 FILLER_43_1419 ();
 sg13g2_fill_2 FILLER_43_1426 ();
 sg13g2_decap_8 FILLER_43_1433 ();
 sg13g2_decap_8 FILLER_43_1466 ();
 sg13g2_decap_8 FILLER_43_1473 ();
 sg13g2_fill_2 FILLER_43_1480 ();
 sg13g2_fill_1 FILLER_43_1482 ();
 sg13g2_fill_2 FILLER_43_1515 ();
 sg13g2_fill_2 FILLER_43_1543 ();
 sg13g2_fill_1 FILLER_43_1545 ();
 sg13g2_fill_2 FILLER_43_1561 ();
 sg13g2_decap_8 FILLER_43_1619 ();
 sg13g2_decap_8 FILLER_43_1626 ();
 sg13g2_fill_2 FILLER_43_1633 ();
 sg13g2_fill_1 FILLER_43_1635 ();
 sg13g2_fill_2 FILLER_43_1640 ();
 sg13g2_fill_1 FILLER_43_1642 ();
 sg13g2_decap_4 FILLER_43_1667 ();
 sg13g2_fill_1 FILLER_43_1671 ();
 sg13g2_fill_2 FILLER_43_1683 ();
 sg13g2_fill_1 FILLER_43_1708 ();
 sg13g2_decap_4 FILLER_43_1713 ();
 sg13g2_fill_2 FILLER_43_1717 ();
 sg13g2_decap_8 FILLER_43_1733 ();
 sg13g2_decap_8 FILLER_43_1740 ();
 sg13g2_decap_4 FILLER_43_1747 ();
 sg13g2_fill_2 FILLER_43_1751 ();
 sg13g2_decap_8 FILLER_43_1766 ();
 sg13g2_decap_4 FILLER_43_1773 ();
 sg13g2_decap_8 FILLER_43_1785 ();
 sg13g2_decap_8 FILLER_43_1792 ();
 sg13g2_decap_8 FILLER_43_1816 ();
 sg13g2_decap_4 FILLER_43_1823 ();
 sg13g2_fill_2 FILLER_43_1853 ();
 sg13g2_fill_2 FILLER_43_1922 ();
 sg13g2_fill_1 FILLER_43_1951 ();
 sg13g2_fill_2 FILLER_43_2050 ();
 sg13g2_fill_1 FILLER_43_2052 ();
 sg13g2_fill_2 FILLER_43_2100 ();
 sg13g2_fill_1 FILLER_43_2146 ();
 sg13g2_fill_1 FILLER_43_2213 ();
 sg13g2_fill_2 FILLER_43_2262 ();
 sg13g2_decap_8 FILLER_43_2307 ();
 sg13g2_fill_2 FILLER_43_2314 ();
 sg13g2_decap_8 FILLER_43_2333 ();
 sg13g2_decap_8 FILLER_43_2340 ();
 sg13g2_decap_4 FILLER_43_2347 ();
 sg13g2_decap_4 FILLER_43_2391 ();
 sg13g2_decap_8 FILLER_43_2399 ();
 sg13g2_fill_2 FILLER_43_2406 ();
 sg13g2_fill_2 FILLER_43_2413 ();
 sg13g2_fill_1 FILLER_43_2415 ();
 sg13g2_fill_2 FILLER_43_2454 ();
 sg13g2_decap_4 FILLER_43_2462 ();
 sg13g2_fill_2 FILLER_43_2466 ();
 sg13g2_decap_4 FILLER_43_2494 ();
 sg13g2_decap_4 FILLER_43_2517 ();
 sg13g2_fill_2 FILLER_43_2563 ();
 sg13g2_decap_8 FILLER_43_2621 ();
 sg13g2_decap_8 FILLER_43_2628 ();
 sg13g2_decap_8 FILLER_43_2635 ();
 sg13g2_decap_8 FILLER_43_2642 ();
 sg13g2_decap_8 FILLER_43_2649 ();
 sg13g2_decap_8 FILLER_43_2656 ();
 sg13g2_decap_8 FILLER_43_2663 ();
 sg13g2_decap_4 FILLER_43_2670 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_476 ();
 sg13g2_decap_8 FILLER_44_483 ();
 sg13g2_decap_8 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_497 ();
 sg13g2_decap_4 FILLER_44_504 ();
 sg13g2_fill_1 FILLER_44_548 ();
 sg13g2_fill_2 FILLER_44_599 ();
 sg13g2_fill_1 FILLER_44_612 ();
 sg13g2_fill_2 FILLER_44_627 ();
 sg13g2_fill_2 FILLER_44_647 ();
 sg13g2_fill_1 FILLER_44_649 ();
 sg13g2_fill_2 FILLER_44_667 ();
 sg13g2_fill_1 FILLER_44_669 ();
 sg13g2_fill_1 FILLER_44_699 ();
 sg13g2_fill_1 FILLER_44_713 ();
 sg13g2_fill_2 FILLER_44_724 ();
 sg13g2_fill_1 FILLER_44_726 ();
 sg13g2_decap_4 FILLER_44_745 ();
 sg13g2_fill_1 FILLER_44_749 ();
 sg13g2_decap_4 FILLER_44_755 ();
 sg13g2_fill_1 FILLER_44_781 ();
 sg13g2_fill_1 FILLER_44_786 ();
 sg13g2_fill_2 FILLER_44_819 ();
 sg13g2_fill_1 FILLER_44_821 ();
 sg13g2_fill_1 FILLER_44_857 ();
 sg13g2_fill_1 FILLER_44_898 ();
 sg13g2_fill_2 FILLER_44_904 ();
 sg13g2_fill_1 FILLER_44_906 ();
 sg13g2_fill_1 FILLER_44_932 ();
 sg13g2_fill_1 FILLER_44_942 ();
 sg13g2_fill_2 FILLER_44_955 ();
 sg13g2_fill_1 FILLER_44_957 ();
 sg13g2_fill_1 FILLER_44_984 ();
 sg13g2_fill_1 FILLER_44_1017 ();
 sg13g2_decap_4 FILLER_44_1042 ();
 sg13g2_fill_1 FILLER_44_1046 ();
 sg13g2_fill_1 FILLER_44_1086 ();
 sg13g2_fill_1 FILLER_44_1101 ();
 sg13g2_fill_2 FILLER_44_1138 ();
 sg13g2_fill_2 FILLER_44_1175 ();
 sg13g2_fill_2 FILLER_44_1203 ();
 sg13g2_fill_1 FILLER_44_1205 ();
 sg13g2_fill_2 FILLER_44_1232 ();
 sg13g2_fill_1 FILLER_44_1234 ();
 sg13g2_decap_8 FILLER_44_1274 ();
 sg13g2_decap_4 FILLER_44_1281 ();
 sg13g2_fill_2 FILLER_44_1285 ();
 sg13g2_fill_1 FILLER_44_1297 ();
 sg13g2_fill_1 FILLER_44_1314 ();
 sg13g2_decap_4 FILLER_44_1341 ();
 sg13g2_fill_1 FILLER_44_1350 ();
 sg13g2_fill_2 FILLER_44_1377 ();
 sg13g2_fill_1 FILLER_44_1379 ();
 sg13g2_decap_4 FILLER_44_1403 ();
 sg13g2_fill_2 FILLER_44_1407 ();
 sg13g2_fill_2 FILLER_44_1452 ();
 sg13g2_fill_2 FILLER_44_1567 ();
 sg13g2_fill_1 FILLER_44_1583 ();
 sg13g2_fill_1 FILLER_44_1628 ();
 sg13g2_fill_1 FILLER_44_1679 ();
 sg13g2_fill_2 FILLER_44_1727 ();
 sg13g2_fill_1 FILLER_44_1750 ();
 sg13g2_decap_8 FILLER_44_1755 ();
 sg13g2_decap_4 FILLER_44_1762 ();
 sg13g2_fill_2 FILLER_44_1766 ();
 sg13g2_decap_8 FILLER_44_1802 ();
 sg13g2_decap_4 FILLER_44_1809 ();
 sg13g2_fill_1 FILLER_44_1813 ();
 sg13g2_fill_2 FILLER_44_1822 ();
 sg13g2_fill_1 FILLER_44_1824 ();
 sg13g2_fill_2 FILLER_44_1851 ();
 sg13g2_fill_2 FILLER_44_1895 ();
 sg13g2_fill_2 FILLER_44_1944 ();
 sg13g2_fill_1 FILLER_44_2015 ();
 sg13g2_decap_8 FILLER_44_2051 ();
 sg13g2_decap_4 FILLER_44_2058 ();
 sg13g2_decap_8 FILLER_44_2101 ();
 sg13g2_fill_1 FILLER_44_2144 ();
 sg13g2_fill_2 FILLER_44_2158 ();
 sg13g2_fill_1 FILLER_44_2160 ();
 sg13g2_fill_1 FILLER_44_2165 ();
 sg13g2_fill_1 FILLER_44_2179 ();
 sg13g2_fill_2 FILLER_44_2215 ();
 sg13g2_fill_2 FILLER_44_2251 ();
 sg13g2_decap_4 FILLER_44_2341 ();
 sg13g2_decap_8 FILLER_44_2349 ();
 sg13g2_decap_4 FILLER_44_2364 ();
 sg13g2_fill_1 FILLER_44_2385 ();
 sg13g2_decap_8 FILLER_44_2410 ();
 sg13g2_decap_4 FILLER_44_2421 ();
 sg13g2_fill_1 FILLER_44_2433 ();
 sg13g2_fill_1 FILLER_44_2442 ();
 sg13g2_fill_1 FILLER_44_2466 ();
 sg13g2_fill_1 FILLER_44_2493 ();
 sg13g2_fill_2 FILLER_44_2520 ();
 sg13g2_fill_1 FILLER_44_2522 ();
 sg13g2_fill_2 FILLER_44_2570 ();
 sg13g2_fill_1 FILLER_44_2572 ();
 sg13g2_fill_2 FILLER_44_2587 ();
 sg13g2_decap_8 FILLER_44_2628 ();
 sg13g2_decap_8 FILLER_44_2635 ();
 sg13g2_decap_8 FILLER_44_2642 ();
 sg13g2_decap_8 FILLER_44_2649 ();
 sg13g2_decap_8 FILLER_44_2656 ();
 sg13g2_decap_8 FILLER_44_2663 ();
 sg13g2_decap_4 FILLER_44_2670 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_decap_8 FILLER_45_476 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_decap_8 FILLER_45_490 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_4 FILLER_45_511 ();
 sg13g2_fill_1 FILLER_45_515 ();
 sg13g2_fill_1 FILLER_45_529 ();
 sg13g2_fill_1 FILLER_45_538 ();
 sg13g2_fill_1 FILLER_45_543 ();
 sg13g2_decap_4 FILLER_45_548 ();
 sg13g2_fill_1 FILLER_45_552 ();
 sg13g2_fill_1 FILLER_45_583 ();
 sg13g2_fill_2 FILLER_45_640 ();
 sg13g2_fill_1 FILLER_45_642 ();
 sg13g2_fill_1 FILLER_45_742 ();
 sg13g2_fill_1 FILLER_45_781 ();
 sg13g2_fill_2 FILLER_45_819 ();
 sg13g2_fill_2 FILLER_45_829 ();
 sg13g2_fill_1 FILLER_45_831 ();
 sg13g2_fill_1 FILLER_45_888 ();
 sg13g2_fill_1 FILLER_45_898 ();
 sg13g2_fill_2 FILLER_45_916 ();
 sg13g2_fill_1 FILLER_45_918 ();
 sg13g2_fill_1 FILLER_45_928 ();
 sg13g2_fill_2 FILLER_45_943 ();
 sg13g2_fill_1 FILLER_45_945 ();
 sg13g2_fill_2 FILLER_45_952 ();
 sg13g2_fill_2 FILLER_45_1027 ();
 sg13g2_fill_2 FILLER_45_1042 ();
 sg13g2_fill_2 FILLER_45_1080 ();
 sg13g2_fill_1 FILLER_45_1174 ();
 sg13g2_fill_2 FILLER_45_1223 ();
 sg13g2_decap_8 FILLER_45_1278 ();
 sg13g2_decap_4 FILLER_45_1285 ();
 sg13g2_fill_2 FILLER_45_1289 ();
 sg13g2_decap_8 FILLER_45_1324 ();
 sg13g2_decap_8 FILLER_45_1331 ();
 sg13g2_decap_8 FILLER_45_1338 ();
 sg13g2_decap_8 FILLER_45_1345 ();
 sg13g2_decap_4 FILLER_45_1352 ();
 sg13g2_fill_1 FILLER_45_1356 ();
 sg13g2_fill_2 FILLER_45_1375 ();
 sg13g2_fill_1 FILLER_45_1377 ();
 sg13g2_fill_1 FILLER_45_1416 ();
 sg13g2_fill_1 FILLER_45_1443 ();
 sg13g2_fill_2 FILLER_45_1506 ();
 sg13g2_decap_4 FILLER_45_1513 ();
 sg13g2_fill_2 FILLER_45_1517 ();
 sg13g2_fill_2 FILLER_45_1532 ();
 sg13g2_fill_2 FILLER_45_1539 ();
 sg13g2_fill_1 FILLER_45_1541 ();
 sg13g2_fill_2 FILLER_45_1551 ();
 sg13g2_fill_1 FILLER_45_1553 ();
 sg13g2_fill_2 FILLER_45_1646 ();
 sg13g2_fill_2 FILLER_45_1678 ();
 sg13g2_fill_2 FILLER_45_1790 ();
 sg13g2_fill_2 FILLER_45_1801 ();
 sg13g2_fill_1 FILLER_45_1803 ();
 sg13g2_fill_1 FILLER_45_1843 ();
 sg13g2_fill_1 FILLER_45_1925 ();
 sg13g2_fill_2 FILLER_45_1971 ();
 sg13g2_decap_8 FILLER_45_2062 ();
 sg13g2_decap_4 FILLER_45_2069 ();
 sg13g2_fill_2 FILLER_45_2073 ();
 sg13g2_decap_4 FILLER_45_2083 ();
 sg13g2_fill_2 FILLER_45_2087 ();
 sg13g2_decap_8 FILLER_45_2102 ();
 sg13g2_decap_8 FILLER_45_2158 ();
 sg13g2_decap_4 FILLER_45_2165 ();
 sg13g2_fill_2 FILLER_45_2169 ();
 sg13g2_fill_2 FILLER_45_2180 ();
 sg13g2_fill_1 FILLER_45_2187 ();
 sg13g2_fill_1 FILLER_45_2197 ();
 sg13g2_fill_2 FILLER_45_2211 ();
 sg13g2_fill_2 FILLER_45_2259 ();
 sg13g2_fill_1 FILLER_45_2261 ();
 sg13g2_fill_2 FILLER_45_2297 ();
 sg13g2_decap_8 FILLER_45_2355 ();
 sg13g2_decap_8 FILLER_45_2362 ();
 sg13g2_fill_2 FILLER_45_2369 ();
 sg13g2_fill_1 FILLER_45_2371 ();
 sg13g2_fill_1 FILLER_45_2377 ();
 sg13g2_fill_2 FILLER_45_2398 ();
 sg13g2_fill_1 FILLER_45_2400 ();
 sg13g2_fill_2 FILLER_45_2427 ();
 sg13g2_fill_1 FILLER_45_2429 ();
 sg13g2_fill_2 FILLER_45_2462 ();
 sg13g2_fill_1 FILLER_45_2464 ();
 sg13g2_decap_8 FILLER_45_2514 ();
 sg13g2_fill_2 FILLER_45_2521 ();
 sg13g2_fill_2 FILLER_45_2542 ();
 sg13g2_fill_2 FILLER_45_2567 ();
 sg13g2_fill_1 FILLER_45_2569 ();
 sg13g2_fill_2 FILLER_45_2579 ();
 sg13g2_fill_1 FILLER_45_2604 ();
 sg13g2_decap_8 FILLER_45_2631 ();
 sg13g2_decap_8 FILLER_45_2638 ();
 sg13g2_decap_8 FILLER_45_2645 ();
 sg13g2_decap_8 FILLER_45_2652 ();
 sg13g2_decap_8 FILLER_45_2659 ();
 sg13g2_decap_8 FILLER_45_2666 ();
 sg13g2_fill_1 FILLER_45_2673 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_4 FILLER_46_504 ();
 sg13g2_fill_2 FILLER_46_508 ();
 sg13g2_fill_2 FILLER_46_513 ();
 sg13g2_fill_1 FILLER_46_515 ();
 sg13g2_fill_1 FILLER_46_524 ();
 sg13g2_fill_2 FILLER_46_533 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_fill_2 FILLER_46_579 ();
 sg13g2_fill_1 FILLER_46_581 ();
 sg13g2_fill_2 FILLER_46_715 ();
 sg13g2_fill_2 FILLER_46_798 ();
 sg13g2_decap_4 FILLER_46_829 ();
 sg13g2_fill_2 FILLER_46_833 ();
 sg13g2_fill_2 FILLER_46_867 ();
 sg13g2_fill_2 FILLER_46_878 ();
 sg13g2_fill_2 FILLER_46_910 ();
 sg13g2_fill_1 FILLER_46_912 ();
 sg13g2_fill_1 FILLER_46_934 ();
 sg13g2_fill_1 FILLER_46_960 ();
 sg13g2_decap_8 FILLER_46_965 ();
 sg13g2_fill_2 FILLER_46_972 ();
 sg13g2_decap_4 FILLER_46_979 ();
 sg13g2_fill_1 FILLER_46_983 ();
 sg13g2_decap_8 FILLER_46_1028 ();
 sg13g2_fill_1 FILLER_46_1035 ();
 sg13g2_fill_1 FILLER_46_1138 ();
 sg13g2_fill_2 FILLER_46_1174 ();
 sg13g2_fill_1 FILLER_46_1176 ();
 sg13g2_fill_1 FILLER_46_1216 ();
 sg13g2_decap_8 FILLER_46_1274 ();
 sg13g2_fill_1 FILLER_46_1281 ();
 sg13g2_fill_1 FILLER_46_1324 ();
 sg13g2_decap_8 FILLER_46_1329 ();
 sg13g2_decap_8 FILLER_46_1336 ();
 sg13g2_decap_8 FILLER_46_1343 ();
 sg13g2_decap_8 FILLER_46_1350 ();
 sg13g2_decap_8 FILLER_46_1357 ();
 sg13g2_decap_8 FILLER_46_1364 ();
 sg13g2_decap_4 FILLER_46_1371 ();
 sg13g2_decap_8 FILLER_46_1379 ();
 sg13g2_fill_2 FILLER_46_1399 ();
 sg13g2_fill_1 FILLER_46_1419 ();
 sg13g2_fill_2 FILLER_46_1465 ();
 sg13g2_decap_4 FILLER_46_1492 ();
 sg13g2_fill_1 FILLER_46_1496 ();
 sg13g2_fill_1 FILLER_46_1502 ();
 sg13g2_decap_4 FILLER_46_1511 ();
 sg13g2_fill_1 FILLER_46_1515 ();
 sg13g2_fill_2 FILLER_46_1623 ();
 sg13g2_fill_1 FILLER_46_1625 ();
 sg13g2_fill_2 FILLER_46_1684 ();
 sg13g2_fill_2 FILLER_46_1698 ();
 sg13g2_fill_1 FILLER_46_1705 ();
 sg13g2_fill_2 FILLER_46_1716 ();
 sg13g2_fill_1 FILLER_46_1744 ();
 sg13g2_fill_2 FILLER_46_1755 ();
 sg13g2_fill_1 FILLER_46_1757 ();
 sg13g2_fill_1 FILLER_46_1763 ();
 sg13g2_fill_2 FILLER_46_1835 ();
 sg13g2_fill_1 FILLER_46_1837 ();
 sg13g2_fill_2 FILLER_46_1852 ();
 sg13g2_fill_1 FILLER_46_1877 ();
 sg13g2_fill_2 FILLER_46_1914 ();
 sg13g2_fill_2 FILLER_46_1925 ();
 sg13g2_fill_1 FILLER_46_2059 ();
 sg13g2_decap_8 FILLER_46_2077 ();
 sg13g2_decap_8 FILLER_46_2084 ();
 sg13g2_decap_8 FILLER_46_2091 ();
 sg13g2_fill_1 FILLER_46_2142 ();
 sg13g2_decap_8 FILLER_46_2178 ();
 sg13g2_fill_1 FILLER_46_2185 ();
 sg13g2_fill_2 FILLER_46_2215 ();
 sg13g2_decap_8 FILLER_46_2254 ();
 sg13g2_decap_4 FILLER_46_2261 ();
 sg13g2_fill_2 FILLER_46_2265 ();
 sg13g2_fill_1 FILLER_46_2298 ();
 sg13g2_fill_2 FILLER_46_2361 ();
 sg13g2_fill_1 FILLER_46_2363 ();
 sg13g2_fill_1 FILLER_46_2393 ();
 sg13g2_fill_2 FILLER_46_2420 ();
 sg13g2_fill_1 FILLER_46_2422 ();
 sg13g2_fill_2 FILLER_46_2449 ();
 sg13g2_decap_4 FILLER_46_2456 ();
 sg13g2_fill_2 FILLER_46_2460 ();
 sg13g2_decap_8 FILLER_46_2501 ();
 sg13g2_decap_8 FILLER_46_2508 ();
 sg13g2_decap_8 FILLER_46_2515 ();
 sg13g2_decap_4 FILLER_46_2522 ();
 sg13g2_fill_2 FILLER_46_2526 ();
 sg13g2_fill_1 FILLER_46_2571 ();
 sg13g2_fill_2 FILLER_46_2584 ();
 sg13g2_decap_8 FILLER_46_2627 ();
 sg13g2_decap_8 FILLER_46_2634 ();
 sg13g2_decap_8 FILLER_46_2641 ();
 sg13g2_decap_8 FILLER_46_2648 ();
 sg13g2_decap_8 FILLER_46_2655 ();
 sg13g2_decap_8 FILLER_46_2662 ();
 sg13g2_decap_4 FILLER_46_2669 ();
 sg13g2_fill_1 FILLER_46_2673 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_fill_2 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_554 ();
 sg13g2_fill_1 FILLER_47_561 ();
 sg13g2_fill_2 FILLER_47_570 ();
 sg13g2_fill_1 FILLER_47_628 ();
 sg13g2_fill_2 FILLER_47_638 ();
 sg13g2_fill_1 FILLER_47_640 ();
 sg13g2_decap_4 FILLER_47_691 ();
 sg13g2_fill_2 FILLER_47_695 ();
 sg13g2_fill_2 FILLER_47_702 ();
 sg13g2_fill_1 FILLER_47_721 ();
 sg13g2_fill_2 FILLER_47_731 ();
 sg13g2_fill_2 FILLER_47_764 ();
 sg13g2_fill_1 FILLER_47_788 ();
 sg13g2_fill_1 FILLER_47_820 ();
 sg13g2_fill_1 FILLER_47_825 ();
 sg13g2_decap_8 FILLER_47_834 ();
 sg13g2_decap_4 FILLER_47_841 ();
 sg13g2_fill_2 FILLER_47_845 ();
 sg13g2_fill_2 FILLER_47_851 ();
 sg13g2_fill_2 FILLER_47_858 ();
 sg13g2_fill_1 FILLER_47_860 ();
 sg13g2_fill_2 FILLER_47_920 ();
 sg13g2_fill_1 FILLER_47_922 ();
 sg13g2_decap_8 FILLER_47_982 ();
 sg13g2_fill_1 FILLER_47_989 ();
 sg13g2_fill_2 FILLER_47_1040 ();
 sg13g2_fill_1 FILLER_47_1099 ();
 sg13g2_fill_2 FILLER_47_1133 ();
 sg13g2_decap_8 FILLER_47_1165 ();
 sg13g2_fill_1 FILLER_47_1172 ();
 sg13g2_fill_2 FILLER_47_1181 ();
 sg13g2_fill_1 FILLER_47_1183 ();
 sg13g2_fill_1 FILLER_47_1189 ();
 sg13g2_fill_2 FILLER_47_1242 ();
 sg13g2_fill_2 FILLER_47_1275 ();
 sg13g2_fill_2 FILLER_47_1338 ();
 sg13g2_fill_2 FILLER_47_1374 ();
 sg13g2_fill_2 FILLER_47_1384 ();
 sg13g2_fill_1 FILLER_47_1386 ();
 sg13g2_fill_2 FILLER_47_1418 ();
 sg13g2_fill_2 FILLER_47_1425 ();
 sg13g2_fill_1 FILLER_47_1427 ();
 sg13g2_fill_2 FILLER_47_1436 ();
 sg13g2_fill_1 FILLER_47_1452 ();
 sg13g2_fill_2 FILLER_47_1512 ();
 sg13g2_fill_1 FILLER_47_1540 ();
 sg13g2_fill_1 FILLER_47_1604 ();
 sg13g2_fill_1 FILLER_47_1643 ();
 sg13g2_fill_2 FILLER_47_1713 ();
 sg13g2_fill_1 FILLER_47_1715 ();
 sg13g2_fill_1 FILLER_47_1725 ();
 sg13g2_fill_1 FILLER_47_1753 ();
 sg13g2_fill_2 FILLER_47_1797 ();
 sg13g2_fill_1 FILLER_47_1799 ();
 sg13g2_fill_1 FILLER_47_1851 ();
 sg13g2_fill_1 FILLER_47_1883 ();
 sg13g2_fill_1 FILLER_47_1973 ();
 sg13g2_fill_1 FILLER_47_1996 ();
 sg13g2_fill_2 FILLER_47_2015 ();
 sg13g2_fill_1 FILLER_47_2052 ();
 sg13g2_decap_4 FILLER_47_2088 ();
 sg13g2_fill_2 FILLER_47_2139 ();
 sg13g2_fill_1 FILLER_47_2141 ();
 sg13g2_fill_2 FILLER_47_2265 ();
 sg13g2_fill_1 FILLER_47_2267 ();
 sg13g2_fill_1 FILLER_47_2286 ();
 sg13g2_fill_1 FILLER_47_2296 ();
 sg13g2_fill_1 FILLER_47_2307 ();
 sg13g2_fill_1 FILLER_47_2318 ();
 sg13g2_fill_2 FILLER_47_2346 ();
 sg13g2_fill_1 FILLER_47_2348 ();
 sg13g2_fill_1 FILLER_47_2408 ();
 sg13g2_fill_2 FILLER_47_2483 ();
 sg13g2_fill_2 FILLER_47_2490 ();
 sg13g2_fill_1 FILLER_47_2492 ();
 sg13g2_fill_1 FILLER_47_2498 ();
 sg13g2_fill_1 FILLER_47_2520 ();
 sg13g2_decap_8 FILLER_47_2525 ();
 sg13g2_fill_2 FILLER_47_2536 ();
 sg13g2_fill_2 FILLER_47_2546 ();
 sg13g2_fill_1 FILLER_47_2548 ();
 sg13g2_fill_1 FILLER_47_2575 ();
 sg13g2_decap_8 FILLER_47_2616 ();
 sg13g2_decap_8 FILLER_47_2623 ();
 sg13g2_decap_8 FILLER_47_2630 ();
 sg13g2_decap_8 FILLER_47_2637 ();
 sg13g2_decap_8 FILLER_47_2644 ();
 sg13g2_decap_8 FILLER_47_2651 ();
 sg13g2_decap_8 FILLER_47_2658 ();
 sg13g2_decap_8 FILLER_47_2665 ();
 sg13g2_fill_2 FILLER_47_2672 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_fill_1 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_4 FILLER_48_469 ();
 sg13g2_fill_2 FILLER_48_473 ();
 sg13g2_decap_8 FILLER_48_480 ();
 sg13g2_decap_8 FILLER_48_487 ();
 sg13g2_decap_8 FILLER_48_494 ();
 sg13g2_decap_8 FILLER_48_501 ();
 sg13g2_decap_4 FILLER_48_508 ();
 sg13g2_fill_2 FILLER_48_549 ();
 sg13g2_decap_8 FILLER_48_565 ();
 sg13g2_decap_4 FILLER_48_576 ();
 sg13g2_fill_2 FILLER_48_580 ();
 sg13g2_fill_1 FILLER_48_634 ();
 sg13g2_fill_2 FILLER_48_644 ();
 sg13g2_fill_1 FILLER_48_646 ();
 sg13g2_fill_2 FILLER_48_669 ();
 sg13g2_fill_2 FILLER_48_686 ();
 sg13g2_fill_1 FILLER_48_688 ();
 sg13g2_fill_2 FILLER_48_706 ();
 sg13g2_fill_1 FILLER_48_716 ();
 sg13g2_fill_2 FILLER_48_747 ();
 sg13g2_fill_2 FILLER_48_769 ();
 sg13g2_fill_1 FILLER_48_797 ();
 sg13g2_decap_8 FILLER_48_824 ();
 sg13g2_decap_8 FILLER_48_831 ();
 sg13g2_fill_2 FILLER_48_874 ();
 sg13g2_fill_1 FILLER_48_876 ();
 sg13g2_fill_2 FILLER_48_902 ();
 sg13g2_fill_1 FILLER_48_904 ();
 sg13g2_fill_1 FILLER_48_912 ();
 sg13g2_fill_2 FILLER_48_998 ();
 sg13g2_decap_8 FILLER_48_1012 ();
 sg13g2_decap_4 FILLER_48_1019 ();
 sg13g2_fill_2 FILLER_48_1023 ();
 sg13g2_fill_1 FILLER_48_1072 ();
 sg13g2_fill_2 FILLER_48_1082 ();
 sg13g2_fill_2 FILLER_48_1157 ();
 sg13g2_fill_1 FILLER_48_1167 ();
 sg13g2_fill_1 FILLER_48_1172 ();
 sg13g2_decap_8 FILLER_48_1177 ();
 sg13g2_decap_4 FILLER_48_1184 ();
 sg13g2_fill_2 FILLER_48_1198 ();
 sg13g2_fill_1 FILLER_48_1212 ();
 sg13g2_decap_4 FILLER_48_1217 ();
 sg13g2_fill_1 FILLER_48_1221 ();
 sg13g2_fill_2 FILLER_48_1279 ();
 sg13g2_decap_4 FILLER_48_1338 ();
 sg13g2_fill_2 FILLER_48_1342 ();
 sg13g2_fill_2 FILLER_48_1389 ();
 sg13g2_fill_1 FILLER_48_1417 ();
 sg13g2_decap_8 FILLER_48_1444 ();
 sg13g2_decap_4 FILLER_48_1451 ();
 sg13g2_fill_2 FILLER_48_1455 ();
 sg13g2_fill_1 FILLER_48_1487 ();
 sg13g2_fill_1 FILLER_48_1538 ();
 sg13g2_fill_2 FILLER_48_1568 ();
 sg13g2_fill_1 FILLER_48_1570 ();
 sg13g2_decap_8 FILLER_48_1631 ();
 sg13g2_fill_2 FILLER_48_1638 ();
 sg13g2_fill_2 FILLER_48_1644 ();
 sg13g2_fill_2 FILLER_48_1650 ();
 sg13g2_fill_1 FILLER_48_1652 ();
 sg13g2_fill_1 FILLER_48_1766 ();
 sg13g2_fill_2 FILLER_48_1809 ();
 sg13g2_fill_1 FILLER_48_1811 ();
 sg13g2_decap_8 FILLER_48_1834 ();
 sg13g2_decap_8 FILLER_48_1841 ();
 sg13g2_decap_8 FILLER_48_1848 ();
 sg13g2_decap_8 FILLER_48_1855 ();
 sg13g2_decap_8 FILLER_48_1866 ();
 sg13g2_decap_4 FILLER_48_1873 ();
 sg13g2_fill_2 FILLER_48_1877 ();
 sg13g2_fill_2 FILLER_48_1910 ();
 sg13g2_fill_1 FILLER_48_1963 ();
 sg13g2_fill_1 FILLER_48_1969 ();
 sg13g2_fill_1 FILLER_48_1975 ();
 sg13g2_fill_1 FILLER_48_2096 ();
 sg13g2_fill_1 FILLER_48_2207 ();
 sg13g2_fill_2 FILLER_48_2217 ();
 sg13g2_fill_1 FILLER_48_2266 ();
 sg13g2_fill_2 FILLER_48_2284 ();
 sg13g2_fill_1 FILLER_48_2286 ();
 sg13g2_fill_2 FILLER_48_2305 ();
 sg13g2_fill_2 FILLER_48_2333 ();
 sg13g2_fill_2 FILLER_48_2401 ();
 sg13g2_fill_2 FILLER_48_2417 ();
 sg13g2_fill_1 FILLER_48_2458 ();
 sg13g2_fill_2 FILLER_48_2472 ();
 sg13g2_fill_1 FILLER_48_2474 ();
 sg13g2_fill_2 FILLER_48_2479 ();
 sg13g2_fill_1 FILLER_48_2525 ();
 sg13g2_fill_2 FILLER_48_2583 ();
 sg13g2_decap_8 FILLER_48_2620 ();
 sg13g2_decap_8 FILLER_48_2627 ();
 sg13g2_decap_8 FILLER_48_2634 ();
 sg13g2_decap_8 FILLER_48_2641 ();
 sg13g2_decap_8 FILLER_48_2648 ();
 sg13g2_decap_8 FILLER_48_2655 ();
 sg13g2_decap_8 FILLER_48_2662 ();
 sg13g2_decap_4 FILLER_48_2669 ();
 sg13g2_fill_1 FILLER_48_2673 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_4 FILLER_49_483 ();
 sg13g2_decap_4 FILLER_49_492 ();
 sg13g2_fill_2 FILLER_49_500 ();
 sg13g2_fill_1 FILLER_49_502 ();
 sg13g2_fill_1 FILLER_49_549 ();
 sg13g2_fill_2 FILLER_49_565 ();
 sg13g2_fill_1 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_576 ();
 sg13g2_fill_1 FILLER_49_603 ();
 sg13g2_fill_2 FILLER_49_617 ();
 sg13g2_fill_1 FILLER_49_619 ();
 sg13g2_fill_2 FILLER_49_681 ();
 sg13g2_fill_1 FILLER_49_732 ();
 sg13g2_fill_1 FILLER_49_737 ();
 sg13g2_fill_2 FILLER_49_781 ();
 sg13g2_fill_1 FILLER_49_788 ();
 sg13g2_fill_1 FILLER_49_802 ();
 sg13g2_decap_8 FILLER_49_816 ();
 sg13g2_fill_1 FILLER_49_823 ();
 sg13g2_fill_1 FILLER_49_891 ();
 sg13g2_fill_1 FILLER_49_931 ();
 sg13g2_fill_1 FILLER_49_955 ();
 sg13g2_fill_2 FILLER_49_1013 ();
 sg13g2_fill_1 FILLER_49_1015 ();
 sg13g2_fill_2 FILLER_49_1047 ();
 sg13g2_fill_1 FILLER_49_1049 ();
 sg13g2_fill_2 FILLER_49_1063 ();
 sg13g2_fill_2 FILLER_49_1073 ();
 sg13g2_fill_1 FILLER_49_1114 ();
 sg13g2_fill_1 FILLER_49_1128 ();
 sg13g2_fill_2 FILLER_49_1160 ();
 sg13g2_fill_1 FILLER_49_1162 ();
 sg13g2_fill_1 FILLER_49_1248 ();
 sg13g2_fill_2 FILLER_49_1259 ();
 sg13g2_decap_8 FILLER_49_1319 ();
 sg13g2_fill_1 FILLER_49_1388 ();
 sg13g2_fill_1 FILLER_49_1415 ();
 sg13g2_fill_1 FILLER_49_1446 ();
 sg13g2_fill_1 FILLER_49_1451 ();
 sg13g2_fill_1 FILLER_49_1465 ();
 sg13g2_decap_4 FILLER_49_1484 ();
 sg13g2_fill_1 FILLER_49_1531 ();
 sg13g2_fill_2 FILLER_49_1544 ();
 sg13g2_fill_2 FILLER_49_1624 ();
 sg13g2_decap_8 FILLER_49_1640 ();
 sg13g2_decap_8 FILLER_49_1647 ();
 sg13g2_fill_2 FILLER_49_1685 ();
 sg13g2_fill_1 FILLER_49_1708 ();
 sg13g2_fill_1 FILLER_49_1722 ();
 sg13g2_fill_1 FILLER_49_1815 ();
 sg13g2_decap_4 FILLER_49_1842 ();
 sg13g2_fill_2 FILLER_49_1846 ();
 sg13g2_fill_2 FILLER_49_1879 ();
 sg13g2_fill_1 FILLER_49_1881 ();
 sg13g2_fill_2 FILLER_49_1899 ();
 sg13g2_fill_1 FILLER_49_1901 ();
 sg13g2_fill_2 FILLER_49_1970 ();
 sg13g2_fill_1 FILLER_49_2043 ();
 sg13g2_fill_1 FILLER_49_2092 ();
 sg13g2_decap_4 FILLER_49_2102 ();
 sg13g2_fill_2 FILLER_49_2106 ();
 sg13g2_fill_2 FILLER_49_2139 ();
 sg13g2_fill_2 FILLER_49_2181 ();
 sg13g2_fill_1 FILLER_49_2209 ();
 sg13g2_decap_4 FILLER_49_2224 ();
 sg13g2_fill_2 FILLER_49_2260 ();
 sg13g2_fill_1 FILLER_49_2262 ();
 sg13g2_fill_2 FILLER_49_2289 ();
 sg13g2_fill_1 FILLER_49_2291 ();
 sg13g2_fill_2 FILLER_49_2348 ();
 sg13g2_fill_1 FILLER_49_2350 ();
 sg13g2_fill_2 FILLER_49_2381 ();
 sg13g2_fill_2 FILLER_49_2388 ();
 sg13g2_fill_1 FILLER_49_2390 ();
 sg13g2_fill_1 FILLER_49_2417 ();
 sg13g2_fill_2 FILLER_49_2427 ();
 sg13g2_fill_2 FILLER_49_2485 ();
 sg13g2_fill_2 FILLER_49_2513 ();
 sg13g2_fill_1 FILLER_49_2515 ();
 sg13g2_fill_2 FILLER_49_2521 ();
 sg13g2_fill_1 FILLER_49_2567 ();
 sg13g2_decap_8 FILLER_49_2620 ();
 sg13g2_decap_8 FILLER_49_2627 ();
 sg13g2_decap_8 FILLER_49_2634 ();
 sg13g2_decap_8 FILLER_49_2641 ();
 sg13g2_decap_8 FILLER_49_2648 ();
 sg13g2_decap_8 FILLER_49_2655 ();
 sg13g2_decap_8 FILLER_49_2662 ();
 sg13g2_decap_4 FILLER_49_2669 ();
 sg13g2_fill_1 FILLER_49_2673 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_203 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_decap_8 FILLER_50_224 ();
 sg13g2_decap_8 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_decap_8 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_259 ();
 sg13g2_decap_8 FILLER_50_266 ();
 sg13g2_decap_8 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_decap_8 FILLER_50_287 ();
 sg13g2_decap_8 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_301 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_315 ();
 sg13g2_decap_8 FILLER_50_322 ();
 sg13g2_decap_8 FILLER_50_329 ();
 sg13g2_decap_8 FILLER_50_336 ();
 sg13g2_decap_8 FILLER_50_343 ();
 sg13g2_decap_8 FILLER_50_350 ();
 sg13g2_decap_8 FILLER_50_357 ();
 sg13g2_decap_8 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_371 ();
 sg13g2_decap_8 FILLER_50_378 ();
 sg13g2_decap_8 FILLER_50_385 ();
 sg13g2_decap_8 FILLER_50_392 ();
 sg13g2_decap_8 FILLER_50_399 ();
 sg13g2_decap_8 FILLER_50_406 ();
 sg13g2_decap_8 FILLER_50_413 ();
 sg13g2_decap_8 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_427 ();
 sg13g2_decap_8 FILLER_50_434 ();
 sg13g2_decap_8 FILLER_50_441 ();
 sg13g2_decap_8 FILLER_50_448 ();
 sg13g2_decap_8 FILLER_50_455 ();
 sg13g2_decap_8 FILLER_50_462 ();
 sg13g2_fill_1 FILLER_50_469 ();
 sg13g2_fill_1 FILLER_50_501 ();
 sg13g2_fill_1 FILLER_50_512 ();
 sg13g2_fill_2 FILLER_50_574 ();
 sg13g2_fill_1 FILLER_50_576 ();
 sg13g2_fill_1 FILLER_50_581 ();
 sg13g2_decap_4 FILLER_50_592 ();
 sg13g2_decap_4 FILLER_50_604 ();
 sg13g2_fill_1 FILLER_50_612 ();
 sg13g2_fill_2 FILLER_50_617 ();
 sg13g2_fill_1 FILLER_50_649 ();
 sg13g2_fill_2 FILLER_50_682 ();
 sg13g2_fill_1 FILLER_50_714 ();
 sg13g2_fill_1 FILLER_50_771 ();
 sg13g2_fill_1 FILLER_50_777 ();
 sg13g2_fill_1 FILLER_50_788 ();
 sg13g2_fill_2 FILLER_50_804 ();
 sg13g2_fill_1 FILLER_50_815 ();
 sg13g2_fill_2 FILLER_50_854 ();
 sg13g2_fill_2 FILLER_50_881 ();
 sg13g2_fill_1 FILLER_50_883 ();
 sg13g2_fill_2 FILLER_50_933 ();
 sg13g2_fill_2 FILLER_50_1013 ();
 sg13g2_fill_1 FILLER_50_1015 ();
 sg13g2_decap_4 FILLER_50_1052 ();
 sg13g2_fill_2 FILLER_50_1069 ();
 sg13g2_decap_4 FILLER_50_1093 ();
 sg13g2_fill_2 FILLER_50_1097 ();
 sg13g2_fill_2 FILLER_50_1102 ();
 sg13g2_fill_1 FILLER_50_1104 ();
 sg13g2_decap_4 FILLER_50_1110 ();
 sg13g2_fill_2 FILLER_50_1114 ();
 sg13g2_decap_8 FILLER_50_1133 ();
 sg13g2_decap_8 FILLER_50_1140 ();
 sg13g2_decap_4 FILLER_50_1147 ();
 sg13g2_fill_2 FILLER_50_1171 ();
 sg13g2_fill_1 FILLER_50_1173 ();
 sg13g2_fill_1 FILLER_50_1203 ();
 sg13g2_fill_1 FILLER_50_1238 ();
 sg13g2_fill_1 FILLER_50_1252 ();
 sg13g2_fill_2 FILLER_50_1273 ();
 sg13g2_decap_8 FILLER_50_1321 ();
 sg13g2_decap_8 FILLER_50_1328 ();
 sg13g2_fill_2 FILLER_50_1335 ();
 sg13g2_fill_1 FILLER_50_1337 ();
 sg13g2_fill_2 FILLER_50_1377 ();
 sg13g2_fill_1 FILLER_50_1443 ();
 sg13g2_fill_1 FILLER_50_1459 ();
 sg13g2_fill_2 FILLER_50_1524 ();
 sg13g2_fill_1 FILLER_50_1526 ();
 sg13g2_fill_2 FILLER_50_1552 ();
 sg13g2_fill_1 FILLER_50_1554 ();
 sg13g2_fill_2 FILLER_50_1595 ();
 sg13g2_fill_1 FILLER_50_1623 ();
 sg13g2_fill_2 FILLER_50_1637 ();
 sg13g2_fill_2 FILLER_50_1665 ();
 sg13g2_fill_1 FILLER_50_1675 ();
 sg13g2_fill_2 FILLER_50_1766 ();
 sg13g2_fill_2 FILLER_50_1774 ();
 sg13g2_fill_1 FILLER_50_1776 ();
 sg13g2_fill_2 FILLER_50_1811 ();
 sg13g2_decap_4 FILLER_50_1839 ();
 sg13g2_fill_2 FILLER_50_1843 ();
 sg13g2_decap_4 FILLER_50_1889 ();
 sg13g2_fill_1 FILLER_50_1942 ();
 sg13g2_fill_2 FILLER_50_1968 ();
 sg13g2_fill_2 FILLER_50_1981 ();
 sg13g2_fill_2 FILLER_50_2058 ();
 sg13g2_fill_1 FILLER_50_2060 ();
 sg13g2_fill_2 FILLER_50_2082 ();
 sg13g2_fill_1 FILLER_50_2097 ();
 sg13g2_fill_2 FILLER_50_2106 ();
 sg13g2_fill_1 FILLER_50_2108 ();
 sg13g2_fill_2 FILLER_50_2117 ();
 sg13g2_fill_2 FILLER_50_2123 ();
 sg13g2_fill_2 FILLER_50_2148 ();
 sg13g2_fill_1 FILLER_50_2150 ();
 sg13g2_fill_1 FILLER_50_2172 ();
 sg13g2_decap_4 FILLER_50_2178 ();
 sg13g2_fill_2 FILLER_50_2216 ();
 sg13g2_fill_1 FILLER_50_2218 ();
 sg13g2_decap_4 FILLER_50_2227 ();
 sg13g2_fill_2 FILLER_50_2247 ();
 sg13g2_fill_1 FILLER_50_2249 ();
 sg13g2_fill_2 FILLER_50_2302 ();
 sg13g2_fill_1 FILLER_50_2338 ();
 sg13g2_fill_2 FILLER_50_2373 ();
 sg13g2_fill_1 FILLER_50_2375 ();
 sg13g2_fill_2 FILLER_50_2385 ();
 sg13g2_fill_1 FILLER_50_2387 ();
 sg13g2_fill_2 FILLER_50_2414 ();
 sg13g2_fill_2 FILLER_50_2459 ();
 sg13g2_fill_1 FILLER_50_2461 ();
 sg13g2_fill_1 FILLER_50_2488 ();
 sg13g2_fill_2 FILLER_50_2538 ();
 sg13g2_fill_1 FILLER_50_2540 ();
 sg13g2_fill_2 FILLER_50_2560 ();
 sg13g2_fill_1 FILLER_50_2562 ();
 sg13g2_fill_1 FILLER_50_2568 ();
 sg13g2_fill_2 FILLER_50_2582 ();
 sg13g2_fill_1 FILLER_50_2584 ();
 sg13g2_fill_1 FILLER_50_2603 ();
 sg13g2_decap_8 FILLER_50_2622 ();
 sg13g2_decap_8 FILLER_50_2629 ();
 sg13g2_decap_8 FILLER_50_2636 ();
 sg13g2_decap_8 FILLER_50_2643 ();
 sg13g2_decap_8 FILLER_50_2650 ();
 sg13g2_decap_8 FILLER_50_2657 ();
 sg13g2_decap_8 FILLER_50_2664 ();
 sg13g2_fill_2 FILLER_50_2671 ();
 sg13g2_fill_1 FILLER_50_2673 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_182 ();
 sg13g2_decap_8 FILLER_51_189 ();
 sg13g2_decap_8 FILLER_51_196 ();
 sg13g2_decap_8 FILLER_51_203 ();
 sg13g2_decap_8 FILLER_51_210 ();
 sg13g2_decap_8 FILLER_51_217 ();
 sg13g2_decap_8 FILLER_51_224 ();
 sg13g2_decap_8 FILLER_51_231 ();
 sg13g2_decap_8 FILLER_51_238 ();
 sg13g2_decap_8 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_252 ();
 sg13g2_decap_8 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_266 ();
 sg13g2_decap_8 FILLER_51_273 ();
 sg13g2_decap_8 FILLER_51_280 ();
 sg13g2_decap_8 FILLER_51_287 ();
 sg13g2_decap_8 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_301 ();
 sg13g2_decap_8 FILLER_51_308 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_decap_8 FILLER_51_322 ();
 sg13g2_decap_8 FILLER_51_329 ();
 sg13g2_decap_8 FILLER_51_336 ();
 sg13g2_decap_8 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_350 ();
 sg13g2_decap_8 FILLER_51_357 ();
 sg13g2_decap_8 FILLER_51_364 ();
 sg13g2_decap_8 FILLER_51_371 ();
 sg13g2_decap_8 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_decap_8 FILLER_51_406 ();
 sg13g2_decap_8 FILLER_51_413 ();
 sg13g2_decap_8 FILLER_51_420 ();
 sg13g2_decap_8 FILLER_51_427 ();
 sg13g2_decap_8 FILLER_51_434 ();
 sg13g2_decap_8 FILLER_51_441 ();
 sg13g2_decap_8 FILLER_51_448 ();
 sg13g2_decap_8 FILLER_51_455 ();
 sg13g2_decap_8 FILLER_51_462 ();
 sg13g2_fill_1 FILLER_51_552 ();
 sg13g2_fill_1 FILLER_51_572 ();
 sg13g2_decap_8 FILLER_51_592 ();
 sg13g2_decap_8 FILLER_51_599 ();
 sg13g2_decap_8 FILLER_51_606 ();
 sg13g2_fill_1 FILLER_51_613 ();
 sg13g2_fill_1 FILLER_51_636 ();
 sg13g2_fill_2 FILLER_51_642 ();
 sg13g2_fill_1 FILLER_51_658 ();
 sg13g2_fill_2 FILLER_51_677 ();
 sg13g2_fill_1 FILLER_51_679 ();
 sg13g2_fill_1 FILLER_51_715 ();
 sg13g2_fill_2 FILLER_51_751 ();
 sg13g2_fill_1 FILLER_51_771 ();
 sg13g2_fill_2 FILLER_51_831 ();
 sg13g2_fill_2 FILLER_51_865 ();
 sg13g2_fill_1 FILLER_51_867 ();
 sg13g2_fill_1 FILLER_51_933 ();
 sg13g2_fill_1 FILLER_51_996 ();
 sg13g2_fill_2 FILLER_51_1010 ();
 sg13g2_fill_2 FILLER_51_1042 ();
 sg13g2_decap_8 FILLER_51_1052 ();
 sg13g2_decap_8 FILLER_51_1059 ();
 sg13g2_decap_8 FILLER_51_1066 ();
 sg13g2_decap_4 FILLER_51_1073 ();
 sg13g2_fill_2 FILLER_51_1077 ();
 sg13g2_decap_8 FILLER_51_1083 ();
 sg13g2_decap_8 FILLER_51_1090 ();
 sg13g2_decap_8 FILLER_51_1097 ();
 sg13g2_decap_4 FILLER_51_1104 ();
 sg13g2_fill_2 FILLER_51_1134 ();
 sg13g2_fill_1 FILLER_51_1136 ();
 sg13g2_fill_1 FILLER_51_1176 ();
 sg13g2_fill_2 FILLER_51_1215 ();
 sg13g2_fill_1 FILLER_51_1221 ();
 sg13g2_fill_2 FILLER_51_1227 ();
 sg13g2_fill_1 FILLER_51_1229 ();
 sg13g2_fill_2 FILLER_51_1271 ();
 sg13g2_decap_4 FILLER_51_1277 ();
 sg13g2_fill_1 FILLER_51_1281 ();
 sg13g2_decap_8 FILLER_51_1318 ();
 sg13g2_fill_2 FILLER_51_1325 ();
 sg13g2_fill_2 FILLER_51_1348 ();
 sg13g2_fill_1 FILLER_51_1350 ();
 sg13g2_fill_2 FILLER_51_1382 ();
 sg13g2_fill_2 FILLER_51_1410 ();
 sg13g2_fill_1 FILLER_51_1412 ();
 sg13g2_decap_4 FILLER_51_1488 ();
 sg13g2_fill_2 FILLER_51_1501 ();
 sg13g2_fill_1 FILLER_51_1503 ();
 sg13g2_fill_2 FILLER_51_1564 ();
 sg13g2_fill_1 FILLER_51_1566 ();
 sg13g2_fill_1 FILLER_51_1577 ();
 sg13g2_fill_1 FILLER_51_1594 ();
 sg13g2_fill_2 FILLER_51_1669 ();
 sg13g2_fill_1 FILLER_51_1671 ();
 sg13g2_fill_1 FILLER_51_1720 ();
 sg13g2_fill_1 FILLER_51_1773 ();
 sg13g2_fill_1 FILLER_51_1782 ();
 sg13g2_decap_8 FILLER_51_1806 ();
 sg13g2_decap_4 FILLER_51_1813 ();
 sg13g2_fill_1 FILLER_51_1817 ();
 sg13g2_fill_2 FILLER_51_1858 ();
 sg13g2_fill_1 FILLER_51_1860 ();
 sg13g2_decap_8 FILLER_51_1883 ();
 sg13g2_fill_2 FILLER_51_1890 ();
 sg13g2_fill_2 FILLER_51_1925 ();
 sg13g2_fill_2 FILLER_51_1953 ();
 sg13g2_fill_2 FILLER_51_1963 ();
 sg13g2_fill_2 FILLER_51_1985 ();
 sg13g2_fill_1 FILLER_51_1991 ();
 sg13g2_fill_1 FILLER_51_2000 ();
 sg13g2_fill_2 FILLER_51_2033 ();
 sg13g2_fill_1 FILLER_51_2047 ();
 sg13g2_fill_2 FILLER_51_2053 ();
 sg13g2_fill_1 FILLER_51_2055 ();
 sg13g2_fill_1 FILLER_51_2061 ();
 sg13g2_fill_1 FILLER_51_2077 ();
 sg13g2_fill_2 FILLER_51_2090 ();
 sg13g2_decap_4 FILLER_51_2101 ();
 sg13g2_fill_2 FILLER_51_2105 ();
 sg13g2_decap_8 FILLER_51_2119 ();
 sg13g2_decap_8 FILLER_51_2126 ();
 sg13g2_fill_1 FILLER_51_2133 ();
 sg13g2_fill_1 FILLER_51_2147 ();
 sg13g2_fill_1 FILLER_51_2161 ();
 sg13g2_fill_2 FILLER_51_2175 ();
 sg13g2_fill_1 FILLER_51_2177 ();
 sg13g2_decap_4 FILLER_51_2183 ();
 sg13g2_fill_2 FILLER_51_2191 ();
 sg13g2_fill_1 FILLER_51_2197 ();
 sg13g2_fill_2 FILLER_51_2215 ();
 sg13g2_fill_2 FILLER_51_2282 ();
 sg13g2_decap_8 FILLER_51_2344 ();
 sg13g2_fill_1 FILLER_51_2351 ();
 sg13g2_fill_2 FILLER_51_2366 ();
 sg13g2_fill_1 FILLER_51_2368 ();
 sg13g2_decap_8 FILLER_51_2382 ();
 sg13g2_decap_8 FILLER_51_2389 ();
 sg13g2_fill_2 FILLER_51_2405 ();
 sg13g2_fill_1 FILLER_51_2407 ();
 sg13g2_fill_1 FILLER_51_2425 ();
 sg13g2_fill_2 FILLER_51_2499 ();
 sg13g2_fill_2 FILLER_51_2529 ();
 sg13g2_decap_8 FILLER_51_2544 ();
 sg13g2_fill_2 FILLER_51_2551 ();
 sg13g2_fill_2 FILLER_51_2557 ();
 sg13g2_fill_1 FILLER_51_2571 ();
 sg13g2_fill_2 FILLER_51_2598 ();
 sg13g2_decap_8 FILLER_51_2608 ();
 sg13g2_decap_8 FILLER_51_2615 ();
 sg13g2_decap_8 FILLER_51_2622 ();
 sg13g2_decap_8 FILLER_51_2629 ();
 sg13g2_decap_8 FILLER_51_2636 ();
 sg13g2_decap_8 FILLER_51_2643 ();
 sg13g2_decap_8 FILLER_51_2650 ();
 sg13g2_decap_8 FILLER_51_2657 ();
 sg13g2_decap_8 FILLER_51_2664 ();
 sg13g2_fill_2 FILLER_51_2671 ();
 sg13g2_fill_1 FILLER_51_2673 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_decap_8 FILLER_52_175 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_196 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_210 ();
 sg13g2_decap_8 FILLER_52_217 ();
 sg13g2_decap_8 FILLER_52_224 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_decap_8 FILLER_52_252 ();
 sg13g2_decap_8 FILLER_52_259 ();
 sg13g2_decap_8 FILLER_52_266 ();
 sg13g2_decap_8 FILLER_52_273 ();
 sg13g2_decap_8 FILLER_52_280 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_294 ();
 sg13g2_decap_8 FILLER_52_301 ();
 sg13g2_decap_8 FILLER_52_308 ();
 sg13g2_decap_8 FILLER_52_315 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_8 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_420 ();
 sg13g2_decap_8 FILLER_52_427 ();
 sg13g2_decap_8 FILLER_52_434 ();
 sg13g2_decap_8 FILLER_52_441 ();
 sg13g2_decap_8 FILLER_52_448 ();
 sg13g2_decap_8 FILLER_52_455 ();
 sg13g2_fill_2 FILLER_52_462 ();
 sg13g2_fill_2 FILLER_52_521 ();
 sg13g2_fill_1 FILLER_52_523 ();
 sg13g2_fill_2 FILLER_52_555 ();
 sg13g2_fill_2 FILLER_52_587 ();
 sg13g2_decap_4 FILLER_52_595 ();
 sg13g2_fill_2 FILLER_52_599 ();
 sg13g2_fill_2 FILLER_52_606 ();
 sg13g2_fill_1 FILLER_52_639 ();
 sg13g2_fill_1 FILLER_52_653 ();
 sg13g2_fill_2 FILLER_52_659 ();
 sg13g2_fill_1 FILLER_52_661 ();
 sg13g2_fill_2 FILLER_52_672 ();
 sg13g2_fill_2 FILLER_52_683 ();
 sg13g2_fill_2 FILLER_52_715 ();
 sg13g2_fill_1 FILLER_52_717 ();
 sg13g2_fill_1 FILLER_52_761 ();
 sg13g2_fill_2 FILLER_52_771 ();
 sg13g2_fill_1 FILLER_52_773 ();
 sg13g2_fill_2 FILLER_52_791 ();
 sg13g2_fill_2 FILLER_52_819 ();
 sg13g2_fill_2 FILLER_52_855 ();
 sg13g2_fill_2 FILLER_52_882 ();
 sg13g2_fill_2 FILLER_52_919 ();
 sg13g2_fill_2 FILLER_52_933 ();
 sg13g2_fill_2 FILLER_52_977 ();
 sg13g2_fill_1 FILLER_52_979 ();
 sg13g2_fill_1 FILLER_52_997 ();
 sg13g2_fill_1 FILLER_52_1010 ();
 sg13g2_fill_2 FILLER_52_1026 ();
 sg13g2_fill_1 FILLER_52_1028 ();
 sg13g2_fill_1 FILLER_52_1033 ();
 sg13g2_decap_8 FILLER_52_1040 ();
 sg13g2_decap_8 FILLER_52_1047 ();
 sg13g2_fill_2 FILLER_52_1058 ();
 sg13g2_decap_8 FILLER_52_1086 ();
 sg13g2_fill_2 FILLER_52_1093 ();
 sg13g2_fill_1 FILLER_52_1095 ();
 sg13g2_fill_2 FILLER_52_1106 ();
 sg13g2_fill_1 FILLER_52_1108 ();
 sg13g2_fill_2 FILLER_52_1160 ();
 sg13g2_fill_1 FILLER_52_1172 ();
 sg13g2_fill_2 FILLER_52_1186 ();
 sg13g2_fill_1 FILLER_52_1192 ();
 sg13g2_fill_2 FILLER_52_1215 ();
 sg13g2_fill_1 FILLER_52_1239 ();
 sg13g2_fill_1 FILLER_52_1279 ();
 sg13g2_fill_2 FILLER_52_1285 ();
 sg13g2_fill_1 FILLER_52_1287 ();
 sg13g2_fill_2 FILLER_52_1303 ();
 sg13g2_fill_1 FILLER_52_1305 ();
 sg13g2_decap_8 FILLER_52_1318 ();
 sg13g2_fill_2 FILLER_52_1325 ();
 sg13g2_fill_1 FILLER_52_1337 ();
 sg13g2_decap_4 FILLER_52_1343 ();
 sg13g2_fill_2 FILLER_52_1347 ();
 sg13g2_fill_2 FILLER_52_1406 ();
 sg13g2_decap_8 FILLER_52_1517 ();
 sg13g2_fill_1 FILLER_52_1536 ();
 sg13g2_fill_1 FILLER_52_1546 ();
 sg13g2_fill_2 FILLER_52_1581 ();
 sg13g2_fill_2 FILLER_52_1600 ();
 sg13g2_fill_1 FILLER_52_1611 ();
 sg13g2_fill_1 FILLER_52_1682 ();
 sg13g2_fill_1 FILLER_52_1739 ();
 sg13g2_fill_2 FILLER_52_1762 ();
 sg13g2_fill_2 FILLER_52_1772 ();
 sg13g2_fill_2 FILLER_52_1797 ();
 sg13g2_fill_1 FILLER_52_1806 ();
 sg13g2_fill_2 FILLER_52_1814 ();
 sg13g2_fill_1 FILLER_52_1816 ();
 sg13g2_fill_2 FILLER_52_1822 ();
 sg13g2_fill_1 FILLER_52_1853 ();
 sg13g2_fill_2 FILLER_52_1875 ();
 sg13g2_fill_2 FILLER_52_1900 ();
 sg13g2_fill_2 FILLER_52_1920 ();
 sg13g2_fill_1 FILLER_52_1922 ();
 sg13g2_fill_1 FILLER_52_1941 ();
 sg13g2_fill_1 FILLER_52_1960 ();
 sg13g2_fill_1 FILLER_52_1992 ();
 sg13g2_fill_2 FILLER_52_2028 ();
 sg13g2_fill_2 FILLER_52_2038 ();
 sg13g2_fill_1 FILLER_52_2049 ();
 sg13g2_fill_2 FILLER_52_2128 ();
 sg13g2_decap_4 FILLER_52_2173 ();
 sg13g2_decap_4 FILLER_52_2182 ();
 sg13g2_fill_1 FILLER_52_2186 ();
 sg13g2_decap_4 FILLER_52_2213 ();
 sg13g2_fill_2 FILLER_52_2217 ();
 sg13g2_fill_1 FILLER_52_2250 ();
 sg13g2_fill_2 FILLER_52_2276 ();
 sg13g2_fill_2 FILLER_52_2334 ();
 sg13g2_fill_1 FILLER_52_2336 ();
 sg13g2_decap_4 FILLER_52_2341 ();
 sg13g2_fill_1 FILLER_52_2345 ();
 sg13g2_decap_8 FILLER_52_2350 ();
 sg13g2_fill_1 FILLER_52_2357 ();
 sg13g2_decap_8 FILLER_52_2371 ();
 sg13g2_fill_1 FILLER_52_2378 ();
 sg13g2_decap_8 FILLER_52_2392 ();
 sg13g2_fill_2 FILLER_52_2399 ();
 sg13g2_fill_2 FILLER_52_2409 ();
 sg13g2_fill_2 FILLER_52_2458 ();
 sg13g2_fill_1 FILLER_52_2460 ();
 sg13g2_fill_2 FILLER_52_2487 ();
 sg13g2_fill_1 FILLER_52_2489 ();
 sg13g2_fill_2 FILLER_52_2512 ();
 sg13g2_fill_1 FILLER_52_2514 ();
 sg13g2_fill_1 FILLER_52_2551 ();
 sg13g2_fill_1 FILLER_52_2578 ();
 sg13g2_decap_8 FILLER_52_2614 ();
 sg13g2_decap_8 FILLER_52_2621 ();
 sg13g2_decap_8 FILLER_52_2628 ();
 sg13g2_decap_8 FILLER_52_2635 ();
 sg13g2_decap_8 FILLER_52_2642 ();
 sg13g2_decap_8 FILLER_52_2649 ();
 sg13g2_decap_8 FILLER_52_2656 ();
 sg13g2_decap_8 FILLER_52_2663 ();
 sg13g2_decap_4 FILLER_52_2670 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_decap_8 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_231 ();
 sg13g2_decap_8 FILLER_53_238 ();
 sg13g2_decap_8 FILLER_53_245 ();
 sg13g2_decap_8 FILLER_53_252 ();
 sg13g2_decap_8 FILLER_53_259 ();
 sg13g2_decap_8 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_decap_8 FILLER_53_280 ();
 sg13g2_decap_8 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_301 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_decap_8 FILLER_53_315 ();
 sg13g2_decap_8 FILLER_53_322 ();
 sg13g2_decap_8 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_336 ();
 sg13g2_decap_8 FILLER_53_343 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_383 ();
 sg13g2_decap_8 FILLER_53_415 ();
 sg13g2_decap_8 FILLER_53_422 ();
 sg13g2_decap_8 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_53_436 ();
 sg13g2_decap_8 FILLER_53_443 ();
 sg13g2_decap_8 FILLER_53_450 ();
 sg13g2_decap_8 FILLER_53_457 ();
 sg13g2_decap_8 FILLER_53_464 ();
 sg13g2_decap_4 FILLER_53_471 ();
 sg13g2_fill_1 FILLER_53_475 ();
 sg13g2_fill_2 FILLER_53_527 ();
 sg13g2_fill_1 FILLER_53_529 ();
 sg13g2_fill_2 FILLER_53_539 ();
 sg13g2_fill_1 FILLER_53_559 ();
 sg13g2_decap_8 FILLER_53_590 ();
 sg13g2_fill_2 FILLER_53_597 ();
 sg13g2_fill_1 FILLER_53_599 ();
 sg13g2_fill_1 FILLER_53_688 ();
 sg13g2_fill_1 FILLER_53_713 ();
 sg13g2_fill_2 FILLER_53_745 ();
 sg13g2_fill_1 FILLER_53_747 ();
 sg13g2_fill_1 FILLER_53_795 ();
 sg13g2_fill_1 FILLER_53_818 ();
 sg13g2_fill_2 FILLER_53_827 ();
 sg13g2_fill_2 FILLER_53_886 ();
 sg13g2_fill_1 FILLER_53_897 ();
 sg13g2_fill_2 FILLER_53_915 ();
 sg13g2_fill_1 FILLER_53_917 ();
 sg13g2_fill_1 FILLER_53_981 ();
 sg13g2_fill_2 FILLER_53_986 ();
 sg13g2_fill_1 FILLER_53_988 ();
 sg13g2_fill_1 FILLER_53_1043 ();
 sg13g2_fill_1 FILLER_53_1070 ();
 sg13g2_fill_1 FILLER_53_1131 ();
 sg13g2_fill_1 FILLER_53_1168 ();
 sg13g2_fill_1 FILLER_53_1241 ();
 sg13g2_fill_1 FILLER_53_1259 ();
 sg13g2_fill_2 FILLER_53_1273 ();
 sg13g2_fill_1 FILLER_53_1275 ();
 sg13g2_fill_2 FILLER_53_1284 ();
 sg13g2_fill_1 FILLER_53_1312 ();
 sg13g2_decap_4 FILLER_53_1320 ();
 sg13g2_fill_2 FILLER_53_1324 ();
 sg13g2_decap_8 FILLER_53_1330 ();
 sg13g2_decap_4 FILLER_53_1337 ();
 sg13g2_fill_1 FILLER_53_1344 ();
 sg13g2_fill_1 FILLER_53_1365 ();
 sg13g2_fill_2 FILLER_53_1373 ();
 sg13g2_fill_2 FILLER_53_1397 ();
 sg13g2_fill_1 FILLER_53_1399 ();
 sg13g2_fill_2 FILLER_53_1435 ();
 sg13g2_fill_1 FILLER_53_1437 ();
 sg13g2_fill_2 FILLER_53_1474 ();
 sg13g2_fill_1 FILLER_53_1476 ();
 sg13g2_decap_8 FILLER_53_1508 ();
 sg13g2_fill_1 FILLER_53_1515 ();
 sg13g2_decap_4 FILLER_53_1521 ();
 sg13g2_fill_1 FILLER_53_1563 ();
 sg13g2_fill_2 FILLER_53_1593 ();
 sg13g2_fill_2 FILLER_53_1689 ();
 sg13g2_fill_1 FILLER_53_1691 ();
 sg13g2_fill_1 FILLER_53_1767 ();
 sg13g2_fill_2 FILLER_53_1834 ();
 sg13g2_fill_1 FILLER_53_1836 ();
 sg13g2_fill_2 FILLER_53_1852 ();
 sg13g2_fill_1 FILLER_53_1880 ();
 sg13g2_fill_1 FILLER_53_1921 ();
 sg13g2_fill_2 FILLER_53_1962 ();
 sg13g2_fill_1 FILLER_53_1964 ();
 sg13g2_fill_2 FILLER_53_1991 ();
 sg13g2_fill_2 FILLER_53_2060 ();
 sg13g2_fill_2 FILLER_53_2123 ();
 sg13g2_fill_2 FILLER_53_2181 ();
 sg13g2_fill_1 FILLER_53_2183 ();
 sg13g2_decap_8 FILLER_53_2214 ();
 sg13g2_fill_1 FILLER_53_2221 ();
 sg13g2_fill_2 FILLER_53_2266 ();
 sg13g2_fill_1 FILLER_53_2278 ();
 sg13g2_fill_2 FILLER_53_2324 ();
 sg13g2_decap_8 FILLER_53_2366 ();
 sg13g2_fill_2 FILLER_53_2470 ();
 sg13g2_fill_2 FILLER_53_2547 ();
 sg13g2_fill_1 FILLER_53_2549 ();
 sg13g2_decap_8 FILLER_53_2624 ();
 sg13g2_decap_8 FILLER_53_2631 ();
 sg13g2_decap_8 FILLER_53_2638 ();
 sg13g2_decap_8 FILLER_53_2645 ();
 sg13g2_decap_8 FILLER_53_2652 ();
 sg13g2_decap_8 FILLER_53_2659 ();
 sg13g2_decap_8 FILLER_53_2666 ();
 sg13g2_fill_1 FILLER_53_2673 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_decap_8 FILLER_54_189 ();
 sg13g2_decap_8 FILLER_54_196 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_decap_8 FILLER_54_210 ();
 sg13g2_decap_8 FILLER_54_217 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_decap_8 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_238 ();
 sg13g2_decap_8 FILLER_54_245 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_259 ();
 sg13g2_decap_8 FILLER_54_266 ();
 sg13g2_decap_8 FILLER_54_273 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_decap_8 FILLER_54_287 ();
 sg13g2_decap_8 FILLER_54_294 ();
 sg13g2_decap_8 FILLER_54_301 ();
 sg13g2_decap_8 FILLER_54_308 ();
 sg13g2_decap_8 FILLER_54_315 ();
 sg13g2_decap_8 FILLER_54_322 ();
 sg13g2_decap_8 FILLER_54_329 ();
 sg13g2_decap_8 FILLER_54_336 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_fill_1 FILLER_54_350 ();
 sg13g2_decap_4 FILLER_54_384 ();
 sg13g2_fill_1 FILLER_54_388 ();
 sg13g2_decap_8 FILLER_54_425 ();
 sg13g2_decap_8 FILLER_54_432 ();
 sg13g2_decap_8 FILLER_54_439 ();
 sg13g2_decap_8 FILLER_54_446 ();
 sg13g2_decap_8 FILLER_54_453 ();
 sg13g2_decap_8 FILLER_54_460 ();
 sg13g2_decap_8 FILLER_54_467 ();
 sg13g2_decap_4 FILLER_54_474 ();
 sg13g2_fill_2 FILLER_54_478 ();
 sg13g2_fill_1 FILLER_54_492 ();
 sg13g2_decap_8 FILLER_54_502 ();
 sg13g2_decap_8 FILLER_54_509 ();
 sg13g2_decap_8 FILLER_54_516 ();
 sg13g2_fill_2 FILLER_54_528 ();
 sg13g2_fill_2 FILLER_54_535 ();
 sg13g2_fill_1 FILLER_54_537 ();
 sg13g2_fill_2 FILLER_54_718 ();
 sg13g2_fill_2 FILLER_54_755 ();
 sg13g2_fill_1 FILLER_54_757 ();
 sg13g2_fill_2 FILLER_54_796 ();
 sg13g2_fill_1 FILLER_54_798 ();
 sg13g2_fill_2 FILLER_54_804 ();
 sg13g2_fill_1 FILLER_54_811 ();
 sg13g2_fill_2 FILLER_54_820 ();
 sg13g2_fill_1 FILLER_54_822 ();
 sg13g2_fill_2 FILLER_54_876 ();
 sg13g2_fill_2 FILLER_54_887 ();
 sg13g2_fill_2 FILLER_54_894 ();
 sg13g2_fill_1 FILLER_54_896 ();
 sg13g2_fill_2 FILLER_54_1014 ();
 sg13g2_fill_2 FILLER_54_1032 ();
 sg13g2_fill_2 FILLER_54_1037 ();
 sg13g2_fill_1 FILLER_54_1047 ();
 sg13g2_fill_2 FILLER_54_1072 ();
 sg13g2_fill_1 FILLER_54_1100 ();
 sg13g2_fill_1 FILLER_54_1109 ();
 sg13g2_fill_2 FILLER_54_1123 ();
 sg13g2_decap_4 FILLER_54_1148 ();
 sg13g2_fill_1 FILLER_54_1178 ();
 sg13g2_fill_2 FILLER_54_1219 ();
 sg13g2_fill_2 FILLER_54_1243 ();
 sg13g2_fill_1 FILLER_54_1248 ();
 sg13g2_fill_2 FILLER_54_1268 ();
 sg13g2_fill_1 FILLER_54_1270 ();
 sg13g2_fill_1 FILLER_54_1340 ();
 sg13g2_fill_1 FILLER_54_1357 ();
 sg13g2_fill_1 FILLER_54_1371 ();
 sg13g2_fill_1 FILLER_54_1387 ();
 sg13g2_fill_1 FILLER_54_1392 ();
 sg13g2_fill_2 FILLER_54_1445 ();
 sg13g2_fill_1 FILLER_54_1447 ();
 sg13g2_fill_2 FILLER_54_1477 ();
 sg13g2_fill_1 FILLER_54_1479 ();
 sg13g2_fill_2 FILLER_54_1485 ();
 sg13g2_fill_2 FILLER_54_1505 ();
 sg13g2_decap_4 FILLER_54_1516 ();
 sg13g2_fill_2 FILLER_54_1534 ();
 sg13g2_fill_1 FILLER_54_1536 ();
 sg13g2_fill_2 FILLER_54_1577 ();
 sg13g2_fill_1 FILLER_54_1618 ();
 sg13g2_fill_2 FILLER_54_1636 ();
 sg13g2_fill_2 FILLER_54_1697 ();
 sg13g2_fill_2 FILLER_54_1739 ();
 sg13g2_fill_2 FILLER_54_1762 ();
 sg13g2_fill_1 FILLER_54_1764 ();
 sg13g2_decap_4 FILLER_54_1794 ();
 sg13g2_fill_2 FILLER_54_1798 ();
 sg13g2_fill_2 FILLER_54_1809 ();
 sg13g2_fill_1 FILLER_54_1837 ();
 sg13g2_fill_2 FILLER_54_1908 ();
 sg13g2_fill_1 FILLER_54_1970 ();
 sg13g2_fill_1 FILLER_54_1980 ();
 sg13g2_fill_2 FILLER_54_2005 ();
 sg13g2_fill_1 FILLER_54_2007 ();
 sg13g2_fill_2 FILLER_54_2026 ();
 sg13g2_fill_1 FILLER_54_2038 ();
 sg13g2_fill_2 FILLER_54_2138 ();
 sg13g2_fill_2 FILLER_54_2184 ();
 sg13g2_fill_2 FILLER_54_2246 ();
 sg13g2_fill_1 FILLER_54_2268 ();
 sg13g2_fill_1 FILLER_54_2283 ();
 sg13g2_fill_2 FILLER_54_2289 ();
 sg13g2_fill_1 FILLER_54_2291 ();
 sg13g2_fill_1 FILLER_54_2297 ();
 sg13g2_fill_1 FILLER_54_2310 ();
 sg13g2_fill_2 FILLER_54_2320 ();
 sg13g2_fill_1 FILLER_54_2414 ();
 sg13g2_fill_1 FILLER_54_2450 ();
 sg13g2_fill_1 FILLER_54_2462 ();
 sg13g2_fill_2 FILLER_54_2515 ();
 sg13g2_fill_1 FILLER_54_2517 ();
 sg13g2_fill_1 FILLER_54_2553 ();
 sg13g2_decap_8 FILLER_54_2627 ();
 sg13g2_decap_8 FILLER_54_2634 ();
 sg13g2_decap_8 FILLER_54_2641 ();
 sg13g2_decap_8 FILLER_54_2648 ();
 sg13g2_decap_8 FILLER_54_2655 ();
 sg13g2_decap_8 FILLER_54_2662 ();
 sg13g2_decap_4 FILLER_54_2669 ();
 sg13g2_fill_1 FILLER_54_2673 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_189 ();
 sg13g2_decap_8 FILLER_55_196 ();
 sg13g2_decap_8 FILLER_55_203 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_224 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_decap_8 FILLER_55_238 ();
 sg13g2_decap_8 FILLER_55_245 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_decap_8 FILLER_55_294 ();
 sg13g2_decap_8 FILLER_55_301 ();
 sg13g2_decap_8 FILLER_55_308 ();
 sg13g2_decap_8 FILLER_55_315 ();
 sg13g2_decap_8 FILLER_55_322 ();
 sg13g2_decap_8 FILLER_55_329 ();
 sg13g2_decap_4 FILLER_55_336 ();
 sg13g2_fill_2 FILLER_55_340 ();
 sg13g2_fill_2 FILLER_55_456 ();
 sg13g2_fill_1 FILLER_55_458 ();
 sg13g2_decap_8 FILLER_55_464 ();
 sg13g2_decap_8 FILLER_55_471 ();
 sg13g2_decap_8 FILLER_55_478 ();
 sg13g2_fill_2 FILLER_55_485 ();
 sg13g2_decap_4 FILLER_55_492 ();
 sg13g2_fill_2 FILLER_55_496 ();
 sg13g2_fill_2 FILLER_55_550 ();
 sg13g2_fill_1 FILLER_55_552 ();
 sg13g2_fill_2 FILLER_55_589 ();
 sg13g2_fill_2 FILLER_55_630 ();
 sg13g2_fill_1 FILLER_55_632 ();
 sg13g2_fill_1 FILLER_55_672 ();
 sg13g2_fill_1 FILLER_55_679 ();
 sg13g2_decap_4 FILLER_55_714 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_fill_2 FILLER_55_785 ();
 sg13g2_fill_1 FILLER_55_787 ();
 sg13g2_fill_2 FILLER_55_832 ();
 sg13g2_fill_2 FILLER_55_870 ();
 sg13g2_fill_1 FILLER_55_872 ();
 sg13g2_fill_2 FILLER_55_912 ();
 sg13g2_fill_1 FILLER_55_914 ();
 sg13g2_fill_2 FILLER_55_928 ();
 sg13g2_fill_2 FILLER_55_952 ();
 sg13g2_fill_2 FILLER_55_962 ();
 sg13g2_fill_1 FILLER_55_999 ();
 sg13g2_fill_1 FILLER_55_1009 ();
 sg13g2_fill_2 FILLER_55_1042 ();
 sg13g2_fill_2 FILLER_55_1074 ();
 sg13g2_fill_1 FILLER_55_1076 ();
 sg13g2_decap_8 FILLER_55_1115 ();
 sg13g2_fill_1 FILLER_55_1122 ();
 sg13g2_decap_8 FILLER_55_1127 ();
 sg13g2_decap_8 FILLER_55_1134 ();
 sg13g2_decap_4 FILLER_55_1141 ();
 sg13g2_fill_2 FILLER_55_1145 ();
 sg13g2_fill_2 FILLER_55_1230 ();
 sg13g2_fill_2 FILLER_55_1283 ();
 sg13g2_fill_1 FILLER_55_1285 ();
 sg13g2_decap_4 FILLER_55_1362 ();
 sg13g2_fill_2 FILLER_55_1405 ();
 sg13g2_fill_2 FILLER_55_1436 ();
 sg13g2_fill_1 FILLER_55_1438 ();
 sg13g2_fill_2 FILLER_55_1466 ();
 sg13g2_fill_1 FILLER_55_1468 ();
 sg13g2_fill_2 FILLER_55_1511 ();
 sg13g2_fill_2 FILLER_55_1523 ();
 sg13g2_fill_1 FILLER_55_1533 ();
 sg13g2_fill_1 FILLER_55_1539 ();
 sg13g2_fill_2 FILLER_55_1561 ();
 sg13g2_fill_2 FILLER_55_1577 ();
 sg13g2_fill_1 FILLER_55_1579 ();
 sg13g2_fill_1 FILLER_55_1629 ();
 sg13g2_fill_2 FILLER_55_1635 ();
 sg13g2_fill_1 FILLER_55_1637 ();
 sg13g2_fill_2 FILLER_55_1642 ();
 sg13g2_fill_1 FILLER_55_1644 ();
 sg13g2_fill_2 FILLER_55_1659 ();
 sg13g2_fill_1 FILLER_55_1661 ();
 sg13g2_fill_2 FILLER_55_1692 ();
 sg13g2_fill_1 FILLER_55_1694 ();
 sg13g2_fill_2 FILLER_55_1699 ();
 sg13g2_fill_1 FILLER_55_1701 ();
 sg13g2_fill_2 FILLER_55_1733 ();
 sg13g2_fill_1 FILLER_55_1735 ();
 sg13g2_fill_2 FILLER_55_1749 ();
 sg13g2_fill_1 FILLER_55_1751 ();
 sg13g2_fill_2 FILLER_55_1764 ();
 sg13g2_fill_1 FILLER_55_1766 ();
 sg13g2_fill_2 FILLER_55_1809 ();
 sg13g2_fill_1 FILLER_55_1811 ();
 sg13g2_fill_2 FILLER_55_1868 ();
 sg13g2_fill_2 FILLER_55_1890 ();
 sg13g2_fill_1 FILLER_55_1892 ();
 sg13g2_fill_2 FILLER_55_1910 ();
 sg13g2_fill_2 FILLER_55_1963 ();
 sg13g2_fill_2 FILLER_55_1970 ();
 sg13g2_fill_1 FILLER_55_1972 ();
 sg13g2_fill_2 FILLER_55_1978 ();
 sg13g2_fill_1 FILLER_55_1989 ();
 sg13g2_fill_2 FILLER_55_2012 ();
 sg13g2_fill_1 FILLER_55_2044 ();
 sg13g2_fill_2 FILLER_55_2054 ();
 sg13g2_fill_1 FILLER_55_2056 ();
 sg13g2_fill_2 FILLER_55_2078 ();
 sg13g2_fill_1 FILLER_55_2080 ();
 sg13g2_fill_1 FILLER_55_2087 ();
 sg13g2_fill_1 FILLER_55_2100 ();
 sg13g2_fill_2 FILLER_55_2129 ();
 sg13g2_fill_2 FILLER_55_2187 ();
 sg13g2_fill_1 FILLER_55_2189 ();
 sg13g2_fill_2 FILLER_55_2195 ();
 sg13g2_fill_2 FILLER_55_2206 ();
 sg13g2_decap_8 FILLER_55_2238 ();
 sg13g2_decap_8 FILLER_55_2245 ();
 sg13g2_decap_4 FILLER_55_2252 ();
 sg13g2_fill_1 FILLER_55_2256 ();
 sg13g2_fill_2 FILLER_55_2262 ();
 sg13g2_fill_2 FILLER_55_2300 ();
 sg13g2_fill_1 FILLER_55_2302 ();
 sg13g2_fill_1 FILLER_55_2308 ();
 sg13g2_fill_1 FILLER_55_2335 ();
 sg13g2_fill_2 FILLER_55_2371 ();
 sg13g2_fill_1 FILLER_55_2425 ();
 sg13g2_fill_2 FILLER_55_2451 ();
 sg13g2_fill_1 FILLER_55_2453 ();
 sg13g2_decap_8 FILLER_55_2466 ();
 sg13g2_fill_2 FILLER_55_2495 ();
 sg13g2_fill_1 FILLER_55_2497 ();
 sg13g2_fill_2 FILLER_55_2558 ();
 sg13g2_decap_8 FILLER_55_2630 ();
 sg13g2_decap_8 FILLER_55_2637 ();
 sg13g2_decap_8 FILLER_55_2644 ();
 sg13g2_decap_8 FILLER_55_2651 ();
 sg13g2_decap_8 FILLER_55_2658 ();
 sg13g2_decap_8 FILLER_55_2665 ();
 sg13g2_fill_2 FILLER_55_2672 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_182 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_decap_8 FILLER_56_196 ();
 sg13g2_decap_8 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_decap_8 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_decap_8 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_252 ();
 sg13g2_decap_8 FILLER_56_259 ();
 sg13g2_decap_8 FILLER_56_266 ();
 sg13g2_decap_8 FILLER_56_273 ();
 sg13g2_decap_8 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_287 ();
 sg13g2_decap_8 FILLER_56_294 ();
 sg13g2_decap_8 FILLER_56_301 ();
 sg13g2_decap_8 FILLER_56_308 ();
 sg13g2_decap_8 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_322 ();
 sg13g2_decap_8 FILLER_56_329 ();
 sg13g2_decap_4 FILLER_56_336 ();
 sg13g2_fill_2 FILLER_56_340 ();
 sg13g2_decap_8 FILLER_56_388 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_462 ();
 sg13g2_fill_1 FILLER_56_469 ();
 sg13g2_decap_8 FILLER_56_477 ();
 sg13g2_decap_8 FILLER_56_489 ();
 sg13g2_decap_8 FILLER_56_496 ();
 sg13g2_fill_1 FILLER_56_503 ();
 sg13g2_decap_8 FILLER_56_517 ();
 sg13g2_decap_8 FILLER_56_524 ();
 sg13g2_fill_2 FILLER_56_531 ();
 sg13g2_fill_1 FILLER_56_533 ();
 sg13g2_fill_2 FILLER_56_546 ();
 sg13g2_decap_8 FILLER_56_590 ();
 sg13g2_fill_2 FILLER_56_597 ();
 sg13g2_fill_1 FILLER_56_599 ();
 sg13g2_fill_1 FILLER_56_617 ();
 sg13g2_fill_2 FILLER_56_623 ();
 sg13g2_fill_1 FILLER_56_625 ();
 sg13g2_fill_1 FILLER_56_647 ();
 sg13g2_decap_8 FILLER_56_714 ();
 sg13g2_decap_4 FILLER_56_721 ();
 sg13g2_fill_2 FILLER_56_725 ();
 sg13g2_fill_2 FILLER_56_732 ();
 sg13g2_fill_1 FILLER_56_734 ();
 sg13g2_fill_2 FILLER_56_748 ();
 sg13g2_fill_1 FILLER_56_750 ();
 sg13g2_fill_2 FILLER_56_786 ();
 sg13g2_fill_2 FILLER_56_792 ();
 sg13g2_fill_2 FILLER_56_824 ();
 sg13g2_fill_2 FILLER_56_838 ();
 sg13g2_fill_1 FILLER_56_840 ();
 sg13g2_fill_1 FILLER_56_863 ();
 sg13g2_fill_1 FILLER_56_1034 ();
 sg13g2_fill_1 FILLER_56_1078 ();
 sg13g2_decap_4 FILLER_56_1118 ();
 sg13g2_fill_1 FILLER_56_1122 ();
 sg13g2_fill_2 FILLER_56_1137 ();
 sg13g2_fill_1 FILLER_56_1139 ();
 sg13g2_fill_2 FILLER_56_1150 ();
 sg13g2_fill_2 FILLER_56_1160 ();
 sg13g2_fill_1 FILLER_56_1166 ();
 sg13g2_fill_1 FILLER_56_1194 ();
 sg13g2_fill_2 FILLER_56_1241 ();
 sg13g2_fill_1 FILLER_56_1243 ();
 sg13g2_fill_1 FILLER_56_1270 ();
 sg13g2_decap_8 FILLER_56_1276 ();
 sg13g2_fill_2 FILLER_56_1283 ();
 sg13g2_decap_8 FILLER_56_1289 ();
 sg13g2_decap_8 FILLER_56_1296 ();
 sg13g2_fill_1 FILLER_56_1303 ();
 sg13g2_fill_1 FILLER_56_1327 ();
 sg13g2_decap_4 FILLER_56_1353 ();
 sg13g2_fill_1 FILLER_56_1357 ();
 sg13g2_decap_4 FILLER_56_1366 ();
 sg13g2_fill_1 FILLER_56_1378 ();
 sg13g2_decap_8 FILLER_56_1387 ();
 sg13g2_fill_2 FILLER_56_1394 ();
 sg13g2_fill_1 FILLER_56_1396 ();
 sg13g2_fill_2 FILLER_56_1409 ();
 sg13g2_fill_1 FILLER_56_1411 ();
 sg13g2_decap_4 FILLER_56_1424 ();
 sg13g2_fill_1 FILLER_56_1428 ();
 sg13g2_decap_8 FILLER_56_1433 ();
 sg13g2_decap_4 FILLER_56_1440 ();
 sg13g2_fill_2 FILLER_56_1531 ();
 sg13g2_decap_4 FILLER_56_1571 ();
 sg13g2_fill_1 FILLER_56_1575 ();
 sg13g2_fill_1 FILLER_56_1580 ();
 sg13g2_fill_2 FILLER_56_1622 ();
 sg13g2_fill_1 FILLER_56_1624 ();
 sg13g2_decap_8 FILLER_56_1709 ();
 sg13g2_fill_2 FILLER_56_1716 ();
 sg13g2_decap_4 FILLER_56_1787 ();
 sg13g2_decap_4 FILLER_56_1794 ();
 sg13g2_fill_2 FILLER_56_1798 ();
 sg13g2_fill_1 FILLER_56_1820 ();
 sg13g2_fill_2 FILLER_56_1918 ();
 sg13g2_fill_1 FILLER_56_1928 ();
 sg13g2_fill_1 FILLER_56_1956 ();
 sg13g2_fill_2 FILLER_56_2004 ();
 sg13g2_decap_8 FILLER_56_2036 ();
 sg13g2_decap_8 FILLER_56_2043 ();
 sg13g2_decap_8 FILLER_56_2054 ();
 sg13g2_decap_8 FILLER_56_2070 ();
 sg13g2_decap_8 FILLER_56_2077 ();
 sg13g2_fill_2 FILLER_56_2084 ();
 sg13g2_fill_1 FILLER_56_2086 ();
 sg13g2_fill_2 FILLER_56_2113 ();
 sg13g2_fill_1 FILLER_56_2115 ();
 sg13g2_fill_1 FILLER_56_2129 ();
 sg13g2_fill_2 FILLER_56_2153 ();
 sg13g2_fill_1 FILLER_56_2155 ();
 sg13g2_fill_2 FILLER_56_2182 ();
 sg13g2_fill_1 FILLER_56_2184 ();
 sg13g2_fill_1 FILLER_56_2194 ();
 sg13g2_fill_2 FILLER_56_2204 ();
 sg13g2_fill_1 FILLER_56_2234 ();
 sg13g2_fill_1 FILLER_56_2274 ();
 sg13g2_fill_2 FILLER_56_2322 ();
 sg13g2_fill_1 FILLER_56_2324 ();
 sg13g2_fill_2 FILLER_56_2355 ();
 sg13g2_decap_4 FILLER_56_2374 ();
 sg13g2_fill_1 FILLER_56_2378 ();
 sg13g2_fill_2 FILLER_56_2388 ();
 sg13g2_fill_1 FILLER_56_2390 ();
 sg13g2_fill_1 FILLER_56_2410 ();
 sg13g2_fill_1 FILLER_56_2450 ();
 sg13g2_fill_1 FILLER_56_2456 ();
 sg13g2_fill_1 FILLER_56_2481 ();
 sg13g2_fill_2 FILLER_56_2487 ();
 sg13g2_fill_1 FILLER_56_2489 ();
 sg13g2_fill_2 FILLER_56_2512 ();
 sg13g2_fill_1 FILLER_56_2545 ();
 sg13g2_decap_8 FILLER_56_2632 ();
 sg13g2_decap_8 FILLER_56_2639 ();
 sg13g2_decap_8 FILLER_56_2646 ();
 sg13g2_decap_8 FILLER_56_2653 ();
 sg13g2_decap_8 FILLER_56_2660 ();
 sg13g2_decap_8 FILLER_56_2667 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_238 ();
 sg13g2_decap_8 FILLER_57_245 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_8 FILLER_57_259 ();
 sg13g2_decap_8 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_decap_8 FILLER_57_294 ();
 sg13g2_decap_8 FILLER_57_301 ();
 sg13g2_decap_8 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_8 FILLER_57_329 ();
 sg13g2_decap_8 FILLER_57_336 ();
 sg13g2_decap_8 FILLER_57_343 ();
 sg13g2_decap_4 FILLER_57_350 ();
 sg13g2_fill_1 FILLER_57_370 ();
 sg13g2_decap_8 FILLER_57_383 ();
 sg13g2_fill_2 FILLER_57_390 ();
 sg13g2_fill_1 FILLER_57_418 ();
 sg13g2_decap_8 FILLER_57_439 ();
 sg13g2_fill_2 FILLER_57_454 ();
 sg13g2_fill_1 FILLER_57_456 ();
 sg13g2_decap_4 FILLER_57_519 ();
 sg13g2_decap_8 FILLER_57_528 ();
 sg13g2_decap_8 FILLER_57_535 ();
 sg13g2_fill_2 FILLER_57_542 ();
 sg13g2_fill_1 FILLER_57_544 ();
 sg13g2_fill_2 FILLER_57_553 ();
 sg13g2_fill_1 FILLER_57_555 ();
 sg13g2_decap_8 FILLER_57_586 ();
 sg13g2_decap_8 FILLER_57_593 ();
 sg13g2_decap_8 FILLER_57_600 ();
 sg13g2_decap_4 FILLER_57_607 ();
 sg13g2_decap_4 FILLER_57_619 ();
 sg13g2_fill_2 FILLER_57_631 ();
 sg13g2_fill_1 FILLER_57_633 ();
 sg13g2_fill_2 FILLER_57_642 ();
 sg13g2_fill_1 FILLER_57_644 ();
 sg13g2_fill_2 FILLER_57_657 ();
 sg13g2_fill_1 FILLER_57_659 ();
 sg13g2_fill_2 FILLER_57_673 ();
 sg13g2_fill_1 FILLER_57_675 ();
 sg13g2_decap_8 FILLER_57_684 ();
 sg13g2_fill_1 FILLER_57_691 ();
 sg13g2_decap_8 FILLER_57_696 ();
 sg13g2_fill_1 FILLER_57_703 ();
 sg13g2_decap_8 FILLER_57_712 ();
 sg13g2_fill_2 FILLER_57_719 ();
 sg13g2_fill_2 FILLER_57_821 ();
 sg13g2_fill_1 FILLER_57_876 ();
 sg13g2_fill_2 FILLER_57_907 ();
 sg13g2_fill_1 FILLER_57_909 ();
 sg13g2_fill_1 FILLER_57_999 ();
 sg13g2_fill_1 FILLER_57_1012 ();
 sg13g2_fill_1 FILLER_57_1023 ();
 sg13g2_fill_1 FILLER_57_1041 ();
 sg13g2_fill_1 FILLER_57_1051 ();
 sg13g2_fill_2 FILLER_57_1111 ();
 sg13g2_fill_1 FILLER_57_1113 ();
 sg13g2_fill_2 FILLER_57_1149 ();
 sg13g2_fill_1 FILLER_57_1186 ();
 sg13g2_fill_2 FILLER_57_1197 ();
 sg13g2_fill_1 FILLER_57_1199 ();
 sg13g2_fill_1 FILLER_57_1210 ();
 sg13g2_fill_1 FILLER_57_1249 ();
 sg13g2_fill_1 FILLER_57_1279 ();
 sg13g2_decap_8 FILLER_57_1290 ();
 sg13g2_decap_8 FILLER_57_1297 ();
 sg13g2_decap_4 FILLER_57_1304 ();
 sg13g2_fill_2 FILLER_57_1313 ();
 sg13g2_fill_1 FILLER_57_1315 ();
 sg13g2_decap_8 FILLER_57_1322 ();
 sg13g2_decap_4 FILLER_57_1329 ();
 sg13g2_fill_1 FILLER_57_1333 ();
 sg13g2_fill_1 FILLER_57_1347 ();
 sg13g2_fill_1 FILLER_57_1352 ();
 sg13g2_decap_8 FILLER_57_1358 ();
 sg13g2_decap_4 FILLER_57_1365 ();
 sg13g2_decap_4 FILLER_57_1382 ();
 sg13g2_fill_1 FILLER_57_1386 ();
 sg13g2_decap_8 FILLER_57_1392 ();
 sg13g2_decap_4 FILLER_57_1399 ();
 sg13g2_fill_2 FILLER_57_1403 ();
 sg13g2_fill_2 FILLER_57_1440 ();
 sg13g2_fill_1 FILLER_57_1472 ();
 sg13g2_decap_4 FILLER_57_1575 ();
 sg13g2_fill_1 FILLER_57_1579 ();
 sg13g2_fill_1 FILLER_57_1588 ();
 sg13g2_fill_1 FILLER_57_1597 ();
 sg13g2_fill_2 FILLER_57_1624 ();
 sg13g2_decap_4 FILLER_57_1630 ();
 sg13g2_fill_2 FILLER_57_1634 ();
 sg13g2_decap_8 FILLER_57_1640 ();
 sg13g2_fill_2 FILLER_57_1647 ();
 sg13g2_fill_1 FILLER_57_1649 ();
 sg13g2_fill_2 FILLER_57_1662 ();
 sg13g2_fill_1 FILLER_57_1664 ();
 sg13g2_fill_1 FILLER_57_1691 ();
 sg13g2_fill_2 FILLER_57_1703 ();
 sg13g2_fill_2 FILLER_57_1717 ();
 sg13g2_fill_1 FILLER_57_1719 ();
 sg13g2_fill_2 FILLER_57_1746 ();
 sg13g2_decap_8 FILLER_57_1791 ();
 sg13g2_fill_2 FILLER_57_1798 ();
 sg13g2_decap_4 FILLER_57_1821 ();
 sg13g2_fill_1 FILLER_57_1825 ();
 sg13g2_fill_2 FILLER_57_1852 ();
 sg13g2_fill_1 FILLER_57_1858 ();
 sg13g2_decap_4 FILLER_57_1906 ();
 sg13g2_fill_2 FILLER_57_1919 ();
 sg13g2_fill_1 FILLER_57_1921 ();
 sg13g2_fill_1 FILLER_57_1963 ();
 sg13g2_fill_2 FILLER_57_1999 ();
 sg13g2_fill_1 FILLER_57_2001 ();
 sg13g2_decap_8 FILLER_57_2028 ();
 sg13g2_fill_1 FILLER_57_2035 ();
 sg13g2_decap_4 FILLER_57_2040 ();
 sg13g2_fill_1 FILLER_57_2044 ();
 sg13g2_fill_2 FILLER_57_2066 ();
 sg13g2_fill_1 FILLER_57_2068 ();
 sg13g2_decap_4 FILLER_57_2082 ();
 sg13g2_fill_2 FILLER_57_2148 ();
 sg13g2_fill_1 FILLER_57_2210 ();
 sg13g2_fill_2 FILLER_57_2241 ();
 sg13g2_fill_2 FILLER_57_2262 ();
 sg13g2_fill_1 FILLER_57_2322 ();
 sg13g2_decap_8 FILLER_57_2361 ();
 sg13g2_decap_8 FILLER_57_2368 ();
 sg13g2_decap_8 FILLER_57_2375 ();
 sg13g2_fill_2 FILLER_57_2382 ();
 sg13g2_fill_1 FILLER_57_2384 ();
 sg13g2_fill_1 FILLER_57_2393 ();
 sg13g2_fill_2 FILLER_57_2457 ();
 sg13g2_fill_1 FILLER_57_2472 ();
 sg13g2_fill_1 FILLER_57_2482 ();
 sg13g2_fill_1 FILLER_57_2488 ();
 sg13g2_fill_1 FILLER_57_2494 ();
 sg13g2_fill_2 FILLER_57_2504 ();
 sg13g2_fill_1 FILLER_57_2506 ();
 sg13g2_fill_2 FILLER_57_2516 ();
 sg13g2_fill_1 FILLER_57_2518 ();
 sg13g2_fill_1 FILLER_57_2609 ();
 sg13g2_decap_8 FILLER_57_2627 ();
 sg13g2_decap_8 FILLER_57_2634 ();
 sg13g2_decap_8 FILLER_57_2641 ();
 sg13g2_decap_8 FILLER_57_2648 ();
 sg13g2_decap_8 FILLER_57_2655 ();
 sg13g2_decap_8 FILLER_57_2662 ();
 sg13g2_decap_4 FILLER_57_2669 ();
 sg13g2_fill_1 FILLER_57_2673 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_decap_8 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_224 ();
 sg13g2_decap_8 FILLER_58_231 ();
 sg13g2_decap_8 FILLER_58_238 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_decap_8 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_266 ();
 sg13g2_decap_8 FILLER_58_273 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_308 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_decap_8 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_343 ();
 sg13g2_decap_4 FILLER_58_350 ();
 sg13g2_fill_2 FILLER_58_354 ();
 sg13g2_decap_8 FILLER_58_379 ();
 sg13g2_fill_2 FILLER_58_386 ();
 sg13g2_fill_1 FILLER_58_388 ();
 sg13g2_decap_4 FILLER_58_415 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_2 FILLER_58_438 ();
 sg13g2_fill_1 FILLER_58_440 ();
 sg13g2_fill_1 FILLER_58_486 ();
 sg13g2_decap_4 FILLER_58_518 ();
 sg13g2_decap_8 FILLER_58_548 ();
 sg13g2_decap_8 FILLER_58_555 ();
 sg13g2_fill_2 FILLER_58_562 ();
 sg13g2_decap_8 FILLER_58_569 ();
 sg13g2_decap_8 FILLER_58_576 ();
 sg13g2_fill_2 FILLER_58_583 ();
 sg13g2_decap_8 FILLER_58_589 ();
 sg13g2_fill_2 FILLER_58_596 ();
 sg13g2_fill_2 FILLER_58_639 ();
 sg13g2_decap_4 FILLER_58_646 ();
 sg13g2_decap_8 FILLER_58_663 ();
 sg13g2_decap_4 FILLER_58_679 ();
 sg13g2_fill_2 FILLER_58_683 ();
 sg13g2_fill_2 FILLER_58_711 ();
 sg13g2_fill_2 FILLER_58_717 ();
 sg13g2_fill_1 FILLER_58_719 ();
 sg13g2_decap_8 FILLER_58_750 ();
 sg13g2_fill_1 FILLER_58_757 ();
 sg13g2_decap_4 FILLER_58_780 ();
 sg13g2_fill_1 FILLER_58_784 ();
 sg13g2_fill_2 FILLER_58_790 ();
 sg13g2_fill_1 FILLER_58_792 ();
 sg13g2_fill_2 FILLER_58_798 ();
 sg13g2_fill_2 FILLER_58_886 ();
 sg13g2_fill_1 FILLER_58_888 ();
 sg13g2_fill_1 FILLER_58_988 ();
 sg13g2_fill_1 FILLER_58_1015 ();
 sg13g2_fill_2 FILLER_58_1020 ();
 sg13g2_fill_2 FILLER_58_1035 ();
 sg13g2_fill_2 FILLER_58_1063 ();
 sg13g2_fill_2 FILLER_58_1179 ();
 sg13g2_fill_2 FILLER_58_1190 ();
 sg13g2_fill_1 FILLER_58_1219 ();
 sg13g2_fill_1 FILLER_58_1225 ();
 sg13g2_fill_2 FILLER_58_1269 ();
 sg13g2_decap_8 FILLER_58_1301 ();
 sg13g2_decap_8 FILLER_58_1308 ();
 sg13g2_decap_8 FILLER_58_1315 ();
 sg13g2_decap_4 FILLER_58_1322 ();
 sg13g2_fill_1 FILLER_58_1362 ();
 sg13g2_fill_1 FILLER_58_1393 ();
 sg13g2_fill_1 FILLER_58_1399 ();
 sg13g2_fill_2 FILLER_58_1408 ();
 sg13g2_fill_1 FILLER_58_1463 ();
 sg13g2_fill_2 FILLER_58_1469 ();
 sg13g2_fill_1 FILLER_58_1471 ();
 sg13g2_fill_2 FILLER_58_1481 ();
 sg13g2_fill_2 FILLER_58_1497 ();
 sg13g2_fill_1 FILLER_58_1518 ();
 sg13g2_fill_2 FILLER_58_1602 ();
 sg13g2_fill_2 FILLER_58_1618 ();
 sg13g2_fill_2 FILLER_58_1633 ();
 sg13g2_fill_2 FILLER_58_1674 ();
 sg13g2_fill_1 FILLER_58_1676 ();
 sg13g2_fill_2 FILLER_58_1718 ();
 sg13g2_fill_2 FILLER_58_1729 ();
 sg13g2_fill_1 FILLER_58_1731 ();
 sg13g2_fill_2 FILLER_58_1743 ();
 sg13g2_fill_1 FILLER_58_1759 ();
 sg13g2_decap_8 FILLER_58_1795 ();
 sg13g2_decap_4 FILLER_58_1802 ();
 sg13g2_fill_1 FILLER_58_1833 ();
 sg13g2_decap_8 FILLER_58_1839 ();
 sg13g2_fill_1 FILLER_58_1846 ();
 sg13g2_decap_8 FILLER_58_1851 ();
 sg13g2_fill_2 FILLER_58_1914 ();
 sg13g2_fill_1 FILLER_58_1916 ();
 sg13g2_fill_2 FILLER_58_2000 ();
 sg13g2_fill_1 FILLER_58_2002 ();
 sg13g2_fill_2 FILLER_58_2038 ();
 sg13g2_decap_4 FILLER_58_2066 ();
 sg13g2_fill_2 FILLER_58_2070 ();
 sg13g2_fill_1 FILLER_58_2088 ();
 sg13g2_fill_2 FILLER_58_2105 ();
 sg13g2_fill_1 FILLER_58_2163 ();
 sg13g2_fill_2 FILLER_58_2292 ();
 sg13g2_fill_1 FILLER_58_2325 ();
 sg13g2_decap_4 FILLER_58_2371 ();
 sg13g2_fill_2 FILLER_58_2375 ();
 sg13g2_fill_2 FILLER_58_2427 ();
 sg13g2_fill_1 FILLER_58_2429 ();
 sg13g2_fill_2 FILLER_58_2452 ();
 sg13g2_fill_1 FILLER_58_2544 ();
 sg13g2_fill_2 FILLER_58_2588 ();
 sg13g2_decap_8 FILLER_58_2620 ();
 sg13g2_decap_8 FILLER_58_2627 ();
 sg13g2_decap_8 FILLER_58_2634 ();
 sg13g2_decap_8 FILLER_58_2641 ();
 sg13g2_decap_8 FILLER_58_2648 ();
 sg13g2_decap_8 FILLER_58_2655 ();
 sg13g2_decap_8 FILLER_58_2662 ();
 sg13g2_decap_4 FILLER_58_2669 ();
 sg13g2_fill_1 FILLER_58_2673 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_decap_8 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_8 FILLER_59_231 ();
 sg13g2_decap_8 FILLER_59_238 ();
 sg13g2_decap_8 FILLER_59_245 ();
 sg13g2_decap_8 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_decap_8 FILLER_59_308 ();
 sg13g2_decap_8 FILLER_59_315 ();
 sg13g2_decap_8 FILLER_59_322 ();
 sg13g2_decap_8 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_decap_4 FILLER_59_350 ();
 sg13g2_fill_1 FILLER_59_354 ();
 sg13g2_decap_8 FILLER_59_390 ();
 sg13g2_decap_4 FILLER_59_397 ();
 sg13g2_decap_8 FILLER_59_409 ();
 sg13g2_decap_8 FILLER_59_416 ();
 sg13g2_decap_8 FILLER_59_433 ();
 sg13g2_fill_1 FILLER_59_440 ();
 sg13g2_decap_4 FILLER_59_449 ();
 sg13g2_fill_1 FILLER_59_453 ();
 sg13g2_decap_8 FILLER_59_485 ();
 sg13g2_decap_4 FILLER_59_492 ();
 sg13g2_decap_8 FILLER_59_553 ();
 sg13g2_fill_2 FILLER_59_560 ();
 sg13g2_fill_1 FILLER_59_592 ();
 sg13g2_fill_1 FILLER_59_633 ();
 sg13g2_fill_2 FILLER_59_643 ();
 sg13g2_fill_1 FILLER_59_645 ();
 sg13g2_fill_2 FILLER_59_654 ();
 sg13g2_fill_1 FILLER_59_656 ();
 sg13g2_fill_2 FILLER_59_668 ();
 sg13g2_fill_2 FILLER_59_690 ();
 sg13g2_fill_1 FILLER_59_701 ();
 sg13g2_fill_1 FILLER_59_741 ();
 sg13g2_decap_8 FILLER_59_755 ();
 sg13g2_fill_2 FILLER_59_762 ();
 sg13g2_fill_1 FILLER_59_764 ();
 sg13g2_fill_1 FILLER_59_769 ();
 sg13g2_fill_2 FILLER_59_775 ();
 sg13g2_fill_1 FILLER_59_817 ();
 sg13g2_fill_2 FILLER_59_826 ();
 sg13g2_fill_2 FILLER_59_875 ();
 sg13g2_fill_1 FILLER_59_881 ();
 sg13g2_fill_2 FILLER_59_913 ();
 sg13g2_fill_1 FILLER_59_945 ();
 sg13g2_fill_2 FILLER_59_1106 ();
 sg13g2_fill_1 FILLER_59_1108 ();
 sg13g2_fill_1 FILLER_59_1166 ();
 sg13g2_fill_2 FILLER_59_1187 ();
 sg13g2_fill_1 FILLER_59_1189 ();
 sg13g2_fill_1 FILLER_59_1221 ();
 sg13g2_fill_1 FILLER_59_1234 ();
 sg13g2_fill_2 FILLER_59_1244 ();
 sg13g2_fill_2 FILLER_59_1263 ();
 sg13g2_fill_1 FILLER_59_1276 ();
 sg13g2_decap_8 FILLER_59_1303 ();
 sg13g2_decap_4 FILLER_59_1310 ();
 sg13g2_fill_1 FILLER_59_1368 ();
 sg13g2_fill_2 FILLER_59_1378 ();
 sg13g2_fill_2 FILLER_59_1385 ();
 sg13g2_fill_2 FILLER_59_1428 ();
 sg13g2_fill_2 FILLER_59_1439 ();
 sg13g2_fill_1 FILLER_59_1521 ();
 sg13g2_fill_1 FILLER_59_1530 ();
 sg13g2_fill_1 FILLER_59_1536 ();
 sg13g2_fill_2 FILLER_59_1547 ();
 sg13g2_fill_2 FILLER_59_1588 ();
 sg13g2_fill_1 FILLER_59_1590 ();
 sg13g2_fill_2 FILLER_59_1674 ();
 sg13g2_fill_1 FILLER_59_1676 ();
 sg13g2_fill_2 FILLER_59_1725 ();
 sg13g2_fill_1 FILLER_59_1727 ();
 sg13g2_fill_1 FILLER_59_1743 ();
 sg13g2_fill_2 FILLER_59_1782 ();
 sg13g2_decap_4 FILLER_59_1810 ();
 sg13g2_fill_1 FILLER_59_1814 ();
 sg13g2_decap_4 FILLER_59_1850 ();
 sg13g2_fill_1 FILLER_59_1854 ();
 sg13g2_fill_1 FILLER_59_1911 ();
 sg13g2_fill_1 FILLER_59_1948 ();
 sg13g2_fill_2 FILLER_59_1984 ();
 sg13g2_fill_1 FILLER_59_1990 ();
 sg13g2_decap_4 FILLER_59_2082 ();
 sg13g2_fill_2 FILLER_59_2086 ();
 sg13g2_fill_2 FILLER_59_2093 ();
 sg13g2_fill_1 FILLER_59_2095 ();
 sg13g2_fill_2 FILLER_59_2100 ();
 sg13g2_fill_2 FILLER_59_2165 ();
 sg13g2_fill_1 FILLER_59_2219 ();
 sg13g2_fill_2 FILLER_59_2229 ();
 sg13g2_fill_2 FILLER_59_2240 ();
 sg13g2_fill_1 FILLER_59_2242 ();
 sg13g2_fill_2 FILLER_59_2282 ();
 sg13g2_fill_2 FILLER_59_2371 ();
 sg13g2_fill_1 FILLER_59_2373 ();
 sg13g2_fill_1 FILLER_59_2404 ();
 sg13g2_fill_1 FILLER_59_2436 ();
 sg13g2_fill_2 FILLER_59_2445 ();
 sg13g2_fill_2 FILLER_59_2546 ();
 sg13g2_fill_1 FILLER_59_2548 ();
 sg13g2_fill_2 FILLER_59_2580 ();
 sg13g2_decap_8 FILLER_59_2613 ();
 sg13g2_decap_8 FILLER_59_2620 ();
 sg13g2_decap_8 FILLER_59_2627 ();
 sg13g2_decap_8 FILLER_59_2634 ();
 sg13g2_decap_8 FILLER_59_2641 ();
 sg13g2_decap_8 FILLER_59_2648 ();
 sg13g2_decap_8 FILLER_59_2655 ();
 sg13g2_decap_8 FILLER_59_2662 ();
 sg13g2_decap_4 FILLER_59_2669 ();
 sg13g2_fill_1 FILLER_59_2673 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_decap_8 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_252 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_decap_8 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_8 FILLER_60_301 ();
 sg13g2_decap_8 FILLER_60_308 ();
 sg13g2_decap_8 FILLER_60_315 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_decap_4 FILLER_60_350 ();
 sg13g2_fill_2 FILLER_60_354 ();
 sg13g2_fill_2 FILLER_60_389 ();
 sg13g2_decap_4 FILLER_60_417 ();
 sg13g2_fill_2 FILLER_60_421 ();
 sg13g2_decap_8 FILLER_60_449 ();
 sg13g2_decap_8 FILLER_60_456 ();
 sg13g2_decap_4 FILLER_60_463 ();
 sg13g2_decap_4 FILLER_60_480 ();
 sg13g2_fill_2 FILLER_60_484 ();
 sg13g2_decap_4 FILLER_60_548 ();
 sg13g2_fill_2 FILLER_60_570 ();
 sg13g2_fill_1 FILLER_60_572 ();
 sg13g2_fill_2 FILLER_60_608 ();
 sg13g2_fill_2 FILLER_60_674 ();
 sg13g2_fill_1 FILLER_60_676 ();
 sg13g2_fill_1 FILLER_60_708 ();
 sg13g2_fill_2 FILLER_60_715 ();
 sg13g2_fill_2 FILLER_60_727 ();
 sg13g2_fill_2 FILLER_60_738 ();
 sg13g2_fill_2 FILLER_60_756 ();
 sg13g2_fill_1 FILLER_60_758 ();
 sg13g2_fill_2 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_807 ();
 sg13g2_decap_4 FILLER_60_814 ();
 sg13g2_fill_1 FILLER_60_818 ();
 sg13g2_decap_8 FILLER_60_827 ();
 sg13g2_fill_1 FILLER_60_834 ();
 sg13g2_decap_4 FILLER_60_858 ();
 sg13g2_fill_1 FILLER_60_866 ();
 sg13g2_fill_2 FILLER_60_876 ();
 sg13g2_decap_4 FILLER_60_882 ();
 sg13g2_fill_2 FILLER_60_911 ();
 sg13g2_fill_2 FILLER_60_922 ();
 sg13g2_fill_2 FILLER_60_964 ();
 sg13g2_fill_1 FILLER_60_966 ();
 sg13g2_fill_2 FILLER_60_977 ();
 sg13g2_fill_1 FILLER_60_1032 ();
 sg13g2_fill_1 FILLER_60_1059 ();
 sg13g2_fill_2 FILLER_60_1082 ();
 sg13g2_fill_1 FILLER_60_1084 ();
 sg13g2_fill_2 FILLER_60_1100 ();
 sg13g2_fill_1 FILLER_60_1111 ();
 sg13g2_fill_2 FILLER_60_1117 ();
 sg13g2_fill_1 FILLER_60_1119 ();
 sg13g2_fill_2 FILLER_60_1138 ();
 sg13g2_fill_1 FILLER_60_1140 ();
 sg13g2_fill_1 FILLER_60_1163 ();
 sg13g2_fill_2 FILLER_60_1202 ();
 sg13g2_fill_1 FILLER_60_1239 ();
 sg13g2_fill_2 FILLER_60_1245 ();
 sg13g2_fill_1 FILLER_60_1304 ();
 sg13g2_fill_2 FILLER_60_1340 ();
 sg13g2_fill_2 FILLER_60_1354 ();
 sg13g2_fill_1 FILLER_60_1356 ();
 sg13g2_fill_2 FILLER_60_1397 ();
 sg13g2_fill_2 FILLER_60_1404 ();
 sg13g2_fill_2 FILLER_60_1411 ();
 sg13g2_fill_1 FILLER_60_1413 ();
 sg13g2_fill_2 FILLER_60_1445 ();
 sg13g2_fill_1 FILLER_60_1635 ();
 sg13g2_fill_1 FILLER_60_1670 ();
 sg13g2_fill_2 FILLER_60_1710 ();
 sg13g2_fill_1 FILLER_60_1712 ();
 sg13g2_fill_1 FILLER_60_1817 ();
 sg13g2_fill_1 FILLER_60_1844 ();
 sg13g2_decap_8 FILLER_60_1853 ();
 sg13g2_fill_2 FILLER_60_1865 ();
 sg13g2_fill_1 FILLER_60_1880 ();
 sg13g2_decap_4 FILLER_60_1898 ();
 sg13g2_fill_2 FILLER_60_1910 ();
 sg13g2_fill_1 FILLER_60_1925 ();
 sg13g2_fill_1 FILLER_60_1960 ();
 sg13g2_decap_4 FILLER_60_1973 ();
 sg13g2_fill_2 FILLER_60_1977 ();
 sg13g2_fill_2 FILLER_60_2018 ();
 sg13g2_fill_2 FILLER_60_2075 ();
 sg13g2_fill_1 FILLER_60_2077 ();
 sg13g2_decap_4 FILLER_60_2089 ();
 sg13g2_fill_2 FILLER_60_2093 ();
 sg13g2_fill_2 FILLER_60_2108 ();
 sg13g2_fill_1 FILLER_60_2110 ();
 sg13g2_fill_1 FILLER_60_2120 ();
 sg13g2_fill_1 FILLER_60_2134 ();
 sg13g2_fill_2 FILLER_60_2165 ();
 sg13g2_fill_1 FILLER_60_2167 ();
 sg13g2_fill_2 FILLER_60_2173 ();
 sg13g2_fill_1 FILLER_60_2175 ();
 sg13g2_fill_2 FILLER_60_2207 ();
 sg13g2_fill_1 FILLER_60_2214 ();
 sg13g2_fill_2 FILLER_60_2240 ();
 sg13g2_fill_1 FILLER_60_2242 ();
 sg13g2_fill_2 FILLER_60_2252 ();
 sg13g2_fill_1 FILLER_60_2254 ();
 sg13g2_fill_1 FILLER_60_2317 ();
 sg13g2_fill_2 FILLER_60_2422 ();
 sg13g2_fill_1 FILLER_60_2424 ();
 sg13g2_fill_2 FILLER_60_2469 ();
 sg13g2_fill_1 FILLER_60_2482 ();
 sg13g2_decap_4 FILLER_60_2544 ();
 sg13g2_fill_2 FILLER_60_2552 ();
 sg13g2_decap_8 FILLER_60_2614 ();
 sg13g2_decap_8 FILLER_60_2621 ();
 sg13g2_decap_8 FILLER_60_2628 ();
 sg13g2_decap_8 FILLER_60_2635 ();
 sg13g2_decap_8 FILLER_60_2642 ();
 sg13g2_decap_8 FILLER_60_2649 ();
 sg13g2_decap_8 FILLER_60_2656 ();
 sg13g2_decap_8 FILLER_60_2663 ();
 sg13g2_decap_4 FILLER_60_2670 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_decap_8 FILLER_61_189 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_decap_8 FILLER_61_224 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_259 ();
 sg13g2_decap_8 FILLER_61_266 ();
 sg13g2_decap_8 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_decap_8 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_322 ();
 sg13g2_decap_8 FILLER_61_329 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_fill_1 FILLER_61_357 ();
 sg13g2_fill_2 FILLER_61_423 ();
 sg13g2_fill_1 FILLER_61_425 ();
 sg13g2_decap_8 FILLER_61_452 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_fill_2 FILLER_61_466 ();
 sg13g2_decap_8 FILLER_61_472 ();
 sg13g2_fill_2 FILLER_61_479 ();
 sg13g2_fill_1 FILLER_61_515 ();
 sg13g2_decap_8 FILLER_61_526 ();
 sg13g2_decap_8 FILLER_61_533 ();
 sg13g2_decap_8 FILLER_61_540 ();
 sg13g2_decap_4 FILLER_61_547 ();
 sg13g2_fill_1 FILLER_61_551 ();
 sg13g2_fill_2 FILLER_61_582 ();
 sg13g2_fill_2 FILLER_61_598 ();
 sg13g2_decap_4 FILLER_61_610 ();
 sg13g2_fill_2 FILLER_61_635 ();
 sg13g2_fill_1 FILLER_61_642 ();
 sg13g2_fill_2 FILLER_61_670 ();
 sg13g2_fill_1 FILLER_61_672 ();
 sg13g2_fill_2 FILLER_61_704 ();
 sg13g2_fill_1 FILLER_61_706 ();
 sg13g2_fill_2 FILLER_61_721 ();
 sg13g2_fill_2 FILLER_61_728 ();
 sg13g2_fill_1 FILLER_61_730 ();
 sg13g2_fill_2 FILLER_61_744 ();
 sg13g2_fill_1 FILLER_61_746 ();
 sg13g2_fill_1 FILLER_61_787 ();
 sg13g2_fill_2 FILLER_61_802 ();
 sg13g2_fill_2 FILLER_61_817 ();
 sg13g2_fill_1 FILLER_61_819 ();
 sg13g2_decap_8 FILLER_61_824 ();
 sg13g2_decap_8 FILLER_61_831 ();
 sg13g2_decap_8 FILLER_61_838 ();
 sg13g2_fill_2 FILLER_61_845 ();
 sg13g2_fill_2 FILLER_61_851 ();
 sg13g2_decap_8 FILLER_61_863 ();
 sg13g2_decap_4 FILLER_61_870 ();
 sg13g2_fill_2 FILLER_61_878 ();
 sg13g2_fill_1 FILLER_61_880 ();
 sg13g2_fill_2 FILLER_61_891 ();
 sg13g2_fill_1 FILLER_61_893 ();
 sg13g2_fill_1 FILLER_61_903 ();
 sg13g2_fill_2 FILLER_61_924 ();
 sg13g2_fill_1 FILLER_61_926 ();
 sg13g2_fill_2 FILLER_61_957 ();
 sg13g2_fill_2 FILLER_61_963 ();
 sg13g2_fill_1 FILLER_61_965 ();
 sg13g2_fill_2 FILLER_61_1024 ();
 sg13g2_fill_1 FILLER_61_1026 ();
 sg13g2_fill_1 FILLER_61_1071 ();
 sg13g2_decap_8 FILLER_61_1082 ();
 sg13g2_fill_2 FILLER_61_1089 ();
 sg13g2_fill_1 FILLER_61_1091 ();
 sg13g2_fill_2 FILLER_61_1123 ();
 sg13g2_fill_2 FILLER_61_1164 ();
 sg13g2_fill_1 FILLER_61_1166 ();
 sg13g2_fill_2 FILLER_61_1193 ();
 sg13g2_fill_1 FILLER_61_1204 ();
 sg13g2_fill_2 FILLER_61_1215 ();
 sg13g2_fill_1 FILLER_61_1233 ();
 sg13g2_fill_1 FILLER_61_1273 ();
 sg13g2_fill_1 FILLER_61_1356 ();
 sg13g2_fill_2 FILLER_61_1399 ();
 sg13g2_fill_1 FILLER_61_1401 ();
 sg13g2_fill_2 FILLER_61_1419 ();
 sg13g2_fill_2 FILLER_61_1434 ();
 sg13g2_fill_2 FILLER_61_1473 ();
 sg13g2_fill_1 FILLER_61_1475 ();
 sg13g2_fill_1 FILLER_61_1555 ();
 sg13g2_fill_1 FILLER_61_1565 ();
 sg13g2_fill_1 FILLER_61_1574 ();
 sg13g2_decap_4 FILLER_61_1604 ();
 sg13g2_fill_1 FILLER_61_1608 ();
 sg13g2_fill_1 FILLER_61_1639 ();
 sg13g2_fill_1 FILLER_61_1658 ();
 sg13g2_fill_1 FILLER_61_1681 ();
 sg13g2_fill_1 FILLER_61_1713 ();
 sg13g2_fill_2 FILLER_61_1758 ();
 sg13g2_fill_2 FILLER_61_1809 ();
 sg13g2_fill_2 FILLER_61_1826 ();
 sg13g2_fill_1 FILLER_61_1828 ();
 sg13g2_decap_8 FILLER_61_1861 ();
 sg13g2_decap_8 FILLER_61_1868 ();
 sg13g2_decap_4 FILLER_61_1875 ();
 sg13g2_fill_1 FILLER_61_1879 ();
 sg13g2_decap_4 FILLER_61_1888 ();
 sg13g2_fill_1 FILLER_61_1892 ();
 sg13g2_fill_1 FILLER_61_1928 ();
 sg13g2_fill_1 FILLER_61_1938 ();
 sg13g2_decap_4 FILLER_61_1979 ();
 sg13g2_fill_2 FILLER_61_1983 ();
 sg13g2_decap_4 FILLER_61_2065 ();
 sg13g2_fill_1 FILLER_61_2069 ();
 sg13g2_fill_2 FILLER_61_2097 ();
 sg13g2_fill_1 FILLER_61_2099 ();
 sg13g2_decap_8 FILLER_61_2120 ();
 sg13g2_decap_4 FILLER_61_2127 ();
 sg13g2_fill_1 FILLER_61_2136 ();
 sg13g2_fill_2 FILLER_61_2180 ();
 sg13g2_fill_1 FILLER_61_2182 ();
 sg13g2_fill_1 FILLER_61_2198 ();
 sg13g2_fill_2 FILLER_61_2217 ();
 sg13g2_decap_4 FILLER_61_2264 ();
 sg13g2_fill_2 FILLER_61_2280 ();
 sg13g2_fill_2 FILLER_61_2304 ();
 sg13g2_fill_2 FILLER_61_2332 ();
 sg13g2_fill_1 FILLER_61_2334 ();
 sg13g2_fill_1 FILLER_61_2370 ();
 sg13g2_fill_1 FILLER_61_2381 ();
 sg13g2_fill_1 FILLER_61_2396 ();
 sg13g2_fill_1 FILLER_61_2437 ();
 sg13g2_decap_8 FILLER_61_2482 ();
 sg13g2_decap_4 FILLER_61_2489 ();
 sg13g2_fill_1 FILLER_61_2493 ();
 sg13g2_decap_4 FILLER_61_2504 ();
 sg13g2_fill_1 FILLER_61_2508 ();
 sg13g2_decap_8 FILLER_61_2513 ();
 sg13g2_fill_2 FILLER_61_2520 ();
 sg13g2_decap_8 FILLER_61_2535 ();
 sg13g2_decap_8 FILLER_61_2542 ();
 sg13g2_decap_8 FILLER_61_2549 ();
 sg13g2_decap_4 FILLER_61_2556 ();
 sg13g2_decap_8 FILLER_61_2605 ();
 sg13g2_decap_8 FILLER_61_2612 ();
 sg13g2_decap_8 FILLER_61_2619 ();
 sg13g2_decap_8 FILLER_61_2626 ();
 sg13g2_decap_8 FILLER_61_2633 ();
 sg13g2_decap_8 FILLER_61_2640 ();
 sg13g2_decap_8 FILLER_61_2647 ();
 sg13g2_decap_8 FILLER_61_2654 ();
 sg13g2_decap_8 FILLER_61_2661 ();
 sg13g2_decap_4 FILLER_61_2668 ();
 sg13g2_fill_2 FILLER_61_2672 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_decap_8 FILLER_62_245 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_280 ();
 sg13g2_decap_8 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_4 FILLER_62_357 ();
 sg13g2_decap_4 FILLER_62_387 ();
 sg13g2_fill_1 FILLER_62_391 ();
 sg13g2_decap_8 FILLER_62_418 ();
 sg13g2_fill_2 FILLER_62_451 ();
 sg13g2_fill_2 FILLER_62_531 ();
 sg13g2_decap_8 FILLER_62_538 ();
 sg13g2_decap_4 FILLER_62_545 ();
 sg13g2_fill_2 FILLER_62_549 ();
 sg13g2_fill_1 FILLER_62_577 ();
 sg13g2_fill_2 FILLER_62_591 ();
 sg13g2_fill_1 FILLER_62_593 ();
 sg13g2_fill_1 FILLER_62_598 ();
 sg13g2_fill_1 FILLER_62_608 ();
 sg13g2_fill_1 FILLER_62_632 ();
 sg13g2_fill_1 FILLER_62_651 ();
 sg13g2_fill_1 FILLER_62_689 ();
 sg13g2_fill_1 FILLER_62_704 ();
 sg13g2_fill_1 FILLER_62_711 ();
 sg13g2_fill_2 FILLER_62_751 ();
 sg13g2_fill_1 FILLER_62_753 ();
 sg13g2_fill_2 FILLER_62_793 ();
 sg13g2_decap_8 FILLER_62_835 ();
 sg13g2_fill_2 FILLER_62_842 ();
 sg13g2_fill_2 FILLER_62_852 ();
 sg13g2_fill_1 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_930 ();
 sg13g2_fill_2 FILLER_62_972 ();
 sg13g2_fill_1 FILLER_62_1000 ();
 sg13g2_fill_2 FILLER_62_1041 ();
 sg13g2_fill_1 FILLER_62_1070 ();
 sg13g2_fill_2 FILLER_62_1080 ();
 sg13g2_fill_2 FILLER_62_1131 ();
 sg13g2_fill_2 FILLER_62_1169 ();
 sg13g2_fill_2 FILLER_62_1273 ();
 sg13g2_fill_2 FILLER_62_1392 ();
 sg13g2_fill_1 FILLER_62_1394 ();
 sg13g2_decap_4 FILLER_62_1404 ();
 sg13g2_fill_2 FILLER_62_1417 ();
 sg13g2_fill_1 FILLER_62_1419 ();
 sg13g2_fill_2 FILLER_62_1429 ();
 sg13g2_fill_2 FILLER_62_1470 ();
 sg13g2_decap_4 FILLER_62_1489 ();
 sg13g2_fill_1 FILLER_62_1493 ();
 sg13g2_fill_1 FILLER_62_1506 ();
 sg13g2_fill_2 FILLER_62_1559 ();
 sg13g2_fill_2 FILLER_62_1628 ();
 sg13g2_fill_2 FILLER_62_1644 ();
 sg13g2_fill_1 FILLER_62_1646 ();
 sg13g2_fill_2 FILLER_62_1682 ();
 sg13g2_fill_2 FILLER_62_1690 ();
 sg13g2_fill_1 FILLER_62_1692 ();
 sg13g2_fill_2 FILLER_62_1721 ();
 sg13g2_fill_1 FILLER_62_1748 ();
 sg13g2_fill_1 FILLER_62_1832 ();
 sg13g2_fill_2 FILLER_62_1855 ();
 sg13g2_fill_1 FILLER_62_1857 ();
 sg13g2_fill_1 FILLER_62_1889 ();
 sg13g2_fill_2 FILLER_62_1979 ();
 sg13g2_fill_2 FILLER_62_2011 ();
 sg13g2_decap_4 FILLER_62_2060 ();
 sg13g2_fill_2 FILLER_62_2116 ();
 sg13g2_fill_1 FILLER_62_2118 ();
 sg13g2_fill_1 FILLER_62_2227 ();
 sg13g2_fill_2 FILLER_62_2259 ();
 sg13g2_fill_1 FILLER_62_2274 ();
 sg13g2_fill_1 FILLER_62_2279 ();
 sg13g2_decap_4 FILLER_62_2284 ();
 sg13g2_fill_2 FILLER_62_2288 ();
 sg13g2_fill_1 FILLER_62_2294 ();
 sg13g2_decap_4 FILLER_62_2321 ();
 sg13g2_fill_1 FILLER_62_2325 ();
 sg13g2_fill_2 FILLER_62_2334 ();
 sg13g2_fill_1 FILLER_62_2336 ();
 sg13g2_decap_8 FILLER_62_2357 ();
 sg13g2_decap_4 FILLER_62_2364 ();
 sg13g2_fill_1 FILLER_62_2368 ();
 sg13g2_fill_2 FILLER_62_2395 ();
 sg13g2_fill_1 FILLER_62_2459 ();
 sg13g2_fill_2 FILLER_62_2473 ();
 sg13g2_fill_1 FILLER_62_2526 ();
 sg13g2_fill_1 FILLER_62_2566 ();
 sg13g2_decap_8 FILLER_62_2598 ();
 sg13g2_decap_8 FILLER_62_2605 ();
 sg13g2_decap_8 FILLER_62_2612 ();
 sg13g2_decap_8 FILLER_62_2619 ();
 sg13g2_decap_8 FILLER_62_2626 ();
 sg13g2_decap_8 FILLER_62_2633 ();
 sg13g2_decap_8 FILLER_62_2640 ();
 sg13g2_decap_8 FILLER_62_2647 ();
 sg13g2_decap_8 FILLER_62_2654 ();
 sg13g2_decap_8 FILLER_62_2661 ();
 sg13g2_decap_4 FILLER_62_2668 ();
 sg13g2_fill_2 FILLER_62_2672 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_266 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_8 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_315 ();
 sg13g2_decap_8 FILLER_63_322 ();
 sg13g2_decap_8 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_fill_2 FILLER_63_364 ();
 sg13g2_fill_1 FILLER_63_366 ();
 sg13g2_decap_8 FILLER_63_380 ();
 sg13g2_decap_8 FILLER_63_387 ();
 sg13g2_decap_8 FILLER_63_394 ();
 sg13g2_decap_8 FILLER_63_401 ();
 sg13g2_decap_4 FILLER_63_408 ();
 sg13g2_fill_2 FILLER_63_412 ();
 sg13g2_fill_2 FILLER_63_450 ();
 sg13g2_decap_8 FILLER_63_491 ();
 sg13g2_fill_2 FILLER_63_498 ();
 sg13g2_decap_4 FILLER_63_525 ();
 sg13g2_decap_8 FILLER_63_544 ();
 sg13g2_decap_4 FILLER_63_551 ();
 sg13g2_fill_2 FILLER_63_581 ();
 sg13g2_fill_1 FILLER_63_583 ();
 sg13g2_fill_1 FILLER_63_607 ();
 sg13g2_fill_2 FILLER_63_618 ();
 sg13g2_fill_2 FILLER_63_672 ();
 sg13g2_fill_1 FILLER_63_674 ();
 sg13g2_fill_1 FILLER_63_740 ();
 sg13g2_fill_1 FILLER_63_767 ();
 sg13g2_fill_2 FILLER_63_791 ();
 sg13g2_fill_2 FILLER_63_817 ();
 sg13g2_fill_2 FILLER_63_833 ();
 sg13g2_fill_1 FILLER_63_835 ();
 sg13g2_fill_2 FILLER_63_857 ();
 sg13g2_fill_1 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_923 ();
 sg13g2_fill_1 FILLER_63_978 ();
 sg13g2_fill_2 FILLER_63_994 ();
 sg13g2_fill_1 FILLER_63_1005 ();
 sg13g2_fill_2 FILLER_63_1078 ();
 sg13g2_fill_1 FILLER_63_1115 ();
 sg13g2_fill_1 FILLER_63_1122 ();
 sg13g2_fill_1 FILLER_63_1157 ();
 sg13g2_fill_1 FILLER_63_1196 ();
 sg13g2_fill_1 FILLER_63_1202 ();
 sg13g2_fill_1 FILLER_63_1209 ();
 sg13g2_fill_2 FILLER_63_1218 ();
 sg13g2_fill_1 FILLER_63_1260 ();
 sg13g2_decap_8 FILLER_63_1297 ();
 sg13g2_fill_1 FILLER_63_1304 ();
 sg13g2_fill_1 FILLER_63_1313 ();
 sg13g2_fill_1 FILLER_63_1342 ();
 sg13g2_decap_4 FILLER_63_1377 ();
 sg13g2_fill_2 FILLER_63_1381 ();
 sg13g2_fill_2 FILLER_63_1387 ();
 sg13g2_fill_2 FILLER_63_1398 ();
 sg13g2_decap_8 FILLER_63_1497 ();
 sg13g2_decap_4 FILLER_63_1504 ();
 sg13g2_fill_2 FILLER_63_1520 ();
 sg13g2_fill_1 FILLER_63_1522 ();
 sg13g2_fill_2 FILLER_63_1561 ();
 sg13g2_fill_1 FILLER_63_1563 ();
 sg13g2_fill_2 FILLER_63_1590 ();
 sg13g2_fill_1 FILLER_63_1592 ();
 sg13g2_fill_2 FILLER_63_1664 ();
 sg13g2_fill_1 FILLER_63_1666 ();
 sg13g2_fill_1 FILLER_63_1680 ();
 sg13g2_fill_2 FILLER_63_1710 ();
 sg13g2_fill_1 FILLER_63_1720 ();
 sg13g2_fill_2 FILLER_63_1739 ();
 sg13g2_fill_1 FILLER_63_1741 ();
 sg13g2_fill_2 FILLER_63_1777 ();
 sg13g2_fill_2 FILLER_63_1787 ();
 sg13g2_fill_1 FILLER_63_1815 ();
 sg13g2_fill_1 FILLER_63_1847 ();
 sg13g2_fill_1 FILLER_63_1911 ();
 sg13g2_fill_2 FILLER_63_1987 ();
 sg13g2_fill_1 FILLER_63_1989 ();
 sg13g2_fill_1 FILLER_63_2005 ();
 sg13g2_fill_2 FILLER_63_2031 ();
 sg13g2_fill_1 FILLER_63_2039 ();
 sg13g2_fill_1 FILLER_63_2066 ();
 sg13g2_fill_2 FILLER_63_2125 ();
 sg13g2_fill_1 FILLER_63_2127 ();
 sg13g2_fill_1 FILLER_63_2173 ();
 sg13g2_fill_2 FILLER_63_2235 ();
 sg13g2_fill_1 FILLER_63_2237 ();
 sg13g2_decap_4 FILLER_63_2274 ();
 sg13g2_decap_4 FILLER_63_2306 ();
 sg13g2_fill_1 FILLER_63_2310 ();
 sg13g2_decap_8 FILLER_63_2316 ();
 sg13g2_decap_8 FILLER_63_2323 ();
 sg13g2_decap_8 FILLER_63_2330 ();
 sg13g2_decap_4 FILLER_63_2341 ();
 sg13g2_decap_8 FILLER_63_2370 ();
 sg13g2_fill_2 FILLER_63_2377 ();
 sg13g2_fill_1 FILLER_63_2379 ();
 sg13g2_fill_1 FILLER_63_2384 ();
 sg13g2_fill_1 FILLER_63_2394 ();
 sg13g2_fill_2 FILLER_63_2424 ();
 sg13g2_fill_1 FILLER_63_2426 ();
 sg13g2_fill_2 FILLER_63_2448 ();
 sg13g2_fill_2 FILLER_63_2455 ();
 sg13g2_fill_1 FILLER_63_2457 ();
 sg13g2_decap_4 FILLER_63_2492 ();
 sg13g2_fill_1 FILLER_63_2496 ();
 sg13g2_decap_8 FILLER_63_2605 ();
 sg13g2_decap_8 FILLER_63_2612 ();
 sg13g2_decap_8 FILLER_63_2619 ();
 sg13g2_decap_8 FILLER_63_2626 ();
 sg13g2_decap_8 FILLER_63_2633 ();
 sg13g2_decap_8 FILLER_63_2640 ();
 sg13g2_decap_8 FILLER_63_2647 ();
 sg13g2_decap_8 FILLER_63_2654 ();
 sg13g2_decap_8 FILLER_63_2661 ();
 sg13g2_decap_4 FILLER_63_2668 ();
 sg13g2_fill_2 FILLER_63_2672 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_decap_8 FILLER_64_175 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_decap_8 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_decap_8 FILLER_64_217 ();
 sg13g2_decap_8 FILLER_64_224 ();
 sg13g2_decap_8 FILLER_64_231 ();
 sg13g2_decap_8 FILLER_64_238 ();
 sg13g2_decap_8 FILLER_64_245 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_decap_8 FILLER_64_280 ();
 sg13g2_decap_8 FILLER_64_287 ();
 sg13g2_decap_8 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_decap_8 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_329 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_fill_1 FILLER_64_357 ();
 sg13g2_decap_4 FILLER_64_389 ();
 sg13g2_fill_1 FILLER_64_419 ();
 sg13g2_decap_8 FILLER_64_448 ();
 sg13g2_decap_8 FILLER_64_455 ();
 sg13g2_fill_2 FILLER_64_470 ();
 sg13g2_decap_8 FILLER_64_482 ();
 sg13g2_decap_8 FILLER_64_489 ();
 sg13g2_decap_8 FILLER_64_496 ();
 sg13g2_decap_4 FILLER_64_503 ();
 sg13g2_decap_8 FILLER_64_522 ();
 sg13g2_fill_2 FILLER_64_529 ();
 sg13g2_fill_1 FILLER_64_587 ();
 sg13g2_fill_2 FILLER_64_597 ();
 sg13g2_fill_1 FILLER_64_678 ();
 sg13g2_fill_2 FILLER_64_692 ();
 sg13g2_fill_1 FILLER_64_694 ();
 sg13g2_fill_2 FILLER_64_723 ();
 sg13g2_fill_1 FILLER_64_748 ();
 sg13g2_fill_2 FILLER_64_775 ();
 sg13g2_fill_1 FILLER_64_777 ();
 sg13g2_fill_1 FILLER_64_809 ();
 sg13g2_fill_1 FILLER_64_849 ();
 sg13g2_fill_2 FILLER_64_885 ();
 sg13g2_fill_1 FILLER_64_887 ();
 sg13g2_fill_1 FILLER_64_905 ();
 sg13g2_fill_2 FILLER_64_910 ();
 sg13g2_fill_2 FILLER_64_921 ();
 sg13g2_fill_1 FILLER_64_973 ();
 sg13g2_fill_1 FILLER_64_989 ();
 sg13g2_fill_1 FILLER_64_1003 ();
 sg13g2_fill_2 FILLER_64_1060 ();
 sg13g2_fill_1 FILLER_64_1062 ();
 sg13g2_fill_1 FILLER_64_1068 ();
 sg13g2_fill_1 FILLER_64_1101 ();
 sg13g2_decap_4 FILLER_64_1153 ();
 sg13g2_fill_1 FILLER_64_1157 ();
 sg13g2_fill_1 FILLER_64_1177 ();
 sg13g2_fill_2 FILLER_64_1254 ();
 sg13g2_decap_8 FILLER_64_1292 ();
 sg13g2_decap_8 FILLER_64_1299 ();
 sg13g2_fill_2 FILLER_64_1306 ();
 sg13g2_fill_1 FILLER_64_1308 ();
 sg13g2_fill_2 FILLER_64_1314 ();
 sg13g2_fill_1 FILLER_64_1316 ();
 sg13g2_fill_2 FILLER_64_1322 ();
 sg13g2_fill_2 FILLER_64_1329 ();
 sg13g2_decap_4 FILLER_64_1387 ();
 sg13g2_fill_1 FILLER_64_1391 ();
 sg13g2_fill_2 FILLER_64_1405 ();
 sg13g2_fill_2 FILLER_64_1420 ();
 sg13g2_fill_2 FILLER_64_1426 ();
 sg13g2_fill_1 FILLER_64_1491 ();
 sg13g2_fill_2 FILLER_64_1500 ();
 sg13g2_fill_1 FILLER_64_1502 ();
 sg13g2_fill_1 FILLER_64_1506 ();
 sg13g2_fill_1 FILLER_64_1525 ();
 sg13g2_decap_8 FILLER_64_1574 ();
 sg13g2_decap_8 FILLER_64_1581 ();
 sg13g2_decap_8 FILLER_64_1588 ();
 sg13g2_fill_2 FILLER_64_1595 ();
 sg13g2_fill_2 FILLER_64_1632 ();
 sg13g2_fill_2 FILLER_64_1674 ();
 sg13g2_fill_1 FILLER_64_1710 ();
 sg13g2_fill_1 FILLER_64_1746 ();
 sg13g2_fill_1 FILLER_64_1855 ();
 sg13g2_fill_2 FILLER_64_1925 ();
 sg13g2_fill_2 FILLER_64_1932 ();
 sg13g2_fill_2 FILLER_64_1977 ();
 sg13g2_fill_1 FILLER_64_1979 ();
 sg13g2_fill_1 FILLER_64_1992 ();
 sg13g2_fill_1 FILLER_64_2016 ();
 sg13g2_decap_4 FILLER_64_2069 ();
 sg13g2_fill_1 FILLER_64_2110 ();
 sg13g2_decap_4 FILLER_64_2170 ();
 sg13g2_fill_1 FILLER_64_2174 ();
 sg13g2_fill_1 FILLER_64_2235 ();
 sg13g2_decap_8 FILLER_64_2288 ();
 sg13g2_fill_2 FILLER_64_2295 ();
 sg13g2_decap_8 FILLER_64_2301 ();
 sg13g2_fill_2 FILLER_64_2334 ();
 sg13g2_fill_1 FILLER_64_2336 ();
 sg13g2_decap_8 FILLER_64_2368 ();
 sg13g2_decap_8 FILLER_64_2375 ();
 sg13g2_decap_8 FILLER_64_2382 ();
 sg13g2_decap_8 FILLER_64_2416 ();
 sg13g2_fill_1 FILLER_64_2437 ();
 sg13g2_decap_4 FILLER_64_2492 ();
 sg13g2_fill_1 FILLER_64_2496 ();
 sg13g2_fill_2 FILLER_64_2516 ();
 sg13g2_fill_1 FILLER_64_2518 ();
 sg13g2_decap_8 FILLER_64_2611 ();
 sg13g2_decap_8 FILLER_64_2618 ();
 sg13g2_decap_8 FILLER_64_2625 ();
 sg13g2_decap_8 FILLER_64_2632 ();
 sg13g2_decap_8 FILLER_64_2639 ();
 sg13g2_decap_8 FILLER_64_2646 ();
 sg13g2_decap_8 FILLER_64_2653 ();
 sg13g2_decap_8 FILLER_64_2660 ();
 sg13g2_decap_8 FILLER_64_2667 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_decap_8 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_266 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_294 ();
 sg13g2_decap_8 FILLER_65_301 ();
 sg13g2_decap_8 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_8 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_4 FILLER_65_350 ();
 sg13g2_fill_2 FILLER_65_354 ();
 sg13g2_fill_2 FILLER_65_395 ();
 sg13g2_fill_1 FILLER_65_397 ();
 sg13g2_decap_8 FILLER_65_403 ();
 sg13g2_decap_8 FILLER_65_415 ();
 sg13g2_decap_4 FILLER_65_422 ();
 sg13g2_decap_8 FILLER_65_457 ();
 sg13g2_fill_2 FILLER_65_464 ();
 sg13g2_fill_1 FILLER_65_466 ();
 sg13g2_decap_4 FILLER_65_492 ();
 sg13g2_fill_2 FILLER_65_496 ();
 sg13g2_decap_8 FILLER_65_524 ();
 sg13g2_fill_1 FILLER_65_531 ();
 sg13g2_decap_4 FILLER_65_558 ();
 sg13g2_fill_1 FILLER_65_588 ();
 sg13g2_fill_2 FILLER_65_647 ();
 sg13g2_fill_1 FILLER_65_649 ();
 sg13g2_fill_2 FILLER_65_665 ();
 sg13g2_fill_2 FILLER_65_709 ();
 sg13g2_fill_1 FILLER_65_711 ();
 sg13g2_fill_2 FILLER_65_747 ();
 sg13g2_fill_1 FILLER_65_769 ();
 sg13g2_fill_2 FILLER_65_790 ();
 sg13g2_fill_1 FILLER_65_792 ();
 sg13g2_fill_1 FILLER_65_819 ();
 sg13g2_decap_8 FILLER_65_824 ();
 sg13g2_fill_2 FILLER_65_831 ();
 sg13g2_fill_1 FILLER_65_833 ();
 sg13g2_decap_8 FILLER_65_842 ();
 sg13g2_fill_1 FILLER_65_858 ();
 sg13g2_fill_1 FILLER_65_897 ();
 sg13g2_fill_2 FILLER_65_910 ();
 sg13g2_decap_8 FILLER_65_920 ();
 sg13g2_fill_2 FILLER_65_927 ();
 sg13g2_fill_1 FILLER_65_929 ();
 sg13g2_fill_1 FILLER_65_935 ();
 sg13g2_fill_2 FILLER_65_953 ();
 sg13g2_fill_2 FILLER_65_963 ();
 sg13g2_fill_1 FILLER_65_965 ();
 sg13g2_fill_2 FILLER_65_972 ();
 sg13g2_fill_1 FILLER_65_974 ();
 sg13g2_decap_4 FILLER_65_979 ();
 sg13g2_fill_2 FILLER_65_1026 ();
 sg13g2_fill_1 FILLER_65_1074 ();
 sg13g2_fill_1 FILLER_65_1084 ();
 sg13g2_fill_2 FILLER_65_1102 ();
 sg13g2_fill_1 FILLER_65_1104 ();
 sg13g2_fill_2 FILLER_65_1141 ();
 sg13g2_fill_2 FILLER_65_1178 ();
 sg13g2_fill_2 FILLER_65_1245 ();
 sg13g2_fill_1 FILLER_65_1251 ();
 sg13g2_fill_1 FILLER_65_1269 ();
 sg13g2_fill_2 FILLER_65_1283 ();
 sg13g2_fill_2 FILLER_65_1389 ();
 sg13g2_fill_1 FILLER_65_1520 ();
 sg13g2_fill_1 FILLER_65_1525 ();
 sg13g2_decap_8 FILLER_65_1534 ();
 sg13g2_fill_2 FILLER_65_1541 ();
 sg13g2_fill_1 FILLER_65_1543 ();
 sg13g2_fill_1 FILLER_65_1548 ();
 sg13g2_fill_2 FILLER_65_1557 ();
 sg13g2_fill_2 FILLER_65_1585 ();
 sg13g2_fill_1 FILLER_65_1587 ();
 sg13g2_decap_8 FILLER_65_1594 ();
 sg13g2_fill_2 FILLER_65_1601 ();
 sg13g2_fill_1 FILLER_65_1603 ();
 sg13g2_fill_2 FILLER_65_1626 ();
 sg13g2_fill_1 FILLER_65_1628 ();
 sg13g2_fill_1 FILLER_65_1651 ();
 sg13g2_decap_4 FILLER_65_1698 ();
 sg13g2_fill_1 FILLER_65_1702 ();
 sg13g2_fill_2 FILLER_65_1756 ();
 sg13g2_fill_1 FILLER_65_1758 ();
 sg13g2_fill_1 FILLER_65_1790 ();
 sg13g2_fill_2 FILLER_65_1830 ();
 sg13g2_fill_1 FILLER_65_1832 ();
 sg13g2_fill_1 FILLER_65_1893 ();
 sg13g2_fill_1 FILLER_65_1902 ();
 sg13g2_fill_1 FILLER_65_1907 ();
 sg13g2_fill_1 FILLER_65_1922 ();
 sg13g2_decap_8 FILLER_65_1976 ();
 sg13g2_decap_4 FILLER_65_1983 ();
 sg13g2_fill_2 FILLER_65_1987 ();
 sg13g2_fill_2 FILLER_65_1994 ();
 sg13g2_fill_1 FILLER_65_1996 ();
 sg13g2_decap_8 FILLER_65_2017 ();
 sg13g2_fill_2 FILLER_65_2084 ();
 sg13g2_fill_1 FILLER_65_2086 ();
 sg13g2_fill_2 FILLER_65_2149 ();
 sg13g2_fill_1 FILLER_65_2151 ();
 sg13g2_fill_1 FILLER_65_2161 ();
 sg13g2_decap_4 FILLER_65_2168 ();
 sg13g2_decap_8 FILLER_65_2176 ();
 sg13g2_fill_2 FILLER_65_2183 ();
 sg13g2_fill_1 FILLER_65_2185 ();
 sg13g2_fill_1 FILLER_65_2194 ();
 sg13g2_fill_2 FILLER_65_2204 ();
 sg13g2_fill_1 FILLER_65_2206 ();
 sg13g2_fill_2 FILLER_65_2236 ();
 sg13g2_fill_1 FILLER_65_2248 ();
 sg13g2_fill_2 FILLER_65_2291 ();
 sg13g2_fill_1 FILLER_65_2293 ();
 sg13g2_fill_1 FILLER_65_2300 ();
 sg13g2_fill_1 FILLER_65_2332 ();
 sg13g2_fill_1 FILLER_65_2377 ();
 sg13g2_fill_2 FILLER_65_2394 ();
 sg13g2_fill_1 FILLER_65_2396 ();
 sg13g2_fill_1 FILLER_65_2407 ();
 sg13g2_fill_2 FILLER_65_2438 ();
 sg13g2_fill_1 FILLER_65_2440 ();
 sg13g2_fill_2 FILLER_65_2451 ();
 sg13g2_decap_4 FILLER_65_2497 ();
 sg13g2_fill_2 FILLER_65_2501 ();
 sg13g2_fill_2 FILLER_65_2513 ();
 sg13g2_fill_2 FILLER_65_2542 ();
 sg13g2_fill_1 FILLER_65_2544 ();
 sg13g2_fill_2 FILLER_65_2558 ();
 sg13g2_fill_1 FILLER_65_2560 ();
 sg13g2_fill_2 FILLER_65_2592 ();
 sg13g2_decap_8 FILLER_65_2612 ();
 sg13g2_decap_8 FILLER_65_2619 ();
 sg13g2_decap_8 FILLER_65_2626 ();
 sg13g2_decap_8 FILLER_65_2633 ();
 sg13g2_decap_8 FILLER_65_2640 ();
 sg13g2_decap_8 FILLER_65_2647 ();
 sg13g2_decap_8 FILLER_65_2654 ();
 sg13g2_decap_8 FILLER_65_2661 ();
 sg13g2_decap_4 FILLER_65_2668 ();
 sg13g2_fill_2 FILLER_65_2672 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_252 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_8 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_decap_8 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_308 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_decap_8 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_decap_8 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_350 ();
 sg13g2_decap_4 FILLER_66_357 ();
 sg13g2_fill_1 FILLER_66_361 ();
 sg13g2_decap_4 FILLER_66_388 ();
 sg13g2_fill_1 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_419 ();
 sg13g2_decap_4 FILLER_66_452 ();
 sg13g2_fill_1 FILLER_66_456 ();
 sg13g2_decap_8 FILLER_66_496 ();
 sg13g2_fill_1 FILLER_66_503 ();
 sg13g2_fill_2 FILLER_66_566 ();
 sg13g2_fill_2 FILLER_66_587 ();
 sg13g2_fill_1 FILLER_66_589 ();
 sg13g2_fill_2 FILLER_66_616 ();
 sg13g2_fill_2 FILLER_66_622 ();
 sg13g2_fill_2 FILLER_66_671 ();
 sg13g2_fill_1 FILLER_66_673 ();
 sg13g2_fill_2 FILLER_66_721 ();
 sg13g2_fill_1 FILLER_66_723 ();
 sg13g2_decap_8 FILLER_66_739 ();
 sg13g2_fill_1 FILLER_66_746 ();
 sg13g2_decap_8 FILLER_66_816 ();
 sg13g2_decap_8 FILLER_66_823 ();
 sg13g2_decap_8 FILLER_66_834 ();
 sg13g2_decap_4 FILLER_66_841 ();
 sg13g2_fill_2 FILLER_66_854 ();
 sg13g2_fill_2 FILLER_66_876 ();
 sg13g2_fill_1 FILLER_66_878 ();
 sg13g2_fill_2 FILLER_66_884 ();
 sg13g2_fill_1 FILLER_66_886 ();
 sg13g2_fill_2 FILLER_66_901 ();
 sg13g2_fill_2 FILLER_66_908 ();
 sg13g2_decap_4 FILLER_66_914 ();
 sg13g2_fill_1 FILLER_66_944 ();
 sg13g2_fill_1 FILLER_66_950 ();
 sg13g2_decap_8 FILLER_66_980 ();
 sg13g2_fill_2 FILLER_66_987 ();
 sg13g2_fill_1 FILLER_66_989 ();
 sg13g2_fill_2 FILLER_66_998 ();
 sg13g2_fill_1 FILLER_66_1018 ();
 sg13g2_fill_1 FILLER_66_1028 ();
 sg13g2_fill_1 FILLER_66_1034 ();
 sg13g2_fill_2 FILLER_66_1038 ();
 sg13g2_fill_1 FILLER_66_1040 ();
 sg13g2_fill_2 FILLER_66_1093 ();
 sg13g2_fill_1 FILLER_66_1130 ();
 sg13g2_fill_2 FILLER_66_1140 ();
 sg13g2_fill_1 FILLER_66_1173 ();
 sg13g2_fill_1 FILLER_66_1201 ();
 sg13g2_decap_8 FILLER_66_1247 ();
 sg13g2_fill_2 FILLER_66_1254 ();
 sg13g2_decap_4 FILLER_66_1260 ();
 sg13g2_decap_8 FILLER_66_1272 ();
 sg13g2_fill_2 FILLER_66_1279 ();
 sg13g2_fill_1 FILLER_66_1281 ();
 sg13g2_fill_2 FILLER_66_1286 ();
 sg13g2_fill_2 FILLER_66_1293 ();
 sg13g2_fill_2 FILLER_66_1304 ();
 sg13g2_fill_1 FILLER_66_1315 ();
 sg13g2_fill_2 FILLER_66_1330 ();
 sg13g2_fill_2 FILLER_66_1394 ();
 sg13g2_fill_1 FILLER_66_1422 ();
 sg13g2_decap_4 FILLER_66_1461 ();
 sg13g2_decap_8 FILLER_66_1497 ();
 sg13g2_fill_2 FILLER_66_1517 ();
 sg13g2_fill_2 FILLER_66_1553 ();
 sg13g2_fill_1 FILLER_66_1555 ();
 sg13g2_fill_1 FILLER_66_1601 ();
 sg13g2_fill_2 FILLER_66_1611 ();
 sg13g2_fill_2 FILLER_66_1676 ();
 sg13g2_fill_1 FILLER_66_1699 ();
 sg13g2_fill_1 FILLER_66_1704 ();
 sg13g2_fill_2 FILLER_66_1713 ();
 sg13g2_fill_2 FILLER_66_1756 ();
 sg13g2_decap_8 FILLER_66_1793 ();
 sg13g2_fill_1 FILLER_66_1800 ();
 sg13g2_fill_2 FILLER_66_1823 ();
 sg13g2_decap_8 FILLER_66_1839 ();
 sg13g2_decap_8 FILLER_66_1846 ();
 sg13g2_fill_2 FILLER_66_1865 ();
 sg13g2_fill_1 FILLER_66_1867 ();
 sg13g2_fill_1 FILLER_66_1903 ();
 sg13g2_fill_1 FILLER_66_1973 ();
 sg13g2_fill_1 FILLER_66_2021 ();
 sg13g2_decap_4 FILLER_66_2067 ();
 sg13g2_fill_1 FILLER_66_2071 ();
 sg13g2_fill_2 FILLER_66_2112 ();
 sg13g2_fill_1 FILLER_66_2114 ();
 sg13g2_fill_2 FILLER_66_2141 ();
 sg13g2_decap_8 FILLER_66_2147 ();
 sg13g2_decap_8 FILLER_66_2154 ();
 sg13g2_fill_1 FILLER_66_2161 ();
 sg13g2_fill_1 FILLER_66_2172 ();
 sg13g2_fill_2 FILLER_66_2189 ();
 sg13g2_fill_1 FILLER_66_2200 ();
 sg13g2_fill_2 FILLER_66_2227 ();
 sg13g2_fill_1 FILLER_66_2229 ();
 sg13g2_fill_2 FILLER_66_2245 ();
 sg13g2_fill_1 FILLER_66_2247 ();
 sg13g2_fill_2 FILLER_66_2256 ();
 sg13g2_fill_1 FILLER_66_2258 ();
 sg13g2_decap_8 FILLER_66_2285 ();
 sg13g2_fill_2 FILLER_66_2292 ();
 sg13g2_fill_2 FILLER_66_2339 ();
 sg13g2_fill_2 FILLER_66_2389 ();
 sg13g2_fill_1 FILLER_66_2478 ();
 sg13g2_fill_2 FILLER_66_2523 ();
 sg13g2_fill_1 FILLER_66_2550 ();
 sg13g2_fill_1 FILLER_66_2559 ();
 sg13g2_decap_8 FILLER_66_2606 ();
 sg13g2_decap_8 FILLER_66_2613 ();
 sg13g2_decap_8 FILLER_66_2620 ();
 sg13g2_decap_8 FILLER_66_2627 ();
 sg13g2_decap_8 FILLER_66_2634 ();
 sg13g2_decap_8 FILLER_66_2641 ();
 sg13g2_decap_8 FILLER_66_2648 ();
 sg13g2_decap_8 FILLER_66_2655 ();
 sg13g2_decap_8 FILLER_66_2662 ();
 sg13g2_decap_4 FILLER_66_2669 ();
 sg13g2_fill_1 FILLER_66_2673 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_decap_8 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_decap_8 FILLER_67_308 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_decap_8 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_350 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_fill_1 FILLER_67_372 ();
 sg13g2_fill_2 FILLER_67_377 ();
 sg13g2_fill_1 FILLER_67_379 ();
 sg13g2_decap_4 FILLER_67_393 ();
 sg13g2_fill_1 FILLER_67_397 ();
 sg13g2_decap_4 FILLER_67_450 ();
 sg13g2_fill_2 FILLER_67_556 ();
 sg13g2_fill_2 FILLER_67_583 ();
 sg13g2_fill_1 FILLER_67_630 ();
 sg13g2_fill_2 FILLER_67_678 ();
 sg13g2_fill_1 FILLER_67_685 ();
 sg13g2_fill_2 FILLER_67_711 ();
 sg13g2_fill_1 FILLER_67_713 ();
 sg13g2_fill_2 FILLER_67_769 ();
 sg13g2_fill_2 FILLER_67_878 ();
 sg13g2_decap_8 FILLER_67_920 ();
 sg13g2_fill_2 FILLER_67_949 ();
 sg13g2_fill_2 FILLER_67_991 ();
 sg13g2_fill_2 FILLER_67_1068 ();
 sg13g2_fill_1 FILLER_67_1088 ();
 sg13g2_fill_1 FILLER_67_1097 ();
 sg13g2_fill_1 FILLER_67_1120 ();
 sg13g2_fill_1 FILLER_67_1126 ();
 sg13g2_fill_2 FILLER_67_1193 ();
 sg13g2_fill_1 FILLER_67_1195 ();
 sg13g2_fill_2 FILLER_67_1200 ();
 sg13g2_decap_4 FILLER_67_1210 ();
 sg13g2_fill_2 FILLER_67_1230 ();
 sg13g2_fill_2 FILLER_67_1246 ();
 sg13g2_fill_2 FILLER_67_1279 ();
 sg13g2_fill_1 FILLER_67_1281 ();
 sg13g2_fill_2 FILLER_67_1326 ();
 sg13g2_fill_1 FILLER_67_1342 ();
 sg13g2_fill_1 FILLER_67_1349 ();
 sg13g2_decap_4 FILLER_67_1355 ();
 sg13g2_fill_1 FILLER_67_1388 ();
 sg13g2_fill_2 FILLER_67_1402 ();
 sg13g2_fill_1 FILLER_67_1404 ();
 sg13g2_fill_1 FILLER_67_1448 ();
 sg13g2_fill_1 FILLER_67_1459 ();
 sg13g2_decap_4 FILLER_67_1465 ();
 sg13g2_fill_2 FILLER_67_1469 ();
 sg13g2_fill_2 FILLER_67_1474 ();
 sg13g2_decap_8 FILLER_67_1489 ();
 sg13g2_decap_4 FILLER_67_1504 ();
 sg13g2_decap_4 FILLER_67_1511 ();
 sg13g2_fill_1 FILLER_67_1550 ();
 sg13g2_fill_2 FILLER_67_1656 ();
 sg13g2_fill_1 FILLER_67_1670 ();
 sg13g2_decap_8 FILLER_67_1690 ();
 sg13g2_fill_2 FILLER_67_1720 ();
 sg13g2_fill_1 FILLER_67_1734 ();
 sg13g2_fill_2 FILLER_67_1779 ();
 sg13g2_fill_1 FILLER_67_1793 ();
 sg13g2_fill_2 FILLER_67_1802 ();
 sg13g2_fill_2 FILLER_67_1810 ();
 sg13g2_decap_8 FILLER_67_1845 ();
 sg13g2_fill_2 FILLER_67_1852 ();
 sg13g2_fill_1 FILLER_67_1894 ();
 sg13g2_fill_2 FILLER_67_1973 ();
 sg13g2_fill_2 FILLER_67_2001 ();
 sg13g2_fill_1 FILLER_67_2003 ();
 sg13g2_fill_2 FILLER_67_2030 ();
 sg13g2_fill_1 FILLER_67_2032 ();
 sg13g2_decap_8 FILLER_67_2064 ();
 sg13g2_fill_2 FILLER_67_2097 ();
 sg13g2_fill_1 FILLER_67_2099 ();
 sg13g2_fill_2 FILLER_67_2182 ();
 sg13g2_fill_1 FILLER_67_2184 ();
 sg13g2_fill_2 FILLER_67_2211 ();
 sg13g2_fill_2 FILLER_67_2227 ();
 sg13g2_fill_1 FILLER_67_2229 ();
 sg13g2_decap_4 FILLER_67_2293 ();
 sg13g2_fill_1 FILLER_67_2297 ();
 sg13g2_decap_4 FILLER_67_2345 ();
 sg13g2_fill_1 FILLER_67_2362 ();
 sg13g2_fill_1 FILLER_67_2376 ();
 sg13g2_fill_1 FILLER_67_2442 ();
 sg13g2_fill_1 FILLER_67_2467 ();
 sg13g2_decap_8 FILLER_67_2498 ();
 sg13g2_fill_1 FILLER_67_2505 ();
 sg13g2_fill_1 FILLER_67_2545 ();
 sg13g2_fill_2 FILLER_67_2555 ();
 sg13g2_fill_1 FILLER_67_2557 ();
 sg13g2_fill_2 FILLER_67_2563 ();
 sg13g2_fill_1 FILLER_67_2565 ();
 sg13g2_fill_1 FILLER_67_2571 ();
 sg13g2_decap_8 FILLER_67_2598 ();
 sg13g2_decap_8 FILLER_67_2605 ();
 sg13g2_decap_8 FILLER_67_2612 ();
 sg13g2_decap_8 FILLER_67_2619 ();
 sg13g2_decap_8 FILLER_67_2626 ();
 sg13g2_decap_8 FILLER_67_2633 ();
 sg13g2_decap_8 FILLER_67_2640 ();
 sg13g2_decap_8 FILLER_67_2647 ();
 sg13g2_decap_8 FILLER_67_2654 ();
 sg13g2_decap_8 FILLER_67_2661 ();
 sg13g2_decap_4 FILLER_67_2668 ();
 sg13g2_fill_2 FILLER_67_2672 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_decap_8 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_decap_8 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_252 ();
 sg13g2_decap_8 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_280 ();
 sg13g2_decap_8 FILLER_68_287 ();
 sg13g2_decap_8 FILLER_68_294 ();
 sg13g2_decap_8 FILLER_68_301 ();
 sg13g2_decap_8 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_315 ();
 sg13g2_decap_8 FILLER_68_322 ();
 sg13g2_decap_8 FILLER_68_329 ();
 sg13g2_decap_8 FILLER_68_336 ();
 sg13g2_decap_8 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_350 ();
 sg13g2_decap_8 FILLER_68_357 ();
 sg13g2_decap_4 FILLER_68_364 ();
 sg13g2_fill_1 FILLER_68_368 ();
 sg13g2_fill_2 FILLER_68_395 ();
 sg13g2_decap_4 FILLER_68_423 ();
 sg13g2_fill_2 FILLER_68_427 ();
 sg13g2_decap_8 FILLER_68_449 ();
 sg13g2_decap_8 FILLER_68_456 ();
 sg13g2_fill_2 FILLER_68_499 ();
 sg13g2_decap_4 FILLER_68_527 ();
 sg13g2_decap_8 FILLER_68_541 ();
 sg13g2_decap_8 FILLER_68_548 ();
 sg13g2_fill_1 FILLER_68_555 ();
 sg13g2_fill_2 FILLER_68_623 ();
 sg13g2_fill_1 FILLER_68_625 ();
 sg13g2_fill_1 FILLER_68_666 ();
 sg13g2_fill_2 FILLER_68_676 ();
 sg13g2_fill_2 FILLER_68_686 ();
 sg13g2_fill_1 FILLER_68_688 ();
 sg13g2_fill_2 FILLER_68_720 ();
 sg13g2_fill_1 FILLER_68_722 ();
 sg13g2_fill_2 FILLER_68_735 ();
 sg13g2_fill_1 FILLER_68_751 ();
 sg13g2_fill_2 FILLER_68_757 ();
 sg13g2_fill_1 FILLER_68_768 ();
 sg13g2_fill_2 FILLER_68_782 ();
 sg13g2_fill_1 FILLER_68_784 ();
 sg13g2_fill_1 FILLER_68_868 ();
 sg13g2_fill_1 FILLER_68_910 ();
 sg13g2_fill_2 FILLER_68_934 ();
 sg13g2_fill_1 FILLER_68_936 ();
 sg13g2_fill_2 FILLER_68_1020 ();
 sg13g2_fill_2 FILLER_68_1027 ();
 sg13g2_fill_2 FILLER_68_1039 ();
 sg13g2_fill_1 FILLER_68_1049 ();
 sg13g2_fill_1 FILLER_68_1088 ();
 sg13g2_fill_2 FILLER_68_1096 ();
 sg13g2_decap_8 FILLER_68_1179 ();
 sg13g2_fill_1 FILLER_68_1186 ();
 sg13g2_fill_2 FILLER_68_1200 ();
 sg13g2_fill_1 FILLER_68_1250 ();
 sg13g2_fill_2 FILLER_68_1287 ();
 sg13g2_fill_1 FILLER_68_1289 ();
 sg13g2_fill_1 FILLER_68_1307 ();
 sg13g2_fill_1 FILLER_68_1352 ();
 sg13g2_fill_2 FILLER_68_1362 ();
 sg13g2_fill_2 FILLER_68_1376 ();
 sg13g2_fill_1 FILLER_68_1391 ();
 sg13g2_decap_8 FILLER_68_1407 ();
 sg13g2_fill_2 FILLER_68_1414 ();
 sg13g2_fill_2 FILLER_68_1420 ();
 sg13g2_fill_2 FILLER_68_1468 ();
 sg13g2_decap_8 FILLER_68_1515 ();
 sg13g2_fill_1 FILLER_68_1522 ();
 sg13g2_fill_2 FILLER_68_1528 ();
 sg13g2_fill_1 FILLER_68_1530 ();
 sg13g2_fill_2 FILLER_68_1542 ();
 sg13g2_fill_2 FILLER_68_1563 ();
 sg13g2_fill_1 FILLER_68_1565 ();
 sg13g2_fill_2 FILLER_68_1688 ();
 sg13g2_fill_2 FILLER_68_1773 ();
 sg13g2_decap_4 FILLER_68_1779 ();
 sg13g2_fill_1 FILLER_68_1783 ();
 sg13g2_fill_1 FILLER_68_1821 ();
 sg13g2_fill_1 FILLER_68_1848 ();
 sg13g2_fill_1 FILLER_68_1881 ();
 sg13g2_fill_1 FILLER_68_1920 ();
 sg13g2_fill_1 FILLER_68_1931 ();
 sg13g2_fill_1 FILLER_68_1984 ();
 sg13g2_decap_8 FILLER_68_2067 ();
 sg13g2_fill_2 FILLER_68_2074 ();
 sg13g2_fill_2 FILLER_68_2092 ();
 sg13g2_fill_1 FILLER_68_2094 ();
 sg13g2_decap_8 FILLER_68_2134 ();
 sg13g2_decap_4 FILLER_68_2141 ();
 sg13g2_fill_1 FILLER_68_2253 ();
 sg13g2_fill_1 FILLER_68_2340 ();
 sg13g2_decap_4 FILLER_68_2381 ();
 sg13g2_fill_2 FILLER_68_2415 ();
 sg13g2_fill_1 FILLER_68_2430 ();
 sg13g2_fill_1 FILLER_68_2444 ();
 sg13g2_fill_2 FILLER_68_2465 ();
 sg13g2_fill_1 FILLER_68_2505 ();
 sg13g2_fill_2 FILLER_68_2537 ();
 sg13g2_fill_1 FILLER_68_2539 ();
 sg13g2_decap_8 FILLER_68_2604 ();
 sg13g2_decap_8 FILLER_68_2611 ();
 sg13g2_decap_8 FILLER_68_2618 ();
 sg13g2_decap_8 FILLER_68_2625 ();
 sg13g2_decap_8 FILLER_68_2632 ();
 sg13g2_decap_8 FILLER_68_2639 ();
 sg13g2_decap_8 FILLER_68_2646 ();
 sg13g2_decap_8 FILLER_68_2653 ();
 sg13g2_decap_8 FILLER_68_2660 ();
 sg13g2_decap_8 FILLER_68_2667 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_decap_8 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_182 ();
 sg13g2_decap_8 FILLER_69_189 ();
 sg13g2_decap_8 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_203 ();
 sg13g2_decap_8 FILLER_69_210 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_decap_8 FILLER_69_238 ();
 sg13g2_decap_8 FILLER_69_245 ();
 sg13g2_decap_8 FILLER_69_252 ();
 sg13g2_decap_8 FILLER_69_259 ();
 sg13g2_decap_8 FILLER_69_266 ();
 sg13g2_decap_8 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_decap_8 FILLER_69_301 ();
 sg13g2_decap_8 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_315 ();
 sg13g2_decap_8 FILLER_69_322 ();
 sg13g2_decap_8 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_336 ();
 sg13g2_decap_8 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_350 ();
 sg13g2_decap_8 FILLER_69_357 ();
 sg13g2_decap_8 FILLER_69_364 ();
 sg13g2_fill_2 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_decap_4 FILLER_69_406 ();
 sg13g2_fill_2 FILLER_69_410 ();
 sg13g2_fill_2 FILLER_69_443 ();
 sg13g2_fill_1 FILLER_69_445 ();
 sg13g2_decap_8 FILLER_69_451 ();
 sg13g2_fill_1 FILLER_69_458 ();
 sg13g2_fill_2 FILLER_69_501 ();
 sg13g2_decap_4 FILLER_69_555 ();
 sg13g2_fill_2 FILLER_69_559 ();
 sg13g2_fill_1 FILLER_69_592 ();
 sg13g2_fill_2 FILLER_69_665 ();
 sg13g2_fill_1 FILLER_69_667 ();
 sg13g2_fill_1 FILLER_69_694 ();
 sg13g2_fill_2 FILLER_69_699 ();
 sg13g2_fill_1 FILLER_69_701 ();
 sg13g2_fill_2 FILLER_69_762 ();
 sg13g2_fill_1 FILLER_69_764 ();
 sg13g2_fill_1 FILLER_69_779 ();
 sg13g2_fill_1 FILLER_69_850 ();
 sg13g2_fill_1 FILLER_69_894 ();
 sg13g2_fill_2 FILLER_69_961 ();
 sg13g2_fill_1 FILLER_69_963 ();
 sg13g2_fill_2 FILLER_69_1037 ();
 sg13g2_fill_1 FILLER_69_1039 ();
 sg13g2_fill_1 FILLER_69_1050 ();
 sg13g2_fill_2 FILLER_69_1115 ();
 sg13g2_decap_4 FILLER_69_1135 ();
 sg13g2_decap_4 FILLER_69_1164 ();
 sg13g2_fill_1 FILLER_69_1168 ();
 sg13g2_decap_8 FILLER_69_1173 ();
 sg13g2_fill_2 FILLER_69_1180 ();
 sg13g2_fill_2 FILLER_69_1217 ();
 sg13g2_fill_1 FILLER_69_1219 ();
 sg13g2_fill_2 FILLER_69_1230 ();
 sg13g2_fill_1 FILLER_69_1232 ();
 sg13g2_fill_1 FILLER_69_1246 ();
 sg13g2_fill_1 FILLER_69_1262 ();
 sg13g2_fill_2 FILLER_69_1272 ();
 sg13g2_fill_1 FILLER_69_1274 ();
 sg13g2_fill_1 FILLER_69_1402 ();
 sg13g2_fill_1 FILLER_69_1494 ();
 sg13g2_fill_2 FILLER_69_1511 ();
 sg13g2_fill_2 FILLER_69_1535 ();
 sg13g2_fill_1 FILLER_69_1541 ();
 sg13g2_fill_2 FILLER_69_1547 ();
 sg13g2_fill_1 FILLER_69_1573 ();
 sg13g2_fill_2 FILLER_69_1601 ();
 sg13g2_fill_1 FILLER_69_1603 ();
 sg13g2_fill_2 FILLER_69_1705 ();
 sg13g2_fill_1 FILLER_69_1728 ();
 sg13g2_fill_1 FILLER_69_1739 ();
 sg13g2_fill_2 FILLER_69_1761 ();
 sg13g2_fill_2 FILLER_69_1775 ();
 sg13g2_fill_1 FILLER_69_1777 ();
 sg13g2_decap_4 FILLER_69_1818 ();
 sg13g2_decap_4 FILLER_69_1865 ();
 sg13g2_fill_2 FILLER_69_1891 ();
 sg13g2_fill_1 FILLER_69_1893 ();
 sg13g2_fill_2 FILLER_69_1907 ();
 sg13g2_fill_1 FILLER_69_1945 ();
 sg13g2_fill_2 FILLER_69_2014 ();
 sg13g2_fill_1 FILLER_69_2016 ();
 sg13g2_fill_2 FILLER_69_2043 ();
 sg13g2_fill_1 FILLER_69_2045 ();
 sg13g2_fill_2 FILLER_69_2080 ();
 sg13g2_fill_2 FILLER_69_2090 ();
 sg13g2_fill_2 FILLER_69_2096 ();
 sg13g2_fill_1 FILLER_69_2098 ();
 sg13g2_fill_1 FILLER_69_2107 ();
 sg13g2_fill_2 FILLER_69_2116 ();
 sg13g2_fill_1 FILLER_69_2227 ();
 sg13g2_fill_1 FILLER_69_2250 ();
 sg13g2_fill_1 FILLER_69_2303 ();
 sg13g2_fill_1 FILLER_69_2334 ();
 sg13g2_fill_2 FILLER_69_2356 ();
 sg13g2_decap_8 FILLER_69_2414 ();
 sg13g2_decap_4 FILLER_69_2421 ();
 sg13g2_fill_2 FILLER_69_2425 ();
 sg13g2_fill_1 FILLER_69_2437 ();
 sg13g2_fill_1 FILLER_69_2443 ();
 sg13g2_fill_1 FILLER_69_2475 ();
 sg13g2_decap_8 FILLER_69_2611 ();
 sg13g2_decap_8 FILLER_69_2618 ();
 sg13g2_decap_8 FILLER_69_2625 ();
 sg13g2_decap_8 FILLER_69_2632 ();
 sg13g2_decap_8 FILLER_69_2639 ();
 sg13g2_decap_8 FILLER_69_2646 ();
 sg13g2_decap_8 FILLER_69_2653 ();
 sg13g2_decap_8 FILLER_69_2660 ();
 sg13g2_decap_8 FILLER_69_2667 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_203 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_decap_8 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_266 ();
 sg13g2_decap_8 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_280 ();
 sg13g2_decap_8 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_301 ();
 sg13g2_decap_8 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_4 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_393 ();
 sg13g2_decap_8 FILLER_70_400 ();
 sg13g2_decap_8 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_70_414 ();
 sg13g2_fill_2 FILLER_70_421 ();
 sg13g2_fill_2 FILLER_70_453 ();
 sg13g2_fill_1 FILLER_70_455 ();
 sg13g2_decap_4 FILLER_70_460 ();
 sg13g2_fill_1 FILLER_70_464 ();
 sg13g2_decap_8 FILLER_70_496 ();
 sg13g2_decap_8 FILLER_70_503 ();
 sg13g2_decap_8 FILLER_70_510 ();
 sg13g2_fill_2 FILLER_70_517 ();
 sg13g2_fill_1 FILLER_70_519 ();
 sg13g2_decap_8 FILLER_70_540 ();
 sg13g2_decap_8 FILLER_70_547 ();
 sg13g2_decap_8 FILLER_70_554 ();
 sg13g2_fill_1 FILLER_70_561 ();
 sg13g2_fill_2 FILLER_70_579 ();
 sg13g2_fill_1 FILLER_70_581 ();
 sg13g2_fill_1 FILLER_70_613 ();
 sg13g2_fill_1 FILLER_70_628 ();
 sg13g2_fill_2 FILLER_70_634 ();
 sg13g2_fill_2 FILLER_70_656 ();
 sg13g2_fill_1 FILLER_70_658 ();
 sg13g2_fill_1 FILLER_70_695 ();
 sg13g2_fill_2 FILLER_70_709 ();
 sg13g2_fill_1 FILLER_70_743 ();
 sg13g2_fill_1 FILLER_70_757 ();
 sg13g2_fill_2 FILLER_70_839 ();
 sg13g2_fill_1 FILLER_70_873 ();
 sg13g2_fill_2 FILLER_70_884 ();
 sg13g2_fill_1 FILLER_70_891 ();
 sg13g2_fill_2 FILLER_70_900 ();
 sg13g2_fill_1 FILLER_70_902 ();
 sg13g2_fill_2 FILLER_70_933 ();
 sg13g2_fill_1 FILLER_70_949 ();
 sg13g2_fill_1 FILLER_70_964 ();
 sg13g2_fill_1 FILLER_70_986 ();
 sg13g2_fill_1 FILLER_70_1008 ();
 sg13g2_fill_1 FILLER_70_1023 ();
 sg13g2_fill_2 FILLER_70_1082 ();
 sg13g2_fill_1 FILLER_70_1095 ();
 sg13g2_decap_8 FILLER_70_1143 ();
 sg13g2_decap_8 FILLER_70_1150 ();
 sg13g2_fill_2 FILLER_70_1157 ();
 sg13g2_fill_2 FILLER_70_1173 ();
 sg13g2_fill_1 FILLER_70_1192 ();
 sg13g2_fill_1 FILLER_70_1203 ();
 sg13g2_fill_1 FILLER_70_1209 ();
 sg13g2_fill_2 FILLER_70_1223 ();
 sg13g2_fill_1 FILLER_70_1225 ();
 sg13g2_fill_1 FILLER_70_1252 ();
 sg13g2_fill_2 FILLER_70_1269 ();
 sg13g2_fill_1 FILLER_70_1271 ();
 sg13g2_fill_2 FILLER_70_1283 ();
 sg13g2_fill_1 FILLER_70_1285 ();
 sg13g2_fill_1 FILLER_70_1290 ();
 sg13g2_fill_2 FILLER_70_1323 ();
 sg13g2_fill_1 FILLER_70_1371 ();
 sg13g2_fill_1 FILLER_70_1378 ();
 sg13g2_fill_2 FILLER_70_1414 ();
 sg13g2_fill_1 FILLER_70_1416 ();
 sg13g2_fill_2 FILLER_70_1443 ();
 sg13g2_fill_2 FILLER_70_1480 ();
 sg13g2_fill_1 FILLER_70_1562 ();
 sg13g2_fill_2 FILLER_70_1576 ();
 sg13g2_fill_2 FILLER_70_1583 ();
 sg13g2_fill_1 FILLER_70_1585 ();
 sg13g2_decap_8 FILLER_70_1603 ();
 sg13g2_decap_4 FILLER_70_1610 ();
 sg13g2_fill_2 FILLER_70_1632 ();
 sg13g2_fill_1 FILLER_70_1634 ();
 sg13g2_fill_2 FILLER_70_1656 ();
 sg13g2_fill_1 FILLER_70_1667 ();
 sg13g2_fill_2 FILLER_70_1682 ();
 sg13g2_fill_2 FILLER_70_1693 ();
 sg13g2_fill_1 FILLER_70_1730 ();
 sg13g2_fill_1 FILLER_70_1771 ();
 sg13g2_fill_2 FILLER_70_1822 ();
 sg13g2_fill_1 FILLER_70_1824 ();
 sg13g2_fill_2 FILLER_70_1858 ();
 sg13g2_fill_2 FILLER_70_1864 ();
 sg13g2_fill_1 FILLER_70_1874 ();
 sg13g2_fill_1 FILLER_70_1889 ();
 sg13g2_fill_1 FILLER_70_1924 ();
 sg13g2_fill_2 FILLER_70_1994 ();
 sg13g2_fill_1 FILLER_70_1996 ();
 sg13g2_fill_2 FILLER_70_2016 ();
 sg13g2_fill_1 FILLER_70_2048 ();
 sg13g2_fill_1 FILLER_70_2061 ();
 sg13g2_decap_4 FILLER_70_2092 ();
 sg13g2_fill_1 FILLER_70_2096 ();
 sg13g2_decap_4 FILLER_70_2102 ();
 sg13g2_fill_2 FILLER_70_2106 ();
 sg13g2_fill_2 FILLER_70_2155 ();
 sg13g2_fill_1 FILLER_70_2157 ();
 sg13g2_fill_1 FILLER_70_2162 ();
 sg13g2_fill_1 FILLER_70_2168 ();
 sg13g2_fill_1 FILLER_70_2205 ();
 sg13g2_fill_1 FILLER_70_2215 ();
 sg13g2_fill_2 FILLER_70_2260 ();
 sg13g2_fill_1 FILLER_70_2297 ();
 sg13g2_fill_2 FILLER_70_2311 ();
 sg13g2_fill_2 FILLER_70_2348 ();
 sg13g2_fill_2 FILLER_70_2380 ();
 sg13g2_fill_1 FILLER_70_2458 ();
 sg13g2_fill_1 FILLER_70_2468 ();
 sg13g2_fill_2 FILLER_70_2508 ();
 sg13g2_fill_2 FILLER_70_2568 ();
 sg13g2_fill_2 FILLER_70_2584 ();
 sg13g2_decap_8 FILLER_70_2616 ();
 sg13g2_decap_8 FILLER_70_2623 ();
 sg13g2_decap_8 FILLER_70_2630 ();
 sg13g2_decap_8 FILLER_70_2637 ();
 sg13g2_decap_8 FILLER_70_2644 ();
 sg13g2_decap_8 FILLER_70_2651 ();
 sg13g2_decap_8 FILLER_70_2658 ();
 sg13g2_decap_8 FILLER_70_2665 ();
 sg13g2_fill_2 FILLER_70_2672 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_245 ();
 sg13g2_decap_8 FILLER_71_252 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_315 ();
 sg13g2_decap_8 FILLER_71_322 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_decap_8 FILLER_71_350 ();
 sg13g2_decap_4 FILLER_71_357 ();
 sg13g2_fill_2 FILLER_71_361 ();
 sg13g2_fill_2 FILLER_71_377 ();
 sg13g2_fill_2 FILLER_71_400 ();
 sg13g2_decap_8 FILLER_71_454 ();
 sg13g2_fill_2 FILLER_71_461 ();
 sg13g2_decap_4 FILLER_71_468 ();
 sg13g2_fill_2 FILLER_71_472 ();
 sg13g2_fill_1 FILLER_71_478 ();
 sg13g2_decap_8 FILLER_71_487 ();
 sg13g2_decap_8 FILLER_71_494 ();
 sg13g2_decap_8 FILLER_71_501 ();
 sg13g2_fill_2 FILLER_71_508 ();
 sg13g2_fill_2 FILLER_71_531 ();
 sg13g2_decap_4 FILLER_71_559 ();
 sg13g2_fill_2 FILLER_71_563 ();
 sg13g2_fill_2 FILLER_71_611 ();
 sg13g2_fill_2 FILLER_71_619 ();
 sg13g2_fill_1 FILLER_71_621 ();
 sg13g2_fill_2 FILLER_71_659 ();
 sg13g2_fill_2 FILLER_71_700 ();
 sg13g2_fill_2 FILLER_71_736 ();
 sg13g2_fill_1 FILLER_71_738 ();
 sg13g2_fill_1 FILLER_71_748 ();
 sg13g2_fill_2 FILLER_71_754 ();
 sg13g2_fill_2 FILLER_71_856 ();
 sg13g2_fill_1 FILLER_71_873 ();
 sg13g2_fill_1 FILLER_71_879 ();
 sg13g2_fill_2 FILLER_71_929 ();
 sg13g2_fill_1 FILLER_71_931 ();
 sg13g2_fill_2 FILLER_71_990 ();
 sg13g2_fill_1 FILLER_71_992 ();
 sg13g2_fill_2 FILLER_71_1019 ();
 sg13g2_fill_2 FILLER_71_1030 ();
 sg13g2_fill_2 FILLER_71_1058 ();
 sg13g2_fill_1 FILLER_71_1069 ();
 sg13g2_fill_2 FILLER_71_1105 ();
 sg13g2_fill_1 FILLER_71_1113 ();
 sg13g2_fill_2 FILLER_71_1128 ();
 sg13g2_fill_1 FILLER_71_1148 ();
 sg13g2_fill_2 FILLER_71_1180 ();
 sg13g2_fill_1 FILLER_71_1182 ();
 sg13g2_fill_2 FILLER_71_1234 ();
 sg13g2_fill_1 FILLER_71_1236 ();
 sg13g2_fill_1 FILLER_71_1289 ();
 sg13g2_fill_1 FILLER_71_1338 ();
 sg13g2_fill_2 FILLER_71_1353 ();
 sg13g2_fill_1 FILLER_71_1355 ();
 sg13g2_fill_1 FILLER_71_1423 ();
 sg13g2_fill_2 FILLER_71_1447 ();
 sg13g2_fill_2 FILLER_71_1476 ();
 sg13g2_fill_1 FILLER_71_1484 ();
 sg13g2_fill_2 FILLER_71_1488 ();
 sg13g2_fill_1 FILLER_71_1490 ();
 sg13g2_fill_1 FILLER_71_1503 ();
 sg13g2_fill_1 FILLER_71_1530 ();
 sg13g2_fill_1 FILLER_71_1581 ();
 sg13g2_decap_8 FILLER_71_1610 ();
 sg13g2_fill_2 FILLER_71_1617 ();
 sg13g2_fill_1 FILLER_71_1636 ();
 sg13g2_fill_2 FILLER_71_1648 ();
 sg13g2_fill_2 FILLER_71_1655 ();
 sg13g2_decap_8 FILLER_71_1694 ();
 sg13g2_fill_2 FILLER_71_1701 ();
 sg13g2_fill_1 FILLER_71_1703 ();
 sg13g2_fill_1 FILLER_71_1729 ();
 sg13g2_fill_1 FILLER_71_1745 ();
 sg13g2_decap_8 FILLER_71_1784 ();
 sg13g2_fill_2 FILLER_71_1803 ();
 sg13g2_decap_8 FILLER_71_1852 ();
 sg13g2_fill_2 FILLER_71_1867 ();
 sg13g2_fill_2 FILLER_71_1872 ();
 sg13g2_fill_2 FILLER_71_1905 ();
 sg13g2_fill_2 FILLER_71_1939 ();
 sg13g2_fill_1 FILLER_71_1994 ();
 sg13g2_fill_2 FILLER_71_2021 ();
 sg13g2_fill_2 FILLER_71_2058 ();
 sg13g2_fill_1 FILLER_71_2060 ();
 sg13g2_fill_1 FILLER_71_2087 ();
 sg13g2_fill_1 FILLER_71_2162 ();
 sg13g2_fill_2 FILLER_71_2171 ();
 sg13g2_fill_1 FILLER_71_2173 ();
 sg13g2_decap_4 FILLER_71_2182 ();
 sg13g2_decap_4 FILLER_71_2190 ();
 sg13g2_fill_2 FILLER_71_2227 ();
 sg13g2_fill_1 FILLER_71_2229 ();
 sg13g2_fill_1 FILLER_71_2239 ();
 sg13g2_fill_2 FILLER_71_2245 ();
 sg13g2_fill_1 FILLER_71_2247 ();
 sg13g2_fill_2 FILLER_71_2277 ();
 sg13g2_fill_1 FILLER_71_2279 ();
 sg13g2_fill_2 FILLER_71_2306 ();
 sg13g2_fill_1 FILLER_71_2308 ();
 sg13g2_fill_2 FILLER_71_2353 ();
 sg13g2_fill_2 FILLER_71_2377 ();
 sg13g2_fill_2 FILLER_71_2502 ();
 sg13g2_fill_2 FILLER_71_2517 ();
 sg13g2_fill_1 FILLER_71_2519 ();
 sg13g2_fill_2 FILLER_71_2541 ();
 sg13g2_fill_1 FILLER_71_2543 ();
 sg13g2_fill_2 FILLER_71_2553 ();
 sg13g2_fill_1 FILLER_71_2559 ();
 sg13g2_decap_8 FILLER_71_2611 ();
 sg13g2_decap_8 FILLER_71_2618 ();
 sg13g2_decap_8 FILLER_71_2625 ();
 sg13g2_decap_8 FILLER_71_2632 ();
 sg13g2_decap_8 FILLER_71_2639 ();
 sg13g2_decap_8 FILLER_71_2646 ();
 sg13g2_decap_8 FILLER_71_2653 ();
 sg13g2_decap_8 FILLER_71_2660 ();
 sg13g2_decap_8 FILLER_71_2667 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_252 ();
 sg13g2_decap_8 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_294 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_8 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_343 ();
 sg13g2_decap_4 FILLER_72_350 ();
 sg13g2_fill_2 FILLER_72_354 ();
 sg13g2_decap_4 FILLER_72_464 ();
 sg13g2_fill_1 FILLER_72_468 ();
 sg13g2_decap_4 FILLER_72_503 ();
 sg13g2_fill_1 FILLER_72_559 ();
 sg13g2_fill_2 FILLER_72_586 ();
 sg13g2_fill_2 FILLER_72_612 ();
 sg13g2_fill_1 FILLER_72_614 ();
 sg13g2_fill_2 FILLER_72_688 ();
 sg13g2_fill_1 FILLER_72_690 ();
 sg13g2_fill_1 FILLER_72_735 ();
 sg13g2_fill_1 FILLER_72_776 ();
 sg13g2_fill_2 FILLER_72_801 ();
 sg13g2_fill_1 FILLER_72_833 ();
 sg13g2_fill_1 FILLER_72_869 ();
 sg13g2_fill_1 FILLER_72_905 ();
 sg13g2_fill_2 FILLER_72_915 ();
 sg13g2_fill_2 FILLER_72_937 ();
 sg13g2_fill_1 FILLER_72_939 ();
 sg13g2_fill_2 FILLER_72_1020 ();
 sg13g2_fill_1 FILLER_72_1022 ();
 sg13g2_fill_2 FILLER_72_1034 ();
 sg13g2_fill_2 FILLER_72_1140 ();
 sg13g2_fill_1 FILLER_72_1142 ();
 sg13g2_fill_2 FILLER_72_1148 ();
 sg13g2_fill_1 FILLER_72_1150 ();
 sg13g2_fill_2 FILLER_72_1182 ();
 sg13g2_fill_1 FILLER_72_1184 ();
 sg13g2_decap_4 FILLER_72_1290 ();
 sg13g2_fill_1 FILLER_72_1308 ();
 sg13g2_fill_2 FILLER_72_1327 ();
 sg13g2_fill_1 FILLER_72_1329 ();
 sg13g2_fill_2 FILLER_72_1365 ();
 sg13g2_fill_2 FILLER_72_1406 ();
 sg13g2_fill_1 FILLER_72_1408 ();
 sg13g2_fill_1 FILLER_72_1453 ();
 sg13g2_fill_2 FILLER_72_1484 ();
 sg13g2_fill_2 FILLER_72_1574 ();
 sg13g2_fill_2 FILLER_72_1611 ();
 sg13g2_fill_1 FILLER_72_1653 ();
 sg13g2_decap_4 FILLER_72_1696 ();
 sg13g2_fill_1 FILLER_72_1700 ();
 sg13g2_fill_2 FILLER_72_1738 ();
 sg13g2_fill_1 FILLER_72_1754 ();
 sg13g2_fill_2 FILLER_72_1812 ();
 sg13g2_fill_2 FILLER_72_2011 ();
 sg13g2_fill_1 FILLER_72_2013 ();
 sg13g2_fill_1 FILLER_72_2069 ();
 sg13g2_fill_2 FILLER_72_2170 ();
 sg13g2_fill_1 FILLER_72_2172 ();
 sg13g2_fill_1 FILLER_72_2212 ();
 sg13g2_fill_2 FILLER_72_2226 ();
 sg13g2_fill_2 FILLER_72_2254 ();
 sg13g2_fill_1 FILLER_72_2256 ();
 sg13g2_fill_1 FILLER_72_2306 ();
 sg13g2_fill_2 FILLER_72_2312 ();
 sg13g2_fill_1 FILLER_72_2319 ();
 sg13g2_fill_2 FILLER_72_2350 ();
 sg13g2_fill_2 FILLER_72_2386 ();
 sg13g2_fill_2 FILLER_72_2427 ();
 sg13g2_decap_4 FILLER_72_2500 ();
 sg13g2_fill_1 FILLER_72_2504 ();
 sg13g2_fill_1 FILLER_72_2572 ();
 sg13g2_decap_8 FILLER_72_2608 ();
 sg13g2_decap_8 FILLER_72_2615 ();
 sg13g2_decap_8 FILLER_72_2622 ();
 sg13g2_decap_8 FILLER_72_2629 ();
 sg13g2_decap_8 FILLER_72_2636 ();
 sg13g2_decap_8 FILLER_72_2643 ();
 sg13g2_decap_8 FILLER_72_2650 ();
 sg13g2_decap_8 FILLER_72_2657 ();
 sg13g2_decap_8 FILLER_72_2664 ();
 sg13g2_fill_2 FILLER_72_2671 ();
 sg13g2_fill_1 FILLER_72_2673 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_8 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_259 ();
 sg13g2_decap_8 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_322 ();
 sg13g2_decap_8 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_fill_2 FILLER_73_357 ();
 sg13g2_decap_4 FILLER_73_504 ();
 sg13g2_decap_8 FILLER_73_554 ();
 sg13g2_fill_2 FILLER_73_561 ();
 sg13g2_fill_1 FILLER_73_602 ();
 sg13g2_fill_2 FILLER_73_711 ();
 sg13g2_fill_2 FILLER_73_745 ();
 sg13g2_fill_2 FILLER_73_791 ();
 sg13g2_fill_1 FILLER_73_793 ();
 sg13g2_fill_1 FILLER_73_803 ();
 sg13g2_fill_2 FILLER_73_848 ();
 sg13g2_fill_2 FILLER_73_941 ();
 sg13g2_fill_2 FILLER_73_954 ();
 sg13g2_fill_1 FILLER_73_982 ();
 sg13g2_fill_2 FILLER_73_1000 ();
 sg13g2_fill_1 FILLER_73_1002 ();
 sg13g2_fill_2 FILLER_73_1025 ();
 sg13g2_fill_1 FILLER_73_1041 ();
 sg13g2_fill_2 FILLER_73_1187 ();
 sg13g2_fill_1 FILLER_73_1258 ();
 sg13g2_decap_4 FILLER_73_1293 ();
 sg13g2_fill_2 FILLER_73_1297 ();
 sg13g2_fill_2 FILLER_73_1312 ();
 sg13g2_fill_1 FILLER_73_1314 ();
 sg13g2_fill_1 FILLER_73_1336 ();
 sg13g2_fill_2 FILLER_73_1397 ();
 sg13g2_fill_1 FILLER_73_1408 ();
 sg13g2_fill_1 FILLER_73_1414 ();
 sg13g2_fill_2 FILLER_73_1423 ();
 sg13g2_fill_2 FILLER_73_1456 ();
 sg13g2_fill_1 FILLER_73_1458 ();
 sg13g2_fill_2 FILLER_73_1560 ();
 sg13g2_fill_1 FILLER_73_1601 ();
 sg13g2_fill_1 FILLER_73_1663 ();
 sg13g2_fill_2 FILLER_73_1724 ();
 sg13g2_fill_2 FILLER_73_1774 ();
 sg13g2_fill_1 FILLER_73_1776 ();
 sg13g2_fill_1 FILLER_73_1847 ();
 sg13g2_fill_2 FILLER_73_1935 ();
 sg13g2_fill_2 FILLER_73_1963 ();
 sg13g2_fill_1 FILLER_73_1965 ();
 sg13g2_fill_2 FILLER_73_1974 ();
 sg13g2_fill_1 FILLER_73_1976 ();
 sg13g2_fill_1 FILLER_73_1981 ();
 sg13g2_fill_2 FILLER_73_2021 ();
 sg13g2_fill_2 FILLER_73_2042 ();
 sg13g2_fill_2 FILLER_73_2105 ();
 sg13g2_fill_2 FILLER_73_2121 ();
 sg13g2_fill_1 FILLER_73_2123 ();
 sg13g2_fill_2 FILLER_73_2156 ();
 sg13g2_fill_2 FILLER_73_2238 ();
 sg13g2_fill_1 FILLER_73_2240 ();
 sg13g2_fill_1 FILLER_73_2246 ();
 sg13g2_fill_1 FILLER_73_2327 ();
 sg13g2_fill_2 FILLER_73_2337 ();
 sg13g2_fill_1 FILLER_73_2339 ();
 sg13g2_fill_2 FILLER_73_2345 ();
 sg13g2_fill_1 FILLER_73_2347 ();
 sg13g2_fill_1 FILLER_73_2399 ();
 sg13g2_fill_2 FILLER_73_2474 ();
 sg13g2_fill_1 FILLER_73_2481 ();
 sg13g2_fill_2 FILLER_73_2499 ();
 sg13g2_fill_2 FILLER_73_2553 ();
 sg13g2_fill_1 FILLER_73_2555 ();
 sg13g2_decap_8 FILLER_73_2603 ();
 sg13g2_decap_8 FILLER_73_2610 ();
 sg13g2_decap_8 FILLER_73_2617 ();
 sg13g2_decap_8 FILLER_73_2624 ();
 sg13g2_decap_8 FILLER_73_2631 ();
 sg13g2_decap_8 FILLER_73_2638 ();
 sg13g2_decap_8 FILLER_73_2645 ();
 sg13g2_decap_8 FILLER_73_2652 ();
 sg13g2_decap_8 FILLER_73_2659 ();
 sg13g2_decap_8 FILLER_73_2666 ();
 sg13g2_fill_1 FILLER_73_2673 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_decap_8 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_266 ();
 sg13g2_decap_8 FILLER_74_273 ();
 sg13g2_decap_8 FILLER_74_280 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_decap_8 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_322 ();
 sg13g2_decap_8 FILLER_74_329 ();
 sg13g2_decap_8 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_fill_2 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_404 ();
 sg13g2_fill_1 FILLER_74_411 ();
 sg13g2_decap_4 FILLER_74_462 ();
 sg13g2_fill_1 FILLER_74_502 ();
 sg13g2_decap_4 FILLER_74_529 ();
 sg13g2_fill_1 FILLER_74_585 ();
 sg13g2_fill_1 FILLER_74_627 ();
 sg13g2_fill_1 FILLER_74_755 ();
 sg13g2_fill_2 FILLER_74_839 ();
 sg13g2_fill_1 FILLER_74_867 ();
 sg13g2_fill_1 FILLER_74_877 ();
 sg13g2_fill_2 FILLER_74_970 ();
 sg13g2_fill_2 FILLER_74_986 ();
 sg13g2_fill_2 FILLER_74_1001 ();
 sg13g2_fill_1 FILLER_74_1021 ();
 sg13g2_fill_2 FILLER_74_1036 ();
 sg13g2_fill_2 FILLER_74_1064 ();
 sg13g2_fill_1 FILLER_74_1066 ();
 sg13g2_fill_2 FILLER_74_1129 ();
 sg13g2_fill_1 FILLER_74_1131 ();
 sg13g2_fill_1 FILLER_74_1215 ();
 sg13g2_fill_2 FILLER_74_1221 ();
 sg13g2_fill_2 FILLER_74_1259 ();
 sg13g2_fill_1 FILLER_74_1261 ();
 sg13g2_fill_1 FILLER_74_1294 ();
 sg13g2_fill_2 FILLER_74_1321 ();
 sg13g2_fill_1 FILLER_74_1323 ();
 sg13g2_fill_2 FILLER_74_1332 ();
 sg13g2_fill_2 FILLER_74_1391 ();
 sg13g2_fill_1 FILLER_74_1393 ();
 sg13g2_fill_2 FILLER_74_1478 ();
 sg13g2_fill_1 FILLER_74_1480 ();
 sg13g2_fill_2 FILLER_74_1513 ();
 sg13g2_decap_4 FILLER_74_1520 ();
 sg13g2_fill_2 FILLER_74_1524 ();
 sg13g2_fill_2 FILLER_74_1538 ();
 sg13g2_fill_2 FILLER_74_1555 ();
 sg13g2_fill_2 FILLER_74_1562 ();
 sg13g2_fill_2 FILLER_74_1604 ();
 sg13g2_fill_2 FILLER_74_1655 ();
 sg13g2_fill_1 FILLER_74_1691 ();
 sg13g2_fill_2 FILLER_74_1774 ();
 sg13g2_fill_1 FILLER_74_1776 ();
 sg13g2_fill_2 FILLER_74_1817 ();
 sg13g2_fill_2 FILLER_74_1859 ();
 sg13g2_fill_1 FILLER_74_1861 ();
 sg13g2_fill_1 FILLER_74_1906 ();
 sg13g2_fill_1 FILLER_74_1911 ();
 sg13g2_fill_1 FILLER_74_1917 ();
 sg13g2_fill_2 FILLER_74_1996 ();
 sg13g2_fill_1 FILLER_74_2064 ();
 sg13g2_fill_1 FILLER_74_2088 ();
 sg13g2_fill_1 FILLER_74_2110 ();
 sg13g2_fill_1 FILLER_74_2116 ();
 sg13g2_fill_2 FILLER_74_2125 ();
 sg13g2_fill_1 FILLER_74_2132 ();
 sg13g2_fill_2 FILLER_74_2245 ();
 sg13g2_fill_2 FILLER_74_2252 ();
 sg13g2_fill_2 FILLER_74_2305 ();
 sg13g2_fill_1 FILLER_74_2307 ();
 sg13g2_fill_2 FILLER_74_2317 ();
 sg13g2_fill_1 FILLER_74_2319 ();
 sg13g2_fill_2 FILLER_74_2348 ();
 sg13g2_fill_1 FILLER_74_2390 ();
 sg13g2_fill_1 FILLER_74_2396 ();
 sg13g2_fill_2 FILLER_74_2401 ();
 sg13g2_fill_2 FILLER_74_2416 ();
 sg13g2_fill_2 FILLER_74_2426 ();
 sg13g2_fill_2 FILLER_74_2506 ();
 sg13g2_fill_2 FILLER_74_2518 ();
 sg13g2_fill_2 FILLER_74_2546 ();
 sg13g2_fill_1 FILLER_74_2548 ();
 sg13g2_decap_8 FILLER_74_2597 ();
 sg13g2_decap_8 FILLER_74_2604 ();
 sg13g2_decap_8 FILLER_74_2611 ();
 sg13g2_decap_8 FILLER_74_2618 ();
 sg13g2_decap_8 FILLER_74_2625 ();
 sg13g2_decap_8 FILLER_74_2632 ();
 sg13g2_decap_8 FILLER_74_2639 ();
 sg13g2_decap_8 FILLER_74_2646 ();
 sg13g2_decap_8 FILLER_74_2653 ();
 sg13g2_decap_8 FILLER_74_2660 ();
 sg13g2_decap_8 FILLER_74_2667 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_336 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_decap_8 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_75_412 ();
 sg13g2_decap_8 FILLER_75_419 ();
 sg13g2_decap_8 FILLER_75_426 ();
 sg13g2_decap_8 FILLER_75_433 ();
 sg13g2_decap_8 FILLER_75_440 ();
 sg13g2_decap_8 FILLER_75_447 ();
 sg13g2_decap_8 FILLER_75_454 ();
 sg13g2_fill_2 FILLER_75_466 ();
 sg13g2_fill_2 FILLER_75_472 ();
 sg13g2_fill_1 FILLER_75_474 ();
 sg13g2_fill_1 FILLER_75_489 ();
 sg13g2_decap_8 FILLER_75_493 ();
 sg13g2_decap_8 FILLER_75_500 ();
 sg13g2_decap_8 FILLER_75_515 ();
 sg13g2_decap_8 FILLER_75_522 ();
 sg13g2_fill_1 FILLER_75_529 ();
 sg13g2_decap_8 FILLER_75_540 ();
 sg13g2_decap_8 FILLER_75_547 ();
 sg13g2_decap_8 FILLER_75_554 ();
 sg13g2_fill_1 FILLER_75_561 ();
 sg13g2_fill_1 FILLER_75_588 ();
 sg13g2_fill_1 FILLER_75_603 ();
 sg13g2_fill_1 FILLER_75_618 ();
 sg13g2_fill_1 FILLER_75_624 ();
 sg13g2_fill_1 FILLER_75_639 ();
 sg13g2_fill_2 FILLER_75_645 ();
 sg13g2_fill_1 FILLER_75_647 ();
 sg13g2_fill_1 FILLER_75_666 ();
 sg13g2_fill_1 FILLER_75_677 ();
 sg13g2_decap_8 FILLER_75_704 ();
 sg13g2_decap_8 FILLER_75_711 ();
 sg13g2_decap_4 FILLER_75_718 ();
 sg13g2_fill_2 FILLER_75_722 ();
 sg13g2_fill_1 FILLER_75_772 ();
 sg13g2_fill_1 FILLER_75_777 ();
 sg13g2_fill_2 FILLER_75_829 ();
 sg13g2_fill_1 FILLER_75_844 ();
 sg13g2_fill_2 FILLER_75_875 ();
 sg13g2_fill_1 FILLER_75_877 ();
 sg13g2_fill_2 FILLER_75_895 ();
 sg13g2_fill_2 FILLER_75_951 ();
 sg13g2_fill_2 FILLER_75_957 ();
 sg13g2_fill_2 FILLER_75_968 ();
 sg13g2_fill_1 FILLER_75_970 ();
 sg13g2_fill_1 FILLER_75_1079 ();
 sg13g2_fill_1 FILLER_75_1088 ();
 sg13g2_fill_1 FILLER_75_1094 ();
 sg13g2_decap_4 FILLER_75_1179 ();
 sg13g2_fill_2 FILLER_75_1183 ();
 sg13g2_fill_1 FILLER_75_1195 ();
 sg13g2_fill_2 FILLER_75_1210 ();
 sg13g2_fill_1 FILLER_75_1212 ();
 sg13g2_decap_8 FILLER_75_1252 ();
 sg13g2_fill_1 FILLER_75_1259 ();
 sg13g2_fill_2 FILLER_75_1265 ();
 sg13g2_fill_2 FILLER_75_1333 ();
 sg13g2_fill_1 FILLER_75_1340 ();
 sg13g2_decap_4 FILLER_75_1355 ();
 sg13g2_fill_1 FILLER_75_1359 ();
 sg13g2_fill_2 FILLER_75_1391 ();
 sg13g2_fill_2 FILLER_75_1423 ();
 sg13g2_fill_1 FILLER_75_1425 ();
 sg13g2_fill_1 FILLER_75_1447 ();
 sg13g2_fill_2 FILLER_75_1457 ();
 sg13g2_fill_1 FILLER_75_1494 ();
 sg13g2_fill_2 FILLER_75_1508 ();
 sg13g2_fill_1 FILLER_75_1515 ();
 sg13g2_fill_1 FILLER_75_1566 ();
 sg13g2_fill_2 FILLER_75_1611 ();
 sg13g2_fill_2 FILLER_75_1630 ();
 sg13g2_fill_1 FILLER_75_1632 ();
 sg13g2_fill_1 FILLER_75_1642 ();
 sg13g2_fill_1 FILLER_75_1656 ();
 sg13g2_fill_2 FILLER_75_1685 ();
 sg13g2_fill_2 FILLER_75_1696 ();
 sg13g2_fill_1 FILLER_75_1698 ();
 sg13g2_fill_2 FILLER_75_1704 ();
 sg13g2_fill_1 FILLER_75_1706 ();
 sg13g2_fill_1 FILLER_75_1734 ();
 sg13g2_fill_1 FILLER_75_1739 ();
 sg13g2_fill_2 FILLER_75_1772 ();
 sg13g2_fill_1 FILLER_75_1818 ();
 sg13g2_fill_2 FILLER_75_1840 ();
 sg13g2_decap_4 FILLER_75_1846 ();
 sg13g2_fill_2 FILLER_75_1850 ();
 sg13g2_decap_8 FILLER_75_1888 ();
 sg13g2_decap_8 FILLER_75_1895 ();
 sg13g2_decap_8 FILLER_75_1902 ();
 sg13g2_decap_8 FILLER_75_1909 ();
 sg13g2_decap_4 FILLER_75_1916 ();
 sg13g2_fill_2 FILLER_75_1920 ();
 sg13g2_fill_1 FILLER_75_1945 ();
 sg13g2_fill_2 FILLER_75_1989 ();
 sg13g2_fill_1 FILLER_75_1991 ();
 sg13g2_fill_2 FILLER_75_2005 ();
 sg13g2_fill_2 FILLER_75_2031 ();
 sg13g2_fill_1 FILLER_75_2033 ();
 sg13g2_fill_1 FILLER_75_2048 ();
 sg13g2_fill_2 FILLER_75_2063 ();
 sg13g2_fill_1 FILLER_75_2065 ();
 sg13g2_fill_2 FILLER_75_2136 ();
 sg13g2_decap_8 FILLER_75_2168 ();
 sg13g2_fill_2 FILLER_75_2180 ();
 sg13g2_fill_1 FILLER_75_2182 ();
 sg13g2_fill_2 FILLER_75_2191 ();
 sg13g2_fill_1 FILLER_75_2193 ();
 sg13g2_fill_1 FILLER_75_2226 ();
 sg13g2_fill_2 FILLER_75_2235 ();
 sg13g2_fill_1 FILLER_75_2262 ();
 sg13g2_decap_4 FILLER_75_2280 ();
 sg13g2_fill_1 FILLER_75_2284 ();
 sg13g2_decap_4 FILLER_75_2289 ();
 sg13g2_fill_2 FILLER_75_2293 ();
 sg13g2_fill_2 FILLER_75_2356 ();
 sg13g2_fill_1 FILLER_75_2358 ();
 sg13g2_fill_2 FILLER_75_2394 ();
 sg13g2_fill_2 FILLER_75_2449 ();
 sg13g2_fill_1 FILLER_75_2451 ();
 sg13g2_fill_1 FILLER_75_2501 ();
 sg13g2_fill_2 FILLER_75_2514 ();
 sg13g2_fill_1 FILLER_75_2516 ();
 sg13g2_decap_8 FILLER_75_2549 ();
 sg13g2_decap_8 FILLER_75_2556 ();
 sg13g2_decap_4 FILLER_75_2563 ();
 sg13g2_fill_2 FILLER_75_2567 ();
 sg13g2_decap_8 FILLER_75_2573 ();
 sg13g2_decap_8 FILLER_75_2580 ();
 sg13g2_decap_8 FILLER_75_2587 ();
 sg13g2_decap_8 FILLER_75_2594 ();
 sg13g2_decap_8 FILLER_75_2601 ();
 sg13g2_decap_8 FILLER_75_2608 ();
 sg13g2_decap_8 FILLER_75_2615 ();
 sg13g2_decap_8 FILLER_75_2622 ();
 sg13g2_decap_8 FILLER_75_2629 ();
 sg13g2_decap_8 FILLER_75_2636 ();
 sg13g2_decap_8 FILLER_75_2643 ();
 sg13g2_decap_8 FILLER_75_2650 ();
 sg13g2_decap_8 FILLER_75_2657 ();
 sg13g2_decap_8 FILLER_75_2664 ();
 sg13g2_fill_2 FILLER_75_2671 ();
 sg13g2_fill_1 FILLER_75_2673 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_8 FILLER_76_427 ();
 sg13g2_fill_2 FILLER_76_434 ();
 sg13g2_decap_4 FILLER_76_444 ();
 sg13g2_fill_1 FILLER_76_448 ();
 sg13g2_fill_1 FILLER_76_465 ();
 sg13g2_fill_1 FILLER_76_471 ();
 sg13g2_decap_8 FILLER_76_483 ();
 sg13g2_fill_1 FILLER_76_490 ();
 sg13g2_decap_4 FILLER_76_501 ();
 sg13g2_fill_2 FILLER_76_505 ();
 sg13g2_decap_4 FILLER_76_517 ();
 sg13g2_fill_1 FILLER_76_521 ();
 sg13g2_decap_8 FILLER_76_548 ();
 sg13g2_decap_4 FILLER_76_555 ();
 sg13g2_fill_1 FILLER_76_559 ();
 sg13g2_fill_1 FILLER_76_603 ();
 sg13g2_fill_2 FILLER_76_609 ();
 sg13g2_fill_1 FILLER_76_611 ();
 sg13g2_fill_2 FILLER_76_675 ();
 sg13g2_fill_2 FILLER_76_686 ();
 sg13g2_decap_8 FILLER_76_705 ();
 sg13g2_decap_8 FILLER_76_712 ();
 sg13g2_fill_1 FILLER_76_719 ();
 sg13g2_fill_1 FILLER_76_724 ();
 sg13g2_fill_1 FILLER_76_746 ();
 sg13g2_fill_1 FILLER_76_751 ();
 sg13g2_decap_4 FILLER_76_760 ();
 sg13g2_fill_2 FILLER_76_764 ();
 sg13g2_decap_8 FILLER_76_821 ();
 sg13g2_fill_1 FILLER_76_828 ();
 sg13g2_fill_1 FILLER_76_837 ();
 sg13g2_fill_1 FILLER_76_850 ();
 sg13g2_fill_2 FILLER_76_872 ();
 sg13g2_fill_1 FILLER_76_874 ();
 sg13g2_fill_2 FILLER_76_913 ();
 sg13g2_fill_1 FILLER_76_915 ();
 sg13g2_fill_2 FILLER_76_955 ();
 sg13g2_fill_1 FILLER_76_957 ();
 sg13g2_fill_2 FILLER_76_963 ();
 sg13g2_fill_1 FILLER_76_1035 ();
 sg13g2_fill_2 FILLER_76_1042 ();
 sg13g2_fill_2 FILLER_76_1076 ();
 sg13g2_fill_1 FILLER_76_1078 ();
 sg13g2_fill_2 FILLER_76_1085 ();
 sg13g2_fill_2 FILLER_76_1112 ();
 sg13g2_fill_1 FILLER_76_1114 ();
 sg13g2_fill_2 FILLER_76_1141 ();
 sg13g2_fill_1 FILLER_76_1143 ();
 sg13g2_fill_1 FILLER_76_1161 ();
 sg13g2_decap_4 FILLER_76_1244 ();
 sg13g2_fill_1 FILLER_76_1248 ();
 sg13g2_fill_2 FILLER_76_1279 ();
 sg13g2_fill_2 FILLER_76_1335 ();
 sg13g2_fill_1 FILLER_76_1337 ();
 sg13g2_fill_1 FILLER_76_1342 ();
 sg13g2_fill_1 FILLER_76_1356 ();
 sg13g2_fill_2 FILLER_76_1366 ();
 sg13g2_fill_1 FILLER_76_1394 ();
 sg13g2_fill_2 FILLER_76_1453 ();
 sg13g2_fill_1 FILLER_76_1455 ();
 sg13g2_fill_1 FILLER_76_1487 ();
 sg13g2_decap_4 FILLER_76_1492 ();
 sg13g2_fill_1 FILLER_76_1496 ();
 sg13g2_fill_2 FILLER_76_1501 ();
 sg13g2_fill_1 FILLER_76_1543 ();
 sg13g2_fill_2 FILLER_76_1595 ();
 sg13g2_fill_1 FILLER_76_1597 ();
 sg13g2_fill_2 FILLER_76_1607 ();
 sg13g2_fill_1 FILLER_76_1609 ();
 sg13g2_fill_1 FILLER_76_1625 ();
 sg13g2_fill_2 FILLER_76_1630 ();
 sg13g2_fill_2 FILLER_76_1657 ();
 sg13g2_fill_1 FILLER_76_1659 ();
 sg13g2_decap_4 FILLER_76_1689 ();
 sg13g2_fill_1 FILLER_76_1723 ();
 sg13g2_fill_2 FILLER_76_1758 ();
 sg13g2_fill_2 FILLER_76_1764 ();
 sg13g2_fill_2 FILLER_76_1813 ();
 sg13g2_fill_1 FILLER_76_1815 ();
 sg13g2_fill_2 FILLER_76_1845 ();
 sg13g2_fill_1 FILLER_76_1847 ();
 sg13g2_fill_2 FILLER_76_1871 ();
 sg13g2_fill_1 FILLER_76_1873 ();
 sg13g2_fill_2 FILLER_76_1891 ();
 sg13g2_fill_2 FILLER_76_1932 ();
 sg13g2_fill_1 FILLER_76_1934 ();
 sg13g2_fill_2 FILLER_76_1989 ();
 sg13g2_fill_1 FILLER_76_1991 ();
 sg13g2_fill_1 FILLER_76_2037 ();
 sg13g2_fill_2 FILLER_76_2059 ();
 sg13g2_fill_2 FILLER_76_2086 ();
 sg13g2_fill_1 FILLER_76_2154 ();
 sg13g2_fill_2 FILLER_76_2164 ();
 sg13g2_fill_1 FILLER_76_2171 ();
 sg13g2_fill_2 FILLER_76_2203 ();
 sg13g2_fill_1 FILLER_76_2205 ();
 sg13g2_fill_1 FILLER_76_2211 ();
 sg13g2_fill_2 FILLER_76_2251 ();
 sg13g2_fill_2 FILLER_76_2266 ();
 sg13g2_fill_1 FILLER_76_2268 ();
 sg13g2_fill_2 FILLER_76_2325 ();
 sg13g2_fill_2 FILLER_76_2391 ();
 sg13g2_fill_1 FILLER_76_2393 ();
 sg13g2_fill_2 FILLER_76_2445 ();
 sg13g2_fill_1 FILLER_76_2447 ();
 sg13g2_decap_8 FILLER_76_2547 ();
 sg13g2_decap_8 FILLER_76_2554 ();
 sg13g2_decap_8 FILLER_76_2561 ();
 sg13g2_decap_8 FILLER_76_2568 ();
 sg13g2_decap_8 FILLER_76_2575 ();
 sg13g2_decap_8 FILLER_76_2582 ();
 sg13g2_decap_8 FILLER_76_2589 ();
 sg13g2_decap_8 FILLER_76_2596 ();
 sg13g2_decap_8 FILLER_76_2603 ();
 sg13g2_decap_8 FILLER_76_2610 ();
 sg13g2_decap_8 FILLER_76_2617 ();
 sg13g2_decap_8 FILLER_76_2624 ();
 sg13g2_decap_8 FILLER_76_2631 ();
 sg13g2_decap_8 FILLER_76_2638 ();
 sg13g2_decap_8 FILLER_76_2645 ();
 sg13g2_decap_8 FILLER_76_2652 ();
 sg13g2_decap_8 FILLER_76_2659 ();
 sg13g2_decap_8 FILLER_76_2666 ();
 sg13g2_fill_1 FILLER_76_2673 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_434 ();
 sg13g2_fill_2 FILLER_77_490 ();
 sg13g2_fill_2 FILLER_77_518 ();
 sg13g2_decap_8 FILLER_77_538 ();
 sg13g2_decap_8 FILLER_77_545 ();
 sg13g2_decap_8 FILLER_77_552 ();
 sg13g2_decap_8 FILLER_77_559 ();
 sg13g2_fill_2 FILLER_77_566 ();
 sg13g2_fill_2 FILLER_77_631 ();
 sg13g2_fill_1 FILLER_77_633 ();
 sg13g2_fill_1 FILLER_77_708 ();
 sg13g2_decap_8 FILLER_77_749 ();
 sg13g2_decap_4 FILLER_77_756 ();
 sg13g2_fill_1 FILLER_77_790 ();
 sg13g2_decap_8 FILLER_77_816 ();
 sg13g2_decap_4 FILLER_77_823 ();
 sg13g2_fill_1 FILLER_77_827 ();
 sg13g2_fill_2 FILLER_77_863 ();
 sg13g2_fill_1 FILLER_77_865 ();
 sg13g2_fill_2 FILLER_77_924 ();
 sg13g2_fill_1 FILLER_77_926 ();
 sg13g2_fill_1 FILLER_77_967 ();
 sg13g2_fill_1 FILLER_77_1016 ();
 sg13g2_fill_1 FILLER_77_1030 ();
 sg13g2_fill_2 FILLER_77_1045 ();
 sg13g2_fill_2 FILLER_77_1052 ();
 sg13g2_fill_1 FILLER_77_1054 ();
 sg13g2_fill_1 FILLER_77_1117 ();
 sg13g2_fill_2 FILLER_77_1136 ();
 sg13g2_fill_1 FILLER_77_1138 ();
 sg13g2_decap_4 FILLER_77_1157 ();
 sg13g2_fill_1 FILLER_77_1161 ();
 sg13g2_fill_2 FILLER_77_1171 ();
 sg13g2_fill_1 FILLER_77_1173 ();
 sg13g2_fill_2 FILLER_77_1200 ();
 sg13g2_fill_2 FILLER_77_1212 ();
 sg13g2_fill_2 FILLER_77_1245 ();
 sg13g2_fill_1 FILLER_77_1303 ();
 sg13g2_fill_1 FILLER_77_1326 ();
 sg13g2_fill_1 FILLER_77_1448 ();
 sg13g2_fill_1 FILLER_77_1497 ();
 sg13g2_fill_2 FILLER_77_1545 ();
 sg13g2_fill_2 FILLER_77_1617 ();
 sg13g2_fill_2 FILLER_77_1645 ();
 sg13g2_fill_1 FILLER_77_1652 ();
 sg13g2_fill_2 FILLER_77_1658 ();
 sg13g2_fill_2 FILLER_77_1686 ();
 sg13g2_fill_2 FILLER_77_1698 ();
 sg13g2_fill_2 FILLER_77_1709 ();
 sg13g2_fill_1 FILLER_77_1711 ();
 sg13g2_decap_8 FILLER_77_1768 ();
 sg13g2_fill_2 FILLER_77_1775 ();
 sg13g2_fill_1 FILLER_77_1781 ();
 sg13g2_fill_1 FILLER_77_1787 ();
 sg13g2_fill_1 FILLER_77_1793 ();
 sg13g2_fill_1 FILLER_77_1804 ();
 sg13g2_fill_2 FILLER_77_1974 ();
 sg13g2_fill_1 FILLER_77_1976 ();
 sg13g2_fill_2 FILLER_77_2008 ();
 sg13g2_fill_1 FILLER_77_2010 ();
 sg13g2_fill_2 FILLER_77_2025 ();
 sg13g2_fill_2 FILLER_77_2083 ();
 sg13g2_fill_1 FILLER_77_2085 ();
 sg13g2_fill_1 FILLER_77_2112 ();
 sg13g2_fill_2 FILLER_77_2153 ();
 sg13g2_fill_1 FILLER_77_2155 ();
 sg13g2_fill_2 FILLER_77_2182 ();
 sg13g2_fill_1 FILLER_77_2184 ();
 sg13g2_fill_2 FILLER_77_2190 ();
 sg13g2_fill_2 FILLER_77_2236 ();
 sg13g2_fill_2 FILLER_77_2285 ();
 sg13g2_fill_2 FILLER_77_2334 ();
 sg13g2_decap_8 FILLER_77_2380 ();
 sg13g2_fill_2 FILLER_77_2387 ();
 sg13g2_fill_2 FILLER_77_2424 ();
 sg13g2_fill_1 FILLER_77_2426 ();
 sg13g2_fill_2 FILLER_77_2475 ();
 sg13g2_fill_2 FILLER_77_2507 ();
 sg13g2_decap_8 FILLER_77_2517 ();
 sg13g2_decap_8 FILLER_77_2524 ();
 sg13g2_decap_8 FILLER_77_2531 ();
 sg13g2_decap_8 FILLER_77_2538 ();
 sg13g2_decap_8 FILLER_77_2545 ();
 sg13g2_decap_8 FILLER_77_2552 ();
 sg13g2_decap_8 FILLER_77_2559 ();
 sg13g2_decap_8 FILLER_77_2566 ();
 sg13g2_decap_8 FILLER_77_2573 ();
 sg13g2_decap_8 FILLER_77_2580 ();
 sg13g2_decap_8 FILLER_77_2587 ();
 sg13g2_decap_8 FILLER_77_2594 ();
 sg13g2_decap_8 FILLER_77_2601 ();
 sg13g2_decap_8 FILLER_77_2608 ();
 sg13g2_decap_8 FILLER_77_2615 ();
 sg13g2_decap_8 FILLER_77_2622 ();
 sg13g2_decap_8 FILLER_77_2629 ();
 sg13g2_decap_8 FILLER_77_2636 ();
 sg13g2_decap_8 FILLER_77_2643 ();
 sg13g2_decap_8 FILLER_77_2650 ();
 sg13g2_decap_8 FILLER_77_2657 ();
 sg13g2_decap_8 FILLER_77_2664 ();
 sg13g2_fill_2 FILLER_77_2671 ();
 sg13g2_fill_1 FILLER_77_2673 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_fill_2 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_532 ();
 sg13g2_decap_8 FILLER_78_539 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_decap_8 FILLER_78_560 ();
 sg13g2_decap_4 FILLER_78_567 ();
 sg13g2_fill_2 FILLER_78_571 ();
 sg13g2_fill_1 FILLER_78_608 ();
 sg13g2_fill_1 FILLER_78_635 ();
 sg13g2_fill_2 FILLER_78_667 ();
 sg13g2_fill_1 FILLER_78_669 ();
 sg13g2_fill_2 FILLER_78_748 ();
 sg13g2_fill_1 FILLER_78_750 ();
 sg13g2_fill_2 FILLER_78_787 ();
 sg13g2_fill_2 FILLER_78_815 ();
 sg13g2_fill_1 FILLER_78_1004 ();
 sg13g2_fill_2 FILLER_78_1169 ();
 sg13g2_fill_2 FILLER_78_1206 ();
 sg13g2_fill_1 FILLER_78_1239 ();
 sg13g2_fill_2 FILLER_78_1292 ();
 sg13g2_fill_1 FILLER_78_1294 ();
 sg13g2_fill_2 FILLER_78_1325 ();
 sg13g2_fill_1 FILLER_78_1327 ();
 sg13g2_fill_1 FILLER_78_1358 ();
 sg13g2_fill_2 FILLER_78_1369 ();
 sg13g2_fill_1 FILLER_78_1371 ();
 sg13g2_fill_1 FILLER_78_1398 ();
 sg13g2_fill_2 FILLER_78_1499 ();
 sg13g2_fill_2 FILLER_78_1614 ();
 sg13g2_fill_2 FILLER_78_1656 ();
 sg13g2_fill_1 FILLER_78_1776 ();
 sg13g2_fill_2 FILLER_78_1807 ();
 sg13g2_fill_2 FILLER_78_1986 ();
 sg13g2_fill_1 FILLER_78_1988 ();
 sg13g2_fill_2 FILLER_78_2046 ();
 sg13g2_fill_1 FILLER_78_2048 ();
 sg13g2_fill_2 FILLER_78_2075 ();
 sg13g2_fill_2 FILLER_78_2113 ();
 sg13g2_fill_1 FILLER_78_2200 ();
 sg13g2_fill_1 FILLER_78_2227 ();
 sg13g2_fill_1 FILLER_78_2285 ();
 sg13g2_fill_2 FILLER_78_2317 ();
 sg13g2_fill_1 FILLER_78_2319 ();
 sg13g2_decap_8 FILLER_78_2372 ();
 sg13g2_decap_8 FILLER_78_2379 ();
 sg13g2_decap_4 FILLER_78_2386 ();
 sg13g2_fill_2 FILLER_78_2435 ();
 sg13g2_fill_2 FILLER_78_2477 ();
 sg13g2_fill_1 FILLER_78_2479 ();
 sg13g2_decap_8 FILLER_78_2515 ();
 sg13g2_decap_8 FILLER_78_2522 ();
 sg13g2_decap_8 FILLER_78_2529 ();
 sg13g2_decap_8 FILLER_78_2536 ();
 sg13g2_decap_8 FILLER_78_2543 ();
 sg13g2_decap_8 FILLER_78_2550 ();
 sg13g2_decap_8 FILLER_78_2557 ();
 sg13g2_decap_8 FILLER_78_2564 ();
 sg13g2_decap_8 FILLER_78_2571 ();
 sg13g2_decap_8 FILLER_78_2578 ();
 sg13g2_decap_8 FILLER_78_2585 ();
 sg13g2_decap_8 FILLER_78_2592 ();
 sg13g2_decap_8 FILLER_78_2599 ();
 sg13g2_decap_8 FILLER_78_2606 ();
 sg13g2_decap_8 FILLER_78_2613 ();
 sg13g2_decap_8 FILLER_78_2620 ();
 sg13g2_decap_8 FILLER_78_2627 ();
 sg13g2_decap_8 FILLER_78_2634 ();
 sg13g2_decap_8 FILLER_78_2641 ();
 sg13g2_decap_8 FILLER_78_2648 ();
 sg13g2_decap_8 FILLER_78_2655 ();
 sg13g2_decap_8 FILLER_78_2662 ();
 sg13g2_decap_4 FILLER_78_2669 ();
 sg13g2_fill_1 FILLER_78_2673 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_4 FILLER_79_266 ();
 sg13g2_fill_2 FILLER_79_270 ();
 sg13g2_fill_2 FILLER_79_285 ();
 sg13g2_fill_1 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_4 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_4 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_341 ();
 sg13g2_decap_4 FILLER_79_348 ();
 sg13g2_decap_8 FILLER_79_365 ();
 sg13g2_decap_8 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_379 ();
 sg13g2_decap_8 FILLER_79_386 ();
 sg13g2_decap_8 FILLER_79_393 ();
 sg13g2_decap_8 FILLER_79_400 ();
 sg13g2_decap_8 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_79_414 ();
 sg13g2_decap_8 FILLER_79_421 ();
 sg13g2_decap_8 FILLER_79_428 ();
 sg13g2_decap_8 FILLER_79_435 ();
 sg13g2_fill_2 FILLER_79_494 ();
 sg13g2_fill_1 FILLER_79_496 ();
 sg13g2_decap_8 FILLER_79_523 ();
 sg13g2_decap_8 FILLER_79_530 ();
 sg13g2_decap_8 FILLER_79_537 ();
 sg13g2_decap_8 FILLER_79_544 ();
 sg13g2_decap_8 FILLER_79_551 ();
 sg13g2_decap_8 FILLER_79_558 ();
 sg13g2_decap_8 FILLER_79_565 ();
 sg13g2_fill_2 FILLER_79_572 ();
 sg13g2_fill_1 FILLER_79_574 ();
 sg13g2_fill_1 FILLER_79_635 ();
 sg13g2_decap_4 FILLER_79_680 ();
 sg13g2_fill_2 FILLER_79_684 ();
 sg13g2_decap_8 FILLER_79_694 ();
 sg13g2_decap_8 FILLER_79_701 ();
 sg13g2_fill_1 FILLER_79_708 ();
 sg13g2_fill_2 FILLER_79_753 ();
 sg13g2_fill_1 FILLER_79_755 ();
 sg13g2_fill_2 FILLER_79_813 ();
 sg13g2_fill_1 FILLER_79_815 ();
 sg13g2_fill_1 FILLER_79_919 ();
 sg13g2_fill_2 FILLER_79_971 ();
 sg13g2_fill_1 FILLER_79_973 ();
 sg13g2_fill_2 FILLER_79_1004 ();
 sg13g2_fill_2 FILLER_79_1036 ();
 sg13g2_fill_1 FILLER_79_1082 ();
 sg13g2_fill_2 FILLER_79_1135 ();
 sg13g2_fill_2 FILLER_79_1193 ();
 sg13g2_fill_2 FILLER_79_1204 ();
 sg13g2_fill_1 FILLER_79_1206 ();
 sg13g2_fill_1 FILLER_79_1233 ();
 sg13g2_fill_2 FILLER_79_1252 ();
 sg13g2_fill_1 FILLER_79_1254 ();
 sg13g2_decap_8 FILLER_79_1285 ();
 sg13g2_decap_8 FILLER_79_1292 ();
 sg13g2_fill_1 FILLER_79_1299 ();
 sg13g2_fill_2 FILLER_79_1357 ();
 sg13g2_decap_4 FILLER_79_1406 ();
 sg13g2_fill_2 FILLER_79_1410 ();
 sg13g2_fill_1 FILLER_79_1447 ();
 sg13g2_fill_1 FILLER_79_1452 ();
 sg13g2_fill_2 FILLER_79_1484 ();
 sg13g2_fill_1 FILLER_79_1486 ();
 sg13g2_fill_1 FILLER_79_1500 ();
 sg13g2_fill_2 FILLER_79_1532 ();
 sg13g2_fill_1 FILLER_79_1534 ();
 sg13g2_fill_2 FILLER_79_1570 ();
 sg13g2_fill_1 FILLER_79_1572 ();
 sg13g2_fill_2 FILLER_79_1651 ();
 sg13g2_fill_1 FILLER_79_1688 ();
 sg13g2_fill_2 FILLER_79_1733 ();
 sg13g2_fill_2 FILLER_79_1770 ();
 sg13g2_fill_1 FILLER_79_1772 ();
 sg13g2_fill_2 FILLER_79_1799 ();
 sg13g2_fill_1 FILLER_79_1801 ();
 sg13g2_fill_2 FILLER_79_1815 ();
 sg13g2_fill_2 FILLER_79_1891 ();
 sg13g2_fill_1 FILLER_79_1893 ();
 sg13g2_fill_2 FILLER_79_2029 ();
 sg13g2_fill_2 FILLER_79_2084 ();
 sg13g2_fill_2 FILLER_79_2112 ();
 sg13g2_fill_2 FILLER_79_2152 ();
 sg13g2_fill_1 FILLER_79_2154 ();
 sg13g2_fill_2 FILLER_79_2198 ();
 sg13g2_fill_1 FILLER_79_2200 ();
 sg13g2_fill_2 FILLER_79_2236 ();
 sg13g2_fill_1 FILLER_79_2296 ();
 sg13g2_decap_8 FILLER_79_2370 ();
 sg13g2_decap_8 FILLER_79_2377 ();
 sg13g2_decap_8 FILLER_79_2384 ();
 sg13g2_decap_4 FILLER_79_2391 ();
 sg13g2_fill_1 FILLER_79_2395 ();
 sg13g2_fill_2 FILLER_79_2405 ();
 sg13g2_fill_2 FILLER_79_2494 ();
 sg13g2_decap_8 FILLER_79_2513 ();
 sg13g2_decap_8 FILLER_79_2520 ();
 sg13g2_decap_8 FILLER_79_2527 ();
 sg13g2_decap_8 FILLER_79_2534 ();
 sg13g2_decap_8 FILLER_79_2541 ();
 sg13g2_decap_8 FILLER_79_2548 ();
 sg13g2_decap_8 FILLER_79_2555 ();
 sg13g2_decap_8 FILLER_79_2562 ();
 sg13g2_decap_8 FILLER_79_2569 ();
 sg13g2_decap_8 FILLER_79_2576 ();
 sg13g2_decap_8 FILLER_79_2583 ();
 sg13g2_decap_8 FILLER_79_2590 ();
 sg13g2_decap_8 FILLER_79_2597 ();
 sg13g2_decap_8 FILLER_79_2604 ();
 sg13g2_decap_8 FILLER_79_2611 ();
 sg13g2_decap_8 FILLER_79_2618 ();
 sg13g2_decap_8 FILLER_79_2625 ();
 sg13g2_decap_8 FILLER_79_2632 ();
 sg13g2_decap_8 FILLER_79_2639 ();
 sg13g2_decap_8 FILLER_79_2646 ();
 sg13g2_decap_8 FILLER_79_2653 ();
 sg13g2_decap_8 FILLER_79_2660 ();
 sg13g2_decap_8 FILLER_79_2667 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_fill_2 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_245 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_423 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_decap_8 FILLER_80_451 ();
 sg13g2_decap_8 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_decap_8 FILLER_80_493 ();
 sg13g2_decap_8 FILLER_80_500 ();
 sg13g2_decap_8 FILLER_80_507 ();
 sg13g2_decap_8 FILLER_80_514 ();
 sg13g2_decap_8 FILLER_80_521 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_fill_1 FILLER_80_570 ();
 sg13g2_fill_2 FILLER_80_626 ();
 sg13g2_fill_1 FILLER_80_628 ();
 sg13g2_fill_1 FILLER_80_647 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_fill_2 FILLER_80_697 ();
 sg13g2_fill_1 FILLER_80_730 ();
 sg13g2_fill_1 FILLER_80_757 ();
 sg13g2_fill_1 FILLER_80_775 ();
 sg13g2_fill_1 FILLER_80_794 ();
 sg13g2_decap_8 FILLER_80_803 ();
 sg13g2_fill_2 FILLER_80_900 ();
 sg13g2_fill_1 FILLER_80_902 ();
 sg13g2_fill_2 FILLER_80_916 ();
 sg13g2_fill_2 FILLER_80_926 ();
 sg13g2_fill_1 FILLER_80_928 ();
 sg13g2_fill_1 FILLER_80_942 ();
 sg13g2_fill_2 FILLER_80_956 ();
 sg13g2_fill_1 FILLER_80_958 ();
 sg13g2_fill_1 FILLER_80_964 ();
 sg13g2_fill_1 FILLER_80_1007 ();
 sg13g2_fill_2 FILLER_80_1024 ();
 sg13g2_fill_1 FILLER_80_1026 ();
 sg13g2_fill_1 FILLER_80_1053 ();
 sg13g2_fill_1 FILLER_80_1063 ();
 sg13g2_fill_2 FILLER_80_1077 ();
 sg13g2_decap_8 FILLER_80_1087 ();
 sg13g2_fill_1 FILLER_80_1094 ();
 sg13g2_fill_2 FILLER_80_1116 ();
 sg13g2_fill_1 FILLER_80_1118 ();
 sg13g2_fill_2 FILLER_80_1131 ();
 sg13g2_fill_2 FILLER_80_1137 ();
 sg13g2_fill_2 FILLER_80_1152 ();
 sg13g2_fill_1 FILLER_80_1154 ();
 sg13g2_fill_2 FILLER_80_1184 ();
 sg13g2_fill_1 FILLER_80_1208 ();
 sg13g2_fill_2 FILLER_80_1235 ();
 sg13g2_fill_1 FILLER_80_1237 ();
 sg13g2_fill_1 FILLER_80_1250 ();
 sg13g2_fill_1 FILLER_80_1259 ();
 sg13g2_fill_1 FILLER_80_1265 ();
 sg13g2_decap_8 FILLER_80_1287 ();
 sg13g2_decap_8 FILLER_80_1294 ();
 sg13g2_fill_2 FILLER_80_1335 ();
 sg13g2_fill_1 FILLER_80_1337 ();
 sg13g2_decap_8 FILLER_80_1346 ();
 sg13g2_decap_4 FILLER_80_1362 ();
 sg13g2_fill_1 FILLER_80_1366 ();
 sg13g2_fill_2 FILLER_80_1375 ();
 sg13g2_fill_2 FILLER_80_1386 ();
 sg13g2_fill_1 FILLER_80_1388 ();
 sg13g2_fill_2 FILLER_80_1406 ();
 sg13g2_decap_8 FILLER_80_1441 ();
 sg13g2_decap_4 FILLER_80_1448 ();
 sg13g2_fill_2 FILLER_80_1452 ();
 sg13g2_fill_1 FILLER_80_1458 ();
 sg13g2_fill_2 FILLER_80_1477 ();
 sg13g2_fill_1 FILLER_80_1496 ();
 sg13g2_fill_2 FILLER_80_1501 ();
 sg13g2_fill_2 FILLER_80_1525 ();
 sg13g2_fill_2 FILLER_80_1553 ();
 sg13g2_fill_1 FILLER_80_1555 ();
 sg13g2_fill_2 FILLER_80_1594 ();
 sg13g2_fill_1 FILLER_80_1596 ();
 sg13g2_fill_2 FILLER_80_1601 ();
 sg13g2_fill_1 FILLER_80_1603 ();
 sg13g2_fill_1 FILLER_80_1630 ();
 sg13g2_fill_1 FILLER_80_1636 ();
 sg13g2_fill_1 FILLER_80_1662 ();
 sg13g2_fill_2 FILLER_80_1689 ();
 sg13g2_fill_1 FILLER_80_1704 ();
 sg13g2_fill_2 FILLER_80_1726 ();
 sg13g2_fill_1 FILLER_80_1728 ();
 sg13g2_fill_2 FILLER_80_1737 ();
 sg13g2_fill_1 FILLER_80_1739 ();
 sg13g2_fill_1 FILLER_80_1823 ();
 sg13g2_fill_1 FILLER_80_1858 ();
 sg13g2_decap_4 FILLER_80_1863 ();
 sg13g2_fill_1 FILLER_80_1880 ();
 sg13g2_fill_1 FILLER_80_1899 ();
 sg13g2_fill_2 FILLER_80_1905 ();
 sg13g2_fill_1 FILLER_80_1907 ();
 sg13g2_fill_2 FILLER_80_1975 ();
 sg13g2_fill_1 FILLER_80_1977 ();
 sg13g2_fill_2 FILLER_80_1982 ();
 sg13g2_fill_1 FILLER_80_1984 ();
 sg13g2_fill_2 FILLER_80_2006 ();
 sg13g2_fill_1 FILLER_80_2008 ();
 sg13g2_fill_2 FILLER_80_2034 ();
 sg13g2_fill_1 FILLER_80_2036 ();
 sg13g2_fill_2 FILLER_80_2042 ();
 sg13g2_fill_1 FILLER_80_2044 ();
 sg13g2_fill_1 FILLER_80_2100 ();
 sg13g2_fill_2 FILLER_80_2127 ();
 sg13g2_fill_1 FILLER_80_2129 ();
 sg13g2_fill_1 FILLER_80_2159 ();
 sg13g2_fill_1 FILLER_80_2168 ();
 sg13g2_fill_2 FILLER_80_2179 ();
 sg13g2_fill_1 FILLER_80_2181 ();
 sg13g2_fill_2 FILLER_80_2204 ();
 sg13g2_fill_2 FILLER_80_2219 ();
 sg13g2_fill_2 FILLER_80_2255 ();
 sg13g2_fill_1 FILLER_80_2286 ();
 sg13g2_decap_4 FILLER_80_2291 ();
 sg13g2_fill_1 FILLER_80_2295 ();
 sg13g2_fill_1 FILLER_80_2300 ();
 sg13g2_fill_2 FILLER_80_2314 ();
 sg13g2_fill_2 FILLER_80_2333 ();
 sg13g2_fill_1 FILLER_80_2335 ();
 sg13g2_decap_8 FILLER_80_2370 ();
 sg13g2_decap_8 FILLER_80_2377 ();
 sg13g2_decap_8 FILLER_80_2384 ();
 sg13g2_decap_4 FILLER_80_2391 ();
 sg13g2_fill_1 FILLER_80_2395 ();
 sg13g2_fill_1 FILLER_80_2404 ();
 sg13g2_fill_2 FILLER_80_2409 ();
 sg13g2_fill_1 FILLER_80_2411 ();
 sg13g2_fill_2 FILLER_80_2460 ();
 sg13g2_fill_1 FILLER_80_2462 ();
 sg13g2_fill_2 FILLER_80_2472 ();
 sg13g2_fill_1 FILLER_80_2474 ();
 sg13g2_decap_8 FILLER_80_2504 ();
 sg13g2_decap_8 FILLER_80_2511 ();
 sg13g2_decap_8 FILLER_80_2518 ();
 sg13g2_decap_8 FILLER_80_2525 ();
 sg13g2_decap_8 FILLER_80_2532 ();
 sg13g2_decap_8 FILLER_80_2539 ();
 sg13g2_decap_8 FILLER_80_2546 ();
 sg13g2_decap_8 FILLER_80_2553 ();
 sg13g2_decap_8 FILLER_80_2560 ();
 sg13g2_decap_8 FILLER_80_2567 ();
 sg13g2_decap_8 FILLER_80_2574 ();
 sg13g2_decap_8 FILLER_80_2581 ();
 sg13g2_decap_8 FILLER_80_2588 ();
 sg13g2_decap_8 FILLER_80_2595 ();
 sg13g2_decap_8 FILLER_80_2602 ();
 sg13g2_decap_8 FILLER_80_2609 ();
 sg13g2_decap_8 FILLER_80_2616 ();
 sg13g2_decap_8 FILLER_80_2623 ();
 sg13g2_decap_8 FILLER_80_2630 ();
 sg13g2_decap_8 FILLER_80_2637 ();
 sg13g2_decap_8 FILLER_80_2644 ();
 sg13g2_decap_8 FILLER_80_2651 ();
 sg13g2_decap_8 FILLER_80_2658 ();
 sg13g2_decap_8 FILLER_80_2665 ();
 sg13g2_fill_2 FILLER_80_2672 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule

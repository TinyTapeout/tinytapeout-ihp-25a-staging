module tt_um_rebeccargb_hardware_utf8 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire clknet_0_clk;
 wire retry;
 wire \u8.empty ;
 wire \u8.hs[0] ;
 wire \u8.hs[1] ;
 wire \u8.hs[2] ;
 wire \u8.hs[3] ;
 wire \u8.hs[4] ;
 wire \u8.hs[5] ;
 wire \u8.ls[0] ;
 wire \u8.ls[1] ;
 wire \u8.ls[2] ;
 wire \u8.ls[3] ;
 wire \u8.ls[4] ;
 wire \u8.ls[5] ;
 wire \u8.ls[6] ;
 wire \u8.ls[7] ;
 wire \u8.ls[8] ;
 wire \u8.ls[9] ;
 wire \u8.rbop[0] ;
 wire \u8.rbop[1] ;
 wire \u8.rbop[2] ;
 wire \u8.rc[16] ;
 wire \u8.rc[17] ;
 wire \u8.rc[18] ;
 wire \u8.rc[19] ;
 wire \u8.rc[20] ;
 wire \u8.rc[21] ;
 wire \u8.rc[22] ;
 wire \u8.rc[23] ;
 wire \u8.rc[24] ;
 wire \u8.rc[25] ;
 wire \u8.rc[26] ;
 wire \u8.rc[27] ;
 wire \u8.rc[28] ;
 wire \u8.rc[29] ;
 wire \u8.rc[30] ;
 wire \u8.rc[31] ;
 wire \u8.rcip[0] ;
 wire \u8.rcip[1] ;
 wire \u8.rcip[2] ;
 wire \u8.rcop[0] ;
 wire \u8.rcop[1] ;
 wire \u8.rcop[2] ;
 wire \u8.ruop[0] ;
 wire \u8.ruop[1] ;
 wire \u8.ruop[2] ;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;

 sg13g2_inv_1 _1259_ (.Y(_0385_),
    .A(\u8.rc[23] ));
 sg13g2_inv_1 _1260_ (.Y(_0386_),
    .A(\u8.rc[22] ));
 sg13g2_inv_1 _1261_ (.Y(_0387_),
    .A(net504));
 sg13g2_inv_1 _1262_ (.Y(_0388_),
    .A(net508));
 sg13g2_inv_1 _1263_ (.Y(_0389_),
    .A(net510));
 sg13g2_inv_1 _1264_ (.Y(_0390_),
    .A(net511));
 sg13g2_inv_2 _1265_ (.Y(_0391_),
    .A(net514));
 sg13g2_inv_1 _1266_ (.Y(_0392_),
    .A(\u8.ruop[2] ));
 sg13g2_inv_1 _1267_ (.Y(_0393_),
    .A(\u8.ruop[0] ));
 sg13g2_inv_1 _1268_ (.Y(_0394_),
    .A(net80));
 sg13g2_inv_1 _1269_ (.Y(_0395_),
    .A(\u8.rcop[1] ));
 sg13g2_inv_1 _1270_ (.Y(_0396_),
    .A(net523));
 sg13g2_inv_2 _1271_ (.Y(_0397_),
    .A(net525));
 sg13g2_inv_1 _1272_ (.Y(_0398_),
    .A(net528));
 sg13g2_inv_2 _1273_ (.Y(_0399_),
    .A(net537));
 sg13g2_inv_2 _1274_ (.Y(_0400_),
    .A(net539));
 sg13g2_inv_2 _1275_ (.Y(_0401_),
    .A(\u8.ls[4] ));
 sg13g2_inv_1 _1276_ (.Y(_0402_),
    .A(\u8.ls[0] ));
 sg13g2_inv_1 _1277_ (.Y(_0403_),
    .A(net548));
 sg13g2_inv_2 _1278_ (.Y(_0404_),
    .A(\u8.rc[27] ));
 sg13g2_inv_2 _1279_ (.Y(_0405_),
    .A(\u8.rc[26] ));
 sg13g2_inv_2 _1280_ (.Y(_0406_),
    .A(net555));
 sg13g2_inv_1 _1281_ (.Y(_0407_),
    .A(net564));
 sg13g2_inv_1 _1282_ (.Y(_0408_),
    .A(net6));
 sg13g2_inv_1 _1283_ (.Y(_0409_),
    .A(_0021_));
 sg13g2_inv_2 _1284_ (.Y(_0410_),
    .A(net545));
 sg13g2_inv_1 _1285_ (.Y(_0411_),
    .A(_0022_));
 sg13g2_inv_2 _1286_ (.Y(_0412_),
    .A(_0024_));
 sg13g2_inv_1 _1287_ (.Y(_0413_),
    .A(_0026_));
 sg13g2_inv_2 _1288_ (.Y(_0414_),
    .A(_0027_));
 sg13g2_inv_1 _1289_ (.Y(_0415_),
    .A(_0028_));
 sg13g2_inv_1 _1290_ (.Y(_0416_),
    .A(net13));
 sg13g2_inv_1 _1291_ (.Y(_0417_),
    .A(net14));
 sg13g2_inv_1 _1292_ (.Y(_0418_),
    .A(net9));
 sg13g2_inv_1 _1293_ (.Y(_0419_),
    .A(net574));
 sg13g2_inv_1 _1294_ (.Y(_0420_),
    .A(net10));
 sg13g2_inv_1 _1295_ (.Y(_0421_),
    .A(_0031_));
 sg13g2_inv_2 _1296_ (.Y(_0422_),
    .A(_0032_));
 sg13g2_inv_1 _1297_ (.Y(_0423_),
    .A(_0033_));
 sg13g2_inv_1 _1298_ (.Y(_0424_),
    .A(net2));
 sg13g2_inv_1 _1299_ (.Y(_0425_),
    .A(net7));
 sg13g2_inv_2 _1300_ (.Y(_0426_),
    .A(_0000_));
 sg13g2_inv_1 _1301_ (.Y(_0427_),
    .A(net8));
 sg13g2_inv_2 _1302_ (.Y(_0428_),
    .A(_0002_));
 sg13g2_inv_2 _1303_ (.Y(_0429_),
    .A(_0008_));
 sg13g2_inv_2 _1304_ (.Y(_0430_),
    .A(_0009_));
 sg13g2_inv_2 _1305_ (.Y(_0431_),
    .A(_0010_));
 sg13g2_inv_1 _1306_ (.Y(_0432_),
    .A(_0013_));
 sg13g2_inv_1 _1307_ (.Y(_0433_),
    .A(_0014_));
 sg13g2_inv_2 _1308_ (.Y(_0434_),
    .A(_0015_));
 sg13g2_inv_1 _1309_ (.Y(_0435_),
    .A(_0019_));
 sg13g2_inv_1 _1310_ (.Y(_0436_),
    .A(_0018_));
 sg13g2_inv_1 _1311_ (.Y(_0437_),
    .A(_0020_));
 sg13g2_nand2_2 _1312_ (.Y(_0438_),
    .A(net549),
    .B(\u8.rc[29] ));
 sg13g2_nor2b_1 _1313_ (.A(\u8.rc[29] ),
    .B_N(\u8.rc[28] ),
    .Y(_0439_));
 sg13g2_and3_1 _1314_ (.X(_0440_),
    .A(net549),
    .B(net553),
    .C(_0439_));
 sg13g2_nand3_1 _1315_ (.B(net553),
    .C(_0439_),
    .A(net549),
    .Y(_0441_));
 sg13g2_nor2_1 _1316_ (.A(_0405_),
    .B(_0406_),
    .Y(_0442_));
 sg13g2_nand2_1 _1317_ (.Y(_0443_),
    .A(net554),
    .B(\u8.rc[25] ));
 sg13g2_nand3_1 _1318_ (.B(\u8.rc[22] ),
    .C(\u8.rc[24] ),
    .A(\u8.rc[23] ),
    .Y(_0444_));
 sg13g2_nor3_1 _1319_ (.A(_0405_),
    .B(net555),
    .C(_0444_),
    .Y(_0445_));
 sg13g2_nand3_1 _1320_ (.B(net509),
    .C(\u8.rc[18] ),
    .A(net505),
    .Y(_0446_));
 sg13g2_and2_1 _1321_ (.A(net514),
    .B(net518),
    .X(_0447_));
 sg13g2_and2_2 _1322_ (.A(net518),
    .B(net520),
    .X(_0448_));
 sg13g2_and3_2 _1323_ (.X(_0449_),
    .A(net514),
    .B(net518),
    .C(net519));
 sg13g2_and2_1 _1324_ (.A(net527),
    .B(net530),
    .X(_0450_));
 sg13g2_and4_1 _1325_ (.A(net524),
    .B(net527),
    .C(net529),
    .D(net532),
    .X(_0451_));
 sg13g2_and2_1 _1326_ (.A(net520),
    .B(net521),
    .X(_0452_));
 sg13g2_a221oi_1 _1327_ (.B2(_0447_),
    .C1(net511),
    .B1(_0452_),
    .A1(_0449_),
    .Y(_0453_),
    .A2(_0451_));
 sg13g2_o21ai_1 _1328_ (.B1(_0387_),
    .Y(_0454_),
    .A1(_0446_),
    .A2(_0453_));
 sg13g2_a21oi_1 _1329_ (.A1(_0445_),
    .A2(_0454_),
    .Y(_0455_),
    .B1(_0442_));
 sg13g2_nand2b_1 _1330_ (.Y(_0456_),
    .B(_0440_),
    .A_N(_0455_));
 sg13g2_o21ai_1 _1331_ (.B1(_0438_),
    .Y(_0457_),
    .A1(_0441_),
    .A2(_0455_));
 sg13g2_nand2_1 _1332_ (.Y(_0458_),
    .A(net551),
    .B(\u8.rc[28] ));
 sg13g2_nand4_1 _1333_ (.B(net551),
    .C(net552),
    .A(net549),
    .Y(_0459_),
    .D(net553));
 sg13g2_or3_1 _1334_ (.A(_0024_),
    .B(_0443_),
    .C(_0459_),
    .X(_0460_));
 sg13g2_nand4_1 _1335_ (.B(\u8.rc[22] ),
    .C(net504),
    .A(\u8.rc[23] ),
    .Y(_0461_),
    .D(\u8.rc[24] ));
 sg13g2_nor3_1 _1336_ (.A(_0443_),
    .B(_0459_),
    .C(_0461_),
    .Y(_0462_));
 sg13g2_nand3_1 _1337_ (.B(net508),
    .C(_0412_),
    .A(net505),
    .Y(_0463_));
 sg13g2_nand3_1 _1338_ (.B(_0462_),
    .C(_0463_),
    .A(net547),
    .Y(_0464_));
 sg13g2_nor2_1 _1339_ (.A(_0444_),
    .B(_0460_),
    .Y(_0465_));
 sg13g2_nor2b_1 _1340_ (.A(_0460_),
    .B_N(_0464_),
    .Y(_0466_));
 sg13g2_nand4_1 _1341_ (.B(net506),
    .C(net509),
    .A(net504),
    .Y(_0467_),
    .D(\u8.rc[18] ));
 sg13g2_and2_1 _1342_ (.A(net511),
    .B(net513),
    .X(_0468_));
 sg13g2_nand2b_1 _1343_ (.Y(_0469_),
    .B(_0468_),
    .A_N(_0467_));
 sg13g2_nand2_1 _1344_ (.Y(_0470_),
    .A(net546),
    .B(net549));
 sg13g2_nor2_1 _1345_ (.A(_0404_),
    .B(_0405_),
    .Y(_0471_));
 sg13g2_nand3_1 _1346_ (.B(net554),
    .C(net555),
    .A(net553),
    .Y(_0472_));
 sg13g2_or2_1 _1347_ (.X(_0473_),
    .B(_0472_),
    .A(_0444_));
 sg13g2_nor3_1 _1348_ (.A(_0444_),
    .B(_0458_),
    .C(_0472_),
    .Y(_0474_));
 sg13g2_nor2b_2 _1349_ (.A(_0470_),
    .B_N(_0474_),
    .Y(_0475_));
 sg13g2_nand2b_2 _1350_ (.Y(_0476_),
    .B(_0475_),
    .A_N(_0469_));
 sg13g2_nand4_1 _1351_ (.B(net508),
    .C(\u8.rc[18] ),
    .A(net505),
    .Y(_0477_),
    .D(net511));
 sg13g2_nor4_2 _1352_ (.A(_0443_),
    .B(_0459_),
    .C(_0461_),
    .Y(_0478_),
    .D(_0477_));
 sg13g2_and2_1 _1353_ (.A(net533),
    .B(net536),
    .X(_0479_));
 sg13g2_and4_1 _1354_ (.A(net547),
    .B(_0451_),
    .C(_0452_),
    .D(_0479_),
    .X(_0480_));
 sg13g2_and3_1 _1355_ (.X(_0481_),
    .A(_0447_),
    .B(_0478_),
    .C(_0480_));
 sg13g2_nand4_1 _1356_ (.B(\u8.ls[3] ),
    .C(net544),
    .A(net542),
    .Y(_0482_),
    .D(\u8.ls[1] ));
 sg13g2_nand2_1 _1357_ (.Y(_0483_),
    .A(\u8.ls[6] ),
    .B(net541));
 sg13g2_nand4_1 _1358_ (.B(net537),
    .C(net539),
    .A(net534),
    .Y(_0484_),
    .D(net541));
 sg13g2_o21ai_1 _1359_ (.B1(net538),
    .Y(_0485_),
    .A1(_0482_),
    .A2(_0484_));
 sg13g2_nand4_1 _1360_ (.B(_0478_),
    .C(_0480_),
    .A(_0447_),
    .Y(_0486_),
    .D(_0485_));
 sg13g2_nand3_1 _1361_ (.B(net524),
    .C(_0448_),
    .A(net521),
    .Y(_0487_));
 sg13g2_nor2_1 _1362_ (.A(_0398_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_nand2_1 _1363_ (.Y(_0489_),
    .A(_0412_),
    .B(_0478_));
 sg13g2_nand4_1 _1364_ (.B(_0412_),
    .C(_0449_),
    .A(net521),
    .Y(_0490_),
    .D(_0478_));
 sg13g2_a21oi_1 _1365_ (.A1(_0486_),
    .A2(_0488_),
    .Y(_0491_),
    .B1(_0490_));
 sg13g2_and4_1 _1366_ (.A(net546),
    .B(net550),
    .C(net551),
    .D(net552),
    .X(_0492_));
 sg13g2_nand4_1 _1367_ (.B(net549),
    .C(net551),
    .A(net546),
    .Y(_0493_),
    .D(net552));
 sg13g2_nor2_1 _1368_ (.A(_0473_),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_o21ai_1 _1369_ (.B1(_0466_),
    .Y(_0495_),
    .A1(_0476_),
    .A2(_0491_));
 sg13g2_nor2_2 _1370_ (.A(_0404_),
    .B(_0493_),
    .Y(_0496_));
 sg13g2_nor3_1 _1371_ (.A(_0404_),
    .B(_0405_),
    .C(_0493_),
    .Y(_0497_));
 sg13g2_a22oi_1 _1372_ (.Y(_0498_),
    .B1(_0495_),
    .B2(_0497_),
    .A2(_0456_),
    .A1(_0438_));
 sg13g2_a21oi_1 _1373_ (.A1(net505),
    .A2(net508),
    .Y(_0499_),
    .B1(net504));
 sg13g2_nor4_1 _1374_ (.A(_0405_),
    .B(net555),
    .C(_0444_),
    .D(_0499_),
    .Y(_0500_));
 sg13g2_o21ai_1 _1375_ (.B1(_0440_),
    .Y(_0501_),
    .A1(_0442_),
    .A2(_0500_));
 sg13g2_nand2_1 _1376_ (.Y(_0502_),
    .A(_0438_),
    .B(_0501_));
 sg13g2_a21oi_2 _1377_ (.B1(_0024_),
    .Y(_0503_),
    .A2(_0501_),
    .A1(_0438_));
 sg13g2_nand2b_1 _1378_ (.Y(_0504_),
    .B(_0448_),
    .A_N(_0029_));
 sg13g2_nor2_1 _1379_ (.A(net522),
    .B(_0397_),
    .Y(_0505_));
 sg13g2_nand2_1 _1380_ (.Y(_0506_),
    .A(_0448_),
    .B(_0505_));
 sg13g2_o21ai_1 _1381_ (.B1(_0450_),
    .Y(_0507_),
    .A1(net531),
    .A2(net533));
 sg13g2_o21ai_1 _1382_ (.B1(_0504_),
    .Y(_0508_),
    .A1(_0506_),
    .A2(_0507_));
 sg13g2_nor2_1 _1383_ (.A(net511),
    .B(_0391_),
    .Y(_0509_));
 sg13g2_and2_1 _1384_ (.A(_0026_),
    .B(_0027_),
    .X(_0510_));
 sg13g2_nand3_1 _1385_ (.B(_0028_),
    .C(_0510_),
    .A(_0025_),
    .Y(_0511_));
 sg13g2_a21oi_1 _1386_ (.A1(_0508_),
    .A2(_0509_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_nand2b_1 _1387_ (.Y(_0513_),
    .B(_0503_),
    .A_N(_0512_));
 sg13g2_o21ai_1 _1388_ (.B1(_0510_),
    .Y(_0514_),
    .A1(net503),
    .A2(_0446_));
 sg13g2_o21ai_1 _1389_ (.B1(_0026_),
    .Y(_0515_),
    .A1(net555),
    .A2(_0444_));
 sg13g2_nand4_1 _1390_ (.B(_0471_),
    .C(_0514_),
    .A(_0439_),
    .Y(_0516_),
    .D(_0515_));
 sg13g2_a21oi_2 _1391_ (.B1(_0470_),
    .Y(_0517_),
    .A2(_0516_),
    .A1(_0025_));
 sg13g2_nor2b_1 _1392_ (.A(_0517_),
    .B_N(_0503_),
    .Y(_0518_));
 sg13g2_inv_1 _1393_ (.Y(_0519_),
    .A(_0518_));
 sg13g2_nor2_1 _1394_ (.A(_0410_),
    .B(_0518_),
    .Y(_0520_));
 sg13g2_o21ai_1 _1395_ (.B1(_0520_),
    .Y(_0521_),
    .A1(_0498_),
    .A2(_0513_));
 sg13g2_or3_1 _1396_ (.A(net529),
    .B(net531),
    .C(net533),
    .X(_0522_));
 sg13g2_nor3_2 _1397_ (.A(net521),
    .B(net524),
    .C(net527),
    .Y(_0523_));
 sg13g2_nor2_1 _1398_ (.A(net518),
    .B(net520),
    .Y(_0524_));
 sg13g2_and2_1 _1399_ (.A(_0523_),
    .B(_0524_),
    .X(_0525_));
 sg13g2_nand3b_1 _1400_ (.B(_0523_),
    .C(_0524_),
    .Y(_0526_),
    .A_N(_0522_));
 sg13g2_nor4_2 _1401_ (.A(_0402_),
    .B(net548),
    .C(_0482_),
    .Y(_0527_),
    .D(_0483_));
 sg13g2_nor4_2 _1402_ (.A(net549),
    .B(net551),
    .C(net552),
    .Y(_0528_),
    .D(net553));
 sg13g2_nor2_1 _1403_ (.A(net512),
    .B(net513),
    .Y(_0529_));
 sg13g2_nor3_2 _1404_ (.A(net510),
    .B(net512),
    .C(net514),
    .Y(_0530_));
 sg13g2_or4_1 _1405_ (.A(net508),
    .B(net510),
    .C(net511),
    .D(net514),
    .X(_0531_));
 sg13g2_nor2_1 _1406_ (.A(net506),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_nor2_1 _1407_ (.A(net555),
    .B(\u8.rc[24] ),
    .Y(_0533_));
 sg13g2_nor3_2 _1408_ (.A(\u8.rc[23] ),
    .B(\u8.rc[22] ),
    .C(net503),
    .Y(_0534_));
 sg13g2_nand3_1 _1409_ (.B(_0533_),
    .C(_0534_),
    .A(_0405_),
    .Y(_0535_));
 sg13g2_nor2_1 _1410_ (.A(net546),
    .B(net554),
    .Y(_0536_));
 sg13g2_and4_1 _1411_ (.A(_0528_),
    .B(_0533_),
    .C(_0534_),
    .D(_0536_),
    .X(_0537_));
 sg13g2_nand4_1 _1412_ (.B(_0533_),
    .C(_0534_),
    .A(_0528_),
    .Y(_0538_),
    .D(_0536_));
 sg13g2_nor3_1 _1413_ (.A(net503),
    .B(net505),
    .C(net508),
    .Y(_0539_));
 sg13g2_nand2_1 _1414_ (.Y(_0540_),
    .A(_0530_),
    .B(_0539_));
 sg13g2_and2_1 _1415_ (.A(_0532_),
    .B(_0537_),
    .X(_0541_));
 sg13g2_nand2_1 _1416_ (.Y(_0542_),
    .A(_0532_),
    .B(_0537_));
 sg13g2_o21ai_1 _1417_ (.B1(_0448_),
    .Y(_0543_),
    .A1(net522),
    .A2(net524));
 sg13g2_a21oi_2 _1418_ (.B1(_0543_),
    .Y(_0544_),
    .A2(_0505_),
    .A1(_0398_));
 sg13g2_nor2_1 _1419_ (.A(net487),
    .B(_0544_),
    .Y(_0545_));
 sg13g2_nor3_1 _1420_ (.A(net506),
    .B(net508),
    .C(net536),
    .Y(_0546_));
 sg13g2_nand4_1 _1421_ (.B(_0528_),
    .C(_0530_),
    .A(_0024_),
    .Y(_0547_),
    .D(_0546_));
 sg13g2_nor4_2 _1422_ (.A(_0526_),
    .B(_0527_),
    .C(_0535_),
    .Y(_0548_),
    .D(_0547_));
 sg13g2_nor2_1 _1423_ (.A(_0487_),
    .B(_0507_),
    .Y(_0549_));
 sg13g2_nand2_1 _1424_ (.Y(_0550_),
    .A(net533),
    .B(_0450_));
 sg13g2_nor2_1 _1425_ (.A(net531),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_nand2_1 _1426_ (.Y(_0552_),
    .A(net537),
    .B(net538));
 sg13g2_nor2_1 _1427_ (.A(net541),
    .B(net542),
    .Y(_0553_));
 sg13g2_o21ai_1 _1428_ (.B1(_0551_),
    .Y(_0554_),
    .A1(_0552_),
    .A2(_0553_));
 sg13g2_a21oi_1 _1429_ (.A1(_0549_),
    .A2(_0554_),
    .Y(_0555_),
    .B1(_0542_));
 sg13g2_nand2_1 _1430_ (.Y(_0556_),
    .A(net537),
    .B(net542));
 sg13g2_o21ai_1 _1431_ (.B1(_0551_),
    .Y(_0557_),
    .A1(_0483_),
    .A2(_0556_));
 sg13g2_a21oi_1 _1432_ (.A1(_0549_),
    .A2(_0557_),
    .Y(_0558_),
    .B1(_0542_));
 sg13g2_nor4_2 _1433_ (.A(_0388_),
    .B(_0389_),
    .C(_0390_),
    .Y(_0559_),
    .D(_0391_));
 sg13g2_nor3_1 _1434_ (.A(net505),
    .B(_0538_),
    .C(_0559_),
    .Y(_0560_));
 sg13g2_inv_1 _1435_ (.Y(_0561_),
    .A(_0560_));
 sg13g2_nand3_1 _1436_ (.B(net531),
    .C(net533),
    .A(net528),
    .Y(_0562_));
 sg13g2_nand3_1 _1437_ (.B(net533),
    .C(_0450_),
    .A(net531),
    .Y(_0563_));
 sg13g2_nor4_2 _1438_ (.A(_0482_),
    .B(_0484_),
    .C(_0487_),
    .Y(_0564_),
    .D(_0563_));
 sg13g2_nor3_1 _1439_ (.A(_0558_),
    .B(_0561_),
    .C(_0564_),
    .Y(_0565_));
 sg13g2_nor2_1 _1440_ (.A(_0555_),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_nor2_1 _1441_ (.A(net528),
    .B(_0522_),
    .Y(_0567_));
 sg13g2_nor4_2 _1442_ (.A(\u8.ls[3] ),
    .B(\u8.ls[2] ),
    .C(\u8.ls[1] ),
    .Y(_0568_),
    .D(\u8.ls[0] ));
 sg13g2_nand4_1 _1443_ (.B(_0400_),
    .C(_0553_),
    .A(_0399_),
    .Y(_0569_),
    .D(_0568_));
 sg13g2_nand4_1 _1444_ (.B(_0397_),
    .C(_0448_),
    .A(net521),
    .Y(_0570_),
    .D(_0567_));
 sg13g2_o21ai_1 _1445_ (.B1(_0504_),
    .Y(_0571_),
    .A1(_0569_),
    .A2(_0570_));
 sg13g2_nor2_2 _1446_ (.A(net487),
    .B(_0571_),
    .Y(_0572_));
 sg13g2_a21oi_1 _1447_ (.A1(_0488_),
    .A2(_0522_),
    .Y(_0573_),
    .B1(net487));
 sg13g2_nor3_1 _1448_ (.A(_0566_),
    .B(_0572_),
    .C(_0573_),
    .Y(_0574_));
 sg13g2_or3_1 _1449_ (.A(_0545_),
    .B(_0548_),
    .C(_0574_),
    .X(_0575_));
 sg13g2_nor4_2 _1450_ (.A(net505),
    .B(_0526_),
    .C(_0531_),
    .Y(_0576_),
    .D(_0538_));
 sg13g2_nor3_1 _1451_ (.A(net537),
    .B(net538),
    .C(net540),
    .Y(_0577_));
 sg13g2_or4_1 _1452_ (.A(net542),
    .B(net543),
    .C(net544),
    .D(\u8.ls[1] ),
    .X(_0578_));
 sg13g2_nor2b_1 _1453_ (.A(net538),
    .B_N(net537),
    .Y(_0579_));
 sg13g2_and4_1 _1454_ (.A(net541),
    .B(_0401_),
    .C(_0568_),
    .D(_0579_),
    .X(_0580_));
 sg13g2_a21oi_1 _1455_ (.A1(_0400_),
    .A2(_0033_),
    .Y(_0581_),
    .B1(_0399_));
 sg13g2_nor3_1 _1456_ (.A(_0548_),
    .B(_0580_),
    .C(_0581_),
    .Y(_0582_));
 sg13g2_o21ai_1 _1457_ (.B1(_0576_),
    .Y(_0583_),
    .A1(_0577_),
    .A2(_0582_));
 sg13g2_nor3_1 _1458_ (.A(\u8.empty ),
    .B(net548),
    .C(net2),
    .Y(_0584_));
 sg13g2_or3_1 _1459_ (.A(\u8.empty ),
    .B(net548),
    .C(net2),
    .X(_0585_));
 sg13g2_nand3_1 _1460_ (.B(_0583_),
    .C(_0584_),
    .A(_0575_),
    .Y(_0586_));
 sg13g2_o21ai_1 _1461_ (.B1(_0586_),
    .Y(uo_out[0]),
    .A1(_0424_),
    .A2(_0521_));
 sg13g2_nand2_1 _1462_ (.Y(_0587_),
    .A(retry),
    .B(net2));
 sg13g2_o21ai_1 _1463_ (.B1(_0587_),
    .Y(uo_out[1]),
    .A1(_0583_),
    .A2(_0585_));
 sg13g2_a21o_1 _1464_ (.A2(_0457_),
    .A1(net546),
    .B1(_0512_),
    .X(_0588_));
 sg13g2_and2_1 _1465_ (.A(_0517_),
    .B(_0588_),
    .X(_0589_));
 sg13g2_nor2_1 _1466_ (.A(net553),
    .B(net554),
    .Y(_0590_));
 sg13g2_nand2_1 _1467_ (.Y(_0591_),
    .A(_0464_),
    .B(_0540_));
 sg13g2_and2_1 _1468_ (.A(net546),
    .B(_0478_),
    .X(_0592_));
 sg13g2_nand2_1 _1469_ (.Y(_0593_),
    .A(_0399_),
    .B(_0567_));
 sg13g2_and3_1 _1470_ (.X(_0594_),
    .A(net524),
    .B(net547),
    .C(_0452_));
 sg13g2_nand4_1 _1471_ (.B(_0478_),
    .C(_0593_),
    .A(_0447_),
    .Y(_0595_),
    .D(_0594_));
 sg13g2_nor3_1 _1472_ (.A(_0469_),
    .B(_0473_),
    .C(_0487_),
    .Y(_0596_));
 sg13g2_and2_1 _1473_ (.A(_0492_),
    .B(_0596_),
    .X(_0597_));
 sg13g2_a22oi_1 _1474_ (.Y(_0598_),
    .B1(_0595_),
    .B2(_0597_),
    .A2(_0525_),
    .A1(_0391_));
 sg13g2_o21ai_1 _1475_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0476_),
    .A2(_0491_));
 sg13g2_a21oi_1 _1476_ (.A1(_0592_),
    .A2(_0599_),
    .Y(_0600_),
    .B1(_0591_));
 sg13g2_nand2b_1 _1477_ (.Y(_0601_),
    .B(_0475_),
    .A_N(_0600_));
 sg13g2_nand2_1 _1478_ (.Y(_0602_),
    .A(net554),
    .B(_0460_));
 sg13g2_nand3_1 _1479_ (.B(_0601_),
    .C(_0602_),
    .A(_0535_),
    .Y(_0603_));
 sg13g2_a21oi_1 _1480_ (.A1(_0496_),
    .A2(_0603_),
    .Y(_0604_),
    .B1(_0590_));
 sg13g2_a21o_1 _1481_ (.A2(_0516_),
    .A1(_0025_),
    .B1(_0493_),
    .X(_0605_));
 sg13g2_o21ai_1 _1482_ (.B1(_0589_),
    .Y(_0606_),
    .A1(_0604_),
    .A2(_0605_));
 sg13g2_a21o_2 _1483_ (.A2(_0531_),
    .A1(net505),
    .B1(_0538_),
    .X(_0607_));
 sg13g2_nand4_1 _1484_ (.B(_0412_),
    .C(net2),
    .A(_0017_),
    .Y(_0608_),
    .D(_0607_));
 sg13g2_a21oi_1 _1485_ (.A1(_0502_),
    .A2(_0606_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_a21o_1 _1486_ (.A2(_0450_),
    .A1(net524),
    .B1(net521),
    .X(_0610_));
 sg13g2_a21oi_2 _1487_ (.B1(net487),
    .Y(_0611_),
    .A2(_0610_),
    .A1(_0448_));
 sg13g2_nor2_1 _1488_ (.A(_0572_),
    .B(_0611_),
    .Y(_0612_));
 sg13g2_o21ai_1 _1489_ (.B1(_0584_),
    .Y(_0613_),
    .A1(net487),
    .A2(_0544_));
 sg13g2_or2_1 _1490_ (.X(_0614_),
    .B(_0613_),
    .A(_0612_));
 sg13g2_nand2b_2 _1491_ (.Y(uo_out[2]),
    .B(_0614_),
    .A_N(_0609_));
 sg13g2_nand2_1 _1492_ (.Y(_0615_),
    .A(_0475_),
    .B(_0540_));
 sg13g2_a21oi_1 _1493_ (.A1(net546),
    .A2(_0598_),
    .Y(_0616_),
    .B1(_0489_));
 sg13g2_o21ai_1 _1494_ (.B1(_0465_),
    .Y(_0617_),
    .A1(_0615_),
    .A2(_0616_));
 sg13g2_a21oi_1 _1495_ (.A1(_0535_),
    .A2(_0617_),
    .Y(_0618_),
    .B1(_0404_));
 sg13g2_nor3_1 _1496_ (.A(_0493_),
    .B(_0590_),
    .C(_0618_),
    .Y(_0619_));
 sg13g2_nand2_2 _1497_ (.Y(_0620_),
    .A(net545),
    .B(_0503_));
 sg13g2_or4_1 _1498_ (.A(_0424_),
    .B(_0605_),
    .C(_0619_),
    .D(_0620_),
    .X(_0621_));
 sg13g2_nand2_1 _1499_ (.Y(_0622_),
    .A(net3),
    .B(_0607_));
 sg13g2_a21oi_1 _1500_ (.A1(net487),
    .A2(_0622_),
    .Y(_0623_),
    .B1(_0611_));
 sg13g2_o21ai_1 _1501_ (.B1(_0621_),
    .Y(uo_out[3]),
    .A1(_0613_),
    .A2(_0623_));
 sg13g2_and3_1 _1502_ (.X(_0624_),
    .A(_0403_),
    .B(net545),
    .C(_0607_));
 sg13g2_nand2_1 _1503_ (.Y(_0625_),
    .A(net2),
    .B(_0624_));
 sg13g2_nor2_1 _1504_ (.A(_0560_),
    .B(_0564_),
    .Y(_0626_));
 sg13g2_a21oi_1 _1505_ (.A1(_0622_),
    .A2(_0626_),
    .Y(_0627_),
    .B1(_0573_));
 sg13g2_nor2_1 _1506_ (.A(_0572_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nand3_1 _1507_ (.B(_0568_),
    .C(_0579_),
    .A(_0553_),
    .Y(_0629_));
 sg13g2_nor2_1 _1508_ (.A(_0021_),
    .B(_0543_),
    .Y(_0630_));
 sg13g2_nor3_1 _1509_ (.A(net529),
    .B(_0506_),
    .C(_0629_),
    .Y(_0631_));
 sg13g2_a21oi_1 _1510_ (.A1(_0629_),
    .A2(_0630_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_o21ai_1 _1511_ (.B1(_0611_),
    .Y(_0633_),
    .A1(_0562_),
    .A2(_0632_));
 sg13g2_o21ai_1 _1512_ (.B1(_0633_),
    .Y(_0634_),
    .A1(_0611_),
    .A2(_0628_));
 sg13g2_o21ai_1 _1513_ (.B1(_0625_),
    .Y(uo_out[4]),
    .A1(_0585_),
    .A2(_0634_));
 sg13g2_a21oi_1 _1514_ (.A1(_0564_),
    .A2(_0622_),
    .Y(_0635_),
    .B1(_0558_));
 sg13g2_nor4_1 _1515_ (.A(_0555_),
    .B(_0572_),
    .C(_0585_),
    .D(_0635_),
    .Y(_0636_));
 sg13g2_a21o_1 _1516_ (.A2(_0624_),
    .A1(net3),
    .B1(retry),
    .X(_0637_));
 sg13g2_a21oi_1 _1517_ (.A1(net2),
    .A2(_0637_),
    .Y(_0638_),
    .B1(_0636_));
 sg13g2_nand3b_1 _1518_ (.B(_0621_),
    .C(_0638_),
    .Y(uo_out[5]),
    .A_N(_0609_));
 sg13g2_nor3_2 _1519_ (.A(_0410_),
    .B(_0541_),
    .C(_0607_),
    .Y(_0639_));
 sg13g2_or3_2 _1520_ (.A(_0410_),
    .B(_0541_),
    .C(_0607_),
    .X(_0640_));
 sg13g2_xnor2_1 _1521_ (.Y(_0641_),
    .A(\u8.ruop[2] ),
    .B(net478));
 sg13g2_a21oi_2 _1522_ (.B1(_0410_),
    .Y(_0642_),
    .A2(net487),
    .A1(_0519_));
 sg13g2_o21ai_1 _1523_ (.B1(net545),
    .Y(_0643_),
    .A1(_0518_),
    .A2(_0541_));
 sg13g2_nor2_1 _1524_ (.A(net515),
    .B(net472),
    .Y(_0644_));
 sg13g2_a21oi_2 _1525_ (.B1(_0620_),
    .Y(_0645_),
    .A2(_0588_),
    .A1(_0517_));
 sg13g2_a21o_2 _1526_ (.A2(_0588_),
    .A1(_0517_),
    .B1(_0620_),
    .X(_0646_));
 sg13g2_a21oi_1 _1527_ (.A1(net515),
    .A2(net472),
    .Y(_0647_),
    .B1(\u8.ruop[0] ));
 sg13g2_a21o_1 _1528_ (.A2(_0647_),
    .A1(_0645_),
    .B1(_0644_),
    .X(_0648_));
 sg13g2_a21oi_1 _1529_ (.A1(net515),
    .A2(net472),
    .Y(_0649_),
    .B1(_0392_));
 sg13g2_o21ai_1 _1530_ (.B1(_0649_),
    .Y(_0650_),
    .A1(_0393_),
    .A2(_0645_));
 sg13g2_and2_1 _1531_ (.A(_0035_),
    .B(net478),
    .X(_0651_));
 sg13g2_a22oi_1 _1532_ (.Y(_0652_),
    .B1(_0650_),
    .B2(_0651_),
    .A2(_0648_),
    .A1(_0641_));
 sg13g2_nand2_1 _1533_ (.Y(_0653_),
    .A(net566),
    .B(_0652_));
 sg13g2_o21ai_1 _1534_ (.B1(_0653_),
    .Y(uo_out[6]),
    .A1(net566),
    .A2(_0640_));
 sg13g2_a22oi_1 _1535_ (.Y(_0654_),
    .B1(_0532_),
    .B2(_0537_),
    .A2(_0478_),
    .A1(net547));
 sg13g2_a22oi_1 _1536_ (.Y(_0655_),
    .B1(_0528_),
    .B2(_0536_),
    .A2(_0492_),
    .A1(net553));
 sg13g2_and2_1 _1537_ (.A(_0021_),
    .B(_0629_),
    .X(_0656_));
 sg13g2_a21oi_2 _1538_ (.B1(_0481_),
    .Y(_0657_),
    .A2(_0656_),
    .A1(_0576_));
 sg13g2_a21o_1 _1539_ (.A2(_0656_),
    .A1(_0576_),
    .B1(_0481_),
    .X(_0658_));
 sg13g2_a21oi_1 _1540_ (.A1(net546),
    .A2(_0493_),
    .Y(_0659_),
    .B1(_0410_));
 sg13g2_o21ai_1 _1541_ (.B1(net545),
    .Y(_0660_),
    .A1(_0403_),
    .A2(_0492_));
 sg13g2_nand2_2 _1542_ (.Y(_0661_),
    .A(_0655_),
    .B(net501));
 sg13g2_o21ai_1 _1543_ (.B1(_0661_),
    .Y(_0662_),
    .A1(_0410_),
    .A2(_0654_));
 sg13g2_and2_2 _1544_ (.A(_0657_),
    .B(_0662_),
    .X(_0663_));
 sg13g2_nand2_1 _1545_ (.Y(_0664_),
    .A(_0657_),
    .B(_0662_));
 sg13g2_nand2_1 _1546_ (.Y(_0665_),
    .A(_0411_),
    .B(_0664_));
 sg13g2_or3_1 _1547_ (.A(_0474_),
    .B(_0537_),
    .C(_0655_),
    .X(_0666_));
 sg13g2_a221oi_1 _1548_ (.B2(_0666_),
    .C1(_0596_),
    .B1(_0654_),
    .A1(_0525_),
    .Y(_0667_),
    .A2(_0541_));
 sg13g2_o21ai_1 _1549_ (.B1(net545),
    .Y(_0668_),
    .A1(_0658_),
    .A2(_0667_));
 sg13g2_nor2_1 _1550_ (.A(\u8.rbop[0] ),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_nor2_1 _1551_ (.A(_0411_),
    .B(_0664_),
    .Y(_0670_));
 sg13g2_nand3_1 _1552_ (.B(_0657_),
    .C(_0662_),
    .A(_0411_),
    .Y(_0671_));
 sg13g2_a21o_1 _1553_ (.A2(_0662_),
    .A1(_0657_),
    .B1(_0411_),
    .X(_0672_));
 sg13g2_and2_1 _1554_ (.A(_0671_),
    .B(_0672_),
    .X(_0673_));
 sg13g2_o21ai_1 _1555_ (.B1(_0665_),
    .Y(_0674_),
    .A1(_0669_),
    .A2(_0673_));
 sg13g2_and2_1 _1556_ (.A(_0654_),
    .B(net499),
    .X(_0675_));
 sg13g2_nand2_2 _1557_ (.Y(_0676_),
    .A(_0654_),
    .B(net500));
 sg13g2_and2_1 _1558_ (.A(_0016_),
    .B(_0675_),
    .X(_0677_));
 sg13g2_nand2b_1 _1559_ (.Y(_0678_),
    .B(_0676_),
    .A_N(_0016_));
 sg13g2_nor2b_1 _1560_ (.A(_0677_),
    .B_N(_0678_),
    .Y(_0679_));
 sg13g2_a221oi_1 _1561_ (.B2(_0674_),
    .C1(_0407_),
    .B1(_0679_),
    .A1(\u8.rbop[2] ),
    .Y(_0680_),
    .A2(_0676_));
 sg13g2_a21oi_2 _1562_ (.B1(_0680_),
    .Y(uo_out[7]),
    .A2(_0661_),
    .A1(_0407_));
 sg13g2_nor2_2 _1563_ (.A(net567),
    .B(net6),
    .Y(_0681_));
 sg13g2_nor2_2 _1564_ (.A(net567),
    .B(net4),
    .Y(_0682_));
 sg13g2_or2_2 _1565_ (.X(_0683_),
    .B(net4),
    .A(net567));
 sg13g2_nor2_2 _1566_ (.A(_0681_),
    .B(net559),
    .Y(_0684_));
 sg13g2_a21oi_2 _1567_ (.B1(net567),
    .Y(_0685_),
    .A2(net6),
    .A1(net4));
 sg13g2_or3_1 _1568_ (.A(net567),
    .B(net5),
    .C(_0685_),
    .X(_0686_));
 sg13g2_o21ai_1 _1569_ (.B1(net1),
    .Y(_0687_),
    .A1(_0640_),
    .A2(_0686_));
 sg13g2_o21ai_1 _1570_ (.B1(_0684_),
    .Y(_0688_),
    .A1(net567),
    .A2(net5));
 sg13g2_and2_1 _1571_ (.A(_0544_),
    .B(_0611_),
    .X(_0689_));
 sg13g2_nor2_1 _1572_ (.A(net472),
    .B(_0645_),
    .Y(_0690_));
 sg13g2_nand2_1 _1573_ (.Y(_0691_),
    .A(_0642_),
    .B(_0646_));
 sg13g2_or3_1 _1574_ (.A(net471),
    .B(_0645_),
    .C(_0686_),
    .X(_0692_));
 sg13g2_o21ai_1 _1575_ (.B1(_0688_),
    .Y(_0693_),
    .A1(_0689_),
    .A2(_0692_));
 sg13g2_nand3_1 _1576_ (.B(net14),
    .C(_0521_),
    .A(_0416_),
    .Y(_0694_));
 sg13g2_nand2_1 _1577_ (.Y(_0695_),
    .A(net4),
    .B(_0681_));
 sg13g2_nor2_2 _1578_ (.A(_0660_),
    .B(_0695_),
    .Y(_0696_));
 sg13g2_nand4_1 _1579_ (.B(net14),
    .C(_0521_),
    .A(_0416_),
    .Y(_0697_),
    .D(_0696_));
 sg13g2_inv_1 _1580_ (.Y(_0698_),
    .A(_0697_));
 sg13g2_a21o_1 _1581_ (.A2(_0698_),
    .A1(_0655_),
    .B1(_0693_),
    .X(_0699_));
 sg13g2_and2_1 _1582_ (.A(_0694_),
    .B(_0696_),
    .X(_0700_));
 sg13g2_or2_1 _1583_ (.X(_0701_),
    .B(\u8.rcip[0] ),
    .A(\u8.rcip[1] ));
 sg13g2_nand2_2 _1584_ (.Y(_0702_),
    .A(net95),
    .B(net125));
 sg13g2_nand2_1 _1585_ (.Y(_0703_),
    .A(_0701_),
    .B(_0702_));
 sg13g2_and2_1 _1586_ (.A(\u8.rcip[2] ),
    .B(net559),
    .X(_0704_));
 sg13g2_nand2_1 _1587_ (.Y(_0705_),
    .A(_0703_),
    .B(_0704_));
 sg13g2_o21ai_1 _1588_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_0023_),
    .A2(_0683_));
 sg13g2_nor2_1 _1589_ (.A(_0661_),
    .B(_0697_),
    .Y(_0707_));
 sg13g2_or4_1 _1590_ (.A(_0693_),
    .B(_0700_),
    .C(_0706_),
    .D(_0707_),
    .X(_0708_));
 sg13g2_nor2_2 _1591_ (.A(_0687_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_o21ai_1 _1592_ (.B1(_0681_),
    .Y(_0710_),
    .A1(net14),
    .A2(net501));
 sg13g2_inv_1 _1593_ (.Y(_0711_),
    .A(_0710_));
 sg13g2_nor2_1 _1594_ (.A(net558),
    .B(_0710_),
    .Y(_0712_));
 sg13g2_nor2_2 _1595_ (.A(_0663_),
    .B(_0675_),
    .Y(_0713_));
 sg13g2_nor2_1 _1596_ (.A(_0655_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_o21ai_1 _1597_ (.B1(_0661_),
    .Y(_0715_),
    .A1(_0663_),
    .A2(_0675_));
 sg13g2_nor2_1 _1598_ (.A(net540),
    .B(_0552_),
    .Y(_0716_));
 sg13g2_nand3_1 _1599_ (.B(_0578_),
    .C(_0716_),
    .A(_0559_),
    .Y(_0717_));
 sg13g2_or4_1 _1600_ (.A(_0476_),
    .B(_0487_),
    .C(_0563_),
    .D(_0717_),
    .X(_0718_));
 sg13g2_a21oi_1 _1601_ (.A1(net510),
    .A2(net474),
    .Y(_0719_),
    .B1(net466));
 sg13g2_and4_2 _1602_ (.A(net545),
    .B(_0657_),
    .C(_0662_),
    .D(_0667_),
    .X(_0720_));
 sg13g2_nand3b_1 _1603_ (.B(_0007_),
    .C(_0523_),
    .Y(_0721_),
    .A_N(net529));
 sg13g2_nand3_1 _1604_ (.B(_0592_),
    .C(_0721_),
    .A(_0430_),
    .Y(_0722_));
 sg13g2_nand3_1 _1605_ (.B(_0662_),
    .C(_0676_),
    .A(_0657_),
    .Y(_0723_));
 sg13g2_nand2b_1 _1606_ (.Y(_0724_),
    .B(_0668_),
    .A_N(_0723_));
 sg13g2_inv_1 _1607_ (.Y(_0725_),
    .A(net468));
 sg13g2_nand3_1 _1608_ (.B(net524),
    .C(_0004_),
    .A(net521),
    .Y(_0726_));
 sg13g2_nand3b_1 _1609_ (.B(_0003_),
    .C(_0577_),
    .Y(_0727_),
    .A_N(net533));
 sg13g2_nand2_1 _1610_ (.Y(_0728_),
    .A(net511),
    .B(_0449_));
 sg13g2_o21ai_1 _1611_ (.B1(_0720_),
    .Y(_0729_),
    .A1(net518),
    .A2(_0722_));
 sg13g2_nor4_1 _1612_ (.A(_0005_),
    .B(_0467_),
    .C(_0726_),
    .D(_0728_),
    .Y(_0730_));
 sg13g2_nand3_1 _1613_ (.B(_0727_),
    .C(_0730_),
    .A(_0494_),
    .Y(_0731_));
 sg13g2_nand4_1 _1614_ (.B(_0668_),
    .C(_0676_),
    .A(_0663_),
    .Y(_0732_),
    .D(_0731_));
 sg13g2_nand2_2 _1615_ (.Y(_0733_),
    .A(_0729_),
    .B(_0732_));
 sg13g2_a22oi_1 _1616_ (.Y(_0734_),
    .B1(_0733_),
    .B2(_0431_),
    .A2(_0723_),
    .A1(net510));
 sg13g2_o21ai_1 _1617_ (.B1(net499),
    .Y(_0735_),
    .A1(_0719_),
    .A2(_0734_));
 sg13g2_and2_2 _1618_ (.A(_0640_),
    .B(net472),
    .X(_0736_));
 sg13g2_nand2_2 _1619_ (.Y(_0737_),
    .A(_0640_),
    .B(net472));
 sg13g2_nor2_2 _1620_ (.A(_0645_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_nand2_2 _1621_ (.Y(_0739_),
    .A(_0646_),
    .B(_0736_));
 sg13g2_o21ai_1 _1622_ (.B1(_0646_),
    .Y(_0740_),
    .A1(_0642_),
    .A2(_0736_));
 sg13g2_nand2b_2 _1623_ (.Y(_0741_),
    .B(_0684_),
    .A_N(_0740_));
 sg13g2_nor2_2 _1624_ (.A(\u8.rcip[2] ),
    .B(_0702_),
    .Y(_0742_));
 sg13g2_or2_2 _1625_ (.X(_0743_),
    .B(_0702_),
    .A(\u8.rcip[2] ));
 sg13g2_nor2_2 _1626_ (.A(_0683_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nand2_1 _1627_ (.Y(_0745_),
    .A(net513),
    .B(net575));
 sg13g2_o21ai_1 _1628_ (.B1(_0745_),
    .Y(_0746_),
    .A1(net575),
    .A2(_0425_));
 sg13g2_a22oi_1 _1629_ (.Y(_0747_),
    .B1(_0744_),
    .B2(_0746_),
    .A2(_0735_),
    .A1(net477));
 sg13g2_nand3_1 _1630_ (.B(_0741_),
    .C(_0747_),
    .A(net454),
    .Y(_0748_));
 sg13g2_o21ai_1 _1631_ (.B1(net587),
    .Y(_0749_),
    .A1(net103),
    .A2(net454));
 sg13g2_nor2b_1 _1632_ (.A(_0749_),
    .B_N(_0748_),
    .Y(_0038_));
 sg13g2_nor2_2 _1633_ (.A(net585),
    .B(net8),
    .Y(_0750_));
 sg13g2_a21oi_1 _1634_ (.A1(_0390_),
    .A2(net579),
    .Y(_0751_),
    .B1(_0750_));
 sg13g2_nor2_1 _1635_ (.A(_0663_),
    .B(_0676_),
    .Y(_0752_));
 sg13g2_nor3_2 _1636_ (.A(_0663_),
    .B(_0668_),
    .C(_0676_),
    .Y(_0753_));
 sg13g2_and2_1 _1637_ (.A(_0715_),
    .B(net473),
    .X(_0754_));
 sg13g2_nor3_1 _1638_ (.A(_0733_),
    .B(_0753_),
    .C(_0754_),
    .Y(_0755_));
 sg13g2_and2_2 _1639_ (.A(_0668_),
    .B(_0752_),
    .X(_0756_));
 sg13g2_nand2_1 _1640_ (.Y(_0757_),
    .A(net509),
    .B(_0756_));
 sg13g2_a21oi_1 _1641_ (.A1(net509),
    .A2(_0756_),
    .Y(_0758_),
    .B1(net498));
 sg13g2_o21ai_1 _1642_ (.B1(_0758_),
    .Y(_0759_),
    .A1(_0011_),
    .A2(_0755_));
 sg13g2_a22oi_1 _1643_ (.Y(_0760_),
    .B1(_0759_),
    .B2(net477),
    .A2(_0751_),
    .A1(_0744_));
 sg13g2_o21ai_1 _1644_ (.B1(net590),
    .Y(_0761_),
    .A1(net92),
    .A2(net455));
 sg13g2_a21oi_1 _1645_ (.A1(net455),
    .A2(_0760_),
    .Y(_0039_),
    .B1(_0761_));
 sg13g2_nor2_2 _1646_ (.A(_0681_),
    .B(_0738_),
    .Y(_0762_));
 sg13g2_a21oi_2 _1647_ (.B1(net558),
    .Y(_0763_),
    .A2(_0762_),
    .A1(_0691_));
 sg13g2_nor2_1 _1648_ (.A(_0417_),
    .B(net501),
    .Y(_0764_));
 sg13g2_nor2b_1 _1649_ (.A(_0764_),
    .B_N(_0681_),
    .Y(_0765_));
 sg13g2_o21ai_1 _1650_ (.B1(_0432_),
    .Y(_0766_),
    .A1(_0733_),
    .A2(_0756_));
 sg13g2_nand2_1 _1651_ (.Y(_0767_),
    .A(net507),
    .B(_0723_));
 sg13g2_o21ai_1 _1652_ (.B1(_0766_),
    .Y(_0768_),
    .A1(_0756_),
    .A2(_0767_));
 sg13g2_and2_1 _1653_ (.A(net507),
    .B(net473),
    .X(_0769_));
 sg13g2_o21ai_1 _1654_ (.B1(_0768_),
    .Y(_0770_),
    .A1(net466),
    .A2(_0769_));
 sg13g2_o21ai_1 _1655_ (.B1(net476),
    .Y(_0771_),
    .A1(net498),
    .A2(_0770_));
 sg13g2_nor2_2 _1656_ (.A(net9),
    .B(net582),
    .Y(_0772_));
 sg13g2_a21oi_1 _1657_ (.A1(_0389_),
    .A2(net578),
    .Y(_0773_),
    .B1(_0772_));
 sg13g2_a22oi_1 _1658_ (.Y(_0774_),
    .B1(_0773_),
    .B2(_0744_),
    .A2(_0771_),
    .A1(_0763_));
 sg13g2_o21ai_1 _1659_ (.B1(net589),
    .Y(_0775_),
    .A1(net554),
    .A2(net454));
 sg13g2_a21oi_1 _1660_ (.A1(net454),
    .A2(_0774_),
    .Y(_0040_),
    .B1(_0775_));
 sg13g2_nor2_2 _1661_ (.A(net582),
    .B(net10),
    .Y(_0776_));
 sg13g2_a21oi_1 _1662_ (.A1(_0388_),
    .A2(net578),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_and2_1 _1663_ (.A(net503),
    .B(net473),
    .X(_0778_));
 sg13g2_o21ai_1 _1664_ (.B1(net499),
    .Y(_0779_),
    .A1(net466),
    .A2(_0778_));
 sg13g2_nand3b_1 _1665_ (.B(_0011_),
    .C(_0530_),
    .Y(_0780_),
    .A_N(net518));
 sg13g2_nand4_1 _1666_ (.B(_0013_),
    .C(_0475_),
    .A(_0414_),
    .Y(_0781_),
    .D(_0780_));
 sg13g2_a21o_1 _1667_ (.A2(_0781_),
    .A1(_0756_),
    .B1(_0733_),
    .X(_0782_));
 sg13g2_a221oi_1 _1668_ (.B2(_0414_),
    .C1(_0715_),
    .B1(_0782_),
    .A1(net503),
    .Y(_0783_),
    .A2(_0753_));
 sg13g2_o21ai_1 _1669_ (.B1(net476),
    .Y(_0784_),
    .A1(_0779_),
    .A2(_0783_));
 sg13g2_a22oi_1 _1670_ (.Y(_0785_),
    .B1(_0784_),
    .B2(_0763_),
    .A2(_0777_),
    .A1(_0744_));
 sg13g2_o21ai_1 _1671_ (.B1(net587),
    .Y(_0786_),
    .A1(net553),
    .A2(net454));
 sg13g2_a21oi_1 _1672_ (.A1(net454),
    .A2(_0785_),
    .Y(_0041_),
    .B1(_0786_));
 sg13g2_or2_1 _1673_ (.X(_0787_),
    .B(_0782_),
    .A(_0753_));
 sg13g2_nand3b_1 _1674_ (.B(_0019_),
    .C(_0534_),
    .Y(_0788_),
    .A_N(net507));
 sg13g2_nand4_1 _1675_ (.B(_0436_),
    .C(_0496_),
    .A(_0406_),
    .Y(_0789_),
    .D(_0788_));
 sg13g2_a21o_1 _1676_ (.A2(_0789_),
    .A1(_0753_),
    .B1(_0715_),
    .X(_0790_));
 sg13g2_a21oi_1 _1677_ (.A1(_0433_),
    .A2(_0787_),
    .Y(_0791_),
    .B1(_0790_));
 sg13g2_and2_1 _1678_ (.A(\u8.rc[22] ),
    .B(net475),
    .X(_0792_));
 sg13g2_o21ai_1 _1679_ (.B1(net500),
    .Y(_0793_),
    .A1(_0714_),
    .A2(_0792_));
 sg13g2_o21ai_1 _1680_ (.B1(net476),
    .Y(_0794_),
    .A1(_0791_),
    .A2(_0793_));
 sg13g2_or2_1 _1681_ (.X(_0795_),
    .B(net11),
    .A(net578));
 sg13g2_mux2_1 _1682_ (.A0(net11),
    .A1(net506),
    .S(net579),
    .X(_0796_));
 sg13g2_a22oi_1 _1683_ (.Y(_0797_),
    .B1(_0796_),
    .B2(_0744_),
    .A2(_0794_),
    .A1(_0763_));
 sg13g2_o21ai_1 _1684_ (.B1(net590),
    .Y(_0798_),
    .A1(net552),
    .A2(net455));
 sg13g2_a21oi_1 _1685_ (.A1(net455),
    .A2(_0797_),
    .Y(_0042_),
    .B1(_0798_));
 sg13g2_a21oi_1 _1686_ (.A1(_0434_),
    .A2(net473),
    .Y(_0799_),
    .B1(net466));
 sg13g2_a21oi_1 _1687_ (.A1(_0434_),
    .A2(_0787_),
    .Y(_0800_),
    .B1(_0790_));
 sg13g2_o21ai_1 _1688_ (.B1(net499),
    .Y(_0801_),
    .A1(_0799_),
    .A2(_0800_));
 sg13g2_nor2_2 _1689_ (.A(net582),
    .B(net12),
    .Y(_0802_));
 sg13g2_a21oi_1 _1690_ (.A1(_0387_),
    .A2(net579),
    .Y(_0803_),
    .B1(_0802_));
 sg13g2_a22oi_1 _1691_ (.Y(_0804_),
    .B1(_0803_),
    .B2(_0744_),
    .A2(_0801_),
    .A1(net477));
 sg13g2_o21ai_1 _1692_ (.B1(net590),
    .Y(_0805_),
    .A1(net551),
    .A2(net455));
 sg13g2_a21oi_1 _1693_ (.A1(net455),
    .A2(_0804_),
    .Y(_0043_),
    .B1(_0805_));
 sg13g2_a21oi_1 _1694_ (.A1(_0435_),
    .A2(_0787_),
    .Y(_0806_),
    .B1(_0790_));
 sg13g2_nand3_1 _1695_ (.B(net499),
    .C(net473),
    .A(\u8.rc[24] ),
    .Y(_0807_));
 sg13g2_and2_1 _1696_ (.A(_0715_),
    .B(_0807_),
    .X(_0808_));
 sg13g2_o21ai_1 _1697_ (.B1(net476),
    .Y(_0809_),
    .A1(_0806_),
    .A2(_0808_));
 sg13g2_nor2_2 _1698_ (.A(net13),
    .B(net582),
    .Y(_0810_));
 sg13g2_a21oi_1 _1699_ (.A1(_0386_),
    .A2(net578),
    .Y(_0811_),
    .B1(_0810_));
 sg13g2_a22oi_1 _1700_ (.Y(_0812_),
    .B1(_0811_),
    .B2(_0744_),
    .A2(_0809_),
    .A1(_0763_));
 sg13g2_o21ai_1 _1701_ (.B1(net587),
    .Y(_0813_),
    .A1(net550),
    .A2(net454));
 sg13g2_a21oi_1 _1702_ (.A1(net454),
    .A2(_0812_),
    .Y(_0044_),
    .B1(_0813_));
 sg13g2_nand3_1 _1703_ (.B(net499),
    .C(net473),
    .A(net555),
    .Y(_0814_));
 sg13g2_and2_1 _1704_ (.A(_0715_),
    .B(_0814_),
    .X(_0815_));
 sg13g2_a21oi_1 _1705_ (.A1(_0413_),
    .A2(_0782_),
    .Y(_0816_),
    .B1(_0790_));
 sg13g2_o21ai_1 _1706_ (.B1(net476),
    .Y(_0817_),
    .A1(_0815_),
    .A2(_0816_));
 sg13g2_nor2_2 _1707_ (.A(net14),
    .B(net581),
    .Y(_0818_));
 sg13g2_a21oi_1 _1708_ (.A1(_0385_),
    .A2(net578),
    .Y(_0819_),
    .B1(_0818_));
 sg13g2_a22oi_1 _1709_ (.Y(_0820_),
    .B1(_0819_),
    .B2(_0744_),
    .A2(_0817_),
    .A1(_0763_));
 sg13g2_o21ai_1 _1710_ (.B1(net590),
    .Y(_0821_),
    .A1(net548),
    .A2(net455));
 sg13g2_a21oi_1 _1711_ (.A1(net455),
    .A2(_0820_),
    .Y(_0045_),
    .B1(_0821_));
 sg13g2_nor2_1 _1712_ (.A(net501),
    .B(_0695_),
    .Y(_0822_));
 sg13g2_and3_1 _1713_ (.X(_0823_),
    .A(_0023_),
    .B(net559),
    .C(_0701_));
 sg13g2_nor2_2 _1714_ (.A(\u8.rcip[2] ),
    .B(_0701_),
    .Y(_0824_));
 sg13g2_nand2_2 _1715_ (.Y(_0825_),
    .A(net559),
    .B(_0824_));
 sg13g2_nand3_1 _1716_ (.B(_0688_),
    .C(_0825_),
    .A(net1),
    .Y(_0826_));
 sg13g2_a21oi_1 _1717_ (.A1(net581),
    .A2(_0034_),
    .Y(_0827_),
    .B1(_0810_));
 sg13g2_o21ai_1 _1718_ (.B1(_0795_),
    .Y(_0828_),
    .A1(net562),
    .A2(_0422_));
 sg13g2_a21oi_1 _1719_ (.A1(net582),
    .A2(_0033_),
    .Y(_0829_),
    .B1(_0802_));
 sg13g2_a21oi_2 _1720_ (.B1(_0776_),
    .Y(_0830_),
    .A2(_0031_),
    .A1(net583));
 sg13g2_nand2b_1 _1721_ (.Y(_0831_),
    .B(_0830_),
    .A_N(_0829_));
 sg13g2_a21oi_2 _1722_ (.B1(_0818_),
    .Y(_0832_),
    .A2(net578),
    .A1(_0021_));
 sg13g2_a21o_1 _1723_ (.A2(net581),
    .A1(_0030_),
    .B1(_0772_),
    .X(_0833_));
 sg13g2_nand2_1 _1724_ (.Y(_0834_),
    .A(_0827_),
    .B(_0832_));
 sg13g2_nor4_1 _1725_ (.A(_0828_),
    .B(_0831_),
    .C(_0833_),
    .D(_0834_),
    .Y(_0835_));
 sg13g2_or2_1 _1726_ (.X(_0836_),
    .B(net486),
    .A(net471));
 sg13g2_a221oi_1 _1727_ (.B2(_0645_),
    .C1(_0736_),
    .B1(_0836_),
    .A1(_0689_),
    .Y(_0837_),
    .A2(net457));
 sg13g2_nor2_1 _1728_ (.A(_0686_),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_nor4_1 _1729_ (.A(_0822_),
    .B(_0823_),
    .C(_0826_),
    .D(_0838_),
    .Y(_0839_));
 sg13g2_a21oi_1 _1730_ (.A1(_0697_),
    .A2(_0839_),
    .Y(_0840_),
    .B1(net77));
 sg13g2_nor2b_1 _1731_ (.A(_0840_),
    .B_N(net591),
    .Y(_0046_));
 sg13g2_nor2_2 _1732_ (.A(_0407_),
    .B(net4),
    .Y(_0841_));
 sg13g2_nand2b_2 _1733_ (.Y(_0842_),
    .B(net565),
    .A_N(net4));
 sg13g2_nand2_1 _1734_ (.Y(_0843_),
    .A(net564),
    .B(_0408_));
 sg13g2_inv_1 _1735_ (.Y(_0844_),
    .A(_0843_));
 sg13g2_nand2b_2 _1736_ (.Y(_0845_),
    .B(_0843_),
    .A_N(_0652_));
 sg13g2_nand2_1 _1737_ (.Y(_0846_),
    .A(\u8.ruop[0] ),
    .B(_0035_));
 sg13g2_nor2_1 _1738_ (.A(net515),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_or2_1 _1739_ (.X(_0848_),
    .B(_0846_),
    .A(net516));
 sg13g2_nand2_1 _1740_ (.Y(_0849_),
    .A(net570),
    .B(_0001_));
 sg13g2_nor2_2 _1741_ (.A(net575),
    .B(_0426_),
    .Y(_0850_));
 sg13g2_a21oi_1 _1742_ (.A1(net575),
    .A2(_0001_),
    .Y(_0851_),
    .B1(_0850_));
 sg13g2_nand2_1 _1743_ (.Y(_0852_),
    .A(_0848_),
    .B(_0851_));
 sg13g2_mux2_1 _1744_ (.A0(_0001_),
    .A1(_0000_),
    .S(net576),
    .X(_0853_));
 sg13g2_o21ai_1 _1745_ (.B1(_0852_),
    .Y(_0854_),
    .A1(net495),
    .A2(_0853_));
 sg13g2_xnor2_1 _1746_ (.Y(_0855_),
    .A(_0431_),
    .B(_0529_));
 sg13g2_nand2_1 _1747_ (.Y(_0856_),
    .A(net561),
    .B(_0855_));
 sg13g2_and2_2 _1748_ (.A(net580),
    .B(_0004_),
    .X(_0857_));
 sg13g2_nor2_1 _1749_ (.A(net495),
    .B(_0857_),
    .Y(_0858_));
 sg13g2_and3_2 _1750_ (.X(_0859_),
    .A(net516),
    .B(\u8.ruop[0] ),
    .C(_0035_));
 sg13g2_nand3_1 _1751_ (.B(\u8.ruop[0] ),
    .C(_0035_),
    .A(net515),
    .Y(_0860_));
 sg13g2_nor2_1 _1752_ (.A(_0853_),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_nand2_2 _1753_ (.Y(_0862_),
    .A(_0392_),
    .B(net516));
 sg13g2_and2_1 _1754_ (.A(net495),
    .B(_0862_),
    .X(_0863_));
 sg13g2_nand2_2 _1755_ (.Y(_0864_),
    .A(net494),
    .B(_0862_));
 sg13g2_and3_1 _1756_ (.X(_0865_),
    .A(net515),
    .B(_0393_),
    .C(_0035_));
 sg13g2_nand3_1 _1757_ (.B(_0393_),
    .C(_0035_),
    .A(net515),
    .Y(_0866_));
 sg13g2_nor2b_1 _1758_ (.A(net575),
    .B_N(_0004_),
    .Y(_0867_));
 sg13g2_a21oi_1 _1759_ (.A1(net573),
    .A2(_0855_),
    .Y(_0868_),
    .B1(_0867_));
 sg13g2_a221oi_1 _1760_ (.B2(_0851_),
    .C1(_0861_),
    .B1(net493),
    .A1(_0856_),
    .Y(_0869_),
    .A2(_0858_));
 sg13g2_nand2_1 _1761_ (.Y(_0870_),
    .A(_0863_),
    .B(_0868_));
 sg13g2_o21ai_1 _1762_ (.B1(_0870_),
    .Y(_0871_),
    .A1(_0863_),
    .A2(_0869_));
 sg13g2_a22oi_1 _1763_ (.Y(_0872_),
    .B1(_0871_),
    .B2(_0639_),
    .A2(net465),
    .A1(_0426_));
 sg13g2_a221oi_1 _1764_ (.B2(_0517_),
    .C1(_0620_),
    .B1(_0588_),
    .A1(_0519_),
    .Y(_0873_),
    .A2(net487));
 sg13g2_mux2_1 _1765_ (.A0(_0001_),
    .A1(_0009_),
    .S(net570),
    .X(_0874_));
 sg13g2_xnor2_1 _1766_ (.Y(_0875_),
    .A(net516),
    .B(net98));
 sg13g2_nand2_2 _1767_ (.Y(_0876_),
    .A(net494),
    .B(_0866_));
 sg13g2_inv_1 _1768_ (.Y(_0877_),
    .A(_0876_));
 sg13g2_o21ai_1 _1769_ (.B1(_0849_),
    .Y(_0878_),
    .A1(net570),
    .A2(_0430_));
 sg13g2_nor2_1 _1770_ (.A(net495),
    .B(_0878_),
    .Y(_0879_));
 sg13g2_a21oi_1 _1771_ (.A1(\u8.ls[0] ),
    .A2(net493),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_o21ai_1 _1772_ (.B1(_0880_),
    .Y(_0881_),
    .A1(_0874_),
    .A2(_0876_));
 sg13g2_a22oi_1 _1773_ (.Y(_0882_),
    .B1(net461),
    .B2(_0881_),
    .A2(_0854_),
    .A1(net459));
 sg13g2_a21oi_1 _1774_ (.A1(_0872_),
    .A2(_0882_),
    .Y(_0883_),
    .B1(_0845_));
 sg13g2_a22oi_1 _1775_ (.Y(_0884_),
    .B1(_0671_),
    .B2(_0672_),
    .A2(_0668_),
    .A1(\u8.rbop[0] ));
 sg13g2_o21ai_1 _1776_ (.B1(_0677_),
    .Y(_0885_),
    .A1(_0670_),
    .A2(_0884_));
 sg13g2_or3_1 _1777_ (.A(_0670_),
    .B(_0677_),
    .C(_0884_),
    .X(_0886_));
 sg13g2_nand3_1 _1778_ (.B(_0885_),
    .C(_0886_),
    .A(_0678_),
    .Y(_0887_));
 sg13g2_xor2_1 _1779_ (.B(_0668_),
    .A(\u8.rbop[0] ),
    .X(_0888_));
 sg13g2_and2_1 _1780_ (.A(_0673_),
    .B(_0888_),
    .X(_0889_));
 sg13g2_or2_2 _1781_ (.X(_0890_),
    .B(_0889_),
    .A(_0885_));
 sg13g2_and4_1 _1782_ (.A(\u8.rbop[0] ),
    .B(_0668_),
    .C(_0671_),
    .D(_0672_),
    .X(_0891_));
 sg13g2_nor2_1 _1783_ (.A(_0884_),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_nand4_1 _1784_ (.B(_0885_),
    .C(_0886_),
    .A(_0678_),
    .Y(_0893_),
    .D(_0892_));
 sg13g2_nand3_1 _1785_ (.B(_0890_),
    .C(_0893_),
    .A(_0426_),
    .Y(_0894_));
 sg13g2_and4_2 _1786_ (.A(_0678_),
    .B(_0885_),
    .C(_0886_),
    .D(_0889_),
    .X(_0895_));
 sg13g2_nor3_1 _1787_ (.A(_0884_),
    .B(_0888_),
    .C(_0891_),
    .Y(_0896_));
 sg13g2_and4_2 _1788_ (.A(_0678_),
    .B(_0885_),
    .C(_0886_),
    .D(_0896_),
    .X(_0897_));
 sg13g2_nor2_1 _1789_ (.A(_0885_),
    .B(_0888_),
    .Y(_0898_));
 sg13g2_nor3_2 _1790_ (.A(_0669_),
    .B(_0673_),
    .C(_0885_),
    .Y(_0899_));
 sg13g2_nor2_1 _1791_ (.A(\u8.rbop[1] ),
    .B(\u8.rbop[0] ),
    .Y(_0900_));
 sg13g2_and2_1 _1792_ (.A(_0016_),
    .B(_0900_),
    .X(_0901_));
 sg13g2_nand2_1 _1793_ (.Y(_0902_),
    .A(_0016_),
    .B(_0900_));
 sg13g2_a22oi_1 _1794_ (.Y(_0903_),
    .B1(_0899_),
    .B2(net510),
    .A2(_0898_),
    .A1(_0435_));
 sg13g2_a22oi_1 _1795_ (.Y(_0904_),
    .B1(_0897_),
    .B2(net526),
    .A2(_0895_),
    .A1(net539));
 sg13g2_nand4_1 _1796_ (.B(net491),
    .C(_0903_),
    .A(_0894_),
    .Y(_0905_),
    .D(_0904_));
 sg13g2_and2_2 _1797_ (.A(_0408_),
    .B(_0680_),
    .X(_0906_));
 sg13g2_nor2_1 _1798_ (.A(_0034_),
    .B(net468),
    .Y(_0907_));
 sg13g2_a221oi_1 _1799_ (.B2(\u8.rc[24] ),
    .C1(_0907_),
    .B1(_0753_),
    .A1(net526),
    .Y(_0908_),
    .A2(_0720_));
 sg13g2_nand4_1 _1800_ (.B(net549),
    .C(net545),
    .A(_0403_),
    .Y(_0909_),
    .D(_0655_));
 sg13g2_a221oi_1 _1801_ (.B2(net510),
    .C1(net491),
    .B1(_0756_),
    .A1(_0426_),
    .Y(_0910_),
    .A2(_0713_));
 sg13g2_nand3_1 _1802_ (.B(_0909_),
    .C(_0910_),
    .A(_0908_),
    .Y(_0911_));
 sg13g2_and3_1 _1803_ (.X(_0912_),
    .A(_0905_),
    .B(_0906_),
    .C(_0911_));
 sg13g2_o21ai_1 _1804_ (.B1(_0842_),
    .Y(_0913_),
    .A1(_0883_),
    .A2(_0912_));
 sg13g2_and3_2 _1805_ (.X(_0914_),
    .A(_0408_),
    .B(_0680_),
    .C(_0842_));
 sg13g2_and3_1 _1806_ (.X(_0915_),
    .A(_0887_),
    .B(_0890_),
    .C(net490));
 sg13g2_nand2_1 _1807_ (.Y(_0916_),
    .A(_0012_),
    .B(_0841_));
 sg13g2_nand3_1 _1808_ (.B(net105),
    .C(_0841_),
    .A(\u8.rcop[0] ),
    .Y(_0917_));
 sg13g2_nor2_1 _1809_ (.A(_0395_),
    .B(net106),
    .Y(_0918_));
 sg13g2_nor3_1 _1810_ (.A(_0394_),
    .B(_0395_),
    .C(_0917_),
    .Y(_0919_));
 sg13g2_nand2b_1 _1811_ (.Y(_0920_),
    .B(net564),
    .A_N(net5));
 sg13g2_nand3_1 _1812_ (.B(_0843_),
    .C(_0920_),
    .A(_0842_),
    .Y(_0921_));
 sg13g2_nand2b_1 _1813_ (.Y(_0922_),
    .B(_0921_),
    .A_N(_0919_));
 sg13g2_a21oi_1 _1814_ (.A1(_0914_),
    .A2(_0915_),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_nand2_1 _1815_ (.Y(_0924_),
    .A(_0866_),
    .B(net460));
 sg13g2_nor2b_1 _1816_ (.A(net515),
    .B_N(_0035_),
    .Y(_0925_));
 sg13g2_a22oi_1 _1817_ (.Y(_0926_),
    .B1(_0925_),
    .B2(_0739_),
    .A2(_0924_),
    .A1(_0740_));
 sg13g2_a21oi_1 _1818_ (.A1(\u8.ruop[2] ),
    .A2(net478),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_a21o_1 _1819_ (.A2(net478),
    .A1(\u8.ruop[2] ),
    .B1(_0926_),
    .X(_0928_));
 sg13g2_nor4_2 _1820_ (.A(_0652_),
    .B(_0841_),
    .C(_0844_),
    .Y(_0929_),
    .D(_0920_));
 sg13g2_or4_1 _1821_ (.A(_0652_),
    .B(_0841_),
    .C(_0844_),
    .D(_0920_),
    .X(_0930_));
 sg13g2_a221oi_1 _1822_ (.B2(_0929_),
    .C1(_0922_),
    .B1(_0928_),
    .A1(_0914_),
    .Y(_0931_),
    .A2(_0915_));
 sg13g2_o21ai_1 _1823_ (.B1(_0923_),
    .Y(_0932_),
    .A1(_0927_),
    .A2(_0930_));
 sg13g2_nor3_1 _1824_ (.A(_0394_),
    .B(\u8.rcop[1] ),
    .C(\u8.rcop[0] ),
    .Y(_0933_));
 sg13g2_nor2_1 _1825_ (.A(_0916_),
    .B(_0933_),
    .Y(_0934_));
 sg13g2_nand3_1 _1826_ (.B(\u8.rcop[0] ),
    .C(_0012_),
    .A(_0395_),
    .Y(_0935_));
 sg13g2_nand3b_1 _1827_ (.B(_0012_),
    .C(\u8.rcop[1] ),
    .Y(_0936_),
    .A_N(\u8.rcop[0] ));
 sg13g2_and3_2 _1828_ (.X(_0937_),
    .A(_0394_),
    .B(\u8.rcop[1] ),
    .C(\u8.rcop[0] ));
 sg13g2_nand3_1 _1829_ (.B(\u8.rcop[1] ),
    .C(\u8.rcop[0] ),
    .A(_0394_),
    .Y(_0938_));
 sg13g2_and3_2 _1830_ (.X(_0939_),
    .A(net489),
    .B(net502),
    .C(_0938_));
 sg13g2_a21oi_1 _1831_ (.A1(net570),
    .A2(_0019_),
    .Y(_0940_),
    .B1(_0850_));
 sg13g2_nor2_1 _1832_ (.A(_0874_),
    .B(net489),
    .Y(_0941_));
 sg13g2_mux2_1 _1833_ (.A0(\u8.rc[24] ),
    .A1(\u8.ls[0] ),
    .S(net571),
    .X(_0942_));
 sg13g2_a221oi_1 _1834_ (.B2(_0937_),
    .C1(_0941_),
    .B1(_0942_),
    .A1(_0939_),
    .Y(_0943_),
    .A2(_0940_));
 sg13g2_o21ai_1 _1835_ (.B1(_0943_),
    .Y(_0944_),
    .A1(_0878_),
    .A2(_0936_));
 sg13g2_a21oi_2 _1836_ (.B1(_0932_),
    .Y(_0945_),
    .A2(_0944_),
    .A1(_0934_));
 sg13g2_and2_1 _1837_ (.A(net1),
    .B(net588),
    .X(_0946_));
 sg13g2_nand2_2 _1838_ (.Y(_0947_),
    .A(net1),
    .B(net588));
 sg13g2_o21ai_1 _1839_ (.B1(net557),
    .Y(_0948_),
    .A1(net90),
    .A2(_0931_));
 sg13g2_a21oi_1 _1840_ (.A1(_0913_),
    .A2(_0945_),
    .Y(_0047_),
    .B1(_0948_));
 sg13g2_mux2_1 _1841_ (.A0(_0003_),
    .A1(_0028_),
    .S(net575),
    .X(_0949_));
 sg13g2_and2_1 _1842_ (.A(net570),
    .B(_0003_),
    .X(_0950_));
 sg13g2_nor2_1 _1843_ (.A(_0415_),
    .B(net570),
    .Y(_0951_));
 sg13g2_nor2_1 _1844_ (.A(_0950_),
    .B(_0951_),
    .Y(_0952_));
 sg13g2_a22oi_1 _1845_ (.Y(_0953_),
    .B1(_0952_),
    .B2(net497),
    .A2(net493),
    .A1(\u8.ls[1] ));
 sg13g2_o21ai_1 _1846_ (.B1(_0953_),
    .Y(_0954_),
    .A1(_0876_),
    .A2(_0949_));
 sg13g2_mux2_1 _1847_ (.A0(_0003_),
    .A1(_0002_),
    .S(net576),
    .X(_0955_));
 sg13g2_nor2_2 _1848_ (.A(net576),
    .B(_0428_),
    .Y(_0956_));
 sg13g2_nor2_1 _1849_ (.A(_0950_),
    .B(_0956_),
    .Y(_0957_));
 sg13g2_nor2_1 _1850_ (.A(net497),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_a21oi_1 _1851_ (.A1(net497),
    .A2(_0955_),
    .Y(_0959_),
    .B1(_0958_));
 sg13g2_nor2b_1 _1852_ (.A(net569),
    .B_N(_0005_),
    .Y(_0960_));
 sg13g2_xor2_1 _1853_ (.B(_0530_),
    .A(_0011_),
    .X(_0961_));
 sg13g2_a21oi_1 _1854_ (.A1(net568),
    .A2(_0961_),
    .Y(_0962_),
    .B1(_0960_));
 sg13g2_nor2_1 _1855_ (.A(_0864_),
    .B(_0962_),
    .Y(_0963_));
 sg13g2_nand2_1 _1856_ (.Y(_0964_),
    .A(net561),
    .B(_0961_));
 sg13g2_and2_2 _1857_ (.A(net579),
    .B(_0005_),
    .X(_0965_));
 sg13g2_nor2_1 _1858_ (.A(net494),
    .B(_0965_),
    .Y(_0966_));
 sg13g2_o21ai_1 _1859_ (.B1(_0864_),
    .Y(_0967_),
    .A1(_0860_),
    .A2(_0955_));
 sg13g2_a221oi_1 _1860_ (.B2(_0966_),
    .C1(_0967_),
    .B1(_0964_),
    .A1(net493),
    .Y(_0968_),
    .A2(_0957_));
 sg13g2_nor3_1 _1861_ (.A(_0640_),
    .B(_0963_),
    .C(_0968_),
    .Y(_0969_));
 sg13g2_a21o_1 _1862_ (.A2(_0954_),
    .A1(net461),
    .B1(_0969_),
    .X(_0970_));
 sg13g2_a221oi_1 _1863_ (.B2(net459),
    .C1(_0970_),
    .B1(_0959_),
    .A1(_0428_),
    .Y(_0971_),
    .A2(net465));
 sg13g2_or3_1 _1864_ (.A(_0652_),
    .B(_0844_),
    .C(_0971_),
    .X(_0972_));
 sg13g2_nand3_1 _1865_ (.B(_0890_),
    .C(_0893_),
    .A(_0428_),
    .Y(_0973_));
 sg13g2_a22oi_1 _1866_ (.Y(_0974_),
    .B1(_0899_),
    .B2(net509),
    .A2(_0898_),
    .A1(_0413_));
 sg13g2_a22oi_1 _1867_ (.Y(_0975_),
    .B1(_0897_),
    .B2(net523),
    .A2(_0895_),
    .A1(net536));
 sg13g2_and4_1 _1868_ (.A(net491),
    .B(_0973_),
    .C(_0974_),
    .D(_0975_),
    .X(_0976_));
 sg13g2_nor2_1 _1869_ (.A(_0021_),
    .B(net468),
    .Y(_0977_));
 sg13g2_a21oi_1 _1870_ (.A1(_0428_),
    .A2(_0713_),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_a22oi_1 _1871_ (.Y(_0979_),
    .B1(_0753_),
    .B2(net555),
    .A2(_0720_),
    .A1(net523));
 sg13g2_nand4_1 _1872_ (.B(_0901_),
    .C(_0978_),
    .A(_0757_),
    .Y(_0980_),
    .D(_0979_));
 sg13g2_nand2_1 _1873_ (.Y(_0981_),
    .A(_0906_),
    .B(_0980_));
 sg13g2_o21ai_1 _1874_ (.B1(_0972_),
    .Y(_0982_),
    .A1(_0976_),
    .A2(_0981_));
 sg13g2_a21oi_1 _1875_ (.A1(_0026_),
    .A2(net570),
    .Y(_0983_),
    .B1(_0956_));
 sg13g2_nor3_1 _1876_ (.A(net502),
    .B(_0950_),
    .C(_0951_),
    .Y(_0984_));
 sg13g2_nand2_2 _1877_ (.Y(_0985_),
    .A(\u8.ls[1] ),
    .B(net584));
 sg13g2_o21ai_1 _1878_ (.B1(_0985_),
    .Y(_0986_),
    .A1(_0406_),
    .A2(net586));
 sg13g2_a221oi_1 _1879_ (.B2(_0937_),
    .C1(_0984_),
    .B1(_0986_),
    .A1(_0939_),
    .Y(_0987_),
    .A2(_0983_));
 sg13g2_o21ai_1 _1880_ (.B1(_0987_),
    .Y(_0988_),
    .A1(_0935_),
    .A2(_0949_));
 sg13g2_a221oi_1 _1881_ (.B2(net481),
    .C1(_0932_),
    .B1(_0988_),
    .A1(_0842_),
    .Y(_0989_),
    .A2(_0982_));
 sg13g2_o21ai_1 _1882_ (.B1(net557),
    .Y(_0990_),
    .A1(net88),
    .A2(net453));
 sg13g2_nor2_1 _1883_ (.A(_0989_),
    .B(_0990_),
    .Y(_0048_));
 sg13g2_a21oi_1 _1884_ (.A1(_0030_),
    .A2(net573),
    .Y(_0991_),
    .B1(_0867_));
 sg13g2_nor2b_2 _1885_ (.A(net576),
    .B_N(_0030_),
    .Y(_0992_));
 sg13g2_nor3_1 _1886_ (.A(net496),
    .B(_0857_),
    .C(_0992_),
    .Y(_0993_));
 sg13g2_a21o_1 _1887_ (.A2(_0991_),
    .A1(net496),
    .B1(_0993_),
    .X(_0994_));
 sg13g2_a21oi_1 _1888_ (.A1(net560),
    .A2(_0010_),
    .Y(_0995_),
    .B1(_0857_));
 sg13g2_a21o_1 _1889_ (.A2(_0010_),
    .A1(net574),
    .B1(_0867_),
    .X(_0996_));
 sg13g2_a22oi_1 _1890_ (.Y(_0997_),
    .B1(_0995_),
    .B2(net496),
    .A2(net492),
    .A1(net544));
 sg13g2_o21ai_1 _1891_ (.B1(_0997_),
    .Y(_0998_),
    .A1(_0876_),
    .A2(_0996_));
 sg13g2_nor2_1 _1892_ (.A(net544),
    .B(net574),
    .Y(_0999_));
 sg13g2_o21ai_1 _1893_ (.B1(_0859_),
    .Y(_1000_),
    .A1(net544),
    .A2(net560));
 sg13g2_o21ai_1 _1894_ (.B1(_1000_),
    .Y(_1001_),
    .A1(_0866_),
    .A2(_0999_));
 sg13g2_nor2_1 _1895_ (.A(net573),
    .B(_0864_),
    .Y(_1002_));
 sg13g2_a21oi_2 _1896_ (.B1(_1002_),
    .Y(_1003_),
    .A2(net496),
    .A1(net573));
 sg13g2_inv_1 _1897_ (.Y(_1004_),
    .A(_1003_));
 sg13g2_a22oi_1 _1898_ (.Y(_1005_),
    .B1(_1004_),
    .B2(net526),
    .A2(_1001_),
    .A1(_0864_));
 sg13g2_nor2_1 _1899_ (.A(_0640_),
    .B(_1005_),
    .Y(_1006_));
 sg13g2_a221oi_1 _1900_ (.B2(net460),
    .C1(_1006_),
    .B1(_0998_),
    .A1(net459),
    .Y(_1007_),
    .A2(_0994_));
 sg13g2_o21ai_1 _1901_ (.B1(_1007_),
    .Y(_1008_),
    .A1(_0030_),
    .A2(_0737_));
 sg13g2_nor2b_1 _1902_ (.A(_0845_),
    .B_N(_1008_),
    .Y(_1009_));
 sg13g2_nand3b_1 _1903_ (.B(_0890_),
    .C(_0893_),
    .Y(_1010_),
    .A_N(_0030_));
 sg13g2_a22oi_1 _1904_ (.Y(_1011_),
    .B1(_0899_),
    .B2(net507),
    .A2(_0898_),
    .A1(_0436_));
 sg13g2_a22oi_1 _1905_ (.Y(_1012_),
    .B1(_0897_),
    .B2(net519),
    .A2(_0895_),
    .A1(net535));
 sg13g2_nand4_1 _1906_ (.B(_1010_),
    .C(_1011_),
    .A(net490),
    .Y(_1013_),
    .D(_1012_));
 sg13g2_nor2_1 _1907_ (.A(_0001_),
    .B(net468),
    .Y(_1014_));
 sg13g2_a21oi_1 _1908_ (.A1(net519),
    .A2(_0720_),
    .Y(_1015_),
    .B1(_1014_));
 sg13g2_a221oi_1 _1909_ (.B2(net507),
    .C1(_0715_),
    .B1(_0756_),
    .A1(net554),
    .Y(_1016_),
    .A2(_0753_));
 sg13g2_a22oi_1 _1910_ (.Y(_1017_),
    .B1(_1015_),
    .B2(_1016_),
    .A2(_0713_),
    .A1(_0030_));
 sg13g2_o21ai_1 _1911_ (.B1(_0906_),
    .Y(_1018_),
    .A1(net491),
    .A2(_1017_));
 sg13g2_nor2b_1 _1912_ (.A(_1018_),
    .B_N(_1013_),
    .Y(_1019_));
 sg13g2_o21ai_1 _1913_ (.B1(_0842_),
    .Y(_1020_),
    .A1(_1009_),
    .A2(_1019_));
 sg13g2_a21oi_1 _1914_ (.A1(net571),
    .A2(_0018_),
    .Y(_1021_),
    .B1(_0992_));
 sg13g2_and2_1 _1915_ (.A(\u8.ls[2] ),
    .B(net583),
    .X(_1022_));
 sg13g2_a21oi_1 _1916_ (.A1(net554),
    .A2(net562),
    .Y(_1023_),
    .B1(_1022_));
 sg13g2_nand2b_1 _1917_ (.Y(_1024_),
    .B(_0995_),
    .A_N(net502));
 sg13g2_o21ai_1 _1918_ (.B1(_1024_),
    .Y(_1025_),
    .A1(net489),
    .A2(_0996_));
 sg13g2_a21oi_1 _1919_ (.A1(_0939_),
    .A2(_1021_),
    .Y(_1026_),
    .B1(_1025_));
 sg13g2_o21ai_1 _1920_ (.B1(_1026_),
    .Y(_1027_),
    .A1(_0938_),
    .A2(_1023_));
 sg13g2_a21oi_1 _1921_ (.A1(net481),
    .A2(_1027_),
    .Y(_1028_),
    .B1(_0932_));
 sg13g2_o21ai_1 _1922_ (.B1(net557),
    .Y(_1029_),
    .A1(net85),
    .A2(net453));
 sg13g2_a21oi_1 _1923_ (.A1(_1020_),
    .A2(_1028_),
    .Y(_0049_),
    .B1(_1029_));
 sg13g2_a21oi_1 _1924_ (.A1(net568),
    .A2(_0031_),
    .Y(_1030_),
    .B1(_0960_));
 sg13g2_nor2_2 _1925_ (.A(net568),
    .B(_0421_),
    .Y(_1031_));
 sg13g2_nor3_1 _1926_ (.A(net496),
    .B(_0965_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_a21o_1 _1927_ (.A2(_1030_),
    .A1(net496),
    .B1(_1032_),
    .X(_1033_));
 sg13g2_nand2_1 _1928_ (.Y(_1034_),
    .A(net543),
    .B(net492));
 sg13g2_o21ai_1 _1929_ (.B1(_1034_),
    .Y(_1035_),
    .A1(net574),
    .A2(_0846_));
 sg13g2_a22oi_1 _1930_ (.Y(_1036_),
    .B1(_0864_),
    .B2(_1035_),
    .A2(_0862_),
    .A1(net523));
 sg13g2_a221oi_1 _1931_ (.B2(net494),
    .C1(net492),
    .B1(_0862_),
    .A1(net543),
    .Y(_1037_),
    .A2(_0859_));
 sg13g2_nand2_2 _1932_ (.Y(_1038_),
    .A(net543),
    .B(net584));
 sg13g2_o21ai_1 _1933_ (.B1(_1036_),
    .Y(_1039_),
    .A1(net560),
    .A2(_1037_));
 sg13g2_a22oi_1 _1934_ (.Y(_1040_),
    .B1(_1039_),
    .B2(net478),
    .A2(net465),
    .A1(_0421_));
 sg13g2_a21oi_1 _1935_ (.A1(net568),
    .A2(_0011_),
    .Y(_1041_),
    .B1(_0960_));
 sg13g2_a21o_1 _1936_ (.A2(_0011_),
    .A1(net560),
    .B1(_0965_),
    .X(_1042_));
 sg13g2_a22oi_1 _1937_ (.Y(_1043_),
    .B1(_0877_),
    .B2(_1041_),
    .A2(net492),
    .A1(net543));
 sg13g2_o21ai_1 _1938_ (.B1(_1043_),
    .Y(_1044_),
    .A1(net494),
    .A2(_1042_));
 sg13g2_a22oi_1 _1939_ (.Y(_1045_),
    .B1(_1044_),
    .B2(net460),
    .A2(_1033_),
    .A1(net459));
 sg13g2_a21oi_1 _1940_ (.A1(_1040_),
    .A2(_1045_),
    .Y(_1046_),
    .B1(_0845_));
 sg13g2_nand3_1 _1941_ (.B(_0890_),
    .C(_0893_),
    .A(_0421_),
    .Y(_1047_));
 sg13g2_a22oi_1 _1942_ (.Y(_1048_),
    .B1(_0899_),
    .B2(net503),
    .A2(_0898_),
    .A1(_0437_));
 sg13g2_a22oi_1 _1943_ (.Y(_1049_),
    .B1(_0897_),
    .B2(net517),
    .A2(_0895_),
    .A1(net532));
 sg13g2_nand4_1 _1944_ (.B(_1047_),
    .C(_1048_),
    .A(net490),
    .Y(_1050_),
    .D(_1049_));
 sg13g2_a22oi_1 _1945_ (.Y(_1051_),
    .B1(_0752_),
    .B2(net503),
    .A2(_0720_),
    .A1(net517));
 sg13g2_nor2_1 _1946_ (.A(_0003_),
    .B(net468),
    .Y(_1052_));
 sg13g2_nor3_1 _1947_ (.A(_0715_),
    .B(_0753_),
    .C(_1052_),
    .Y(_1053_));
 sg13g2_a22oi_1 _1948_ (.Y(_1054_),
    .B1(_1051_),
    .B2(_1053_),
    .A2(_0713_),
    .A1(_0031_));
 sg13g2_o21ai_1 _1949_ (.B1(_0906_),
    .Y(_1055_),
    .A1(net490),
    .A2(_1054_));
 sg13g2_nor2b_1 _1950_ (.A(_1055_),
    .B_N(_1050_),
    .Y(_1056_));
 sg13g2_o21ai_1 _1951_ (.B1(_0842_),
    .Y(_1057_),
    .A1(_1046_),
    .A2(_1056_));
 sg13g2_a21oi_1 _1952_ (.A1(net568),
    .A2(_0020_),
    .Y(_1058_),
    .B1(_1031_));
 sg13g2_nor2b_1 _1953_ (.A(net489),
    .B_N(_1041_),
    .Y(_1059_));
 sg13g2_o21ai_1 _1954_ (.B1(_1038_),
    .Y(_1060_),
    .A1(_0404_),
    .A2(net579));
 sg13g2_a221oi_1 _1955_ (.B2(_0937_),
    .C1(_1059_),
    .B1(_1060_),
    .A1(_0939_),
    .Y(_1061_),
    .A2(_1058_));
 sg13g2_o21ai_1 _1956_ (.B1(_1061_),
    .Y(_1062_),
    .A1(net502),
    .A2(_1042_));
 sg13g2_a21oi_1 _1957_ (.A1(net481),
    .A2(_1062_),
    .Y(_1063_),
    .B1(_0932_));
 sg13g2_o21ai_1 _1958_ (.B1(net556),
    .Y(_1064_),
    .A1(net87),
    .A2(net453));
 sg13g2_a21oi_1 _1959_ (.A1(_1057_),
    .A2(_1063_),
    .Y(_0050_),
    .B1(_1064_));
 sg13g2_nand3_1 _1960_ (.B(_0890_),
    .C(_0893_),
    .A(_0422_),
    .Y(_1065_));
 sg13g2_nor3_1 _1961_ (.A(\u8.rc[31] ),
    .B(_0885_),
    .C(_0888_),
    .Y(_1066_));
 sg13g2_a22oi_1 _1962_ (.Y(_1067_),
    .B1(_1066_),
    .B2(net552),
    .A2(_0899_),
    .A1(\u8.rc[22] ));
 sg13g2_a22oi_1 _1963_ (.Y(_1068_),
    .B1(_0897_),
    .B2(net513),
    .A2(_0895_),
    .A1(net530));
 sg13g2_nand4_1 _1964_ (.B(_1065_),
    .C(_1067_),
    .A(net490),
    .Y(_1069_),
    .D(_1068_));
 sg13g2_a21oi_1 _1965_ (.A1(_0422_),
    .A2(_0664_),
    .Y(_1070_),
    .B1(net490));
 sg13g2_nor2_1 _1966_ (.A(_0004_),
    .B(net468),
    .Y(_1071_));
 sg13g2_a21oi_1 _1967_ (.A1(net513),
    .A2(_0720_),
    .Y(_1072_),
    .B1(_1071_));
 sg13g2_nand3_1 _1968_ (.B(_1070_),
    .C(_1072_),
    .A(_0676_),
    .Y(_1073_));
 sg13g2_and3_1 _1969_ (.X(_1074_),
    .A(_0906_),
    .B(_1069_),
    .C(_1073_));
 sg13g2_nor2_1 _1970_ (.A(net578),
    .B(_0006_),
    .Y(_1075_));
 sg13g2_a21oi_2 _1971_ (.B1(_1075_),
    .Y(_1076_),
    .A2(_0432_),
    .A1(net579));
 sg13g2_nand2_1 _1972_ (.Y(_1077_),
    .A(net578),
    .B(_0006_));
 sg13g2_o21ai_1 _1973_ (.B1(_1077_),
    .Y(_1078_),
    .A1(net579),
    .A2(_0432_));
 sg13g2_nor2_1 _1974_ (.A(net495),
    .B(_1078_),
    .Y(_1079_));
 sg13g2_a21oi_1 _1975_ (.A1(net542),
    .A2(net493),
    .Y(_1080_),
    .B1(_1079_));
 sg13g2_o21ai_1 _1976_ (.B1(_1080_),
    .Y(_1081_),
    .A1(_0876_),
    .A2(_1076_));
 sg13g2_nand2_2 _1977_ (.Y(_1082_),
    .A(\u8.ls[4] ),
    .B(net584));
 sg13g2_mux4_1 _1978_ (.S0(net580),
    .A0(_0397_),
    .A1(_0401_),
    .A2(_0032_),
    .A3(_0006_),
    .S1(net495),
    .X(_1083_));
 sg13g2_nor3_1 _1979_ (.A(net519),
    .B(net573),
    .C(_0864_),
    .Y(_1084_));
 sg13g2_nand2_1 _1980_ (.Y(_1085_),
    .A(_0401_),
    .B(net575));
 sg13g2_nand2_1 _1981_ (.Y(_1086_),
    .A(_0401_),
    .B(net560));
 sg13g2_a22oi_1 _1982_ (.Y(_1087_),
    .B1(_1086_),
    .B2(net493),
    .A2(_1085_),
    .A1(_0859_));
 sg13g2_o21ai_1 _1983_ (.B1(_0862_),
    .Y(_1088_),
    .A1(net519),
    .A2(_1003_));
 sg13g2_o21ai_1 _1984_ (.B1(_1088_),
    .Y(_1089_),
    .A1(_1084_),
    .A2(_1087_));
 sg13g2_a22oi_1 _1985_ (.Y(_1090_),
    .B1(_1089_),
    .B2(net478),
    .A2(_1081_),
    .A1(net461));
 sg13g2_o21ai_1 _1986_ (.B1(_1090_),
    .Y(_1091_),
    .A1(net456),
    .A2(_1083_));
 sg13g2_a21oi_1 _1987_ (.A1(_0422_),
    .A2(net465),
    .Y(_1092_),
    .B1(_1091_));
 sg13g2_nor2_1 _1988_ (.A(_0845_),
    .B(_1092_),
    .Y(_1093_));
 sg13g2_o21ai_1 _1989_ (.B1(_0842_),
    .Y(_1094_),
    .A1(_1074_),
    .A2(_1093_));
 sg13g2_nand2_1 _1990_ (.Y(_1095_),
    .A(net552),
    .B(net561));
 sg13g2_a21o_1 _1991_ (.A2(_1095_),
    .A1(_1082_),
    .B1(_0938_),
    .X(_1096_));
 sg13g2_o21ai_1 _1992_ (.B1(_1096_),
    .Y(_1097_),
    .A1(net489),
    .A2(_1076_));
 sg13g2_nand2b_1 _1993_ (.Y(_1098_),
    .B(net571),
    .A_N(net552));
 sg13g2_nand3_1 _1994_ (.B(_1086_),
    .C(_1098_),
    .A(_0939_),
    .Y(_1099_));
 sg13g2_o21ai_1 _1995_ (.B1(_1099_),
    .Y(_1100_),
    .A1(net502),
    .A2(_1078_));
 sg13g2_o21ai_1 _1996_ (.B1(net481),
    .Y(_1101_),
    .A1(_1097_),
    .A2(_1100_));
 sg13g2_and2_1 _1997_ (.A(net453),
    .B(_1101_),
    .X(_1102_));
 sg13g2_o21ai_1 _1998_ (.B1(net557),
    .Y(_1103_),
    .A1(net79),
    .A2(net453));
 sg13g2_a21oi_1 _1999_ (.A1(_1094_),
    .A2(_1102_),
    .Y(_0051_),
    .B1(_1103_));
 sg13g2_nand3_1 _2000_ (.B(_0890_),
    .C(_0893_),
    .A(_0423_),
    .Y(_1104_));
 sg13g2_a22oi_1 _2001_ (.Y(_1105_),
    .B1(_1066_),
    .B2(net551),
    .A2(_0899_),
    .A1(\u8.rc[23] ));
 sg13g2_a22oi_1 _2002_ (.Y(_1106_),
    .B1(_0897_),
    .B2(net512),
    .A2(_0895_),
    .A1(net528));
 sg13g2_nand4_1 _2003_ (.B(_1104_),
    .C(_1105_),
    .A(net491),
    .Y(_1107_),
    .D(_1106_));
 sg13g2_a22oi_1 _2004_ (.Y(_1108_),
    .B1(_0725_),
    .B2(_0005_),
    .A2(_0713_),
    .A1(_0033_));
 sg13g2_o21ai_1 _2005_ (.B1(_0906_),
    .Y(_1109_),
    .A1(net490),
    .A2(_1108_));
 sg13g2_nor2b_1 _2006_ (.A(_1109_),
    .B_N(_1107_),
    .Y(_1110_));
 sg13g2_nor2b_1 _2007_ (.A(net582),
    .B_N(net540),
    .Y(_1111_));
 sg13g2_nor2_1 _2008_ (.A(_0396_),
    .B(net562),
    .Y(_1112_));
 sg13g2_or3_1 _2009_ (.A(net497),
    .B(_1111_),
    .C(_1112_),
    .X(_1113_));
 sg13g2_nor2b_1 _2010_ (.A(net581),
    .B_N(_0029_),
    .Y(_1114_));
 sg13g2_a21oi_1 _2011_ (.A1(net580),
    .A2(_0033_),
    .Y(_1115_),
    .B1(_1114_));
 sg13g2_o21ai_1 _2012_ (.B1(_1113_),
    .Y(_1116_),
    .A1(net495),
    .A2(_1115_));
 sg13g2_a21o_1 _2013_ (.A2(net580),
    .A1(_0027_),
    .B1(_1114_),
    .X(_1117_));
 sg13g2_nand2_1 _2014_ (.Y(_1118_),
    .A(_0029_),
    .B(net581));
 sg13g2_o21ai_1 _2015_ (.B1(_1118_),
    .Y(_1119_),
    .A1(_0414_),
    .A2(net581));
 sg13g2_inv_1 _2016_ (.Y(_1120_),
    .A(_1119_));
 sg13g2_a22oi_1 _2017_ (.Y(_1121_),
    .B1(_1120_),
    .B2(net497),
    .A2(net493),
    .A1(net540));
 sg13g2_o21ai_1 _2018_ (.B1(_1121_),
    .Y(_1122_),
    .A1(_0876_),
    .A2(_1117_));
 sg13g2_nand2b_1 _2019_ (.Y(_1123_),
    .B(net517),
    .A_N(_1003_));
 sg13g2_and2_2 _2020_ (.A(net540),
    .B(net580),
    .X(_1124_));
 sg13g2_a22oi_1 _2021_ (.Y(_1125_),
    .B1(_1124_),
    .B2(_0859_),
    .A2(_1111_),
    .A1(net493));
 sg13g2_o21ai_1 _2022_ (.B1(_1123_),
    .Y(_1126_),
    .A1(_0863_),
    .A2(_1125_));
 sg13g2_a22oi_1 _2023_ (.Y(_1127_),
    .B1(_1126_),
    .B2(net478),
    .A2(_1122_),
    .A1(net461));
 sg13g2_o21ai_1 _2024_ (.B1(_1127_),
    .Y(_1128_),
    .A1(net456),
    .A2(_1116_));
 sg13g2_a21oi_1 _2025_ (.A1(_0423_),
    .A2(net465),
    .Y(_1129_),
    .B1(_1128_));
 sg13g2_nor2_1 _2026_ (.A(_0845_),
    .B(_1129_),
    .Y(_1130_));
 sg13g2_o21ai_1 _2027_ (.B1(_0842_),
    .Y(_1131_),
    .A1(_1110_),
    .A2(_1130_));
 sg13g2_nand2_1 _2028_ (.Y(_1132_),
    .A(net561),
    .B(_0423_));
 sg13g2_o21ai_1 _2029_ (.B1(_1132_),
    .Y(_1133_),
    .A1(_0025_),
    .A2(net561));
 sg13g2_or2_1 _2030_ (.X(_1134_),
    .B(_1117_),
    .A(net489));
 sg13g2_a21o_1 _2031_ (.A2(net561),
    .A1(net551),
    .B1(_1124_),
    .X(_1135_));
 sg13g2_o21ai_1 _2032_ (.B1(_1134_),
    .Y(_1136_),
    .A1(net502),
    .A2(_1119_));
 sg13g2_a22oi_1 _2033_ (.Y(_1137_),
    .B1(_1135_),
    .B2(_0937_),
    .A2(_1133_),
    .A1(_0939_));
 sg13g2_nand2b_1 _2034_ (.Y(_1138_),
    .B(_1137_),
    .A_N(_1136_));
 sg13g2_a21oi_1 _2035_ (.A1(net481),
    .A2(_1138_),
    .Y(_1139_),
    .B1(_0932_));
 sg13g2_o21ai_1 _2036_ (.B1(net556),
    .Y(_1140_),
    .A1(net86),
    .A2(_0931_));
 sg13g2_a21oi_1 _2037_ (.A1(_1131_),
    .A2(_1139_),
    .Y(_0052_),
    .B1(_1140_));
 sg13g2_and2_1 _2038_ (.A(_0034_),
    .B(net465),
    .X(_1141_));
 sg13g2_nor2b_1 _2039_ (.A(net580),
    .B_N(_0007_),
    .Y(_1142_));
 sg13g2_a21oi_1 _2040_ (.A1(net575),
    .A2(_0034_),
    .Y(_1143_),
    .B1(_1142_));
 sg13g2_nand2_2 _2041_ (.Y(_1144_),
    .A(net580),
    .B(_0007_));
 sg13g2_nor2b_2 _2042_ (.A(net582),
    .B_N(_0034_),
    .Y(_1145_));
 sg13g2_nor2_1 _2043_ (.A(net497),
    .B(_1145_),
    .Y(_1146_));
 sg13g2_a22oi_1 _2044_ (.Y(_1147_),
    .B1(_1144_),
    .B2(_1146_),
    .A2(_1143_),
    .A1(net497));
 sg13g2_a21o_1 _2045_ (.A2(_0014_),
    .A1(net571),
    .B1(_1142_),
    .X(_1148_));
 sg13g2_nand2_1 _2046_ (.Y(_1149_),
    .A(net560),
    .B(_0014_));
 sg13g2_and2_1 _2047_ (.A(_1144_),
    .B(_1149_),
    .X(_1150_));
 sg13g2_a22oi_1 _2048_ (.Y(_1151_),
    .B1(_1150_),
    .B2(net496),
    .A2(net492),
    .A1(net539));
 sg13g2_o21ai_1 _2049_ (.B1(_1151_),
    .Y(_1152_),
    .A1(_0876_),
    .A2(_1148_));
 sg13g2_nand2_1 _2050_ (.Y(_1153_),
    .A(_0400_),
    .B(net573));
 sg13g2_o21ai_1 _2051_ (.B1(net492),
    .Y(_1154_),
    .A1(net539),
    .A2(net573));
 sg13g2_a22oi_1 _2052_ (.Y(_1155_),
    .B1(_0859_),
    .B2(_1153_),
    .A2(net496),
    .A1(_0745_));
 sg13g2_nand3_1 _2053_ (.B(_1154_),
    .C(_1155_),
    .A(_0864_),
    .Y(_1156_));
 sg13g2_a21oi_1 _2054_ (.A1(net513),
    .A2(_1002_),
    .Y(_1157_),
    .B1(_0640_));
 sg13g2_o21ai_1 _2055_ (.B1(_0737_),
    .Y(_1158_),
    .A1(net456),
    .A2(_1147_));
 sg13g2_a221oi_1 _2056_ (.B2(_1157_),
    .C1(_1158_),
    .B1(_1156_),
    .A1(net460),
    .Y(_1159_),
    .A2(_1152_));
 sg13g2_nor4_1 _2057_ (.A(_0841_),
    .B(_0845_),
    .C(_1141_),
    .D(_1159_),
    .Y(_1160_));
 sg13g2_a21oi_1 _2058_ (.A1(_0400_),
    .A2(_0713_),
    .Y(_1161_),
    .B1(net490));
 sg13g2_nand2_1 _2059_ (.Y(_1162_),
    .A(_0914_),
    .B(_1161_));
 sg13g2_mux2_1 _2060_ (.A0(net539),
    .A1(net550),
    .S(net568),
    .X(_1163_));
 sg13g2_nand2b_1 _2061_ (.Y(_1164_),
    .B(_1150_),
    .A_N(net502));
 sg13g2_mux2_1 _2062_ (.A0(net550),
    .A1(net539),
    .S(net568),
    .X(_1165_));
 sg13g2_o21ai_1 _2063_ (.B1(_1164_),
    .Y(_1166_),
    .A1(net489),
    .A2(_1148_));
 sg13g2_a221oi_1 _2064_ (.B2(_0937_),
    .C1(_1166_),
    .B1(_1165_),
    .A1(_0939_),
    .Y(_1167_),
    .A2(_1163_));
 sg13g2_nor2b_1 _2065_ (.A(_1167_),
    .B_N(net481),
    .Y(_1168_));
 sg13g2_nor3_1 _2066_ (.A(_0932_),
    .B(_1160_),
    .C(_1168_),
    .Y(_1169_));
 sg13g2_o21ai_1 _2067_ (.B1(net556),
    .Y(_1170_),
    .A1(net97),
    .A2(net453));
 sg13g2_a21oi_1 _2068_ (.A1(_1162_),
    .A2(_1169_),
    .Y(_0053_),
    .B1(_1170_));
 sg13g2_nor2_2 _2069_ (.A(_0409_),
    .B(net569),
    .Y(_1171_));
 sg13g2_a21oi_1 _2070_ (.A1(_0024_),
    .A2(net569),
    .Y(_1172_),
    .B1(_1171_));
 sg13g2_nor2_1 _2071_ (.A(_0399_),
    .B(net562),
    .Y(_1173_));
 sg13g2_a21oi_1 _2072_ (.A1(\u8.rc[31] ),
    .A2(net560),
    .Y(_1174_),
    .B1(_1173_));
 sg13g2_nand2_1 _2073_ (.Y(_1175_),
    .A(net570),
    .B(_0008_));
 sg13g2_o21ai_1 _2074_ (.B1(_1175_),
    .Y(_1176_),
    .A1(net571),
    .A2(_0434_));
 sg13g2_or2_1 _2075_ (.X(_1177_),
    .B(_1176_),
    .A(net502));
 sg13g2_nand2_1 _2076_ (.Y(_1178_),
    .A(net572),
    .B(_0015_));
 sg13g2_o21ai_1 _2077_ (.B1(_1178_),
    .Y(_1179_),
    .A1(net572),
    .A2(_0429_));
 sg13g2_o21ai_1 _2078_ (.B1(_1177_),
    .Y(_1180_),
    .A1(net489),
    .A2(_1179_));
 sg13g2_a21oi_1 _2079_ (.A1(_0939_),
    .A2(_1172_),
    .Y(_1181_),
    .B1(_1180_));
 sg13g2_o21ai_1 _2080_ (.B1(_1181_),
    .Y(_1182_),
    .A1(_0938_),
    .A2(_1174_));
 sg13g2_nand3_1 _2081_ (.B(_0713_),
    .C(_0901_),
    .A(_0021_),
    .Y(_1183_));
 sg13g2_mux4_1 _2082_ (.S0(net569),
    .A0(net517),
    .A1(net536),
    .A2(_0409_),
    .A3(_0429_),
    .S1(net494),
    .X(_1184_));
 sg13g2_nor2_1 _2083_ (.A(_0468_),
    .B(_0529_),
    .Y(_1185_));
 sg13g2_a21oi_1 _2084_ (.A1(net568),
    .A2(_1185_),
    .Y(_1186_),
    .B1(net494));
 sg13g2_nand2_1 _2085_ (.Y(_1187_),
    .A(_0399_),
    .B(net560));
 sg13g2_nand2_1 _2086_ (.Y(_1188_),
    .A(_0399_),
    .B(net573));
 sg13g2_a221oi_1 _2087_ (.B2(_0859_),
    .C1(_1186_),
    .B1(_1188_),
    .A1(net492),
    .Y(_0092_),
    .A2(_1187_));
 sg13g2_a22oi_1 _2088_ (.Y(_0093_),
    .B1(_0092_),
    .B2(_0864_),
    .A2(_1185_),
    .A1(_1002_));
 sg13g2_a21oi_1 _2089_ (.A1(net478),
    .A2(_0093_),
    .Y(_0094_),
    .B1(net465));
 sg13g2_nor2_1 _2090_ (.A(net494),
    .B(_1176_),
    .Y(_0095_));
 sg13g2_a21oi_1 _2091_ (.A1(net536),
    .A2(net492),
    .Y(_0096_),
    .B1(_0095_));
 sg13g2_o21ai_1 _2092_ (.B1(_0096_),
    .Y(_0097_),
    .A1(_0876_),
    .A2(_1179_));
 sg13g2_a22oi_1 _2093_ (.Y(_0098_),
    .B1(_0097_),
    .B2(net460),
    .A2(_1184_),
    .A1(net459));
 sg13g2_a221oi_1 _2094_ (.B2(_0098_),
    .C1(_0841_),
    .B1(_0094_),
    .A1(_0021_),
    .Y(_0099_),
    .A2(net465));
 sg13g2_nor2b_1 _2095_ (.A(_0845_),
    .B_N(_0099_),
    .Y(_0100_));
 sg13g2_a221oi_1 _2096_ (.B2(_0914_),
    .C1(_0100_),
    .B1(_1183_),
    .A1(net481),
    .Y(_0101_),
    .A2(_1182_));
 sg13g2_o21ai_1 _2097_ (.B1(net556),
    .Y(_0102_),
    .A1(net89),
    .A2(net453));
 sg13g2_a21oi_1 _2098_ (.A1(net453),
    .A2(_0101_),
    .Y(_0054_),
    .B1(_0102_));
 sg13g2_nor2_2 _2099_ (.A(_0683_),
    .B(_0824_),
    .Y(_0103_));
 sg13g2_o21ai_1 _2100_ (.B1(net559),
    .Y(_0104_),
    .A1(\u8.rcip[2] ),
    .A2(_0701_));
 sg13g2_nand3_1 _2101_ (.B(_0688_),
    .C(_0104_),
    .A(net1),
    .Y(_0105_));
 sg13g2_nor2_1 _2102_ (.A(_0696_),
    .B(_0105_),
    .Y(_0106_));
 sg13g2_nor2_2 _2103_ (.A(_0685_),
    .B(_0738_),
    .Y(_0107_));
 sg13g2_nand2_2 _2104_ (.Y(_0108_),
    .A(_0684_),
    .B(_0739_));
 sg13g2_o21ai_1 _2105_ (.B1(_0106_),
    .Y(_0109_),
    .A1(_0686_),
    .A2(_0738_));
 sg13g2_nand2_1 _2106_ (.Y(_0110_),
    .A(net78),
    .B(_0109_));
 sg13g2_nand2_1 _2107_ (.Y(_0055_),
    .A(net592),
    .B(_0110_));
 sg13g2_nand3_1 _2108_ (.B(_0742_),
    .C(_0823_),
    .A(net563),
    .Y(_0111_));
 sg13g2_nand2b_1 _2109_ (.Y(_0112_),
    .B(_0111_),
    .A_N(_0687_));
 sg13g2_nand2_1 _2110_ (.Y(_0113_),
    .A(\u8.rcip[1] ),
    .B(_0023_));
 sg13g2_nor2_1 _2111_ (.A(\u8.rcip[0] ),
    .B(_0113_),
    .Y(_0114_));
 sg13g2_or2_1 _2112_ (.X(_0115_),
    .B(_0113_),
    .A(\u8.rcip[0] ));
 sg13g2_nor3_1 _2113_ (.A(net584),
    .B(_0683_),
    .C(_0115_),
    .Y(_0116_));
 sg13g2_nor3_1 _2114_ (.A(_0708_),
    .B(_0112_),
    .C(_0116_),
    .Y(_0117_));
 sg13g2_nand2b_2 _2115_ (.Y(_0118_),
    .B(_0825_),
    .A_N(_0763_));
 sg13g2_a21oi_1 _2116_ (.A1(net576),
    .A2(_0425_),
    .Y(_0119_),
    .B1(_0850_));
 sg13g2_nor2_2 _2117_ (.A(_0742_),
    .B(_0114_),
    .Y(_0120_));
 sg13g2_nand2_1 _2118_ (.Y(_0121_),
    .A(_0743_),
    .B(_0115_));
 sg13g2_a21oi_2 _2119_ (.B1(_0104_),
    .Y(_0122_),
    .A2(net480),
    .A1(net562));
 sg13g2_nand2_1 _2120_ (.Y(_0123_),
    .A(net483),
    .B(_0119_));
 sg13g2_o21ai_1 _2121_ (.B1(_0123_),
    .Y(_0124_),
    .A1(_0001_),
    .A2(net483));
 sg13g2_a22oi_1 _2122_ (.Y(_0125_),
    .B1(_0124_),
    .B2(net460),
    .A2(_0119_),
    .A1(net470));
 sg13g2_nor2_1 _2123_ (.A(_0108_),
    .B(_0125_),
    .Y(_0126_));
 sg13g2_a221oi_1 _2124_ (.B2(_0122_),
    .C1(_0126_),
    .B1(_0119_),
    .A1(net7),
    .Y(_0127_),
    .A2(_0118_));
 sg13g2_o21ai_1 _2125_ (.B1(net588),
    .Y(_0128_),
    .A1(net120),
    .A2(net447));
 sg13g2_a21oi_1 _2126_ (.A1(net448),
    .A2(_0127_),
    .Y(_0056_),
    .B1(_0128_));
 sg13g2_a21oi_1 _2127_ (.A1(net582),
    .A2(_0427_),
    .Y(_0129_),
    .B1(_0956_));
 sg13g2_nand2_1 _2128_ (.Y(_0130_),
    .A(net482),
    .B(_0129_));
 sg13g2_o21ai_1 _2129_ (.B1(_0130_),
    .Y(_0131_),
    .A1(_0003_),
    .A2(net482));
 sg13g2_a22oi_1 _2130_ (.Y(_0132_),
    .B1(_0131_),
    .B2(net462),
    .A2(_0129_),
    .A1(net470));
 sg13g2_nor2_1 _2131_ (.A(_0108_),
    .B(_0132_),
    .Y(_0133_));
 sg13g2_a221oi_1 _2132_ (.B2(_0129_),
    .C1(_0133_),
    .B1(_0122_),
    .A1(net8),
    .Y(_0134_),
    .A2(_0118_));
 sg13g2_o21ai_1 _2133_ (.B1(net589),
    .Y(_0135_),
    .A1(net117),
    .A2(net447));
 sg13g2_a21oi_1 _2134_ (.A1(net449),
    .A2(_0134_),
    .Y(_0057_),
    .B1(_0135_));
 sg13g2_a21oi_1 _2135_ (.A1(_0418_),
    .A2(net576),
    .Y(_0136_),
    .B1(_0992_));
 sg13g2_nand2_1 _2136_ (.Y(_0137_),
    .A(net482),
    .B(_0136_));
 sg13g2_o21ai_1 _2137_ (.B1(_0137_),
    .Y(_0138_),
    .A1(_0004_),
    .A2(net482));
 sg13g2_a22oi_1 _2138_ (.Y(_0139_),
    .B1(_0138_),
    .B2(net460),
    .A2(_0136_),
    .A1(net472));
 sg13g2_nor2_1 _2139_ (.A(_0108_),
    .B(_0139_),
    .Y(_0140_));
 sg13g2_a221oi_1 _2140_ (.B2(_0136_),
    .C1(_0140_),
    .B1(_0122_),
    .A1(net9),
    .Y(_0141_),
    .A2(_0118_));
 sg13g2_o21ai_1 _2141_ (.B1(net588),
    .Y(_0142_),
    .A1(net544),
    .A2(net447));
 sg13g2_a21oi_1 _2142_ (.A1(net447),
    .A2(_0141_),
    .Y(_0058_),
    .B1(_0142_));
 sg13g2_a21oi_1 _2143_ (.A1(net576),
    .A2(_0420_),
    .Y(_0143_),
    .B1(_1031_));
 sg13g2_nand2_1 _2144_ (.Y(_0144_),
    .A(net482),
    .B(_0143_));
 sg13g2_o21ai_1 _2145_ (.B1(_0144_),
    .Y(_0145_),
    .A1(_0005_),
    .A2(net482));
 sg13g2_a22oi_1 _2146_ (.Y(_0146_),
    .B1(_0145_),
    .B2(net460),
    .A2(_0143_),
    .A1(net472));
 sg13g2_nor2_1 _2147_ (.A(_0108_),
    .B(_0146_),
    .Y(_0147_));
 sg13g2_a221oi_1 _2148_ (.B2(_0143_),
    .C1(_0147_),
    .B1(_0122_),
    .A1(net10),
    .Y(_0148_),
    .A2(_0118_));
 sg13g2_o21ai_1 _2149_ (.B1(net588),
    .Y(_0149_),
    .A1(net543),
    .A2(net447));
 sg13g2_a21oi_1 _2150_ (.A1(net447),
    .A2(_0148_),
    .Y(_0059_),
    .B1(_0149_));
 sg13g2_nor2_1 _2151_ (.A(net562),
    .B(net11),
    .Y(_0150_));
 sg13g2_a21oi_1 _2152_ (.A1(net562),
    .A2(_0032_),
    .Y(_0151_),
    .B1(_0150_));
 sg13g2_nand2_1 _2153_ (.Y(_0152_),
    .A(net483),
    .B(_0151_));
 sg13g2_o21ai_1 _2154_ (.B1(_0152_),
    .Y(_0153_),
    .A1(_0006_),
    .A2(net483));
 sg13g2_a22oi_1 _2155_ (.Y(_0154_),
    .B1(_0153_),
    .B2(net462),
    .A2(_0151_),
    .A1(net470));
 sg13g2_nor2_1 _2156_ (.A(_0108_),
    .B(_0154_),
    .Y(_0155_));
 sg13g2_a221oi_1 _2157_ (.B2(_0151_),
    .C1(_0155_),
    .B1(_0122_),
    .A1(net11),
    .Y(_0156_),
    .A2(_0118_));
 sg13g2_o21ai_1 _2158_ (.B1(net588),
    .Y(_0157_),
    .A1(net542),
    .A2(net449));
 sg13g2_a21oi_1 _2159_ (.A1(net449),
    .A2(_0156_),
    .Y(_0060_),
    .B1(_0157_));
 sg13g2_a21o_1 _2160_ (.A2(net12),
    .A1(net583),
    .B1(_1111_),
    .X(_0158_));
 sg13g2_nand2_1 _2161_ (.Y(_0159_),
    .A(net483),
    .B(_0158_));
 sg13g2_o21ai_1 _2162_ (.B1(_0159_),
    .Y(_0160_),
    .A1(_0029_),
    .A2(net483));
 sg13g2_a22oi_1 _2163_ (.Y(_0161_),
    .B1(_0160_),
    .B2(net462),
    .A2(_0158_),
    .A1(net470));
 sg13g2_nor2_1 _2164_ (.A(_0108_),
    .B(_0161_),
    .Y(_0162_));
 sg13g2_a221oi_1 _2165_ (.B2(_0158_),
    .C1(_0162_),
    .B1(_0122_),
    .A1(net12),
    .Y(_0163_),
    .A2(_0118_));
 sg13g2_o21ai_1 _2166_ (.B1(net588),
    .Y(_0164_),
    .A1(net540),
    .A2(net449));
 sg13g2_a21oi_1 _2167_ (.A1(net449),
    .A2(_0163_),
    .Y(_0061_),
    .B1(_0164_));
 sg13g2_nand2_1 _2168_ (.Y(_0165_),
    .A(_0741_),
    .B(_0825_));
 sg13g2_o21ai_1 _2169_ (.B1(net13),
    .Y(_0166_),
    .A1(_0822_),
    .A2(_0165_));
 sg13g2_a21oi_2 _2170_ (.B1(_1145_),
    .Y(_0167_),
    .A2(net585),
    .A1(_0416_));
 sg13g2_a22oi_1 _2171_ (.Y(_0168_),
    .B1(_0122_),
    .B2(_0167_),
    .A2(_0696_),
    .A1(\u8.ls[0] ));
 sg13g2_nand2_1 _2172_ (.Y(_0169_),
    .A(net486),
    .B(_0167_));
 sg13g2_o21ai_1 _2173_ (.B1(_0169_),
    .Y(_0170_),
    .A1(_0007_),
    .A2(net486));
 sg13g2_a22oi_1 _2174_ (.Y(_0171_),
    .B1(_0170_),
    .B2(net463),
    .A2(_0167_),
    .A1(net471));
 sg13g2_nand2b_1 _2175_ (.Y(_0172_),
    .B(_0107_),
    .A_N(_0171_));
 sg13g2_nand4_1 _2176_ (.B(_0166_),
    .C(_0168_),
    .A(net449),
    .Y(_0173_),
    .D(_0172_));
 sg13g2_o21ai_1 _2177_ (.B1(net592),
    .Y(_0174_),
    .A1(net538),
    .A2(net449));
 sg13g2_nor2b_1 _2178_ (.A(_0174_),
    .B_N(_0173_),
    .Y(_0062_));
 sg13g2_a21oi_2 _2179_ (.B1(_1171_),
    .Y(_0175_),
    .A2(net580),
    .A1(_0417_));
 sg13g2_o21ai_1 _2180_ (.B1(net477),
    .Y(_0176_),
    .A1(\u8.ls[1] ),
    .A2(_0660_));
 sg13g2_nand2_1 _2181_ (.Y(_0177_),
    .A(net482),
    .B(_0175_));
 sg13g2_o21ai_1 _2182_ (.B1(_0177_),
    .Y(_0178_),
    .A1(_0008_),
    .A2(net482));
 sg13g2_a22oi_1 _2183_ (.Y(_0179_),
    .B1(_0178_),
    .B2(net462),
    .A2(_0175_),
    .A1(net471));
 sg13g2_o21ai_1 _2184_ (.B1(_0176_),
    .Y(_0180_),
    .A1(_0108_),
    .A2(_0179_));
 sg13g2_a221oi_1 _2185_ (.B2(_0122_),
    .C1(_0180_),
    .B1(_0175_),
    .A1(net14),
    .Y(_0181_),
    .A2(_0165_));
 sg13g2_o21ai_1 _2186_ (.B1(net588),
    .Y(_0182_),
    .A1(net536),
    .A2(net447));
 sg13g2_a21oi_1 _2187_ (.A1(net447),
    .A2(_0181_),
    .Y(_0063_),
    .B1(_0182_));
 sg13g2_nor2_1 _2188_ (.A(net584),
    .B(net7),
    .Y(_0183_));
 sg13g2_a21oi_2 _2189_ (.B1(_0183_),
    .Y(_0184_),
    .A2(_0000_),
    .A1(net584));
 sg13g2_a21oi_1 _2190_ (.A1(\u8.ls[0] ),
    .A2(net584),
    .Y(_0185_),
    .B1(_0120_));
 sg13g2_o21ai_1 _2191_ (.B1(_0103_),
    .Y(_0186_),
    .A1(net480),
    .A2(_0184_));
 sg13g2_nor2_1 _2192_ (.A(_0185_),
    .B(_0186_),
    .Y(_0187_));
 sg13g2_o21ai_1 _2193_ (.B1(net463),
    .Y(_0188_),
    .A1(_0009_),
    .A2(net485));
 sg13g2_a21oi_1 _2194_ (.A1(net485),
    .A2(_0184_),
    .Y(_0189_),
    .B1(_0188_));
 sg13g2_nand2_1 _2195_ (.Y(_0190_),
    .A(_0402_),
    .B(net458));
 sg13g2_o21ai_1 _2196_ (.B1(_0190_),
    .Y(_0191_),
    .A1(_0642_),
    .A2(_0184_));
 sg13g2_o21ai_1 _2197_ (.B1(_0762_),
    .Y(_0192_),
    .A1(_0189_),
    .A2(_0191_));
 sg13g2_nand2_1 _2198_ (.Y(_0193_),
    .A(net544),
    .B(net501));
 sg13g2_a21oi_1 _2199_ (.A1(_0765_),
    .A2(_0193_),
    .Y(_0194_),
    .B1(_0682_));
 sg13g2_a21oi_1 _2200_ (.A1(_0192_),
    .A2(_0194_),
    .Y(_0195_),
    .B1(_0187_));
 sg13g2_o21ai_1 _2201_ (.B1(net591),
    .Y(_0196_),
    .A1(net533),
    .A2(net450));
 sg13g2_a21oi_1 _2202_ (.A1(net450),
    .A2(_0195_),
    .Y(_0064_),
    .B1(_0196_));
 sg13g2_a21oi_2 _2203_ (.B1(_0750_),
    .Y(_0197_),
    .A2(_0002_),
    .A1(net585));
 sg13g2_o21ai_1 _2204_ (.B1(_0107_),
    .Y(_0198_),
    .A1(_0642_),
    .A2(_0197_));
 sg13g2_o21ai_1 _2205_ (.B1(net463),
    .Y(_0199_),
    .A1(_0028_),
    .A2(net486));
 sg13g2_a21oi_1 _2206_ (.A1(net486),
    .A2(_0197_),
    .Y(_0200_),
    .B1(_0199_));
 sg13g2_nor2_1 _2207_ (.A(\u8.ls[1] ),
    .B(net456),
    .Y(_0201_));
 sg13g2_or3_1 _2208_ (.A(_0198_),
    .B(_0200_),
    .C(_0201_),
    .X(_0202_));
 sg13g2_a21oi_1 _2209_ (.A1(_0985_),
    .A2(net479),
    .Y(_0203_),
    .B1(_0104_));
 sg13g2_o21ai_1 _2210_ (.B1(_0203_),
    .Y(_0204_),
    .A1(net479),
    .A2(_0197_));
 sg13g2_o21ai_1 _2211_ (.B1(_0712_),
    .Y(_0205_),
    .A1(net543),
    .A2(_0660_));
 sg13g2_nand4_1 _2212_ (.B(_0202_),
    .C(_0204_),
    .A(net452),
    .Y(_0206_),
    .D(_0205_));
 sg13g2_o21ai_1 _2213_ (.B1(net592),
    .Y(_0207_),
    .A1(net531),
    .A2(net451));
 sg13g2_nor2b_1 _2214_ (.A(_0207_),
    .B_N(_0206_),
    .Y(_0065_));
 sg13g2_nand2_1 _2215_ (.Y(_0208_),
    .A(_1022_),
    .B(net479));
 sg13g2_o21ai_1 _2216_ (.B1(_0208_),
    .Y(_0209_),
    .A1(_0833_),
    .A2(net479));
 sg13g2_nand2_1 _2217_ (.Y(_0210_),
    .A(_0001_),
    .B(net484));
 sg13g2_o21ai_1 _2218_ (.B1(_0210_),
    .Y(_0211_),
    .A1(_0431_),
    .A2(net484));
 sg13g2_a22oi_1 _2219_ (.Y(_0212_),
    .B1(net462),
    .B2(_0211_),
    .A2(_0833_),
    .A1(net470));
 sg13g2_o21ai_1 _2220_ (.B1(_0212_),
    .Y(_0213_),
    .A1(net544),
    .A2(net456));
 sg13g2_nand2_1 _2221_ (.Y(_0214_),
    .A(net542),
    .B(net501));
 sg13g2_a22oi_1 _2222_ (.Y(_0215_),
    .B1(_0214_),
    .B2(net476),
    .A2(_0213_),
    .A1(_0762_));
 sg13g2_a22oi_1 _2223_ (.Y(_0216_),
    .B1(_0215_),
    .B2(_0683_),
    .A2(_0209_),
    .A1(_0103_));
 sg13g2_o21ai_1 _2224_ (.B1(net591),
    .Y(_0217_),
    .A1(net529),
    .A2(net450));
 sg13g2_a21oi_1 _2225_ (.A1(net450),
    .A2(_0216_),
    .Y(_0066_),
    .B1(_0217_));
 sg13g2_nand2_1 _2226_ (.Y(_0218_),
    .A(net543),
    .B(net457));
 sg13g2_nand2b_1 _2227_ (.Y(_0219_),
    .B(net485),
    .A_N(_0003_));
 sg13g2_o21ai_1 _2228_ (.B1(_0219_),
    .Y(_0220_),
    .A1(_0011_),
    .A2(net485));
 sg13g2_a22oi_1 _2229_ (.Y(_0221_),
    .B1(net463),
    .B2(_0220_),
    .A2(_0830_),
    .A1(net471));
 sg13g2_nand3_1 _2230_ (.B(_0218_),
    .C(_0221_),
    .A(_0739_),
    .Y(_0222_));
 sg13g2_o21ai_1 _2231_ (.B1(_0103_),
    .Y(_0223_),
    .A1(_0830_),
    .A2(net480));
 sg13g2_a21oi_1 _2232_ (.A1(_1038_),
    .A2(net480),
    .Y(_0224_),
    .B1(_0223_));
 sg13g2_a21oi_1 _2233_ (.A1(net540),
    .A2(net469),
    .Y(_0225_),
    .B1(net498));
 sg13g2_o21ai_1 _2234_ (.B1(_0225_),
    .Y(_0226_),
    .A1(_0033_),
    .A2(net469));
 sg13g2_a221oi_1 _2235_ (.B2(net477),
    .C1(_0224_),
    .B1(_0226_),
    .A1(_0684_),
    .Y(_0227_),
    .A2(_0222_));
 sg13g2_o21ai_1 _2236_ (.B1(net591),
    .Y(_0228_),
    .A1(net527),
    .A2(net450));
 sg13g2_a21oi_1 _2237_ (.A1(net450),
    .A2(_0227_),
    .Y(_0067_),
    .B1(_0228_));
 sg13g2_nand2b_1 _2238_ (.Y(_0229_),
    .B(net485),
    .A_N(_0004_));
 sg13g2_o21ai_1 _2239_ (.B1(_0229_),
    .Y(_0230_),
    .A1(_0013_),
    .A2(net485));
 sg13g2_o21ai_1 _2240_ (.B1(_0739_),
    .Y(_0231_),
    .A1(_0642_),
    .A2(_0828_));
 sg13g2_a221oi_1 _2241_ (.B2(_0230_),
    .C1(_0231_),
    .B1(net463),
    .A1(net542),
    .Y(_0232_),
    .A2(net457));
 sg13g2_nor2_1 _2242_ (.A(_0685_),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nand2_1 _2243_ (.Y(_0234_),
    .A(_0828_),
    .B(_0120_));
 sg13g2_a21oi_1 _2244_ (.A1(_1082_),
    .A2(net479),
    .Y(_0235_),
    .B1(_0104_));
 sg13g2_a21oi_1 _2245_ (.A1(net538),
    .A2(net475),
    .Y(_0236_),
    .B1(net467));
 sg13g2_a21oi_1 _2246_ (.A1(net538),
    .A2(net469),
    .Y(_0237_),
    .B1(_0907_));
 sg13g2_o21ai_1 _2247_ (.B1(net501),
    .Y(_0238_),
    .A1(_0236_),
    .A2(_0237_));
 sg13g2_a221oi_1 _2248_ (.B2(net477),
    .C1(_0233_),
    .B1(_0238_),
    .A1(_0234_),
    .Y(_0239_),
    .A2(_0235_));
 sg13g2_o21ai_1 _2249_ (.B1(net591),
    .Y(_0240_),
    .A1(net524),
    .A2(net451));
 sg13g2_a21oi_1 _2250_ (.A1(net451),
    .A2(_0239_),
    .Y(_0068_),
    .B1(_0240_));
 sg13g2_nand2_1 _2251_ (.Y(_0241_),
    .A(net540),
    .B(net458));
 sg13g2_nor2_1 _2252_ (.A(_0414_),
    .B(net483),
    .Y(_0242_));
 sg13g2_a21oi_1 _2253_ (.A1(_0005_),
    .A2(net486),
    .Y(_0243_),
    .B1(_0242_));
 sg13g2_a22oi_1 _2254_ (.Y(_0244_),
    .B1(net462),
    .B2(_0243_),
    .A2(_0829_),
    .A1(net470));
 sg13g2_a21o_1 _2255_ (.A2(_0244_),
    .A1(_0241_),
    .B1(_0108_),
    .X(_0245_));
 sg13g2_mux2_1 _2256_ (.A0(_0829_),
    .A1(_1124_),
    .S(net479),
    .X(_0246_));
 sg13g2_a21oi_1 _2257_ (.A1(net536),
    .A2(net468),
    .Y(_0247_),
    .B1(_0977_));
 sg13g2_nand3_1 _2258_ (.B(net499),
    .C(net474),
    .A(net536),
    .Y(_0248_));
 sg13g2_a21oi_1 _2259_ (.A1(_0715_),
    .A2(_0248_),
    .Y(_0249_),
    .B1(_0247_));
 sg13g2_nor2_1 _2260_ (.A(_0764_),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_o21ai_1 _2261_ (.B1(_0245_),
    .Y(_0251_),
    .A1(_0695_),
    .A2(_0250_));
 sg13g2_a21oi_1 _2262_ (.A1(_0103_),
    .A2(_0246_),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_o21ai_1 _2263_ (.B1(net592),
    .Y(_0253_),
    .A1(net521),
    .A2(net451));
 sg13g2_a21oi_1 _2264_ (.A1(net451),
    .A2(_0252_),
    .Y(_0069_),
    .B1(_0253_));
 sg13g2_nor2_1 _2265_ (.A(_0433_),
    .B(net484),
    .Y(_0254_));
 sg13g2_a21oi_1 _2266_ (.A1(_0006_),
    .A2(net484),
    .Y(_0255_),
    .B1(_0254_));
 sg13g2_a221oi_1 _2267_ (.B2(_0255_),
    .C1(_0738_),
    .B1(net462),
    .A1(net470),
    .Y(_0256_),
    .A2(_0827_));
 sg13g2_o21ai_1 _2268_ (.B1(_0256_),
    .Y(_0257_),
    .A1(_0400_),
    .A2(net456));
 sg13g2_a21oi_1 _2269_ (.A1(net538),
    .A2(net581),
    .Y(_0258_),
    .B1(_0120_));
 sg13g2_o21ai_1 _2270_ (.B1(_0103_),
    .Y(_0259_),
    .A1(_0827_),
    .A2(net479));
 sg13g2_nor2_1 _2271_ (.A(_0258_),
    .B(_0259_),
    .Y(_0260_));
 sg13g2_a21oi_1 _2272_ (.A1(net535),
    .A2(net474),
    .Y(_0261_),
    .B1(net466));
 sg13g2_a21oi_1 _2273_ (.A1(net535),
    .A2(net469),
    .Y(_0262_),
    .B1(_1014_));
 sg13g2_o21ai_1 _2274_ (.B1(net499),
    .Y(_0263_),
    .A1(_0261_),
    .A2(_0262_));
 sg13g2_a221oi_1 _2275_ (.B2(net477),
    .C1(_0260_),
    .B1(_0263_),
    .A1(_0684_),
    .Y(_0264_),
    .A2(_0257_));
 sg13g2_o21ai_1 _2276_ (.B1(net590),
    .Y(_0265_),
    .A1(net520),
    .A2(net450));
 sg13g2_a21oi_1 _2277_ (.A1(net450),
    .A2(_0264_),
    .Y(_0070_),
    .B1(_0265_));
 sg13g2_nor2_1 _2278_ (.A(_0434_),
    .B(net484),
    .Y(_0266_));
 sg13g2_a21oi_1 _2279_ (.A1(_0029_),
    .A2(net484),
    .Y(_0267_),
    .B1(_0266_));
 sg13g2_a221oi_1 _2280_ (.B2(_0267_),
    .C1(_0738_),
    .B1(net462),
    .A1(net470),
    .Y(_0268_),
    .A2(_0832_));
 sg13g2_o21ai_1 _2281_ (.B1(_0268_),
    .Y(_0269_),
    .A1(_0399_),
    .A2(net456));
 sg13g2_a21oi_1 _2282_ (.A1(net532),
    .A2(net474),
    .Y(_0270_),
    .B1(net466));
 sg13g2_a21oi_1 _2283_ (.A1(net532),
    .A2(net468),
    .Y(_0271_),
    .B1(_1052_));
 sg13g2_o21ai_1 _2284_ (.B1(net500),
    .Y(_0272_),
    .A1(_0270_),
    .A2(_0271_));
 sg13g2_nor2_1 _2285_ (.A(_1173_),
    .B(_0120_),
    .Y(_0273_));
 sg13g2_o21ai_1 _2286_ (.B1(_0103_),
    .Y(_0274_),
    .A1(_0832_),
    .A2(net479));
 sg13g2_nor2_1 _2287_ (.A(_0273_),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_a221oi_1 _2288_ (.B2(net477),
    .C1(_0275_),
    .B1(_0272_),
    .A1(_0684_),
    .Y(_0276_),
    .A2(_0269_));
 sg13g2_o21ai_1 _2289_ (.B1(net587),
    .Y(_0277_),
    .A1(net517),
    .A2(net448));
 sg13g2_a21oi_1 _2290_ (.A1(net448),
    .A2(_0276_),
    .Y(_0071_),
    .B1(_0277_));
 sg13g2_o21ai_1 _2291_ (.B1(net559),
    .Y(_0278_),
    .A1(_0023_),
    .A2(_0824_));
 sg13g2_nor2b_1 _2292_ (.A(_0278_),
    .B_N(net1),
    .Y(_0279_));
 sg13g2_and2_1 _2293_ (.A(net101),
    .B(_0279_),
    .X(_0280_));
 sg13g2_o21ai_1 _2294_ (.B1(net591),
    .Y(_0281_),
    .A1(net101),
    .A2(_0279_));
 sg13g2_nor2_1 _2295_ (.A(_0280_),
    .B(_0281_),
    .Y(_0072_));
 sg13g2_nor2b_1 _2296_ (.A(_0702_),
    .B_N(_0279_),
    .Y(_0282_));
 sg13g2_o21ai_1 _2297_ (.B1(net591),
    .Y(_0283_),
    .A1(net95),
    .A2(_0280_));
 sg13g2_nor2_1 _2298_ (.A(_0282_),
    .B(net96),
    .Y(_0073_));
 sg13g2_o21ai_1 _2299_ (.B1(net591),
    .Y(_0284_),
    .A1(net93),
    .A2(_0282_));
 sg13g2_a21oi_1 _2300_ (.A1(net93),
    .A2(_0282_),
    .Y(_0074_),
    .B1(_0284_));
 sg13g2_a22oi_1 _2301_ (.Y(_0285_),
    .B1(net481),
    .B2(net69),
    .A2(_0916_),
    .A1(\u8.rcop[0] ));
 sg13g2_nor2_1 _2302_ (.A(_0947_),
    .B(net70),
    .Y(_0075_));
 sg13g2_a21oi_1 _2303_ (.A1(_0395_),
    .A2(net106),
    .Y(_0286_),
    .B1(_0947_));
 sg13g2_nor2b_1 _2304_ (.A(_0918_),
    .B_N(net107),
    .Y(_0076_));
 sg13g2_o21ai_1 _2305_ (.B1(net556),
    .Y(_0287_),
    .A1(net80),
    .A2(_0918_));
 sg13g2_nor2_1 _2306_ (.A(_0919_),
    .B(net81),
    .Y(_0077_));
 sg13g2_xnor2_1 _2307_ (.Y(_0288_),
    .A(net102),
    .B(_0914_));
 sg13g2_nor2_1 _2308_ (.A(_0947_),
    .B(_0288_),
    .Y(_0078_));
 sg13g2_a21oi_1 _2309_ (.A1(\u8.rbop[0] ),
    .A2(_0914_),
    .Y(_0289_),
    .B1(net75));
 sg13g2_and3_1 _2310_ (.X(_0290_),
    .A(net75),
    .B(\u8.rbop[0] ),
    .C(_0914_));
 sg13g2_nor3_1 _2311_ (.A(_0947_),
    .B(net76),
    .C(_0290_),
    .Y(_0079_));
 sg13g2_a21oi_1 _2312_ (.A1(_0901_),
    .A2(_0914_),
    .Y(_0291_),
    .B1(_0947_));
 sg13g2_o21ai_1 _2313_ (.B1(_0291_),
    .Y(_0292_),
    .A1(net73),
    .A2(_0290_));
 sg13g2_a21oi_1 _2314_ (.A1(net73),
    .A2(_0290_),
    .Y(_0080_),
    .B1(_0292_));
 sg13g2_o21ai_1 _2315_ (.B1(net556),
    .Y(_0293_),
    .A1(net71),
    .A2(_0930_));
 sg13g2_a21oi_1 _2316_ (.A1(_0393_),
    .A2(_0930_),
    .Y(_0081_),
    .B1(_0293_));
 sg13g2_o21ai_1 _2317_ (.B1(net556),
    .Y(_0294_),
    .A1(net516),
    .A2(_0929_));
 sg13g2_a21oi_1 _2318_ (.A1(net99),
    .A2(_0929_),
    .Y(_0082_),
    .B1(_0294_));
 sg13g2_and3_1 _2319_ (.X(_0295_),
    .A(net516),
    .B(\u8.ruop[0] ),
    .C(_0929_));
 sg13g2_o21ai_1 _2320_ (.B1(net556),
    .Y(_0296_),
    .A1(net83),
    .A2(_0295_));
 sg13g2_a21oi_1 _2321_ (.A1(net83),
    .A2(_0295_),
    .Y(_0083_),
    .B1(_0296_));
 sg13g2_nor4_2 _2322_ (.A(_0699_),
    .B(_0700_),
    .C(_0704_),
    .Y(_0297_),
    .D(_0112_));
 sg13g2_and2_1 _2323_ (.A(net485),
    .B(net463),
    .X(_0298_));
 sg13g2_nand2_1 _2324_ (.Y(_0299_),
    .A(net485),
    .B(net463));
 sg13g2_a21oi_1 _2325_ (.A1(net534),
    .A2(net457),
    .Y(_0300_),
    .B1(_0738_));
 sg13g2_o21ai_1 _2326_ (.B1(_0300_),
    .Y(_0301_),
    .A1(net520),
    .A2(_0299_));
 sg13g2_nor2_2 _2327_ (.A(net562),
    .B(_0743_),
    .Y(_0302_));
 sg13g2_a21oi_1 _2328_ (.A1(net584),
    .A2(_0001_),
    .Y(_0303_),
    .B1(_0183_));
 sg13g2_a22oi_1 _2329_ (.Y(_0304_),
    .B1(_0303_),
    .B2(net488),
    .A2(_0302_),
    .A1(net534));
 sg13g2_nor2_1 _2330_ (.A(_0683_),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_a21oi_1 _2331_ (.A1(net529),
    .A2(net475),
    .Y(_0306_),
    .B1(net467));
 sg13g2_a21oi_1 _2332_ (.A1(net530),
    .A2(net469),
    .Y(_0307_),
    .B1(_1071_));
 sg13g2_o21ai_1 _2333_ (.B1(net500),
    .Y(_0308_),
    .A1(_0306_),
    .A2(_0307_));
 sg13g2_a221oi_1 _2334_ (.B2(_0712_),
    .C1(_0305_),
    .B1(_0308_),
    .A1(_0684_),
    .Y(_0309_),
    .A2(_0301_));
 sg13g2_o21ai_1 _2335_ (.B1(net593),
    .Y(_0310_),
    .A1(net514),
    .A2(net446));
 sg13g2_a21oi_1 _2336_ (.A1(net446),
    .A2(_0309_),
    .Y(_0084_),
    .B1(_0310_));
 sg13g2_nor2_1 _2337_ (.A(_0750_),
    .B(_0950_),
    .Y(_0311_));
 sg13g2_a22oi_1 _2338_ (.Y(_0312_),
    .B1(_0311_),
    .B2(net488),
    .A2(_0302_),
    .A1(net531));
 sg13g2_nand2_1 _2339_ (.Y(_0313_),
    .A(net531),
    .B(net457));
 sg13g2_or2_1 _2340_ (.X(_0314_),
    .B(_0524_),
    .A(_0448_));
 sg13g2_o21ai_1 _2341_ (.B1(_0313_),
    .Y(_0315_),
    .A1(_0299_),
    .A2(_0314_));
 sg13g2_a21oi_1 _2342_ (.A1(net527),
    .A2(net475),
    .Y(_0316_),
    .B1(net467));
 sg13g2_nor2_1 _2343_ (.A(_0005_),
    .B(_0732_),
    .Y(_0317_));
 sg13g2_a21oi_1 _2344_ (.A1(net527),
    .A2(_0724_),
    .Y(_0318_),
    .B1(_0317_));
 sg13g2_o21ai_1 _2345_ (.B1(net500),
    .Y(_0319_),
    .A1(_0316_),
    .A2(_0318_));
 sg13g2_a221oi_1 _2346_ (.B2(_0711_),
    .C1(net558),
    .B1(_0319_),
    .A1(_0762_),
    .Y(_0320_),
    .A2(_0315_));
 sg13g2_a21o_1 _2347_ (.A2(_0312_),
    .A1(net559),
    .B1(_0320_),
    .X(_0321_));
 sg13g2_o21ai_1 _2348_ (.B1(net590),
    .Y(_0322_),
    .A1(net511),
    .A2(net446));
 sg13g2_a21oi_1 _2349_ (.A1(net446),
    .A2(_0321_),
    .Y(_0085_),
    .B1(_0322_));
 sg13g2_xnor2_1 _2350_ (.Y(_0323_),
    .A(_0391_),
    .B(_0448_));
 sg13g2_a22oi_1 _2351_ (.Y(_0324_),
    .B1(_0298_),
    .B2(_0323_),
    .A2(net457),
    .A1(net529));
 sg13g2_nand2_2 _2352_ (.Y(_0325_),
    .A(_0683_),
    .B(net476));
 sg13g2_nor2_1 _2353_ (.A(_0006_),
    .B(_0732_),
    .Y(_0326_));
 sg13g2_a21oi_1 _2354_ (.A1(net525),
    .A2(_0724_),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_a21oi_1 _2355_ (.A1(net525),
    .A2(net475),
    .Y(_0328_),
    .B1(net467));
 sg13g2_nor3_1 _2356_ (.A(net498),
    .B(_0327_),
    .C(_0328_),
    .Y(_0329_));
 sg13g2_nor2_1 _2357_ (.A(_0772_),
    .B(_0857_),
    .Y(_0330_));
 sg13g2_a22oi_1 _2358_ (.Y(_0331_),
    .B1(_0330_),
    .B2(net488),
    .A2(_0302_),
    .A1(net529));
 sg13g2_a22oi_1 _2359_ (.Y(_0332_),
    .B1(_0331_),
    .B2(net558),
    .A2(_0324_),
    .A1(_0107_));
 sg13g2_o21ai_1 _2360_ (.B1(_0332_),
    .Y(_0333_),
    .A1(_0325_),
    .A2(_0329_));
 sg13g2_o21ai_1 _2361_ (.B1(net587),
    .Y(_0334_),
    .A1(net510),
    .A2(net445));
 sg13g2_a21oi_1 _2362_ (.A1(net445),
    .A2(_0333_),
    .Y(_0086_),
    .B1(_0334_));
 sg13g2_xnor2_1 _2363_ (.Y(_0335_),
    .A(_0028_),
    .B(_0449_));
 sg13g2_a22oi_1 _2364_ (.Y(_0336_),
    .B1(_0298_),
    .B2(_0335_),
    .A2(net457),
    .A1(net527));
 sg13g2_nor2_1 _2365_ (.A(_0029_),
    .B(_0732_),
    .Y(_0337_));
 sg13g2_a21oi_1 _2366_ (.A1(net522),
    .A2(net469),
    .Y(_0338_),
    .B1(_0337_));
 sg13g2_a21oi_1 _2367_ (.A1(net522),
    .A2(net475),
    .Y(_0339_),
    .B1(net467));
 sg13g2_nor3_1 _2368_ (.A(net498),
    .B(_0338_),
    .C(_0339_),
    .Y(_0340_));
 sg13g2_nor2_1 _2369_ (.A(_0776_),
    .B(_0965_),
    .Y(_0341_));
 sg13g2_a22oi_1 _2370_ (.Y(_0342_),
    .B1(_0341_),
    .B2(net488),
    .A2(_0302_),
    .A1(net527));
 sg13g2_a22oi_1 _2371_ (.Y(_0343_),
    .B1(_0342_),
    .B2(net558),
    .A2(_0336_),
    .A1(_0107_));
 sg13g2_o21ai_1 _2372_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0325_),
    .A2(_0340_));
 sg13g2_o21ai_1 _2373_ (.B1(net590),
    .Y(_0345_),
    .A1(net508),
    .A2(net446));
 sg13g2_a21oi_1 _2374_ (.A1(net446),
    .A2(_0344_),
    .Y(_0087_),
    .B1(_0345_));
 sg13g2_nor2b_1 _2375_ (.A(_0728_),
    .B_N(net486),
    .Y(_0346_));
 sg13g2_a22oi_1 _2376_ (.Y(_0347_),
    .B1(_0346_),
    .B2(_0642_),
    .A2(net457),
    .A1(net525));
 sg13g2_nor2_1 _2377_ (.A(_0007_),
    .B(_0732_),
    .Y(_0348_));
 sg13g2_a21oi_1 _2378_ (.A1(net519),
    .A2(net469),
    .Y(_0349_),
    .B1(_0348_));
 sg13g2_a21oi_1 _2379_ (.A1(net519),
    .A2(net475),
    .Y(_0350_),
    .B1(net467));
 sg13g2_nor3_1 _2380_ (.A(net498),
    .B(_0349_),
    .C(_0350_),
    .Y(_0351_));
 sg13g2_nand3_1 _2381_ (.B(_1077_),
    .C(net488),
    .A(_0795_),
    .Y(_0352_));
 sg13g2_a21oi_1 _2382_ (.A1(net525),
    .A2(_0302_),
    .Y(_0353_),
    .B1(_0683_));
 sg13g2_a22oi_1 _2383_ (.Y(_0354_),
    .B1(_0352_),
    .B2(_0353_),
    .A2(_0347_),
    .A1(_0107_));
 sg13g2_o21ai_1 _2384_ (.B1(_0354_),
    .Y(_0355_),
    .A1(_0325_),
    .A2(_0351_));
 sg13g2_o21ai_1 _2385_ (.B1(net590),
    .Y(_0356_),
    .A1(net506),
    .A2(net446));
 sg13g2_a21oi_1 _2386_ (.A1(net446),
    .A2(_0355_),
    .Y(_0088_),
    .B1(_0356_));
 sg13g2_a22oi_1 _2387_ (.Y(_0357_),
    .B1(_0733_),
    .B2(_0429_),
    .A2(_0723_),
    .A1(net517));
 sg13g2_a21oi_1 _2388_ (.A1(net517),
    .A2(net473),
    .Y(_0358_),
    .B1(net466));
 sg13g2_nor3_1 _2389_ (.A(net498),
    .B(_0357_),
    .C(_0358_),
    .Y(_0359_));
 sg13g2_nor2b_1 _2390_ (.A(_0802_),
    .B_N(_1118_),
    .Y(_0360_));
 sg13g2_a22oi_1 _2391_ (.Y(_0361_),
    .B1(net488),
    .B2(_0360_),
    .A2(_1112_),
    .A1(_0742_));
 sg13g2_nand2b_1 _2392_ (.Y(_0362_),
    .B(net458),
    .A_N(_0029_));
 sg13g2_a22oi_1 _2393_ (.Y(_0363_),
    .B1(_0362_),
    .B2(_0684_),
    .A2(_0361_),
    .A1(_0682_));
 sg13g2_o21ai_1 _2394_ (.B1(_0363_),
    .Y(_0364_),
    .A1(_0325_),
    .A2(_0359_));
 sg13g2_o21ai_1 _2395_ (.B1(net587),
    .Y(_0365_),
    .A1(net503),
    .A2(net445));
 sg13g2_a21oi_1 _2396_ (.A1(net445),
    .A2(_0364_),
    .Y(_0089_),
    .B1(_0365_));
 sg13g2_nor2b_1 _2397_ (.A(_0810_),
    .B_N(_1144_),
    .Y(_0366_));
 sg13g2_a22oi_1 _2398_ (.Y(_0367_),
    .B1(_0366_),
    .B2(net488),
    .A2(_0302_),
    .A1(net519));
 sg13g2_a22oi_1 _2399_ (.Y(_0368_),
    .B1(_0733_),
    .B2(_0430_),
    .A2(_0723_),
    .A1(net513));
 sg13g2_and2_1 _2400_ (.A(net513),
    .B(net474),
    .X(_0369_));
 sg13g2_o21ai_1 _2401_ (.B1(net500),
    .Y(_0370_),
    .A1(net467),
    .A2(_0369_));
 sg13g2_o21ai_1 _2402_ (.B1(net476),
    .Y(_0371_),
    .A1(_0368_),
    .A2(_0370_));
 sg13g2_o21ai_1 _2403_ (.B1(_0762_),
    .Y(_0372_),
    .A1(_0007_),
    .A2(net456));
 sg13g2_a21oi_1 _2404_ (.A1(_0371_),
    .A2(_0372_),
    .Y(_0373_),
    .B1(net558));
 sg13g2_a21o_1 _2405_ (.A2(_0367_),
    .A1(net558),
    .B1(_0373_),
    .X(_0374_));
 sg13g2_o21ai_1 _2406_ (.B1(net587),
    .Y(_0375_),
    .A1(net109),
    .A2(net445));
 sg13g2_a21oi_1 _2407_ (.A1(net445),
    .A2(_0374_),
    .Y(_0090_),
    .B1(_0375_));
 sg13g2_a22oi_1 _2408_ (.Y(_0376_),
    .B1(_0733_),
    .B2(_0415_),
    .A2(_0723_),
    .A1(net512));
 sg13g2_a21oi_1 _2409_ (.A1(net512),
    .A2(net473),
    .Y(_0377_),
    .B1(net466));
 sg13g2_nor3_1 _2410_ (.A(net498),
    .B(_0376_),
    .C(_0377_),
    .Y(_0378_));
 sg13g2_nor2b_1 _2411_ (.A(_0818_),
    .B_N(_1175_),
    .Y(_0379_));
 sg13g2_a22oi_1 _2412_ (.Y(_0380_),
    .B1(_0379_),
    .B2(net488),
    .A2(_0302_),
    .A1(net517));
 sg13g2_nand2_1 _2413_ (.Y(_0381_),
    .A(_0429_),
    .B(net458));
 sg13g2_a22oi_1 _2414_ (.Y(_0382_),
    .B1(_0381_),
    .B2(_0107_),
    .A2(_0380_),
    .A1(net558));
 sg13g2_o21ai_1 _2415_ (.B1(_0382_),
    .Y(_0383_),
    .A1(_0325_),
    .A2(_0378_));
 sg13g2_o21ai_1 _2416_ (.B1(net587),
    .Y(_0384_),
    .A1(net104),
    .A2(net445));
 sg13g2_a21oi_1 _2417_ (.A1(net445),
    .A2(_0383_),
    .Y(_0091_),
    .B1(_0384_));
 sg13g2_dfrbp_1 _2418_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net41),
    .D(_0038_),
    .Q_N(_0019_),
    .Q(\u8.rc[24] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net30),
    .D(_0039_),
    .Q_N(_0026_),
    .Q(\u8.rc[25] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net28),
    .D(_0040_),
    .Q_N(_0018_),
    .Q(\u8.rc[26] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net26),
    .D(_0041_),
    .Q_N(_0020_),
    .Q(\u8.rc[27] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net24),
    .D(_0042_),
    .Q_N(_1204_),
    .Q(\u8.rc[28] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net22),
    .D(_0043_),
    .Q_N(_0025_),
    .Q(\u8.rc[29] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net20),
    .D(_0044_),
    .Q_N(_1203_),
    .Q(\u8.rc[30] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net18),
    .D(_0045_),
    .Q_N(_0024_),
    .Q(\u8.rc[31] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net16),
    .D(_0046_),
    .Q_N(_1202_),
    .Q(retry));
 sg13g2_dfrbp_1 _2427_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net68),
    .D(net91),
    .Q_N(_1201_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _2428_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net66),
    .D(_0048_),
    .Q_N(_1200_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _2429_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net64),
    .D(_0049_),
    .Q_N(_1199_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _2430_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net62),
    .D(_0050_),
    .Q_N(_1198_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net60),
    .D(_0051_),
    .Q_N(_1197_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net58),
    .D(_0052_),
    .Q_N(_1196_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net56),
    .D(_0053_),
    .Q_N(_1195_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net54),
    .D(_0054_),
    .Q_N(_1194_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net52),
    .D(_0055_),
    .Q_N(_0017_),
    .Q(\u8.empty ));
 sg13g2_dfrbp_1 _2436_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net50),
    .D(_0056_),
    .Q_N(_0000_),
    .Q(\u8.ls[0] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net48),
    .D(_0057_),
    .Q_N(_0002_),
    .Q(\u8.ls[1] ));
 sg13g2_dfrbp_1 _2438_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net46),
    .D(_0058_),
    .Q_N(_0030_),
    .Q(\u8.ls[2] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net44),
    .D(_0059_),
    .Q_N(_0031_),
    .Q(\u8.ls[3] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net42),
    .D(_0060_),
    .Q_N(_0032_),
    .Q(\u8.ls[4] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net40),
    .D(_0061_),
    .Q_N(_0033_),
    .Q(\u8.ls[5] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net38),
    .D(_0062_),
    .Q_N(_0034_),
    .Q(\u8.ls[6] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net36),
    .D(_0063_),
    .Q_N(_0021_),
    .Q(\u8.ls[7] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net34),
    .D(_0064_),
    .Q_N(_0001_),
    .Q(\u8.ls[8] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net32),
    .D(_0065_),
    .Q_N(_0003_),
    .Q(\u8.ls[9] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net29),
    .D(_0066_),
    .Q_N(_0004_),
    .Q(\u8.hs[0] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net25),
    .D(_0067_),
    .Q_N(_0005_),
    .Q(\u8.hs[1] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net21),
    .D(_0068_),
    .Q_N(_0006_),
    .Q(\u8.hs[2] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net17),
    .D(_0069_),
    .Q_N(_0029_),
    .Q(\u8.hs[3] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net67),
    .D(_0070_),
    .Q_N(_0007_),
    .Q(\u8.hs[4] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net63),
    .D(_0071_),
    .Q_N(_0008_),
    .Q(\u8.hs[5] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net59),
    .D(_0072_),
    .Q_N(_1193_),
    .Q(\u8.rcip[0] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net55),
    .D(_0073_),
    .Q_N(_1192_),
    .Q(\u8.rcip[1] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net51),
    .D(net94),
    .Q_N(_0023_),
    .Q(\u8.rcip[2] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net47),
    .D(_0075_),
    .Q_N(_0037_),
    .Q(\u8.rcop[0] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net43),
    .D(net108),
    .Q_N(_1191_),
    .Q(\u8.rcop[1] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net39),
    .D(net82),
    .Q_N(_0012_),
    .Q(\u8.rcop[2] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net35),
    .D(_0078_),
    .Q_N(_1190_),
    .Q(\u8.rbop[0] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net31),
    .D(_0079_),
    .Q_N(_0022_),
    .Q(\u8.rbop[1] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net23),
    .D(net74),
    .Q_N(_0016_),
    .Q(\u8.rbop[2] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net15),
    .D(net72),
    .Q_N(_0036_),
    .Q(\u8.ruop[0] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net61),
    .D(net100),
    .Q_N(_1189_),
    .Q(\u8.ruop[1] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net53),
    .D(net84),
    .Q_N(_0035_),
    .Q(\u8.ruop[2] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net45),
    .D(_0084_),
    .Q_N(_0009_),
    .Q(\u8.rc[16] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net37),
    .D(_0085_),
    .Q_N(_0028_),
    .Q(\u8.rc[17] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net27),
    .D(_0086_),
    .Q_N(_0010_),
    .Q(\u8.rc[18] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net65),
    .D(_0087_),
    .Q_N(_0011_),
    .Q(\u8.rc[19] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net49),
    .D(_0088_),
    .Q_N(_0013_),
    .Q(\u8.rc[20] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net33),
    .D(_0089_),
    .Q_N(_0027_),
    .Q(\u8.rc[21] ));
 sg13g2_dfrbp_1 _2470_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net57),
    .D(_0090_),
    .Q_N(_0014_),
    .Q(\u8.rc[22] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net19),
    .D(_0091_),
    .Q_N(_0015_),
    .Q(\u8.rc[23] ));
 sg13g2_tiehi _2426__16 (.L_HI(net16));
 sg13g2_tiehi _2449__17 (.L_HI(net17));
 sg13g2_tiehi _2425__18 (.L_HI(net18));
 sg13g2_tiehi _2471__19 (.L_HI(net19));
 sg13g2_tiehi _2424__20 (.L_HI(net20));
 sg13g2_tiehi _2448__21 (.L_HI(net21));
 sg13g2_tiehi _2423__22 (.L_HI(net22));
 sg13g2_tiehi _2460__23 (.L_HI(net23));
 sg13g2_tiehi _2422__24 (.L_HI(net24));
 sg13g2_tiehi _2447__25 (.L_HI(net25));
 sg13g2_tiehi _2421__26 (.L_HI(net26));
 sg13g2_tiehi _2466__27 (.L_HI(net27));
 sg13g2_tiehi _2420__28 (.L_HI(net28));
 sg13g2_tiehi _2446__29 (.L_HI(net29));
 sg13g2_tiehi _2419__30 (.L_HI(net30));
 sg13g2_tiehi _2459__31 (.L_HI(net31));
 sg13g2_tiehi _2445__32 (.L_HI(net32));
 sg13g2_tiehi _2469__33 (.L_HI(net33));
 sg13g2_tiehi _2444__34 (.L_HI(net34));
 sg13g2_tiehi _2458__35 (.L_HI(net35));
 sg13g2_tiehi _2443__36 (.L_HI(net36));
 sg13g2_tiehi _2465__37 (.L_HI(net37));
 sg13g2_tiehi _2442__38 (.L_HI(net38));
 sg13g2_tiehi _2457__39 (.L_HI(net39));
 sg13g2_tiehi _2441__40 (.L_HI(net40));
 sg13g2_tiehi _2418__41 (.L_HI(net41));
 sg13g2_tiehi _2440__42 (.L_HI(net42));
 sg13g2_tiehi _2456__43 (.L_HI(net43));
 sg13g2_tiehi _2439__44 (.L_HI(net44));
 sg13g2_tiehi _2464__45 (.L_HI(net45));
 sg13g2_tiehi _2438__46 (.L_HI(net46));
 sg13g2_tiehi _2455__47 (.L_HI(net47));
 sg13g2_tiehi _2437__48 (.L_HI(net48));
 sg13g2_tiehi _2468__49 (.L_HI(net49));
 sg13g2_tiehi _2436__50 (.L_HI(net50));
 sg13g2_tiehi _2454__51 (.L_HI(net51));
 sg13g2_tiehi _2435__52 (.L_HI(net52));
 sg13g2_tiehi _2463__53 (.L_HI(net53));
 sg13g2_tiehi _2434__54 (.L_HI(net54));
 sg13g2_tiehi _2453__55 (.L_HI(net55));
 sg13g2_tiehi _2433__56 (.L_HI(net56));
 sg13g2_tiehi _2470__57 (.L_HI(net57));
 sg13g2_tiehi _2432__58 (.L_HI(net58));
 sg13g2_tiehi _2452__59 (.L_HI(net59));
 sg13g2_tiehi _2431__60 (.L_HI(net60));
 sg13g2_tiehi _2462__61 (.L_HI(net61));
 sg13g2_tiehi _2430__62 (.L_HI(net62));
 sg13g2_tiehi _2451__63 (.L_HI(net63));
 sg13g2_tiehi _2429__64 (.L_HI(net64));
 sg13g2_tiehi _2467__65 (.L_HI(net65));
 sg13g2_tiehi _2428__66 (.L_HI(net66));
 sg13g2_tiehi _2450__67 (.L_HI(net67));
 sg13g2_tiehi _2427__68 (.L_HI(net68));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _2526_ (.A(net565),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2527_ (.A(net565),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2528_ (.A(net565),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2529_ (.A(net564),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2530_ (.A(net564),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2531_ (.A(net564),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2532_ (.A(net564),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2533_ (.A(net564),
    .X(uio_oe[7]));
 sg13g2_buf_2 fanout445 (.A(_0297_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_0297_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net452),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(net452),
    .X(net450));
 sg13g2_buf_1 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_1 fanout452 (.A(_0117_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_0931_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_0709_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_0709_),
    .X(net455));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(_0691_));
 sg13g2_buf_2 fanout457 (.A(net458),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_0690_),
    .X(net459));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(net464));
 sg13g2_buf_1 fanout461 (.A(net464),
    .X(net461));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(net464));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_0873_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_0736_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net467),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_0714_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(net469),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_0724_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net471),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_0643_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_0643_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_0718_),
    .X(net475));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(_0765_));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(_0712_));
 sg13g2_buf_2 fanout478 (.A(_0639_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_0121_),
    .X(net479));
 sg13g2_buf_1 fanout480 (.A(_0121_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_0934_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net483),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_0835_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_0835_),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(_0542_));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(_0114_));
 sg13g2_buf_2 fanout489 (.A(_0935_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_0902_),
    .X(net490));
 sg13g2_buf_1 fanout491 (.A(_0902_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_0865_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_0865_),
    .X(net493));
 sg13g2_buf_4 fanout494 (.X(net494),
    .A(net495));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(_0848_));
 sg13g2_buf_2 fanout496 (.A(_0847_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_0847_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_0660_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(_0659_));
 sg13g2_buf_2 fanout502 (.A(_0936_),
    .X(net502));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(net110));
 sg13g2_buf_1 fanout504 (.A(\u8.rc[21] ),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(\u8.rc[20] ),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(\u8.rc[19] ),
    .X(net509));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(\u8.rc[18] ));
 sg13g2_buf_2 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_4 fanout512 (.X(net512),
    .A(\u8.rc[17] ));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(\u8.rc[16] ));
 sg13g2_buf_2 fanout514 (.A(net111),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(\u8.ruop[1] ),
    .X(net516));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net112));
 sg13g2_buf_2 fanout518 (.A(\u8.hs[5] ),
    .X(net518));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(\u8.hs[4] ));
 sg13g2_buf_2 fanout520 (.A(net115),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net523),
    .X(net522));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(\u8.hs[3] ));
 sg13g2_buf_2 fanout524 (.A(net525),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(\u8.hs[2] ));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(net528));
 sg13g2_buf_2 fanout528 (.A(\u8.hs[1] ),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(\u8.hs[0] ),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(\u8.ls[9] ),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_1 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(\u8.ls[8] ),
    .X(net535));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net119));
 sg13g2_buf_2 fanout537 (.A(\u8.ls[7] ),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(net539),
    .X(net538));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(\u8.ls[6] ));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net113));
 sg13g2_buf_1 fanout541 (.A(\u8.ls[5] ),
    .X(net541));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(net124));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(net123));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(\u8.ls[2] ));
 sg13g2_buf_2 fanout545 (.A(_0017_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(\u8.rc[31] ));
 sg13g2_buf_2 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net114),
    .X(net550));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(net121));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(net116));
 sg13g2_buf_2 fanout553 (.A(net122),
    .X(net553));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(net118));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(\u8.rc[25] ));
 sg13g2_buf_2 fanout556 (.A(_0946_),
    .X(net556));
 sg13g2_buf_1 fanout557 (.A(_0946_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_0682_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net563),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net563),
    .X(net561));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(net563));
 sg13g2_buf_2 fanout563 (.A(_0419_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net566),
    .X(net564));
 sg13g2_buf_1 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_1 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(ui_in[4]));
 sg13g2_buf_2 fanout568 (.A(net572),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(net572),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net577),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net577),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net577),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net586),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net586),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net583),
    .X(net581));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(net583));
 sg13g2_buf_2 fanout583 (.A(net585),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(ui_in[3]),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net589),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net593),
    .X(net589));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(net593));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(rst_n),
    .X(net593));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[5]));
 sg13g2_buf_2 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_buf_2 input14 (.A(uio_in[7]),
    .X(net14));
 sg13g2_tiehi _2461__15 (.L_HI(net15));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0037_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0285_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0036_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0081_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u8.rbop[2] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0080_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold7 (.A(\u8.rbop[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0289_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold9 (.A(retry),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u8.empty ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold11 (.A(uio_out[4]),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u8.rcop[2] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0287_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0077_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u8.ruop[2] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0083_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold17 (.A(uio_out[2]),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold18 (.A(uio_out[5]),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold19 (.A(uio_out[3]),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold20 (.A(uio_out[1]),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold21 (.A(uio_out[7]),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold22 (.A(uio_out[0]),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0047_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u8.rc[25] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u8.rcip[2] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0074_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u8.rcip[1] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0283_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold29 (.A(uio_out[6]),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold30 (.A(\u8.ruop[0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0875_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0082_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u8.rcip[0] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u8.rbop[0] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u8.rc[24] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u8.rc[23] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0012_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0917_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0286_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0076_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u8.rc[22] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u8.rc[21] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u8.rc[16] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold44 (.A(\u8.hs[5] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u8.ls[5] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold46 (.A(\u8.rc[30] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u8.hs[4] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u8.rc[28] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u8.ls[1] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u8.rc[26] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u8.ls[7] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u8.ls[0] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u8.rc[29] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u8.rc[27] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u8.ls[3] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u8.ls[4] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u8.rcip[0] ),
    .X(net125));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_fill_2 FILLER_7_231 ();
 sg13g2_fill_1 FILLER_7_233 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_4 FILLER_8_147 ();
 sg13g2_fill_2 FILLER_8_164 ();
 sg13g2_decap_8 FILLER_8_171 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_189 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_decap_4 FILLER_8_228 ();
 sg13g2_fill_1 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_290 ();
 sg13g2_decap_4 FILLER_8_297 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_decap_4 FILLER_9_202 ();
 sg13g2_fill_1 FILLER_9_228 ();
 sg13g2_decap_4 FILLER_9_244 ();
 sg13g2_decap_4 FILLER_9_256 ();
 sg13g2_fill_1 FILLER_9_267 ();
 sg13g2_fill_2 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_285 ();
 sg13g2_fill_2 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_fill_1 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_4 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_1 FILLER_10_166 ();
 sg13g2_fill_2 FILLER_10_172 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_fill_2 FILLER_10_189 ();
 sg13g2_fill_1 FILLER_10_191 ();
 sg13g2_fill_2 FILLER_10_202 ();
 sg13g2_decap_4 FILLER_10_209 ();
 sg13g2_fill_1 FILLER_10_213 ();
 sg13g2_fill_1 FILLER_10_227 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_fill_1 FILLER_10_240 ();
 sg13g2_fill_2 FILLER_10_246 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_decap_4 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_286 ();
 sg13g2_fill_2 FILLER_10_303 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_4 FILLER_10_349 ();
 sg13g2_fill_2 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_4 FILLER_11_105 ();
 sg13g2_decap_4 FILLER_11_135 ();
 sg13g2_fill_2 FILLER_11_139 ();
 sg13g2_fill_1 FILLER_11_145 ();
 sg13g2_fill_2 FILLER_11_172 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_185 ();
 sg13g2_fill_1 FILLER_11_187 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_fill_2 FILLER_11_238 ();
 sg13g2_fill_1 FILLER_11_270 ();
 sg13g2_fill_2 FILLER_11_285 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_fill_1 FILLER_11_320 ();
 sg13g2_decap_4 FILLER_11_339 ();
 sg13g2_fill_1 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_fill_1 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_117 ();
 sg13g2_fill_1 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_124 ();
 sg13g2_decap_4 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_161 ();
 sg13g2_decap_4 FILLER_12_185 ();
 sg13g2_decap_4 FILLER_12_203 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_fill_2 FILLER_12_212 ();
 sg13g2_fill_2 FILLER_12_227 ();
 sg13g2_fill_2 FILLER_12_238 ();
 sg13g2_fill_2 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_261 ();
 sg13g2_decap_4 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_272 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_279 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_fill_2 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_338 ();
 sg13g2_decap_4 FILLER_12_355 ();
 sg13g2_fill_1 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_4 FILLER_12_383 ();
 sg13g2_fill_2 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_2 FILLER_13_138 ();
 sg13g2_fill_2 FILLER_13_146 ();
 sg13g2_fill_2 FILLER_13_174 ();
 sg13g2_fill_1 FILLER_13_176 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_decap_4 FILLER_13_255 ();
 sg13g2_fill_2 FILLER_13_259 ();
 sg13g2_decap_4 FILLER_13_266 ();
 sg13g2_fill_1 FILLER_13_270 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_decap_4 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_343 ();
 sg13g2_fill_2 FILLER_13_389 ();
 sg13g2_fill_1 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_4 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_107 ();
 sg13g2_fill_2 FILLER_14_114 ();
 sg13g2_fill_1 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_decap_4 FILLER_14_176 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_220 ();
 sg13g2_decap_8 FILLER_14_227 ();
 sg13g2_fill_2 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_273 ();
 sg13g2_fill_2 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_283 ();
 sg13g2_fill_1 FILLER_14_297 ();
 sg13g2_fill_2 FILLER_14_317 ();
 sg13g2_fill_1 FILLER_14_319 ();
 sg13g2_decap_4 FILLER_14_339 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_fill_1 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_4 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_4 FILLER_15_88 ();
 sg13g2_decap_4 FILLER_15_118 ();
 sg13g2_fill_2 FILLER_15_122 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_192 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_2 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_229 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_fill_2 FILLER_15_307 ();
 sg13g2_decap_4 FILLER_15_317 ();
 sg13g2_decap_4 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_fill_2 FILLER_15_360 ();
 sg13g2_fill_1 FILLER_15_370 ();
 sg13g2_fill_1 FILLER_15_377 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_4 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_decap_4 FILLER_16_87 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_106 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_155 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_fill_2 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_335 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_4 FILLER_16_358 ();
 sg13g2_fill_2 FILLER_16_362 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_4 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_32 ();
 sg13g2_decap_8 FILLER_17_37 ();
 sg13g2_fill_2 FILLER_17_44 ();
 sg13g2_fill_1 FILLER_17_46 ();
 sg13g2_fill_1 FILLER_17_50 ();
 sg13g2_fill_1 FILLER_17_81 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_decap_4 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_148 ();
 sg13g2_decap_4 FILLER_17_158 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_decap_4 FILLER_17_222 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_232 ();
 sg13g2_decap_8 FILLER_17_239 ();
 sg13g2_decap_4 FILLER_17_246 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_fill_1 FILLER_17_264 ();
 sg13g2_fill_1 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_decap_4 FILLER_17_295 ();
 sg13g2_decap_4 FILLER_17_317 ();
 sg13g2_fill_1 FILLER_17_346 ();
 sg13g2_decap_4 FILLER_17_355 ();
 sg13g2_fill_1 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_376 ();
 sg13g2_fill_2 FILLER_17_393 ();
 sg13g2_fill_1 FILLER_17_395 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_68 ();
 sg13g2_decap_8 FILLER_18_94 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_135 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_decap_4 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_189 ();
 sg13g2_fill_1 FILLER_18_191 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_4 FILLER_18_280 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_decap_4 FILLER_18_305 ();
 sg13g2_decap_4 FILLER_18_314 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_decap_4 FILLER_18_365 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_fill_2 FILLER_18_388 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_11 ();
 sg13g2_fill_2 FILLER_19_25 ();
 sg13g2_fill_1 FILLER_19_27 ();
 sg13g2_fill_1 FILLER_19_33 ();
 sg13g2_fill_2 FILLER_19_41 ();
 sg13g2_fill_1 FILLER_19_43 ();
 sg13g2_fill_2 FILLER_19_58 ();
 sg13g2_decap_8 FILLER_19_65 ();
 sg13g2_fill_2 FILLER_19_85 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_fill_2 FILLER_19_118 ();
 sg13g2_fill_2 FILLER_19_131 ();
 sg13g2_decap_8 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_192 ();
 sg13g2_decap_4 FILLER_19_199 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_decap_4 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_fill_1 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_decap_4 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_340 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_350 ();
 sg13g2_decap_4 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_fill_2 FILLER_19_394 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_2 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_fill_1 FILLER_20_51 ();
 sg13g2_fill_2 FILLER_20_57 ();
 sg13g2_fill_1 FILLER_20_59 ();
 sg13g2_fill_2 FILLER_20_72 ();
 sg13g2_decap_8 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_fill_1 FILLER_20_196 ();
 sg13g2_decap_4 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_fill_2 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_4 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_fill_2 FILLER_20_361 ();
 sg13g2_fill_1 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_decap_4 FILLER_21_59 ();
 sg13g2_decap_8 FILLER_21_97 ();
 sg13g2_decap_8 FILLER_21_104 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_160 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_192 ();
 sg13g2_fill_2 FILLER_21_199 ();
 sg13g2_fill_1 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_214 ();
 sg13g2_decap_4 FILLER_21_220 ();
 sg13g2_fill_2 FILLER_21_224 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_decap_4 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_decap_4 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_decap_4 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_29 ();
 sg13g2_fill_1 FILLER_22_31 ();
 sg13g2_fill_2 FILLER_22_62 ();
 sg13g2_decap_4 FILLER_22_83 ();
 sg13g2_decap_8 FILLER_22_99 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_decap_4 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_148 ();
 sg13g2_decap_4 FILLER_22_155 ();
 sg13g2_fill_2 FILLER_22_163 ();
 sg13g2_fill_1 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_fill_2 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_decap_4 FILLER_22_191 ();
 sg13g2_fill_1 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_decap_8 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_226 ();
 sg13g2_decap_4 FILLER_22_233 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_287 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_decap_4 FILLER_22_359 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_51 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_decap_4 FILLER_23_58 ();
 sg13g2_fill_2 FILLER_23_62 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_2 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_fill_2 FILLER_23_146 ();
 sg13g2_fill_1 FILLER_23_163 ();
 sg13g2_fill_2 FILLER_23_169 ();
 sg13g2_fill_1 FILLER_23_175 ();
 sg13g2_fill_2 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_fill_2 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_286 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_fill_2 FILLER_23_295 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_decap_4 FILLER_23_334 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_369 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_fill_2 FILLER_24_38 ();
 sg13g2_fill_1 FILLER_24_40 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_fill_2 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_129 ();
 sg13g2_fill_2 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_169 ();
 sg13g2_fill_1 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_296 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_4 FILLER_24_394 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_16 ();
 sg13g2_fill_1 FILLER_25_22 ();
 sg13g2_fill_2 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_61 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_178 ();
 sg13g2_decap_8 FILLER_25_198 ();
 sg13g2_decap_4 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_decap_4 FILLER_25_295 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_2 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_fill_2 FILLER_26_66 ();
 sg13g2_fill_2 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_decap_4 FILLER_26_92 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_fill_2 FILLER_26_151 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_decap_4 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_213 ();
 sg13g2_fill_2 FILLER_26_219 ();
 sg13g2_decap_4 FILLER_26_226 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_decap_4 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_283 ();
 sg13g2_decap_4 FILLER_26_299 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_4 FILLER_26_344 ();
 sg13g2_decap_4 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_369 ();
 sg13g2_fill_2 FILLER_26_375 ();
 sg13g2_fill_1 FILLER_26_377 ();
 sg13g2_fill_1 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_26_397 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_43 ();
 sg13g2_fill_1 FILLER_27_55 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_decap_4 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_129 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_fill_2 FILLER_27_141 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_174 ();
 sg13g2_decap_8 FILLER_27_181 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_decap_4 FILLER_27_193 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_decap_8 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_277 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_307 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_4 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_decap_4 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_160 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_190 ();
 sg13g2_decap_4 FILLER_28_199 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_fill_2 FILLER_28_229 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_237 ();
 sg13g2_fill_2 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_fill_2 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_2 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_fill_1 FILLER_28_379 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_19 ();
 sg13g2_fill_1 FILLER_29_61 ();
 sg13g2_fill_2 FILLER_29_68 ();
 sg13g2_fill_1 FILLER_29_86 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_fill_2 FILLER_29_113 ();
 sg13g2_fill_1 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_134 ();
 sg13g2_decap_4 FILLER_29_149 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_4 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_193 ();
 sg13g2_fill_2 FILLER_29_200 ();
 sg13g2_decap_4 FILLER_29_207 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_233 ();
 sg13g2_decap_4 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_decap_4 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_decap_4 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_fill_2 FILLER_29_396 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_6 ();
 sg13g2_fill_1 FILLER_30_33 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_83 ();
 sg13g2_fill_1 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_fill_2 FILLER_30_143 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_decap_4 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_decap_4 FILLER_30_349 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_31_40 ();
 sg13g2_decap_4 FILLER_31_58 ();
 sg13g2_fill_2 FILLER_31_62 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_127 ();
 sg13g2_decap_4 FILLER_31_135 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_decap_4 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_decap_8 FILLER_31_208 ();
 sg13g2_fill_2 FILLER_31_215 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_386 ();
 sg13g2_fill_1 FILLER_31_388 ();
 sg13g2_fill_1 FILLER_31_397 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_87 ();
 sg13g2_fill_2 FILLER_32_94 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_32_352 ();
 sg13g2_fill_1 FILLER_32_366 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_27 ();
 sg13g2_fill_2 FILLER_33_65 ();
 sg13g2_fill_2 FILLER_33_86 ();
 sg13g2_decap_8 FILLER_33_92 ();
 sg13g2_fill_2 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_decap_4 FILLER_33_129 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_decap_4 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_4 FILLER_33_282 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_fill_1 FILLER_34_52 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_fill_2 FILLER_34_69 ();
 sg13g2_fill_1 FILLER_34_71 ();
 sg13g2_decap_4 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_154 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_2 FILLER_34_203 ();
 sg13g2_decap_4 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_decap_4 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_295 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_15 ();
 sg13g2_decap_4 FILLER_35_92 ();
 sg13g2_fill_2 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_107 ();
 sg13g2_fill_2 FILLER_35_129 ();
 sg13g2_fill_2 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_fill_2 FILLER_35_144 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_179 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_fill_1 FILLER_35_358 ();
 sg13g2_fill_2 FILLER_35_363 ();
 sg13g2_fill_2 FILLER_35_383 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_58 ();
 sg13g2_fill_2 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_65 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_fill_1 FILLER_36_81 ();
 sg13g2_decap_4 FILLER_36_113 ();
 sg13g2_fill_1 FILLER_36_117 ();
 sg13g2_fill_1 FILLER_36_131 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_4 FILLER_36_142 ();
 sg13g2_fill_2 FILLER_36_146 ();
 sg13g2_decap_4 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_fill_2 FILLER_36_219 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_239 ();
 sg13g2_decap_4 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_1 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_305 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_16 ();
 sg13g2_fill_1 FILLER_37_48 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_150 ();
 sg13g2_fill_1 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_166 ();
 sg13g2_decap_4 FILLER_37_198 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_210 ();
 sg13g2_fill_1 FILLER_37_221 ();
 sg13g2_decap_4 FILLER_37_227 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_271 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_327 ();
 sg13g2_fill_2 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_191 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_2 FILLER_38_378 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
endmodule

module tt_um_a1k0n_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire audio;
 wire hsync;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire \vgademo.a_cos[0] ;
 wire \vgademo.a_cos[10] ;
 wire \vgademo.a_cos[11] ;
 wire \vgademo.a_cos[12] ;
 wire \vgademo.a_cos[13] ;
 wire \vgademo.a_cos[14] ;
 wire \vgademo.a_cos[1] ;
 wire \vgademo.a_cos[2] ;
 wire \vgademo.a_cos[3] ;
 wire \vgademo.a_cos[4] ;
 wire \vgademo.a_cos[5] ;
 wire \vgademo.a_cos[6] ;
 wire \vgademo.a_cos[7] ;
 wire \vgademo.a_cos[8] ;
 wire \vgademo.a_cos[9] ;
 wire \vgademo.a_scrolly[10] ;
 wire \vgademo.a_scrolly[11] ;
 wire \vgademo.a_scrolly[12] ;
 wire \vgademo.a_scrolly[13] ;
 wire \vgademo.a_scrolly[3] ;
 wire \vgademo.a_scrolly[4] ;
 wire \vgademo.a_scrolly[5] ;
 wire \vgademo.a_scrolly[6] ;
 wire \vgademo.a_scrolly[7] ;
 wire \vgademo.a_scrolly[8] ;
 wire \vgademo.a_scrolly[9] ;
 wire \vgademo.a_sin[0] ;
 wire \vgademo.a_sin[10] ;
 wire \vgademo.a_sin[11] ;
 wire \vgademo.a_sin[12] ;
 wire \vgademo.a_sin[13] ;
 wire \vgademo.a_sin[14] ;
 wire \vgademo.a_sin[1] ;
 wire \vgademo.a_sin[2] ;
 wire \vgademo.a_sin[3] ;
 wire \vgademo.a_sin[4] ;
 wire \vgademo.a_sin[5] ;
 wire \vgademo.a_sin[6] ;
 wire \vgademo.a_sin[7] ;
 wire \vgademo.a_sin[8] ;
 wire \vgademo.a_sin[9] ;
 wire \vgademo.audio_beat_out[0] ;
 wire \vgademo.audio_beat_out[1] ;
 wire \vgademo.audio_beat_out[2] ;
 wire \vgademo.audio_beat_out[3] ;
 wire \vgademo.audio_beat_out[4] ;
 wire \vgademo.audio_kick_frames[0] ;
 wire \vgademo.audio_kick_frames[1] ;
 wire \vgademo.audio_kick_frames[2] ;
 wire \vgademo.audio_snare_frames[0] ;
 wire \vgademo.audio_snare_frames[1] ;
 wire \vgademo.audio_snare_frames[2] ;
 wire \vgademo.audio_snare_frames[3] ;
 wire \vgademo.audio_songpos[0] ;
 wire \vgademo.audio_songpos[1] ;
 wire \vgademo.audio_songpos[2] ;
 wire \vgademo.audio_songpos[3] ;
 wire \vgademo.audio_songpos[4] ;
 wire \vgademo.audio_songpos[5] ;
 wire \vgademo.audio_songpos[6] ;
 wire \vgademo.audio_songpos[7] ;
 wire \vgademo.b_cos[0] ;
 wire \vgademo.b_cos[10] ;
 wire \vgademo.b_cos[11] ;
 wire \vgademo.b_cos[1] ;
 wire \vgademo.b_cos[2] ;
 wire \vgademo.b_cos[3] ;
 wire \vgademo.b_cos[4] ;
 wire \vgademo.b_cos[5] ;
 wire \vgademo.b_cos[6] ;
 wire \vgademo.b_cos[7] ;
 wire \vgademo.b_cos[8] ;
 wire \vgademo.b_cos[9] ;
 wire \vgademo.b_sin[0] ;
 wire \vgademo.b_sin[10] ;
 wire \vgademo.b_sin[11] ;
 wire \vgademo.b_sin[1] ;
 wire \vgademo.b_sin[2] ;
 wire \vgademo.b_sin[3] ;
 wire \vgademo.b_sin[4] ;
 wire \vgademo.b_sin[5] ;
 wire \vgademo.b_sin[6] ;
 wire \vgademo.b_sin[7] ;
 wire \vgademo.b_sin[8] ;
 wire \vgademo.b_sin[9] ;
 wire \vgademo.bayer_j[0] ;
 wire \vgademo.bayer_j[1] ;
 wire \vgademo.h_count[0] ;
 wire \vgademo.h_count[10] ;
 wire \vgademo.h_count[1] ;
 wire \vgademo.h_count[2] ;
 wire \vgademo.h_count[3] ;
 wire \vgademo.h_count[4] ;
 wire \vgademo.h_count[5] ;
 wire \vgademo.h_count[6] ;
 wire \vgademo.h_count[7] ;
 wire \vgademo.h_count[8] ;
 wire \vgademo.h_count[9] ;
 wire \vgademo.linelfsr[0] ;
 wire \vgademo.linelfsr[10] ;
 wire \vgademo.linelfsr[11] ;
 wire \vgademo.linelfsr[12] ;
 wire \vgademo.linelfsr[1] ;
 wire \vgademo.linelfsr[2] ;
 wire \vgademo.linelfsr[3] ;
 wire \vgademo.linelfsr[4] ;
 wire \vgademo.linelfsr[5] ;
 wire \vgademo.linelfsr[6] ;
 wire \vgademo.linelfsr[7] ;
 wire \vgademo.linelfsr[8] ;
 wire \vgademo.linelfsr[9] ;
 wire \vgademo.plane_du[0] ;
 wire \vgademo.plane_du[10] ;
 wire \vgademo.plane_du[1] ;
 wire \vgademo.plane_du[2] ;
 wire \vgademo.plane_du[3] ;
 wire \vgademo.plane_du[4] ;
 wire \vgademo.plane_du[5] ;
 wire \vgademo.plane_du[6] ;
 wire \vgademo.plane_du[7] ;
 wire \vgademo.plane_du[8] ;
 wire \vgademo.plane_du[9] ;
 wire \vgademo.plane_dx[0] ;
 wire \vgademo.plane_dx[1] ;
 wire \vgademo.plane_dx[2] ;
 wire \vgademo.plane_dx[3] ;
 wire \vgademo.plane_dx_div.d[16] ;
 wire \vgademo.plane_dx_div.d[17] ;
 wire \vgademo.plane_dx_div.d[18] ;
 wire \vgademo.plane_dx_div.d[19] ;
 wire \vgademo.plane_dx_div.d[20] ;
 wire \vgademo.plane_dx_div.d[21] ;
 wire \vgademo.plane_dx_div.d[22] ;
 wire \vgademo.plane_dx_div.d[23] ;
 wire \vgademo.plane_dx_div.d[24] ;
 wire \vgademo.plane_dx_div.i[0] ;
 wire \vgademo.plane_dx_div.i[1] ;
 wire \vgademo.plane_dx_div.i[2] ;
 wire \vgademo.plane_dx_div.i[3] ;
 wire \vgademo.plane_dx_div.q[3] ;
 wire \vgademo.plane_dx_div.q[4] ;
 wire \vgademo.plane_dx_div.q[5] ;
 wire \vgademo.plane_dx_div.q[6] ;
 wire \vgademo.plane_dx_div.q[7] ;
 wire \vgademo.plane_dx_div.q[8] ;
 wire \vgademo.plane_dx_div.q[9] ;
 wire \vgademo.plane_dx_div.r[16] ;
 wire \vgademo.plane_dx_div.r[17] ;
 wire \vgademo.plane_dx_div.r[18] ;
 wire \vgademo.plane_dx_div.r[19] ;
 wire \vgademo.plane_dx_div.r[20] ;
 wire \vgademo.plane_dx_div.r[21] ;
 wire \vgademo.plane_dx_div.r[22] ;
 wire \vgademo.plane_dx_div.r[23] ;
 wire \vgademo.plane_dx_div.r[24] ;
 wire \vgademo.plane_dx_div.r[25] ;
 wire \vgademo.plane_u[0] ;
 wire \vgademo.plane_u[10] ;
 wire \vgademo.plane_u[11] ;
 wire \vgademo.plane_u[12] ;
 wire \vgademo.plane_u[13] ;
 wire \vgademo.plane_u[14] ;
 wire \vgademo.plane_u[15] ;
 wire \vgademo.plane_u[16] ;
 wire \vgademo.plane_u[17] ;
 wire \vgademo.plane_u[18] ;
 wire \vgademo.plane_u[19] ;
 wire \vgademo.plane_u[1] ;
 wire \vgademo.plane_u[20] ;
 wire \vgademo.plane_u[21] ;
 wire \vgademo.plane_u[2] ;
 wire \vgademo.plane_u[3] ;
 wire \vgademo.plane_u[4] ;
 wire \vgademo.plane_u[5] ;
 wire \vgademo.plane_u[6] ;
 wire \vgademo.plane_u[7] ;
 wire \vgademo.plane_u[8] ;
 wire \vgademo.plane_u[9] ;
 wire \vgademo.scanline_audio_sample[0] ;
 wire \vgademo.scanline_audio_sample[1] ;
 wire \vgademo.scanline_audio_sample[2] ;
 wire \vgademo.scanline_audio_sample[3] ;
 wire \vgademo.scanline_audio_sample[4] ;
 wire \vgademo.scanline_audio_sample[5] ;
 wire \vgademo.scanline_audio_sample[6] ;
 wire \vgademo.soundtrack.noise_lfsr[0] ;
 wire \vgademo.soundtrack.noise_lfsr[10] ;
 wire \vgademo.soundtrack.noise_lfsr[11] ;
 wire \vgademo.soundtrack.noise_lfsr[12] ;
 wire \vgademo.soundtrack.noise_lfsr[13] ;
 wire \vgademo.soundtrack.noise_lfsr[14] ;
 wire \vgademo.soundtrack.noise_lfsr[1] ;
 wire \vgademo.soundtrack.noise_lfsr[2] ;
 wire \vgademo.soundtrack.noise_lfsr[3] ;
 wire \vgademo.soundtrack.noise_lfsr[4] ;
 wire \vgademo.soundtrack.noise_lfsr[5] ;
 wire \vgademo.soundtrack.noise_lfsr[6] ;
 wire \vgademo.soundtrack.noise_lfsr[7] ;
 wire \vgademo.soundtrack.noise_lfsr[8] ;
 wire \vgademo.soundtrack.noise_lfsr[9] ;
 wire \vgademo.soundtrack.pulse_osc_p[0] ;
 wire \vgademo.soundtrack.pulse_osc_p[10] ;
 wire \vgademo.soundtrack.pulse_osc_p[11] ;
 wire \vgademo.soundtrack.pulse_osc_p[12] ;
 wire \vgademo.soundtrack.pulse_osc_p[13] ;
 wire \vgademo.soundtrack.pulse_osc_p[1] ;
 wire \vgademo.soundtrack.pulse_osc_p[2] ;
 wire \vgademo.soundtrack.pulse_osc_p[3] ;
 wire \vgademo.soundtrack.pulse_osc_p[4] ;
 wire \vgademo.soundtrack.pulse_osc_p[5] ;
 wire \vgademo.soundtrack.pulse_osc_p[6] ;
 wire \vgademo.soundtrack.pulse_osc_p[7] ;
 wire \vgademo.soundtrack.pulse_osc_p[8] ;
 wire \vgademo.soundtrack.pulse_osc_p[9] ;
 wire \vgademo.soundtrack.pulse_vol[0] ;
 wire \vgademo.soundtrack.pulse_vol[1] ;
 wire \vgademo.soundtrack.pulse_vol[2] ;
 wire \vgademo.soundtrack.pulse_vol[3] ;
 wire \vgademo.soundtrack.sample_div[0] ;
 wire \vgademo.soundtrack.sample_div[1] ;
 wire \vgademo.soundtrack.sample_div[2] ;
 wire \vgademo.soundtrack.sample_div[3] ;
 wire \vgademo.soundtrack.sample_div[4] ;
 wire \vgademo.soundtrack.sample_div[5] ;
 wire \vgademo.soundtrack.sample_div[6] ;
 wire \vgademo.soundtrack.sample_div[7] ;
 wire \vgademo.soundtrack.sample_div[8] ;
 wire \vgademo.soundtrack.sample_div[9] ;
 wire \vgademo.soundtrack.sample_div_[0] ;
 wire \vgademo.soundtrack.sample_div_[1] ;
 wire \vgademo.soundtrack.sample_div_[2] ;
 wire \vgademo.soundtrack.sample_div_[3] ;
 wire \vgademo.soundtrack.sample_div_[4] ;
 wire \vgademo.soundtrack.sample_div_[5] ;
 wire \vgademo.soundtrack.sample_div_[6] ;
 wire \vgademo.soundtrack.sample_div_[7] ;
 wire \vgademo.soundtrack.sample_div_[8] ;
 wire \vgademo.soundtrack.sample_div_[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[9] ;
 wire \vgademo.soundtrack.tick_div[0] ;
 wire \vgademo.soundtrack.tick_div[1] ;
 wire \vgademo.soundtrack.tick_div[2] ;
 wire \vgademo.soundtrack.tick_div[3] ;
 wire \vgademo.soundtrack.tick_div[4] ;
 wire \vgademo.soundtrack.tick_div[5] ;
 wire \vgademo.soundtrack.tick_div[6] ;
 wire \vgademo.soundtrack.tick_div[7] ;
 wire \vgademo.soundtrack.tick_div_[0] ;
 wire \vgademo.soundtrack.tri_osc_i[0] ;
 wire \vgademo.soundtrack.tri_osc_i[1] ;
 wire \vgademo.soundtrack.tri_osc_i[2] ;
 wire \vgademo.soundtrack.tri_osc_i[3] ;
 wire \vgademo.soundtrack.tri_osc_i[4] ;
 wire \vgademo.soundtrack.tri_osc_i[5] ;
 wire \vgademo.soundtrack.tri_osc_i[6] ;
 wire \vgademo.soundtrack.tri_osc_i[7] ;
 wire \vgademo.soundtrack.tri_osc_i[8] ;
 wire \vgademo.soundtrack.tri_osc_p[0] ;
 wire \vgademo.soundtrack.tri_osc_p[10] ;
 wire \vgademo.soundtrack.tri_osc_p[11] ;
 wire \vgademo.soundtrack.tri_osc_p[12] ;
 wire \vgademo.soundtrack.tri_osc_p[13] ;
 wire \vgademo.soundtrack.tri_osc_p[14] ;
 wire \vgademo.soundtrack.tri_osc_p[15] ;
 wire \vgademo.soundtrack.tri_osc_p[1] ;
 wire \vgademo.soundtrack.tri_osc_p[2] ;
 wire \vgademo.soundtrack.tri_osc_p[3] ;
 wire \vgademo.soundtrack.tri_osc_p[4] ;
 wire \vgademo.soundtrack.tri_osc_p[5] ;
 wire \vgademo.soundtrack.tri_osc_p[6] ;
 wire \vgademo.soundtrack.tri_osc_p[7] ;
 wire \vgademo.soundtrack.tri_osc_p[8] ;
 wire \vgademo.soundtrack.tri_osc_p[9] ;
 wire \vgademo.v_count[2] ;
 wire \vgademo.v_count[3] ;
 wire \vgademo.v_count[4] ;
 wire \vgademo.v_count[5] ;
 wire \vgademo.v_count[6] ;
 wire \vgademo.v_count[7] ;
 wire \vgademo.v_count[8] ;
 wire \vgademo.v_count[9] ;
 wire \vgademo.vsync ;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;

 sg13g2_inv_1 _3726_ (.Y(_3079_),
    .A(net211));
 sg13g2_inv_1 _3727_ (.Y(_3080_),
    .A(net213));
 sg13g2_inv_1 _3728_ (.Y(_3081_),
    .A(net172));
 sg13g2_inv_1 _3729_ (.Y(_3082_),
    .A(net355));
 sg13g2_inv_1 _3730_ (.Y(_3083_),
    .A(\vgademo.plane_dx[3] ));
 sg13g2_inv_1 _3731_ (.Y(_3084_),
    .A(\vgademo.plane_dx[2] ));
 sg13g2_inv_1 _3732_ (.Y(_3085_),
    .A(net1040));
 sg13g2_inv_1 _3733_ (.Y(_3086_),
    .A(net564));
 sg13g2_inv_1 _3734_ (.Y(_3087_),
    .A(net373));
 sg13g2_inv_1 _3735_ (.Y(_3088_),
    .A(\vgademo.linelfsr[10] ));
 sg13g2_inv_1 _3736_ (.Y(_3089_),
    .A(\vgademo.linelfsr[2] ));
 sg13g2_inv_1 _3737_ (.Y(_3090_),
    .A(net1062));
 sg13g2_inv_1 _3738_ (.Y(_3091_),
    .A(net433));
 sg13g2_inv_1 _3739_ (.Y(_3092_),
    .A(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_inv_1 _3740_ (.Y(_3093_),
    .A(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_inv_1 _3741_ (.Y(_3094_),
    .A(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_inv_2 _3742_ (.Y(_3095_),
    .A(net1047));
 sg13g2_inv_1 _3743_ (.Y(_3096_),
    .A(net1052));
 sg13g2_inv_2 _3744_ (.Y(_3097_),
    .A(net1057));
 sg13g2_inv_1 _3745_ (.Y(_3098_),
    .A(net1045));
 sg13g2_inv_1 _3746_ (.Y(_3099_),
    .A(net1042));
 sg13g2_inv_2 _3747_ (.Y(_3100_),
    .A(net415));
 sg13g2_inv_1 _3748_ (.Y(_3101_),
    .A(\vgademo.bayer_j[0] ));
 sg13g2_inv_1 _3749_ (.Y(_3102_),
    .A(\vgademo.v_count[3] ));
 sg13g2_inv_1 _3750_ (.Y(_3103_),
    .A(net965));
 sg13g2_inv_1 _3751_ (.Y(_3104_),
    .A(\vgademo.v_count[4] ));
 sg13g2_inv_1 _3752_ (.Y(_3105_),
    .A(\vgademo.v_count[7] ));
 sg13g2_inv_1 _3753_ (.Y(_3106_),
    .A(net1003));
 sg13g2_inv_1 _3754_ (.Y(_3107_),
    .A(net1001));
 sg13g2_inv_1 _3755_ (.Y(_3108_),
    .A(net1002));
 sg13g2_inv_2 _3756_ (.Y(_3109_),
    .A(\vgademo.h_count[5] ));
 sg13g2_inv_2 _3757_ (.Y(_3110_),
    .A(\vgademo.h_count[7] ));
 sg13g2_inv_1 _3758_ (.Y(_3111_),
    .A(\vgademo.h_count[9] ));
 sg13g2_inv_1 _3759_ (.Y(_3112_),
    .A(\vgademo.a_scrolly[13] ));
 sg13g2_inv_2 _3760_ (.Y(_3113_),
    .A(\vgademo.a_scrolly[11] ));
 sg13g2_inv_2 _3761_ (.Y(_3114_),
    .A(net970));
 sg13g2_inv_1 _3762_ (.Y(_3115_),
    .A(_0065_));
 sg13g2_inv_2 _3763_ (.Y(_3116_),
    .A(net976));
 sg13g2_inv_4 _3764_ (.A(net979),
    .Y(_3117_));
 sg13g2_inv_2 _3765_ (.Y(_3118_),
    .A(net981));
 sg13g2_inv_2 _3766_ (.Y(_3119_),
    .A(_0066_));
 sg13g2_inv_1 _3767_ (.Y(_3120_),
    .A(net517));
 sg13g2_inv_1 _3768_ (.Y(_3121_),
    .A(_0072_));
 sg13g2_inv_1 _3769_ (.Y(_3122_),
    .A(\vgademo.plane_dx_div.r[20] ));
 sg13g2_inv_1 _3770_ (.Y(_3123_),
    .A(_0017_));
 sg13g2_inv_1 _3771_ (.Y(_3124_),
    .A(_0019_));
 sg13g2_inv_1 _3772_ (.Y(_3125_),
    .A(_0021_));
 sg13g2_inv_1 _3773_ (.Y(_3126_),
    .A(net336));
 sg13g2_inv_1 _3774_ (.Y(_3127_),
    .A(net274));
 sg13g2_inv_1 _3775_ (.Y(_3128_),
    .A(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_inv_1 _3776_ (.Y(_3129_),
    .A(net598));
 sg13g2_inv_1 _3777_ (.Y(_3130_),
    .A(net594));
 sg13g2_inv_1 _3778_ (.Y(_3131_),
    .A(net587));
 sg13g2_inv_1 _3779_ (.Y(_3132_),
    .A(net1012));
 sg13g2_inv_1 _3780_ (.Y(_3133_),
    .A(net1008));
 sg13g2_inv_4 _3781_ (.A(net1015),
    .Y(_3134_));
 sg13g2_inv_1 _3782_ (.Y(_3135_),
    .A(\vgademo.b_sin[7] ));
 sg13g2_inv_1 _3783_ (.Y(_3136_),
    .A(net436));
 sg13g2_inv_1 _3784_ (.Y(_3137_),
    .A(\vgademo.b_sin[8] ));
 sg13g2_inv_1 _3785_ (.Y(_3138_),
    .A(net505));
 sg13g2_inv_1 _3786_ (.Y(_3139_),
    .A(\vgademo.b_sin[9] ));
 sg13g2_inv_1 _3787_ (.Y(_3140_),
    .A(\vgademo.b_sin[10] ));
 sg13g2_inv_1 _3788_ (.Y(_3141_),
    .A(net525));
 sg13g2_inv_1 _3789_ (.Y(_3142_),
    .A(net952));
 sg13g2_inv_1 _3790_ (.Y(_3143_),
    .A(net567));
 sg13g2_inv_2 _3791_ (.Y(_3144_),
    .A(net450));
 sg13g2_inv_1 _3792_ (.Y(_3145_),
    .A(\vgademo.b_cos[7] ));
 sg13g2_inv_1 _3793_ (.Y(_3146_),
    .A(net488));
 sg13g2_inv_2 _3794_ (.Y(_3147_),
    .A(net957));
 sg13g2_inv_2 _3795_ (.Y(_3148_),
    .A(net956));
 sg13g2_inv_1 _3796_ (.Y(_3149_),
    .A(net479));
 sg13g2_inv_1 _3797_ (.Y(_3150_),
    .A(net382));
 sg13g2_inv_1 _3798_ (.Y(_3151_),
    .A(net349));
 sg13g2_inv_1 _3799_ (.Y(_3152_),
    .A(net509));
 sg13g2_inv_1 _3800_ (.Y(_3153_),
    .A(\vgademo.a_sin[11] ));
 sg13g2_inv_1 _3801_ (.Y(_3154_),
    .A(\vgademo.a_sin[13] ));
 sg13g2_inv_2 _3802_ (.Y(_3155_),
    .A(net960));
 sg13g2_inv_1 _3803_ (.Y(_3156_),
    .A(net376));
 sg13g2_inv_1 _3804_ (.Y(_3157_),
    .A(net381));
 sg13g2_inv_1 _3805_ (.Y(_3158_),
    .A(\vgademo.plane_du[3] ));
 sg13g2_inv_1 _3806_ (.Y(_3159_),
    .A(net290));
 sg13g2_inv_1 _3807_ (.Y(_3160_),
    .A(_0023_));
 sg13g2_inv_1 _3808_ (.Y(_3161_),
    .A(net357));
 sg13g2_inv_1 _3809_ (.Y(_3162_),
    .A(net377));
 sg13g2_inv_1 _3810_ (.Y(_3163_),
    .A(\vgademo.plane_du[7] ));
 sg13g2_inv_1 _3811_ (.Y(_3164_),
    .A(net289));
 sg13g2_inv_1 _3812_ (.Y(_3165_),
    .A(net399));
 sg13g2_inv_1 _3813_ (.Y(_3166_),
    .A(net404));
 sg13g2_inv_1 _3814_ (.Y(_3167_),
    .A(net282));
 sg13g2_inv_1 _3815_ (.Y(_3168_),
    .A(net420));
 sg13g2_inv_1 _3816_ (.Y(_3169_),
    .A(_0028_));
 sg13g2_inv_1 _3817_ (.Y(_3170_),
    .A(net406));
 sg13g2_inv_1 _3818_ (.Y(_3171_),
    .A(net540));
 sg13g2_inv_1 _3819_ (.Y(_3172_),
    .A(net448));
 sg13g2_inv_1 _3820_ (.Y(_3173_),
    .A(net335));
 sg13g2_inv_1 _3821_ (.Y(_3174_),
    .A(net446));
 sg13g2_inv_1 _3822_ (.Y(_3175_),
    .A(_0033_));
 sg13g2_inv_1 _3823_ (.Y(_3176_),
    .A(net256));
 sg13g2_inv_1 _3824_ (.Y(_3177_),
    .A(\vgademo.linelfsr[5] ));
 sg13g2_inv_1 _3825_ (.Y(_3178_),
    .A(\vgademo.soundtrack.pulse_osc_p[13] ));
 sg13g2_inv_1 _3826_ (.Y(_3179_),
    .A(net369));
 sg13g2_inv_1 _3827_ (.Y(_3180_),
    .A(net424));
 sg13g2_inv_1 _3828_ (.Y(_3181_),
    .A(net428));
 sg13g2_inv_1 _3829_ (.Y(_3182_),
    .A(net398));
 sg13g2_inv_1 _3830_ (.Y(_3183_),
    .A(net316));
 sg13g2_inv_1 _3831_ (.Y(_3184_),
    .A(net265));
 sg13g2_inv_1 _3832_ (.Y(_3185_),
    .A(net328));
 sg13g2_inv_1 _3833_ (.Y(_3186_),
    .A(net321));
 sg13g2_inv_1 _3834_ (.Y(_3187_),
    .A(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_inv_1 _3835_ (.Y(_3188_),
    .A(net425));
 sg13g2_inv_1 _3836_ (.Y(_3189_),
    .A(net575));
 sg13g2_inv_1 _3837_ (.Y(_3190_),
    .A(net396));
 sg13g2_inv_1 _3838_ (.Y(_3191_),
    .A(_0048_));
 sg13g2_inv_1 _3839_ (.Y(_3192_),
    .A(_0050_));
 sg13g2_nand2_1 _3840_ (.Y(_3193_),
    .A(\vgademo.h_count[7] ),
    .B(net996));
 sg13g2_nand4_1 _3841_ (.B(net999),
    .C(\vgademo.h_count[7] ),
    .A(\vgademo.h_count[5] ),
    .Y(_3194_),
    .D(net996));
 sg13g2_inv_1 _3842_ (.Y(_3195_),
    .A(_3194_));
 sg13g2_nor4_2 _3843_ (.A(net1003),
    .B(net1005),
    .C(net1001),
    .Y(_3196_),
    .D(_3108_));
 sg13g2_nor2_1 _3844_ (.A(\vgademo.h_count[9] ),
    .B(net995),
    .Y(_3197_));
 sg13g2_and4_2 _3845_ (.A(\vgademo.h_count[8] ),
    .B(_3195_),
    .C(_3196_),
    .D(_3197_),
    .X(_3198_));
 sg13g2_nand4_1 _3846_ (.B(_3195_),
    .C(_3196_),
    .A(\vgademo.h_count[8] ),
    .Y(_3199_),
    .D(_3197_));
 sg13g2_nor2_1 _3847_ (.A(net1005),
    .B(net941),
    .Y(_0000_));
 sg13g2_nand2_2 _3848_ (.Y(_3200_),
    .A(net1004),
    .B(net1005));
 sg13g2_xor2_1 _3849_ (.B(net1005),
    .A(net1003),
    .X(_0002_));
 sg13g2_and2_1 _3850_ (.A(net477),
    .B(_3200_),
    .X(_3201_));
 sg13g2_nor2_1 _3851_ (.A(net477),
    .B(_3200_),
    .Y(_3202_));
 sg13g2_nor3_1 _3852_ (.A(net941),
    .B(net478),
    .C(_3202_),
    .Y(_0003_));
 sg13g2_xor2_1 _3853_ (.B(_3202_),
    .A(net366),
    .X(_3203_));
 sg13g2_nor2_1 _3854_ (.A(net941),
    .B(net367),
    .Y(_0004_));
 sg13g2_nor3_2 _3855_ (.A(_3107_),
    .B(_3108_),
    .C(_3200_),
    .Y(_3204_));
 sg13g2_nand2_1 _3856_ (.Y(_3205_),
    .A(net998),
    .B(_3204_));
 sg13g2_o21ai_1 _3857_ (.B1(net940),
    .Y(_3206_),
    .A1(net998),
    .A2(_3204_));
 sg13g2_nor2b_1 _3858_ (.A(_3206_),
    .B_N(_3205_),
    .Y(_0005_));
 sg13g2_o21ai_1 _3859_ (.B1(net940),
    .Y(_3207_),
    .A1(net293),
    .A2(_3205_));
 sg13g2_a21oi_1 _3860_ (.A1(net293),
    .A2(_3205_),
    .Y(_0006_),
    .B1(_3207_));
 sg13g2_nand3_1 _3861_ (.B(net999),
    .C(_3204_),
    .A(\vgademo.h_count[5] ),
    .Y(_3208_));
 sg13g2_nor2_1 _3862_ (.A(net589),
    .B(_3208_),
    .Y(_3209_));
 sg13g2_a21oi_1 _3863_ (.A1(net589),
    .A2(_3208_),
    .Y(_3210_),
    .B1(net941));
 sg13g2_nor2b_1 _3864_ (.A(net590),
    .B_N(_3210_),
    .Y(_0007_));
 sg13g2_nor3_1 _3865_ (.A(_0036_),
    .B(net555),
    .C(_3208_),
    .Y(_3211_));
 sg13g2_nor2b_1 _3866_ (.A(_3209_),
    .B_N(net555),
    .Y(_3212_));
 sg13g2_nor3_1 _3867_ (.A(net941),
    .B(_3211_),
    .C(net556),
    .Y(_0008_));
 sg13g2_or2_1 _3868_ (.X(_3213_),
    .B(_3208_),
    .A(_3193_));
 sg13g2_nor2_1 _3869_ (.A(net577),
    .B(_3213_),
    .Y(_3214_));
 sg13g2_a21oi_1 _3870_ (.A1(net577),
    .A2(_3213_),
    .Y(_3215_),
    .B1(net941));
 sg13g2_nor2b_1 _3871_ (.A(_3214_),
    .B_N(_3215_),
    .Y(_0009_));
 sg13g2_o21ai_1 _3872_ (.B1(net940),
    .Y(_3216_),
    .A1(_3176_),
    .A2(_3214_));
 sg13g2_a21oi_1 _3873_ (.A1(_3176_),
    .A2(_3214_),
    .Y(_0010_),
    .B1(_3216_));
 sg13g2_nand2_1 _3874_ (.Y(_3217_),
    .A(\vgademo.h_count[9] ),
    .B(\vgademo.h_count[8] ));
 sg13g2_or2_1 _3875_ (.X(_3218_),
    .B(_3217_),
    .A(_3213_));
 sg13g2_a21oi_1 _3876_ (.A1(net995),
    .A2(_3218_),
    .Y(_3219_),
    .B1(net941));
 sg13g2_o21ai_1 _3877_ (.B1(_3219_),
    .Y(_3220_),
    .A1(net995),
    .A2(_3218_));
 sg13g2_inv_1 _3878_ (.Y(_0001_),
    .A(_3220_));
 sg13g2_nand2_2 _3879_ (.Y(_3221_),
    .A(\vgademo.v_count[7] ),
    .B(\vgademo.v_count[6] ));
 sg13g2_nor2_1 _3880_ (.A(\vgademo.v_count[8] ),
    .B(\vgademo.v_count[9] ),
    .Y(_3222_));
 sg13g2_nor3_1 _3881_ (.A(_0063_),
    .B(_3221_),
    .C(_3222_),
    .Y(_3223_));
 sg13g2_nand2b_1 _3882_ (.Y(_3224_),
    .B(\vgademo.v_count[8] ),
    .A_N(\vgademo.v_count[9] ));
 sg13g2_nor4_2 _3883_ (.A(_3103_),
    .B(net562),
    .C(_3221_),
    .Y(_3225_),
    .D(_3224_));
 sg13g2_o21ai_1 _3884_ (.B1(_3225_),
    .Y(_3226_),
    .A1(_3101_),
    .A2(_3223_));
 sg13g2_or4_1 _3885_ (.A(_3100_),
    .B(_3102_),
    .C(net968),
    .D(_3226_),
    .X(_0012_));
 sg13g2_nor2_2 _3886_ (.A(\vgademo.h_count[9] ),
    .B(\vgademo.h_count[8] ),
    .Y(_3227_));
 sg13g2_nand2_1 _3887_ (.Y(_3228_),
    .A(_3194_),
    .B(_3227_));
 sg13g2_nand3_1 _3888_ (.B(_3108_),
    .C(_3200_),
    .A(_3107_),
    .Y(_3229_));
 sg13g2_nor3_1 _3889_ (.A(_3109_),
    .B(net999),
    .C(_3193_),
    .Y(_3230_));
 sg13g2_a22oi_1 _3890_ (.Y(_3231_),
    .B1(_3229_),
    .B2(_3230_),
    .A2(_3228_),
    .A1(\vgademo.h_count[10] ));
 sg13g2_nor2_1 _3891_ (.A(net1004),
    .B(net1002),
    .Y(_3232_));
 sg13g2_nand2_1 _3892_ (.Y(_3233_),
    .A(net1001),
    .B(net999));
 sg13g2_nor2_1 _3893_ (.A(net997),
    .B(net996),
    .Y(_3234_));
 sg13g2_o21ai_1 _3894_ (.B1(_3234_),
    .Y(_3235_),
    .A1(_3232_),
    .A2(_3233_));
 sg13g2_nand3_1 _3895_ (.B(\vgademo.h_count[8] ),
    .C(_3235_),
    .A(\vgademo.h_count[7] ),
    .Y(_3236_));
 sg13g2_nor2b_1 _3896_ (.A(\vgademo.h_count[9] ),
    .B_N(\vgademo.h_count[10] ),
    .Y(_3237_));
 sg13g2_nor3_2 _3897_ (.A(\vgademo.h_count[9] ),
    .B(\vgademo.h_count[8] ),
    .C(_0061_),
    .Y(_3238_));
 sg13g2_nor3_1 _3898_ (.A(net1001),
    .B(net1002),
    .C(\vgademo.h_count[10] ),
    .Y(_3239_));
 sg13g2_a22oi_1 _3899_ (.Y(_3240_),
    .B1(_3238_),
    .B2(_3239_),
    .A2(_3237_),
    .A1(_3236_));
 sg13g2_or2_2 _3900_ (.X(_0011_),
    .B(_3240_),
    .A(_3231_));
 sg13g2_nand2b_1 _3901_ (.Y(_3241_),
    .B(net1010),
    .A_N(net1011));
 sg13g2_nor2_1 _3902_ (.A(_3099_),
    .B(net1041),
    .Y(_3242_));
 sg13g2_nand2b_1 _3903_ (.Y(_3243_),
    .B(net1042),
    .A_N(net1041));
 sg13g2_nor2_2 _3904_ (.A(net1049),
    .B(net1045),
    .Y(_3244_));
 sg13g2_nand2_2 _3905_ (.Y(_3245_),
    .A(_3095_),
    .B(net946));
 sg13g2_o21ai_1 _3906_ (.B1(net1053),
    .Y(_3246_),
    .A1(net1059),
    .A2(net1055));
 sg13g2_nand2_1 _3907_ (.Y(_3247_),
    .A(_3244_),
    .B(_3246_));
 sg13g2_nand2b_1 _3908_ (.Y(_3248_),
    .B(net1048),
    .A_N(net1044));
 sg13g2_nor2b_1 _3909_ (.A(net1059),
    .B_N(net1053),
    .Y(_3249_));
 sg13g2_nand2b_2 _3910_ (.Y(_3250_),
    .B(net1052),
    .A_N(net1058));
 sg13g2_nor2b_1 _3911_ (.A(net1055),
    .B_N(net1063),
    .Y(_3251_));
 sg13g2_a21oi_1 _3912_ (.A1(_3249_),
    .A2(_3251_),
    .Y(_3252_),
    .B1(_3248_));
 sg13g2_nor2_1 _3913_ (.A(net1063),
    .B(net1059),
    .Y(_3253_));
 sg13g2_or2_1 _3914_ (.X(_3254_),
    .B(net1059),
    .A(net1063));
 sg13g2_nor2_2 _3915_ (.A(net1053),
    .B(net1055),
    .Y(_3255_));
 sg13g2_or2_2 _3916_ (.X(_3256_),
    .B(net1057),
    .A(net1054));
 sg13g2_nor2_1 _3917_ (.A(net1049),
    .B(_3255_),
    .Y(_3257_));
 sg13g2_o21ai_1 _3918_ (.B1(_3254_),
    .Y(_3258_),
    .A1(net1047),
    .A2(_3255_));
 sg13g2_o21ai_1 _3919_ (.B1(_3247_),
    .Y(_3259_),
    .A1(_3252_),
    .A2(_3258_));
 sg13g2_and2_1 _3920_ (.A(_3242_),
    .B(_3259_),
    .X(_3260_));
 sg13g2_and2_1 _3921_ (.A(net1058),
    .B(net1056),
    .X(_3261_));
 sg13g2_nand2_2 _3922_ (.Y(_3262_),
    .A(net1060),
    .B(net1056));
 sg13g2_nand2_1 _3923_ (.Y(_3263_),
    .A(net949),
    .B(net1058));
 sg13g2_nor2_1 _3924_ (.A(net949),
    .B(_3096_),
    .Y(_3264_));
 sg13g2_nand2_1 _3925_ (.Y(_3265_),
    .A(net1051),
    .B(_3262_));
 sg13g2_o21ai_1 _3926_ (.B1(net1053),
    .Y(_3266_),
    .A1(net1062),
    .A2(_3262_));
 sg13g2_and2_2 _3927_ (.A(net1063),
    .B(net1059),
    .X(_3267_));
 sg13g2_xor2_1 _3928_ (.B(net1061),
    .A(net1062),
    .X(_3268_));
 sg13g2_xnor2_1 _3929_ (.Y(_3269_),
    .A(net1062),
    .B(net1060));
 sg13g2_nor2_1 _3930_ (.A(net949),
    .B(net1058),
    .Y(_3270_));
 sg13g2_nor2_1 _3931_ (.A(net1056),
    .B(_3268_),
    .Y(_3271_));
 sg13g2_a221oi_1 _3932_ (.B2(_3097_),
    .C1(_3096_),
    .B1(_3269_),
    .A1(net949),
    .Y(_3272_),
    .A2(_3261_));
 sg13g2_nor2_1 _3933_ (.A(_3256_),
    .B(_3268_),
    .Y(_3273_));
 sg13g2_nand2_1 _3934_ (.Y(_3274_),
    .A(net1056),
    .B(_3269_));
 sg13g2_o21ai_1 _3935_ (.B1(net948),
    .Y(_3275_),
    .A1(_3097_),
    .A2(_3268_));
 sg13g2_a221oi_1 _3936_ (.B2(_3275_),
    .C1(net1048),
    .B1(_3266_),
    .A1(_3097_),
    .Y(_3276_),
    .A2(_3263_));
 sg13g2_o21ai_1 _3937_ (.B1(net1050),
    .Y(_3277_),
    .A1(_3272_),
    .A2(_3273_));
 sg13g2_nand3b_1 _3938_ (.B(_3277_),
    .C(net1044),
    .Y(_3278_),
    .A_N(_3276_));
 sg13g2_nor2b_2 _3939_ (.A(net1056),
    .B_N(net1058),
    .Y(_3279_));
 sg13g2_nand2_2 _3940_ (.Y(_3280_),
    .A(net1058),
    .B(_3097_));
 sg13g2_a21o_1 _3941_ (.A2(_3279_),
    .A1(net1051),
    .B1(net949),
    .X(_3281_));
 sg13g2_nor2_1 _3942_ (.A(net1063),
    .B(net1055),
    .Y(_3282_));
 sg13g2_nand2b_2 _3943_ (.Y(_3283_),
    .B(net1059),
    .A_N(net1053));
 sg13g2_a21oi_1 _3944_ (.A1(net1053),
    .A2(_3282_),
    .Y(_3284_),
    .B1(_3253_));
 sg13g2_a21oi_1 _3945_ (.A1(_3281_),
    .A2(_3284_),
    .Y(_3285_),
    .B1(_3248_));
 sg13g2_mux2_1 _3946_ (.A0(net1055),
    .A1(net1059),
    .S(net1063),
    .X(_3286_));
 sg13g2_a21oi_1 _3947_ (.A1(_3283_),
    .A2(_3286_),
    .Y(_3287_),
    .B1(_3255_));
 sg13g2_and2_2 _3948_ (.A(net1042),
    .B(net1041),
    .X(_3288_));
 sg13g2_o21ai_1 _3949_ (.B1(_3288_),
    .Y(_3289_),
    .A1(_3245_),
    .A2(_3287_));
 sg13g2_nor2_1 _3950_ (.A(_3285_),
    .B(_3289_),
    .Y(_3290_));
 sg13g2_a21o_1 _3951_ (.A2(_3290_),
    .A1(_3278_),
    .B1(_3260_),
    .X(_3291_));
 sg13g2_a221oi_1 _3952_ (.B2(_3290_),
    .C1(_3178_),
    .B1(_3278_),
    .A1(_3242_),
    .Y(_3292_),
    .A2(_3259_));
 sg13g2_a21o_2 _3953_ (.A2(_3291_),
    .A1(\vgademo.soundtrack.pulse_osc_p[12] ),
    .B1(_3292_),
    .X(_3293_));
 sg13g2_a21oi_2 _3954_ (.B1(_3292_),
    .Y(_3294_),
    .A2(_3291_),
    .A1(\vgademo.soundtrack.pulse_osc_p[12] ));
 sg13g2_nor2_1 _3955_ (.A(_3132_),
    .B(_3293_),
    .Y(_3295_));
 sg13g2_nand2_1 _3956_ (.Y(_3296_),
    .A(net1012),
    .B(_3294_));
 sg13g2_a21oi_2 _3957_ (.B1(_3241_),
    .Y(_3297_),
    .A2(_3294_),
    .A1(net1012));
 sg13g2_mux2_1 _3958_ (.A0(\vgademo.soundtrack.noise_lfsr[10] ),
    .A1(\vgademo.soundtrack.noise_lfsr[11] ),
    .S(net1025),
    .X(_3298_));
 sg13g2_nand2_1 _3959_ (.Y(_3299_),
    .A(net1021),
    .B(_3298_));
 sg13g2_nand2b_1 _3960_ (.Y(_3300_),
    .B(net1027),
    .A_N(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_o21ai_1 _3961_ (.B1(_3300_),
    .Y(_3301_),
    .A1(\vgademo.soundtrack.noise_lfsr[8] ),
    .A2(net1026));
 sg13g2_o21ai_1 _3962_ (.B1(_3299_),
    .Y(_3302_),
    .A1(net1021),
    .A2(_3301_));
 sg13g2_nand2b_1 _3963_ (.Y(_3303_),
    .B(\vgademo.soundtrack.noise_lfsr[12] ),
    .A_N(net1025));
 sg13g2_nor2_1 _3964_ (.A(net1024),
    .B(_3303_),
    .Y(_3304_));
 sg13g2_mux2_2 _3965_ (.A0(_3302_),
    .A1(_3304_),
    .S(net1018),
    .X(_3305_));
 sg13g2_nor2_1 _3966_ (.A(net1026),
    .B(_0040_),
    .Y(_3306_));
 sg13g2_a21oi_1 _3967_ (.A1(net1026),
    .A2(\vgademo.soundtrack.noise_lfsr[5] ),
    .Y(_3307_),
    .B1(_3306_));
 sg13g2_nor2_1 _3968_ (.A(net1020),
    .B(_3307_),
    .Y(_3308_));
 sg13g2_mux2_1 _3969_ (.A0(\vgademo.soundtrack.noise_lfsr[6] ),
    .A1(\vgademo.soundtrack.noise_lfsr[7] ),
    .S(net1027),
    .X(_3309_));
 sg13g2_a21oi_1 _3970_ (.A1(net1021),
    .A2(_3309_),
    .Y(_3310_),
    .B1(_3308_));
 sg13g2_mux2_1 _3971_ (.A0(\vgademo.soundtrack.noise_lfsr[2] ),
    .A1(\vgademo.soundtrack.noise_lfsr[3] ),
    .S(net1025),
    .X(_3311_));
 sg13g2_nand2_1 _3972_ (.Y(_3312_),
    .A(net1020),
    .B(_3311_));
 sg13g2_nand2b_1 _3973_ (.Y(_3313_),
    .B(net1026),
    .A_N(\vgademo.soundtrack.noise_lfsr[1] ));
 sg13g2_o21ai_1 _3974_ (.B1(_3313_),
    .Y(_3314_),
    .A1(net1026),
    .A2(\vgademo.soundtrack.noise_lfsr[0] ));
 sg13g2_o21ai_1 _3975_ (.B1(_3312_),
    .Y(_3315_),
    .A1(net1020),
    .A2(_3314_));
 sg13g2_nand2_1 _3976_ (.Y(_3316_),
    .A(net1013),
    .B(_3305_));
 sg13g2_a21oi_1 _3977_ (.A1(net1017),
    .A2(_3310_),
    .Y(_3317_),
    .B1(net1014));
 sg13g2_o21ai_1 _3978_ (.B1(_3317_),
    .Y(_3318_),
    .A1(net1016),
    .A2(_3315_));
 sg13g2_nand2_1 _3979_ (.Y(_3319_),
    .A(_3316_),
    .B(_3318_));
 sg13g2_nand3_1 _3980_ (.B(_3297_),
    .C(_3319_),
    .A(net1008),
    .Y(_3320_));
 sg13g2_a21oi_1 _3981_ (.A1(net1008),
    .A2(_3297_),
    .Y(_3321_),
    .B1(_3319_));
 sg13g2_a21o_1 _3982_ (.A2(_3297_),
    .A1(net1008),
    .B1(_3319_),
    .X(_3322_));
 sg13g2_and2_1 _3983_ (.A(_3320_),
    .B(_3322_),
    .X(_3323_));
 sg13g2_xnor2_1 _3984_ (.Y(_3324_),
    .A(net1007),
    .B(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_xnor2_1 _3985_ (.Y(_3325_),
    .A(_3323_),
    .B(_3324_));
 sg13g2_nand2_1 _3986_ (.Y(_3326_),
    .A(net228),
    .B(_3325_));
 sg13g2_xor2_1 _3987_ (.B(_3325_),
    .A(net228),
    .X(\vgademo.soundtrack.sigma_delta_accum_[0] ));
 sg13g2_o21ai_1 _3988_ (.B1(_3320_),
    .Y(_3327_),
    .A1(_3321_),
    .A2(_3324_));
 sg13g2_and2_1 _3989_ (.A(net1011),
    .B(net1010),
    .X(_3328_));
 sg13g2_nand2_1 _3990_ (.Y(_3329_),
    .A(net1011),
    .B(net1010));
 sg13g2_nor2_1 _3991_ (.A(_3133_),
    .B(_3329_),
    .Y(_3330_));
 sg13g2_xnor2_1 _3992_ (.Y(_3331_),
    .A(net1009),
    .B(_3328_));
 sg13g2_nor2_1 _3993_ (.A(net1011),
    .B(net1010),
    .Y(_3332_));
 sg13g2_or2_2 _3994_ (.X(_3333_),
    .B(_3332_),
    .A(_3328_));
 sg13g2_inv_1 _3995_ (.Y(_3334_),
    .A(_3333_));
 sg13g2_and2_1 _3996_ (.A(net1011),
    .B(net1012),
    .X(_3335_));
 sg13g2_nor2_1 _3997_ (.A(net1011),
    .B(net1012),
    .Y(_3336_));
 sg13g2_nor2_1 _3998_ (.A(_3335_),
    .B(_3336_),
    .Y(_3337_));
 sg13g2_a221oi_1 _3999_ (.B2(_3291_),
    .C1(_3292_),
    .B1(\vgademo.soundtrack.pulse_osc_p[12] ),
    .A1(\vgademo.soundtrack.pulse_vol[1] ),
    .Y(_3338_),
    .A2(\vgademo.soundtrack.pulse_vol[0] ));
 sg13g2_or2_2 _4000_ (.X(_3339_),
    .B(_3338_),
    .A(_3337_));
 sg13g2_nor4_2 _4001_ (.A(_3331_),
    .B(_3333_),
    .C(_3337_),
    .Y(_3340_),
    .D(_3338_));
 sg13g2_nor2b_1 _4002_ (.A(net1027),
    .B_N(\vgademo.soundtrack.noise_lfsr[5] ),
    .Y(_3341_));
 sg13g2_a21oi_1 _4003_ (.A1(\vgademo.soundtrack.noise_lfsr[6] ),
    .A2(net1027),
    .Y(_3342_),
    .B1(_3341_));
 sg13g2_mux2_1 _4004_ (.A0(\vgademo.soundtrack.noise_lfsr[7] ),
    .A1(\vgademo.soundtrack.noise_lfsr[8] ),
    .S(net1027),
    .X(_3343_));
 sg13g2_nand2_1 _4005_ (.Y(_3344_),
    .A(net1022),
    .B(_3343_));
 sg13g2_o21ai_1 _4006_ (.B1(_3344_),
    .Y(_3345_),
    .A1(net1022),
    .A2(_3342_));
 sg13g2_nor2_1 _4007_ (.A(\vgademo.soundtrack.noise_lfsr[3] ),
    .B(net1025),
    .Y(_3346_));
 sg13g2_a21oi_1 _4008_ (.A1(net1025),
    .A2(_0040_),
    .Y(_3347_),
    .B1(_3346_));
 sg13g2_nand2b_1 _4009_ (.Y(_3348_),
    .B(net1025),
    .A_N(\vgademo.soundtrack.noise_lfsr[2] ));
 sg13g2_o21ai_1 _4010_ (.B1(_3348_),
    .Y(_3349_),
    .A1(\vgademo.soundtrack.noise_lfsr[1] ),
    .A2(net1025));
 sg13g2_nor2b_1 _4011_ (.A(net1026),
    .B_N(\vgademo.soundtrack.noise_lfsr[9] ),
    .Y(_3350_));
 sg13g2_a21oi_1 _4012_ (.A1(net1026),
    .A2(\vgademo.soundtrack.noise_lfsr[10] ),
    .Y(_3351_),
    .B1(_3350_));
 sg13g2_mux2_1 _4013_ (.A0(\vgademo.soundtrack.noise_lfsr[11] ),
    .A1(\vgademo.soundtrack.noise_lfsr[12] ),
    .S(net1025),
    .X(_3352_));
 sg13g2_nand2_1 _4014_ (.Y(_3353_),
    .A(net1020),
    .B(_3352_));
 sg13g2_o21ai_1 _4015_ (.B1(_3353_),
    .Y(_3354_),
    .A1(net1021),
    .A2(_3351_));
 sg13g2_nor2b_2 _4016_ (.A(net1016),
    .B_N(_3354_),
    .Y(_3355_));
 sg13g2_a21oi_1 _4017_ (.A1(net1020),
    .A2(_3347_),
    .Y(_3356_),
    .B1(net1016));
 sg13g2_o21ai_1 _4018_ (.B1(_3356_),
    .Y(_3357_),
    .A1(net1021),
    .A2(_3349_));
 sg13g2_nor2b_1 _4019_ (.A(_3345_),
    .B_N(net1017),
    .Y(_3358_));
 sg13g2_nor2_1 _4020_ (.A(net1014),
    .B(_3358_),
    .Y(_3359_));
 sg13g2_a22oi_1 _4021_ (.Y(_3360_),
    .B1(_3357_),
    .B2(_3359_),
    .A2(_3355_),
    .A1(net1014));
 sg13g2_or4_1 _4022_ (.A(_3331_),
    .B(_3333_),
    .C(_3339_),
    .D(_3360_),
    .X(_3361_));
 sg13g2_xor2_1 _4023_ (.B(_3360_),
    .A(_3340_),
    .X(_3362_));
 sg13g2_xnor2_1 _4024_ (.Y(_3363_),
    .A(net1007),
    .B(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_xnor2_1 _4025_ (.Y(_3364_),
    .A(_3362_),
    .B(_3363_));
 sg13g2_nor2b_1 _4026_ (.A(_3364_),
    .B_N(_3327_),
    .Y(_3365_));
 sg13g2_xor2_1 _4027_ (.B(_3364_),
    .A(_3327_),
    .X(_3366_));
 sg13g2_or2_1 _4028_ (.X(_3367_),
    .B(_3366_),
    .A(_3182_));
 sg13g2_xnor2_1 _4029_ (.Y(_3368_),
    .A(_3182_),
    .B(_3366_));
 sg13g2_xor2_1 _4030_ (.B(_3368_),
    .A(_3326_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[1] ));
 sg13g2_o21ai_1 _4031_ (.B1(_3367_),
    .Y(_3369_),
    .A1(_3326_),
    .A2(_3368_));
 sg13g2_o21ai_1 _4032_ (.B1(_3361_),
    .Y(_3370_),
    .A1(_3362_),
    .A2(_3363_));
 sg13g2_nor2b_1 _4033_ (.A(net1010),
    .B_N(net1011),
    .Y(_3371_));
 sg13g2_o21ai_1 _4034_ (.B1(_3371_),
    .Y(_3372_),
    .A1(_3132_),
    .A2(_3293_));
 sg13g2_nor2_1 _4035_ (.A(net1022),
    .B(_3309_),
    .Y(_3373_));
 sg13g2_a21oi_1 _4036_ (.A1(net1022),
    .A2(_3301_),
    .Y(_3374_),
    .B1(_3373_));
 sg13g2_or2_1 _4037_ (.X(_3375_),
    .B(_3311_),
    .A(net1020));
 sg13g2_a21oi_1 _4038_ (.A1(net1020),
    .A2(_3307_),
    .Y(_3376_),
    .B1(net1016));
 sg13g2_a221oi_1 _4039_ (.B2(_3376_),
    .C1(net1013),
    .B1(_3375_),
    .A1(net1016),
    .Y(_3377_),
    .A2(_3374_));
 sg13g2_nor2_1 _4040_ (.A(net1023),
    .B(_3298_),
    .Y(_3378_));
 sg13g2_a21oi_2 _4041_ (.B1(_3378_),
    .Y(_3379_),
    .A2(_3303_),
    .A1(net1023));
 sg13g2_inv_1 _4042_ (.Y(_3380_),
    .A(_3379_));
 sg13g2_nand2b_2 _4043_ (.Y(_3381_),
    .B(_3379_),
    .A_N(net1017));
 sg13g2_a21oi_2 _4044_ (.B1(_3377_),
    .Y(_3382_),
    .A2(_3381_),
    .A1(net1013));
 sg13g2_inv_1 _4045_ (.Y(_3383_),
    .A(_3382_));
 sg13g2_nand4_1 _4046_ (.B(_3296_),
    .C(_3371_),
    .A(net1008),
    .Y(_3384_),
    .D(_3382_));
 sg13g2_o21ai_1 _4047_ (.B1(_3383_),
    .Y(_0365_),
    .A1(_3133_),
    .A2(_3372_));
 sg13g2_xor2_1 _4048_ (.B(\vgademo.soundtrack.tri_osc_p[3] ),
    .A(net1007),
    .X(_0366_));
 sg13g2_nand3_1 _4049_ (.B(_0365_),
    .C(_0366_),
    .A(_3384_),
    .Y(_0367_));
 sg13g2_a21o_1 _4050_ (.A2(_0365_),
    .A1(_3384_),
    .B1(_0366_),
    .X(_0368_));
 sg13g2_and3_1 _4051_ (.X(_0369_),
    .A(_3370_),
    .B(_0367_),
    .C(_0368_));
 sg13g2_nand3_1 _4052_ (.B(_0367_),
    .C(_0368_),
    .A(_3370_),
    .Y(_0370_));
 sg13g2_a21o_1 _4053_ (.A2(_0368_),
    .A1(_0367_),
    .B1(_3370_),
    .X(_0371_));
 sg13g2_and3_1 _4054_ (.X(_0372_),
    .A(_3365_),
    .B(_0370_),
    .C(_0371_));
 sg13g2_a21oi_1 _4055_ (.A1(_0370_),
    .A2(_0371_),
    .Y(_0373_),
    .B1(_3365_));
 sg13g2_nor3_1 _4056_ (.A(_3183_),
    .B(_0372_),
    .C(_0373_),
    .Y(_0374_));
 sg13g2_o21ai_1 _4057_ (.B1(_3183_),
    .Y(_0375_),
    .A1(_0372_),
    .A2(_0373_));
 sg13g2_nand2b_1 _4058_ (.Y(_0376_),
    .B(_0375_),
    .A_N(_0374_));
 sg13g2_xnor2_1 _4059_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .A(_3369_),
    .B(_0376_));
 sg13g2_a21oi_1 _4060_ (.A1(_3369_),
    .A2(_0375_),
    .Y(_0377_),
    .B1(_0374_));
 sg13g2_a21oi_1 _4061_ (.A1(_3365_),
    .A2(_0371_),
    .Y(_0378_),
    .B1(_0369_));
 sg13g2_nand2_1 _4062_ (.Y(_0379_),
    .A(_3384_),
    .B(_0367_));
 sg13g2_nor3_1 _4063_ (.A(net1010),
    .B(_3335_),
    .C(_3336_),
    .Y(_0380_));
 sg13g2_o21ai_1 _4064_ (.B1(_0380_),
    .Y(_0381_),
    .A1(net1012),
    .A2(_3293_));
 sg13g2_nor2_1 _4065_ (.A(_3331_),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_nor2_1 _4066_ (.A(net1020),
    .B(_3343_),
    .Y(_0383_));
 sg13g2_a21oi_1 _4067_ (.A1(net1021),
    .A2(_3351_),
    .Y(_0384_),
    .B1(_0383_));
 sg13g2_nand2b_1 _4068_ (.Y(_0385_),
    .B(_3352_),
    .A_N(net1023));
 sg13g2_or2_2 _4069_ (.X(_0386_),
    .B(_0385_),
    .A(net1017));
 sg13g2_or2_1 _4070_ (.X(_0387_),
    .B(_3347_),
    .A(net1021));
 sg13g2_a21oi_1 _4071_ (.A1(net1022),
    .A2(_3342_),
    .Y(_0388_),
    .B1(net1016));
 sg13g2_a221oi_1 _4072_ (.B2(_0388_),
    .C1(net1013),
    .B1(_0387_),
    .A1(net1016),
    .Y(_0389_),
    .A2(_0384_));
 sg13g2_a21oi_2 _4073_ (.B1(_0389_),
    .Y(_0390_),
    .A2(_0386_),
    .A1(net1013));
 sg13g2_and2_1 _4074_ (.A(_0382_),
    .B(_0390_),
    .X(_0391_));
 sg13g2_xor2_1 _4075_ (.B(_0390_),
    .A(_0382_),
    .X(_0392_));
 sg13g2_xor2_1 _4076_ (.B(\vgademo.soundtrack.tri_osc_p[4] ),
    .A(net1007),
    .X(_0393_));
 sg13g2_xor2_1 _4077_ (.B(_0393_),
    .A(_0392_),
    .X(_0394_));
 sg13g2_nand2_1 _4078_ (.Y(_0395_),
    .A(_0379_),
    .B(_0394_));
 sg13g2_xnor2_1 _4079_ (.Y(_0396_),
    .A(_0379_),
    .B(_0394_));
 sg13g2_xor2_1 _4080_ (.B(_0396_),
    .A(_0378_),
    .X(_0397_));
 sg13g2_xnor2_1 _4081_ (.Y(_0398_),
    .A(\vgademo.soundtrack.sigma_delta_accum[3] ),
    .B(_0397_));
 sg13g2_nor2_1 _4082_ (.A(_0377_),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_xor2_1 _4083_ (.B(_0398_),
    .A(_0377_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[3] ));
 sg13g2_a21oi_1 _4084_ (.A1(\vgademo.soundtrack.sigma_delta_accum[3] ),
    .A2(_0397_),
    .Y(_0400_),
    .B1(_0399_));
 sg13g2_o21ai_1 _4085_ (.B1(_0395_),
    .Y(_0401_),
    .A1(_0378_),
    .A2(_0396_));
 sg13g2_a21oi_1 _4086_ (.A1(_0392_),
    .A2(_0393_),
    .Y(_0402_),
    .B1(_0391_));
 sg13g2_nand3_1 _4087_ (.B(_3296_),
    .C(_3332_),
    .A(net1008),
    .Y(_0403_));
 sg13g2_or2_1 _4088_ (.X(_0404_),
    .B(_3310_),
    .A(net1018));
 sg13g2_a21oi_1 _4089_ (.A1(net1018),
    .A2(_3302_),
    .Y(_0405_),
    .B1(net1013));
 sg13g2_nand2b_2 _4090_ (.Y(_0406_),
    .B(_3304_),
    .A_N(net1018));
 sg13g2_a22oi_1 _4091_ (.Y(_0407_),
    .B1(_0406_),
    .B2(net1013),
    .A2(_0405_),
    .A1(_0404_));
 sg13g2_nand2b_1 _4092_ (.Y(_0408_),
    .B(_0407_),
    .A_N(_0403_));
 sg13g2_xnor2_1 _4093_ (.Y(_0409_),
    .A(_0403_),
    .B(_0407_));
 sg13g2_inv_1 _4094_ (.Y(_0410_),
    .A(_0409_));
 sg13g2_xnor2_1 _4095_ (.Y(_0411_),
    .A(net1007),
    .B(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_xnor2_1 _4096_ (.Y(_0412_),
    .A(_0409_),
    .B(_0411_));
 sg13g2_nand2b_1 _4097_ (.Y(_0413_),
    .B(_0412_),
    .A_N(_0402_));
 sg13g2_xnor2_1 _4098_ (.Y(_0414_),
    .A(_0402_),
    .B(_0412_));
 sg13g2_nand2_1 _4099_ (.Y(_0415_),
    .A(_0401_),
    .B(_0414_));
 sg13g2_xor2_1 _4100_ (.B(_0414_),
    .A(_0401_),
    .X(_0416_));
 sg13g2_nand2_1 _4101_ (.Y(_0417_),
    .A(net550),
    .B(_0416_));
 sg13g2_xnor2_1 _4102_ (.Y(_0418_),
    .A(net550),
    .B(_0416_));
 sg13g2_xor2_1 _4103_ (.B(_0418_),
    .A(_0400_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[4] ));
 sg13g2_o21ai_1 _4104_ (.B1(_0417_),
    .Y(_0419_),
    .A1(_0400_),
    .A2(_0418_));
 sg13g2_and2_1 _4105_ (.A(_0413_),
    .B(_0415_),
    .X(_0420_));
 sg13g2_o21ai_1 _4106_ (.B1(_0408_),
    .Y(_0421_),
    .A1(_0410_),
    .A2(_0411_));
 sg13g2_nor3_1 _4107_ (.A(_3331_),
    .B(_3334_),
    .C(_3339_),
    .Y(_0422_));
 sg13g2_inv_1 _4108_ (.Y(_0423_),
    .A(_0422_));
 sg13g2_mux2_1 _4109_ (.A0(_3345_),
    .A1(_3354_),
    .S(net1016),
    .X(_0424_));
 sg13g2_nand2_1 _4110_ (.Y(_0425_),
    .A(_3134_),
    .B(_0424_));
 sg13g2_xor2_1 _4111_ (.B(_0425_),
    .A(_0422_),
    .X(_0426_));
 sg13g2_xor2_1 _4112_ (.B(\vgademo.soundtrack.tri_osc_p[6] ),
    .A(net1007),
    .X(_0427_));
 sg13g2_nand2b_1 _4113_ (.Y(_0428_),
    .B(_0427_),
    .A_N(_0426_));
 sg13g2_xnor2_1 _4114_ (.Y(_0429_),
    .A(_0426_),
    .B(_0427_));
 sg13g2_nand2_1 _4115_ (.Y(_0430_),
    .A(_0421_),
    .B(_0429_));
 sg13g2_xnor2_1 _4116_ (.Y(_0431_),
    .A(_0421_),
    .B(_0429_));
 sg13g2_xor2_1 _4117_ (.B(_0431_),
    .A(_0420_),
    .X(_0432_));
 sg13g2_and2_1 _4118_ (.A(\vgademo.soundtrack.sigma_delta_accum[5] ),
    .B(_0432_),
    .X(_0433_));
 sg13g2_xor2_1 _4119_ (.B(_0432_),
    .A(net566),
    .X(_0434_));
 sg13g2_xor2_1 _4120_ (.B(_0434_),
    .A(_0419_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[5] ));
 sg13g2_a21oi_1 _4121_ (.A1(_0419_),
    .A2(_0434_),
    .Y(_0435_),
    .B1(_0433_));
 sg13g2_o21ai_1 _4122_ (.B1(_0430_),
    .Y(_0436_),
    .A1(_0420_),
    .A2(_0431_));
 sg13g2_o21ai_1 _4123_ (.B1(_0428_),
    .Y(_0437_),
    .A1(_0423_),
    .A2(_0425_));
 sg13g2_nor3_1 _4124_ (.A(net1009),
    .B(_3295_),
    .C(_3329_),
    .Y(_0438_));
 sg13g2_a21oi_1 _4125_ (.A1(net1017),
    .A2(_3380_),
    .Y(_0439_),
    .B1(net1013));
 sg13g2_o21ai_1 _4126_ (.B1(_0439_),
    .Y(_0440_),
    .A1(net1017),
    .A2(_3374_));
 sg13g2_or4_1 _4127_ (.A(net1008),
    .B(_3295_),
    .C(_3329_),
    .D(_0440_),
    .X(_0441_));
 sg13g2_xor2_1 _4128_ (.B(_0440_),
    .A(_0438_),
    .X(_0442_));
 sg13g2_xnor2_1 _4129_ (.Y(_0443_),
    .A(net1007),
    .B(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_xnor2_1 _4130_ (.Y(_0444_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_nor2b_1 _4131_ (.A(_0444_),
    .B_N(_0437_),
    .Y(_0445_));
 sg13g2_xor2_1 _4132_ (.B(_0444_),
    .A(_0437_),
    .X(_0446_));
 sg13g2_inv_1 _4133_ (.Y(_0447_),
    .A(_0446_));
 sg13g2_xnor2_1 _4134_ (.Y(_0448_),
    .A(_0436_),
    .B(_0446_));
 sg13g2_nand2_1 _4135_ (.Y(_0449_),
    .A(\vgademo.soundtrack.sigma_delta_accum[6] ),
    .B(_0448_));
 sg13g2_xnor2_1 _4136_ (.Y(_0450_),
    .A(net546),
    .B(_0448_));
 sg13g2_xor2_1 _4137_ (.B(_0450_),
    .A(_0435_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[6] ));
 sg13g2_o21ai_1 _4138_ (.B1(_0449_),
    .Y(_0451_),
    .A1(_0435_),
    .A2(_0450_));
 sg13g2_a21oi_1 _4139_ (.A1(_0436_),
    .A2(_0447_),
    .Y(_0452_),
    .B1(_0445_));
 sg13g2_o21ai_1 _4140_ (.B1(_0441_),
    .Y(_0453_),
    .A1(_0442_),
    .A2(_0443_));
 sg13g2_o21ai_1 _4141_ (.B1(_3134_),
    .Y(_0454_),
    .A1(net1017),
    .A2(_0384_));
 sg13g2_a21oi_2 _4142_ (.B1(_0454_),
    .Y(_0455_),
    .A2(_0385_),
    .A1(net1017));
 sg13g2_nor2_1 _4143_ (.A(net1009),
    .B(_3241_),
    .Y(_0456_));
 sg13g2_nor3_1 _4144_ (.A(net1012),
    .B(net1009),
    .C(_3329_),
    .Y(_0457_));
 sg13g2_a22oi_1 _4145_ (.Y(_0458_),
    .B1(_0457_),
    .B2(_3293_),
    .A2(_0456_),
    .A1(net1012));
 sg13g2_nor2b_1 _4146_ (.A(_0458_),
    .B_N(_0455_),
    .Y(_0459_));
 sg13g2_xnor2_1 _4147_ (.Y(_0460_),
    .A(_0455_),
    .B(_0458_));
 sg13g2_xnor2_1 _4148_ (.Y(_0461_),
    .A(net1007),
    .B(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_inv_1 _4149_ (.Y(_0462_),
    .A(_0461_));
 sg13g2_xnor2_1 _4150_ (.Y(_0463_),
    .A(_0460_),
    .B(_0461_));
 sg13g2_nand2_1 _4151_ (.Y(_0464_),
    .A(_0453_),
    .B(_0463_));
 sg13g2_xnor2_1 _4152_ (.Y(_0465_),
    .A(_0453_),
    .B(_0463_));
 sg13g2_xor2_1 _4153_ (.B(_0465_),
    .A(_0452_),
    .X(_0466_));
 sg13g2_xnor2_1 _4154_ (.Y(_0467_),
    .A(net502),
    .B(_0466_));
 sg13g2_nor2b_1 _4155_ (.A(_0467_),
    .B_N(_0451_),
    .Y(_0468_));
 sg13g2_xnor2_1 _4156_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[7] ),
    .A(_0451_),
    .B(_0467_));
 sg13g2_a21oi_1 _4157_ (.A1(net502),
    .A2(_0466_),
    .Y(_0469_),
    .B1(_0468_));
 sg13g2_o21ai_1 _4158_ (.B1(_0464_),
    .Y(_0470_),
    .A1(_0452_),
    .A2(_0465_));
 sg13g2_a21oi_1 _4159_ (.A1(_0460_),
    .A2(_0462_),
    .Y(_0471_),
    .B1(_0459_));
 sg13g2_and2_1 _4160_ (.A(_3133_),
    .B(_3297_),
    .X(_0472_));
 sg13g2_and2_1 _4161_ (.A(_3134_),
    .B(_3305_),
    .X(_0473_));
 sg13g2_nand2_1 _4162_ (.Y(_0474_),
    .A(_0472_),
    .B(_0473_));
 sg13g2_xnor2_1 _4163_ (.Y(_0475_),
    .A(_0472_),
    .B(_0473_));
 sg13g2_xnor2_1 _4164_ (.Y(_0476_),
    .A(net1006),
    .B(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_xnor2_1 _4165_ (.Y(_0477_),
    .A(_0475_),
    .B(_0476_));
 sg13g2_nor2_1 _4166_ (.A(_0471_),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_xor2_1 _4167_ (.B(_0477_),
    .A(_0471_),
    .X(_0479_));
 sg13g2_xor2_1 _4168_ (.B(_0479_),
    .A(_0470_),
    .X(_0480_));
 sg13g2_nand2_1 _4169_ (.Y(_0481_),
    .A(net514),
    .B(_0480_));
 sg13g2_xnor2_1 _4170_ (.Y(_0482_),
    .A(net514),
    .B(_0480_));
 sg13g2_xor2_1 _4171_ (.B(_0482_),
    .A(_0469_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[8] ));
 sg13g2_o21ai_1 _4172_ (.B1(_0481_),
    .Y(_0483_),
    .A1(_0469_),
    .A2(_0482_));
 sg13g2_a21oi_1 _4173_ (.A1(_0470_),
    .A2(_0479_),
    .Y(_0484_),
    .B1(_0478_));
 sg13g2_o21ai_1 _4174_ (.B1(_0474_),
    .Y(_0485_),
    .A1(_0475_),
    .A2(_0476_));
 sg13g2_nor3_2 _4175_ (.A(net1008),
    .B(_3333_),
    .C(_3339_),
    .Y(_0486_));
 sg13g2_nand2_1 _4176_ (.Y(_0487_),
    .A(_3134_),
    .B(_3355_));
 sg13g2_nand3_1 _4177_ (.B(_3355_),
    .C(_0486_),
    .A(_3134_),
    .Y(_0488_));
 sg13g2_xor2_1 _4178_ (.B(_0487_),
    .A(_0486_),
    .X(_0489_));
 sg13g2_xnor2_1 _4179_ (.Y(_0490_),
    .A(net1006),
    .B(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_xnor2_1 _4180_ (.Y(_0491_),
    .A(_0489_),
    .B(_0490_));
 sg13g2_nand2b_1 _4181_ (.Y(_0492_),
    .B(_0485_),
    .A_N(_0491_));
 sg13g2_xor2_1 _4182_ (.B(_0491_),
    .A(_0485_),
    .X(_0493_));
 sg13g2_xor2_1 _4183_ (.B(_0493_),
    .A(_0484_),
    .X(_0494_));
 sg13g2_xnor2_1 _4184_ (.Y(_0495_),
    .A(net520),
    .B(_0494_));
 sg13g2_nor2b_1 _4185_ (.A(_0495_),
    .B_N(_0483_),
    .Y(_0496_));
 sg13g2_xnor2_1 _4186_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .A(_0483_),
    .B(_0495_));
 sg13g2_a21o_1 _4187_ (.A2(_0494_),
    .A1(net520),
    .B1(_0496_),
    .X(_0497_));
 sg13g2_o21ai_1 _4188_ (.B1(_0492_),
    .Y(_0498_),
    .A1(_0484_),
    .A2(_0493_));
 sg13g2_o21ai_1 _4189_ (.B1(_0488_),
    .Y(_0499_),
    .A1(_0489_),
    .A2(_0490_));
 sg13g2_nor2_1 _4190_ (.A(net1009),
    .B(_3372_),
    .Y(_0500_));
 sg13g2_nor2_1 _4191_ (.A(net1015),
    .B(_3381_),
    .Y(_0501_));
 sg13g2_xnor2_1 _4192_ (.Y(_0502_),
    .A(_0500_),
    .B(_0501_));
 sg13g2_xor2_1 _4193_ (.B(\vgademo.soundtrack.tri_osc_p[11] ),
    .A(net1006),
    .X(_0503_));
 sg13g2_nor2b_1 _4194_ (.A(_0502_),
    .B_N(_0503_),
    .Y(_0504_));
 sg13g2_xnor2_1 _4195_ (.Y(_0505_),
    .A(_0502_),
    .B(_0503_));
 sg13g2_xnor2_1 _4196_ (.Y(_0506_),
    .A(_0499_),
    .B(_0505_));
 sg13g2_nor2b_1 _4197_ (.A(_0506_),
    .B_N(_0498_),
    .Y(_0507_));
 sg13g2_xnor2_1 _4198_ (.Y(_0508_),
    .A(_0498_),
    .B(_0506_));
 sg13g2_xnor2_1 _4199_ (.Y(_0509_),
    .A(net533),
    .B(_0508_));
 sg13g2_nor2b_1 _4200_ (.A(_0509_),
    .B_N(_0497_),
    .Y(_0510_));
 sg13g2_xnor2_1 _4201_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .A(_0497_),
    .B(_0509_));
 sg13g2_a21o_1 _4202_ (.A2(_0508_),
    .A1(\vgademo.soundtrack.sigma_delta_accum[10] ),
    .B1(_0510_),
    .X(_0511_));
 sg13g2_a21oi_1 _4203_ (.A1(_0499_),
    .A2(_0505_),
    .Y(_0512_),
    .B1(_0507_));
 sg13g2_a21o_1 _4204_ (.A2(_0501_),
    .A1(_0500_),
    .B1(_0504_),
    .X(_0513_));
 sg13g2_nand2b_1 _4205_ (.Y(_0514_),
    .B(_3331_),
    .A_N(_0381_));
 sg13g2_nor2_1 _4206_ (.A(net1015),
    .B(_0386_),
    .Y(_0515_));
 sg13g2_nor2b_1 _4207_ (.A(_0514_),
    .B_N(_0515_),
    .Y(_0516_));
 sg13g2_xnor2_1 _4208_ (.Y(_0517_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_xor2_1 _4209_ (.B(\vgademo.soundtrack.tri_osc_p[12] ),
    .A(net1006),
    .X(_0518_));
 sg13g2_xor2_1 _4210_ (.B(_0518_),
    .A(_0517_),
    .X(_0519_));
 sg13g2_nand2_1 _4211_ (.Y(_0520_),
    .A(_0513_),
    .B(_0519_));
 sg13g2_xnor2_1 _4212_ (.Y(_0521_),
    .A(_0513_),
    .B(_0519_));
 sg13g2_xor2_1 _4213_ (.B(_0521_),
    .A(_0512_),
    .X(_0522_));
 sg13g2_xnor2_1 _4214_ (.Y(_0523_),
    .A(net529),
    .B(_0522_));
 sg13g2_nor2b_1 _4215_ (.A(_0523_),
    .B_N(_0511_),
    .Y(_0524_));
 sg13g2_xnor2_1 _4216_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .A(_0511_),
    .B(_0523_));
 sg13g2_a21o_1 _4217_ (.A2(_0522_),
    .A1(\vgademo.soundtrack.sigma_delta_accum[11] ),
    .B1(_0524_),
    .X(_0525_));
 sg13g2_o21ai_1 _4218_ (.B1(_0520_),
    .Y(_0526_),
    .A1(_0512_),
    .A2(_0521_));
 sg13g2_a21oi_1 _4219_ (.A1(_0517_),
    .A2(_0518_),
    .Y(_0527_),
    .B1(_0516_));
 sg13g2_nor4_2 _4220_ (.A(net1011),
    .B(net1010),
    .C(net1009),
    .Y(_0528_),
    .D(_3295_));
 sg13g2_nor2_1 _4221_ (.A(net1015),
    .B(_0406_),
    .Y(_0529_));
 sg13g2_nand2_1 _4222_ (.Y(_0530_),
    .A(_0528_),
    .B(_0529_));
 sg13g2_xnor2_1 _4223_ (.Y(_0531_),
    .A(_0528_),
    .B(_0529_));
 sg13g2_xor2_1 _4224_ (.B(\vgademo.soundtrack.tri_osc_p[13] ),
    .A(net1006),
    .X(_0532_));
 sg13g2_inv_1 _4225_ (.Y(_0533_),
    .A(_0532_));
 sg13g2_xnor2_1 _4226_ (.Y(_0534_),
    .A(_0531_),
    .B(_0532_));
 sg13g2_nor2b_1 _4227_ (.A(_0527_),
    .B_N(_0534_),
    .Y(_0535_));
 sg13g2_nand2b_1 _4228_ (.Y(_0536_),
    .B(_0527_),
    .A_N(_0534_));
 sg13g2_nand2b_1 _4229_ (.Y(_0537_),
    .B(_0536_),
    .A_N(_0535_));
 sg13g2_xnor2_1 _4230_ (.Y(_0538_),
    .A(_0526_),
    .B(_0537_));
 sg13g2_xnor2_1 _4231_ (.Y(_0539_),
    .A(net522),
    .B(_0538_));
 sg13g2_nor2b_1 _4232_ (.A(_0539_),
    .B_N(_0525_),
    .Y(_0540_));
 sg13g2_xnor2_1 _4233_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .A(_0525_),
    .B(_0539_));
 sg13g2_a21o_1 _4234_ (.A2(_0538_),
    .A1(\vgademo.soundtrack.sigma_delta_accum[12] ),
    .B1(_0540_),
    .X(_0541_));
 sg13g2_a21o_1 _4235_ (.A2(_0536_),
    .A1(_0526_),
    .B1(_0535_),
    .X(_0542_));
 sg13g2_o21ai_1 _4236_ (.B1(_0530_),
    .Y(_0543_),
    .A1(_0531_),
    .A2(_0533_));
 sg13g2_inv_1 _4237_ (.Y(_0544_),
    .A(_0543_));
 sg13g2_nor4_2 _4238_ (.A(\vgademo.soundtrack.pulse_vol[1] ),
    .B(\vgademo.soundtrack.pulse_vol[2] ),
    .C(net1009),
    .Y(_0545_),
    .D(_3339_));
 sg13g2_nand2b_1 _4239_ (.Y(_0546_),
    .B(net369),
    .A_N(net1006));
 sg13g2_xnor2_1 _4240_ (.Y(_0547_),
    .A(\vgademo.soundtrack.tri_osc_p[14] ),
    .B(net1006));
 sg13g2_nand2b_1 _4241_ (.Y(_0548_),
    .B(_0547_),
    .A_N(_0545_));
 sg13g2_xnor2_1 _4242_ (.Y(_0549_),
    .A(_0545_),
    .B(_0547_));
 sg13g2_xnor2_1 _4243_ (.Y(_0550_),
    .A(_0543_),
    .B(_0549_));
 sg13g2_nand2_1 _4244_ (.Y(_0551_),
    .A(_0542_),
    .B(_0550_));
 sg13g2_xor2_1 _4245_ (.B(_0550_),
    .A(_0542_),
    .X(_0552_));
 sg13g2_xnor2_1 _4246_ (.Y(_0553_),
    .A(net512),
    .B(_0552_));
 sg13g2_nor2b_1 _4247_ (.A(_0553_),
    .B_N(_0541_),
    .Y(_0554_));
 sg13g2_xnor2_1 _4248_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .A(_0541_),
    .B(_0553_));
 sg13g2_a21o_1 _4249_ (.A2(_0552_),
    .A1(net512),
    .B1(_0554_),
    .X(_0555_));
 sg13g2_o21ai_1 _4250_ (.B1(_0551_),
    .Y(_0556_),
    .A1(_0544_),
    .A2(_0549_));
 sg13g2_or2_2 _4251_ (.X(_0557_),
    .B(_0556_),
    .A(_0548_));
 sg13g2_xnor2_1 _4252_ (.Y(_0558_),
    .A(_0548_),
    .B(_0556_));
 sg13g2_and2_1 _4253_ (.A(net572),
    .B(_0558_),
    .X(_0559_));
 sg13g2_xor2_1 _4254_ (.B(_0558_),
    .A(net572),
    .X(_0560_));
 sg13g2_xor2_1 _4255_ (.B(_0560_),
    .A(_0555_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[14] ));
 sg13g2_a21o_1 _4256_ (.A2(_0560_),
    .A1(_0555_),
    .B1(_0559_),
    .X(_0561_));
 sg13g2_and2_1 _4257_ (.A(\vgademo.soundtrack.sigma_delta_accum[15] ),
    .B(_0557_),
    .X(_0562_));
 sg13g2_xor2_1 _4258_ (.B(_0557_),
    .A(net582),
    .X(_0563_));
 sg13g2_xor2_1 _4259_ (.B(_0563_),
    .A(_0561_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[15] ));
 sg13g2_xor2_1 _4260_ (.B(\vgademo.soundtrack.sample_div[1] ),
    .A(net220),
    .X(\vgademo.soundtrack.sample_div_[1] ));
 sg13g2_nand3_1 _4261_ (.B(net471),
    .C(\vgademo.soundtrack.sample_div[1] ),
    .A(net220),
    .Y(_0564_));
 sg13g2_a21o_1 _4262_ (.A2(\vgademo.soundtrack.sample_div[1] ),
    .A1(net220),
    .B1(net471),
    .X(_0565_));
 sg13g2_and2_1 _4263_ (.A(_0564_),
    .B(net472),
    .X(\vgademo.soundtrack.sample_div_[2] ));
 sg13g2_nor2_1 _4264_ (.A(_3093_),
    .B(_0564_),
    .Y(_0566_));
 sg13g2_xnor2_1 _4265_ (.Y(\vgademo.soundtrack.sample_div_[3] ),
    .A(net245),
    .B(_0564_));
 sg13g2_and2_1 _4266_ (.A(net205),
    .B(_0566_),
    .X(_0567_));
 sg13g2_xor2_1 _4267_ (.B(_0566_),
    .A(net205),
    .X(\vgademo.soundtrack.sample_div_[4] ));
 sg13g2_xor2_1 _4268_ (.B(_0567_),
    .A(net269),
    .X(\vgademo.soundtrack.sample_div_[5] ));
 sg13g2_nand3_1 _4269_ (.B(net269),
    .C(_0567_),
    .A(net466),
    .Y(_0568_));
 sg13g2_a21o_1 _4270_ (.A2(_0567_),
    .A1(net269),
    .B1(net466),
    .X(_0569_));
 sg13g2_and2_1 _4271_ (.A(_0568_),
    .B(_0569_),
    .X(\vgademo.soundtrack.sample_div_[6] ));
 sg13g2_nor2_1 _4272_ (.A(_3092_),
    .B(_0568_),
    .Y(_0570_));
 sg13g2_xnor2_1 _4273_ (.Y(\vgademo.soundtrack.sample_div_[7] ),
    .A(net238),
    .B(_0568_));
 sg13g2_and2_1 _4274_ (.A(net207),
    .B(_0570_),
    .X(_0571_));
 sg13g2_xor2_1 _4275_ (.B(_0570_),
    .A(net207),
    .X(\vgademo.soundtrack.sample_div_[8] ));
 sg13g2_and2_1 _4276_ (.A(\vgademo.soundtrack.sample_div[9] ),
    .B(_0571_),
    .X(_0572_));
 sg13g2_nand2_1 _4277_ (.Y(_0573_),
    .A(\vgademo.soundtrack.sample_div[9] ),
    .B(_0571_));
 sg13g2_xor2_1 _4278_ (.B(_0571_),
    .A(net268),
    .X(\vgademo.soundtrack.sample_div_[9] ));
 sg13g2_nor3_1 _4279_ (.A(net997),
    .B(net998),
    .C(_3193_),
    .Y(_0574_));
 sg13g2_and2_1 _4280_ (.A(_3196_),
    .B(_0574_),
    .X(_0575_));
 sg13g2_and2_1 _4281_ (.A(_3238_),
    .B(_0575_),
    .X(_0576_));
 sg13g2_nand2_1 _4282_ (.Y(_0577_),
    .A(_3238_),
    .B(_0575_));
 sg13g2_and2_1 _4283_ (.A(net1092),
    .B(net938),
    .X(_0578_));
 sg13g2_nand2_1 _4284_ (.Y(_0579_),
    .A(net1091),
    .B(net938));
 sg13g2_nor2_1 _4285_ (.A(net926),
    .B(net917),
    .Y(_0580_));
 sg13g2_nor3_1 _4286_ (.A(net963),
    .B(net964),
    .C(\vgademo.v_count[8] ),
    .Y(_0581_));
 sg13g2_nand2_1 _4287_ (.Y(_0582_),
    .A(\vgademo.v_count[3] ),
    .B(net968));
 sg13g2_inv_1 _4288_ (.Y(_0583_),
    .A(_0582_));
 sg13g2_nor4_1 _4289_ (.A(net415),
    .B(net969),
    .C(net965),
    .D(net967),
    .Y(_0584_));
 sg13g2_nand4_1 _4290_ (.B(_0581_),
    .C(_0583_),
    .A(net962),
    .Y(_0585_),
    .D(_0584_));
 sg13g2_nor3_1 _4291_ (.A(net539),
    .B(net969),
    .C(net967),
    .Y(_0586_));
 sg13g2_nor2_1 _4292_ (.A(net965),
    .B(_0582_),
    .Y(_0587_));
 sg13g2_nand4_1 _4293_ (.B(_0581_),
    .C(_0586_),
    .A(net962),
    .Y(_0588_),
    .D(_0587_));
 sg13g2_nor2_1 _4294_ (.A(net938),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_nor2_1 _4295_ (.A(net939),
    .B(_0585_),
    .Y(_0590_));
 sg13g2_or2_1 _4296_ (.X(_0591_),
    .B(_0585_),
    .A(net939));
 sg13g2_a21o_2 _4297_ (.A2(net912),
    .A1(net1091),
    .B1(net891),
    .X(_0592_));
 sg13g2_a21oi_1 _4298_ (.A1(net1064),
    .A2(net884),
    .Y(_0593_),
    .B1(net201));
 sg13g2_o21ai_1 _4299_ (.B1(net885),
    .Y(_0594_),
    .A1(net1066),
    .A2(net922));
 sg13g2_a21o_1 _4300_ (.A2(net1064),
    .A1(net1066),
    .B1(net921),
    .X(_0595_));
 sg13g2_a21oi_1 _4301_ (.A1(net884),
    .A2(_0595_),
    .Y(_0111_),
    .B1(net202));
 sg13g2_nor2_1 _4302_ (.A(net1064),
    .B(net882),
    .Y(_0596_));
 sg13g2_nor2_1 _4303_ (.A(net506),
    .B(net921),
    .Y(_0597_));
 sg13g2_a21oi_1 _4304_ (.A1(net882),
    .A2(_0597_),
    .Y(_0112_),
    .B1(_0596_));
 sg13g2_nand3_1 _4305_ (.B(net932),
    .C(net883),
    .A(net326),
    .Y(_0598_));
 sg13g2_o21ai_1 _4306_ (.B1(_0598_),
    .Y(_0113_),
    .A1(_3089_),
    .A2(net882));
 sg13g2_nor2_1 _4307_ (.A(net326),
    .B(net882),
    .Y(_0599_));
 sg13g2_xor2_1 _4308_ (.B(net348),
    .A(net1067),
    .X(_0600_));
 sg13g2_nor2_1 _4309_ (.A(net921),
    .B(_0600_),
    .Y(_0601_));
 sg13g2_a21oi_1 _4310_ (.A1(net883),
    .A2(_0601_),
    .Y(_0114_),
    .B1(_0599_));
 sg13g2_nor2_1 _4311_ (.A(net348),
    .B(net882),
    .Y(_0602_));
 sg13g2_xor2_1 _4312_ (.B(net302),
    .A(net1067),
    .X(_0603_));
 sg13g2_nor2_1 _4313_ (.A(net921),
    .B(_0603_),
    .Y(_0604_));
 sg13g2_a21oi_1 _4314_ (.A1(net882),
    .A2(_0604_),
    .Y(_0115_),
    .B1(_0602_));
 sg13g2_nor2_1 _4315_ (.A(net302),
    .B(net882),
    .Y(_0605_));
 sg13g2_nor2_1 _4316_ (.A(\vgademo.linelfsr[6] ),
    .B(net921),
    .Y(_0606_));
 sg13g2_a21oi_1 _4317_ (.A1(net882),
    .A2(_0606_),
    .Y(_0116_),
    .B1(_0605_));
 sg13g2_nor2_1 _4318_ (.A(net374),
    .B(net883),
    .Y(_0607_));
 sg13g2_xor2_1 _4319_ (.B(\vgademo.linelfsr[7] ),
    .A(net1067),
    .X(_0608_));
 sg13g2_nor2_1 _4320_ (.A(net921),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_a21oi_1 _4321_ (.A1(net883),
    .A2(_0609_),
    .Y(_0117_),
    .B1(_0607_));
 sg13g2_nor2_1 _4322_ (.A(net426),
    .B(net883),
    .Y(_0610_));
 sg13g2_nor2_1 _4323_ (.A(\vgademo.linelfsr[8] ),
    .B(net922),
    .Y(_0611_));
 sg13g2_a21oi_1 _4324_ (.A1(net883),
    .A2(_0611_),
    .Y(_0118_),
    .B1(_0610_));
 sg13g2_xnor2_1 _4325_ (.Y(_0612_),
    .A(net1066),
    .B(net402));
 sg13g2_o21ai_1 _4326_ (.B1(net884),
    .Y(_0613_),
    .A1(net922),
    .A2(_0612_));
 sg13g2_o21ai_1 _4327_ (.B1(_0613_),
    .Y(_0614_),
    .A1(net493),
    .A2(net884));
 sg13g2_inv_1 _4328_ (.Y(_0119_),
    .A(_0614_));
 sg13g2_nor2_1 _4329_ (.A(net402),
    .B(net884),
    .Y(_0615_));
 sg13g2_nor2_1 _4330_ (.A(\vgademo.linelfsr[10] ),
    .B(net921),
    .Y(_0616_));
 sg13g2_a21oi_1 _4331_ (.A1(net884),
    .A2(_0616_),
    .Y(_0120_),
    .B1(_0615_));
 sg13g2_nand3_1 _4332_ (.B(net932),
    .C(net884),
    .A(net310),
    .Y(_0617_));
 sg13g2_o21ai_1 _4333_ (.B1(_0617_),
    .Y(_0121_),
    .A1(_3088_),
    .A2(net885));
 sg13g2_nor2_1 _4334_ (.A(net310),
    .B(net885),
    .Y(_0618_));
 sg13g2_nor2_1 _4335_ (.A(net373),
    .B(net921),
    .Y(_0619_));
 sg13g2_a21oi_1 _4336_ (.A1(net885),
    .A2(_0619_),
    .Y(_0122_),
    .B1(_0618_));
 sg13g2_o21ai_1 _4337_ (.B1(_0594_),
    .Y(_0123_),
    .A1(_3087_),
    .A2(net884));
 sg13g2_nand3_1 _4338_ (.B(net482),
    .C(net872),
    .A(\vgademo.soundtrack.tick_div[0] ),
    .Y(_0620_));
 sg13g2_nand4_1 _4339_ (.B(\vgademo.soundtrack.tick_div[2] ),
    .C(\vgademo.soundtrack.tick_div[1] ),
    .A(\vgademo.soundtrack.tick_div[0] ),
    .Y(_0621_),
    .D(net872));
 sg13g2_nor2_1 _4340_ (.A(_3094_),
    .B(_0621_),
    .Y(_0622_));
 sg13g2_and2_1 _4341_ (.A(net216),
    .B(_0622_),
    .X(_0623_));
 sg13g2_and3_2 _4342_ (.X(_0624_),
    .A(net198),
    .B(net263),
    .C(_0623_));
 sg13g2_and2_1 _4343_ (.A(net599),
    .B(_0624_),
    .X(_0625_));
 sg13g2_nand2_1 _4344_ (.Y(_0626_),
    .A(net270),
    .B(_0624_));
 sg13g2_or2_1 _4345_ (.X(_0627_),
    .B(\vgademo.audio_beat_out[0] ),
    .A(\vgademo.audio_beat_out[1] ));
 sg13g2_nor4_2 _4346_ (.A(\vgademo.audio_beat_out[3] ),
    .B(\vgademo.audio_beat_out[2] ),
    .C(\vgademo.audio_beat_out[4] ),
    .Y(_0628_),
    .D(_0627_));
 sg13g2_or4_2 _4347_ (.A(\vgademo.audio_beat_out[3] ),
    .B(\vgademo.audio_beat_out[2] ),
    .C(\vgademo.audio_beat_out[4] ),
    .D(_0627_),
    .X(_0629_));
 sg13g2_nand2_1 _4348_ (.Y(_0630_),
    .A(_0625_),
    .B(net945));
 sg13g2_nand3_1 _4349_ (.B(net851),
    .C(net945),
    .A(_3090_),
    .Y(_0631_));
 sg13g2_mux2_1 _4350_ (.A0(net1063),
    .A1(net275),
    .S(net849),
    .X(_0124_));
 sg13g2_nand2_1 _4351_ (.Y(_0632_),
    .A(net203),
    .B(net850));
 sg13g2_o21ai_1 _4352_ (.B1(_0632_),
    .Y(_0125_),
    .A1(_3268_),
    .A2(net850));
 sg13g2_nor2_2 _4353_ (.A(net949),
    .B(_3262_),
    .Y(_0633_));
 sg13g2_nand2_2 _4354_ (.Y(_0634_),
    .A(net1055),
    .B(_3267_));
 sg13g2_nor2_1 _4355_ (.A(net1057),
    .B(_3267_),
    .Y(_0635_));
 sg13g2_nor2_1 _4356_ (.A(_0633_),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_nand2_1 _4357_ (.Y(_0637_),
    .A(net196),
    .B(net849));
 sg13g2_o21ai_1 _4358_ (.B1(_0637_),
    .Y(_0126_),
    .A1(net850),
    .A2(_0636_));
 sg13g2_nand2_1 _4359_ (.Y(_0638_),
    .A(net1062),
    .B(net948));
 sg13g2_xnor2_1 _4360_ (.Y(_0639_),
    .A(net1054),
    .B(_0633_));
 sg13g2_mux2_1 _4361_ (.A0(_0639_),
    .A1(net277),
    .S(net849),
    .X(_0127_));
 sg13g2_nand2_1 _4362_ (.Y(_0640_),
    .A(net1049),
    .B(net1052));
 sg13g2_nor2_2 _4363_ (.A(_0634_),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_nand2_1 _4364_ (.Y(_0642_),
    .A(net1052),
    .B(net1056));
 sg13g2_a21oi_2 _4365_ (.B1(net1050),
    .Y(_0643_),
    .A2(_0633_),
    .A1(net1051));
 sg13g2_nor2_1 _4366_ (.A(_0641_),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_nand2_1 _4367_ (.Y(_0645_),
    .A(net190),
    .B(net850));
 sg13g2_o21ai_1 _4368_ (.B1(_0645_),
    .Y(_0128_),
    .A1(net850),
    .A2(net904));
 sg13g2_nand3_1 _4369_ (.B(net1053),
    .C(net1043),
    .A(net1047),
    .Y(_0646_));
 sg13g2_xnor2_1 _4370_ (.Y(_0647_),
    .A(net946),
    .B(_0641_));
 sg13g2_nand2_1 _4371_ (.Y(_0648_),
    .A(net193),
    .B(net849));
 sg13g2_o21ai_1 _4372_ (.B1(_0648_),
    .Y(_0129_),
    .A1(net849),
    .A2(_0647_));
 sg13g2_nand3_1 _4373_ (.B(net1042),
    .C(_0641_),
    .A(net1044),
    .Y(_0649_));
 sg13g2_o21ai_1 _4374_ (.B1(_3099_),
    .Y(_0650_),
    .A1(_0634_),
    .A2(_0646_));
 sg13g2_nand2_1 _4375_ (.Y(_0651_),
    .A(_0649_),
    .B(_0650_));
 sg13g2_mux2_1 _4376_ (.A0(_0651_),
    .A1(net273),
    .S(net849),
    .X(_0130_));
 sg13g2_xnor2_1 _4377_ (.Y(_0652_),
    .A(net1041),
    .B(_0649_));
 sg13g2_nand2_1 _4378_ (.Y(_0653_),
    .A(net191),
    .B(net849));
 sg13g2_o21ai_1 _4379_ (.B1(_0653_),
    .Y(_0131_),
    .A1(net849),
    .A2(_0652_));
 sg13g2_nor2_1 _4380_ (.A(\vgademo.plane_dx_div.i[1] ),
    .B(net332),
    .Y(_0654_));
 sg13g2_nor4_2 _4381_ (.A(\vgademo.plane_dx_div.i[3] ),
    .B(\vgademo.plane_dx_div.i[2] ),
    .C(\vgademo.plane_dx_div.i[1] ),
    .Y(_0655_),
    .D(net332));
 sg13g2_nand3_1 _4382_ (.B(net998),
    .C(\vgademo.h_count[7] ),
    .A(net997),
    .Y(_0656_));
 sg13g2_nor2_2 _4383_ (.A(net996),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_nand3_1 _4384_ (.B(_3238_),
    .C(_0657_),
    .A(_3196_),
    .Y(_0658_));
 sg13g2_and3_1 _4385_ (.X(_0659_),
    .A(_3196_),
    .B(_3238_),
    .C(_0657_));
 sg13g2_nand3_1 _4386_ (.B(_3238_),
    .C(_0657_),
    .A(_3196_),
    .Y(_0660_));
 sg13g2_nor2_1 _4387_ (.A(_0655_),
    .B(net936),
    .Y(_0661_));
 sg13g2_and2_1 _4388_ (.A(_0655_),
    .B(net937),
    .X(_0662_));
 sg13g2_nand2_2 _4389_ (.Y(_0663_),
    .A(_0655_),
    .B(net937));
 sg13g2_a22oi_1 _4390_ (.Y(_0132_),
    .B1(net901),
    .B2(_3085_),
    .A2(net903),
    .A1(_3086_));
 sg13g2_a22oi_1 _4391_ (.Y(_0664_),
    .B1(net901),
    .B2(net510),
    .A2(net903),
    .A1(net1040));
 sg13g2_inv_1 _4392_ (.Y(_0133_),
    .A(net511));
 sg13g2_a22oi_1 _4393_ (.Y(_0665_),
    .B1(net901),
    .B2(net553),
    .A2(net903),
    .A1(net510));
 sg13g2_inv_1 _4394_ (.Y(_0134_),
    .A(_0665_));
 sg13g2_a22oi_1 _4395_ (.Y(_0666_),
    .B1(net901),
    .B2(net209),
    .A2(net903),
    .A1(\vgademo.plane_dx[3] ));
 sg13g2_inv_1 _4396_ (.Y(_0135_),
    .A(net210));
 sg13g2_a22oi_1 _4397_ (.Y(_0667_),
    .B1(net900),
    .B2(net1037),
    .A2(net902),
    .A1(net209));
 sg13g2_inv_1 _4398_ (.Y(_0136_),
    .A(_0667_));
 sg13g2_a22oi_1 _4399_ (.Y(_0668_),
    .B1(net901),
    .B2(net392),
    .A2(net903),
    .A1(net1037));
 sg13g2_inv_1 _4400_ (.Y(_0137_),
    .A(_0668_));
 sg13g2_a22oi_1 _4401_ (.Y(_0669_),
    .B1(net900),
    .B2(net1034),
    .A2(net902),
    .A1(net1036));
 sg13g2_inv_1 _4402_ (.Y(_0138_),
    .A(_0669_));
 sg13g2_a22oi_1 _4403_ (.Y(_0670_),
    .B1(net900),
    .B2(net1033),
    .A2(net902),
    .A1(net1034));
 sg13g2_inv_1 _4404_ (.Y(_0139_),
    .A(_0670_));
 sg13g2_a22oi_1 _4405_ (.Y(_0671_),
    .B1(net900),
    .B2(net1032),
    .A2(net903),
    .A1(net355));
 sg13g2_inv_1 _4406_ (.Y(_0140_),
    .A(net356));
 sg13g2_a22oi_1 _4407_ (.Y(_0672_),
    .B1(net900),
    .B2(net1030),
    .A2(net902),
    .A1(net1032));
 sg13g2_inv_1 _4408_ (.Y(_0141_),
    .A(_0672_));
 sg13g2_o21ai_1 _4409_ (.B1(_0660_),
    .Y(_0142_),
    .A1(_3081_),
    .A2(_0655_));
 sg13g2_and2_1 _4410_ (.A(\vgademo.plane_dx_div.i[1] ),
    .B(net332),
    .X(_0673_));
 sg13g2_nor3_1 _4411_ (.A(net333),
    .B(net936),
    .C(_0673_),
    .Y(_0143_));
 sg13g2_nand2_1 _4412_ (.Y(_0674_),
    .A(net451),
    .B(_0673_));
 sg13g2_o21ai_1 _4413_ (.B1(_0660_),
    .Y(_0675_),
    .A1(net451),
    .A2(_0673_));
 sg13g2_nor2b_1 _4414_ (.A(net452),
    .B_N(_0674_),
    .Y(_0144_));
 sg13g2_xor2_1 _4415_ (.B(_0674_),
    .A(net418),
    .X(_0676_));
 sg13g2_nor2_1 _4416_ (.A(net936),
    .B(net419),
    .Y(_0145_));
 sg13g2_nor2_2 _4417_ (.A(_0626_),
    .B(net945),
    .Y(_0677_));
 sg13g2_nand2_2 _4418_ (.Y(_0678_),
    .A(net851),
    .B(_0629_));
 sg13g2_nor2_1 _4419_ (.A(net322),
    .B(_0677_),
    .Y(_0679_));
 sg13g2_a21oi_1 _4420_ (.A1(net322),
    .A2(net851),
    .Y(_0146_),
    .B1(_0679_));
 sg13g2_and3_1 _4421_ (.X(_0680_),
    .A(net371),
    .B(net322),
    .C(net851));
 sg13g2_nand3_1 _4422_ (.B(net322),
    .C(net851),
    .A(net371),
    .Y(_0681_));
 sg13g2_a21oi_1 _4423_ (.A1(net322),
    .A2(net851),
    .Y(_0682_),
    .B1(net371));
 sg13g2_o21ai_1 _4424_ (.B1(_0631_),
    .Y(_0147_),
    .A1(_0680_),
    .A2(_0682_));
 sg13g2_nor2_1 _4425_ (.A(net353),
    .B(_0681_),
    .Y(_0683_));
 sg13g2_o21ai_1 _4426_ (.B1(net850),
    .Y(_0684_),
    .A1(net353),
    .A2(_0681_));
 sg13g2_nor2_1 _4427_ (.A(net353),
    .B(_0626_),
    .Y(_0685_));
 sg13g2_a21oi_1 _4428_ (.A1(net1029),
    .A2(_0626_),
    .Y(_0686_),
    .B1(_0685_));
 sg13g2_a21oi_1 _4429_ (.A1(_0681_),
    .A2(_0686_),
    .Y(_0148_),
    .B1(_0684_));
 sg13g2_o21ai_1 _4430_ (.B1(_0631_),
    .Y(_0687_),
    .A1(\vgademo.audio_beat_out[3] ),
    .A2(_0684_));
 sg13g2_a21oi_1 _4431_ (.A1(\vgademo.audio_beat_out[3] ),
    .A2(_0683_),
    .Y(_0149_),
    .B1(_0687_));
 sg13g2_nand3_1 _4432_ (.B(net1029),
    .C(_0680_),
    .A(\vgademo.audio_beat_out[3] ),
    .Y(_0688_));
 sg13g2_xor2_1 _4433_ (.B(_0688_),
    .A(net490),
    .X(_0689_));
 sg13g2_nand2_1 _4434_ (.Y(_0150_),
    .A(_0631_),
    .B(net491));
 sg13g2_nand2_1 _4435_ (.Y(_0690_),
    .A(net948),
    .B(_3261_));
 sg13g2_o21ai_1 _4436_ (.B1(net1046),
    .Y(_0691_),
    .A1(net1062),
    .A2(_0690_));
 sg13g2_a21oi_1 _4437_ (.A1(net1050),
    .A2(_0691_),
    .Y(_0692_),
    .B1(_3267_));
 sg13g2_nor2_1 _4438_ (.A(net1051),
    .B(_3267_),
    .Y(_0693_));
 sg13g2_a21oi_1 _4439_ (.A1(_3262_),
    .A2(_0693_),
    .Y(_0694_),
    .B1(_0647_));
 sg13g2_o21ai_1 _4440_ (.B1(_0694_),
    .Y(_0695_),
    .A1(_3271_),
    .A2(_0639_));
 sg13g2_nor2_1 _4441_ (.A(net947),
    .B(\vgademo.audio_songpos[6] ),
    .Y(_0696_));
 sg13g2_nor3_1 _4442_ (.A(_0641_),
    .B(_0643_),
    .C(_0696_),
    .Y(_0697_));
 sg13g2_a21oi_1 _4443_ (.A1(_0695_),
    .A2(_0697_),
    .Y(_0698_),
    .B1(_0692_));
 sg13g2_o21ai_1 _4444_ (.B1(net851),
    .Y(_0699_),
    .A1(_0629_),
    .A2(_0698_));
 sg13g2_nor2_1 _4445_ (.A(\vgademo.audio_kick_frames[0] ),
    .B(net368),
    .Y(_0700_));
 sg13g2_and2_1 _4446_ (.A(_0060_),
    .B(_0700_),
    .X(_0701_));
 sg13g2_nand2_1 _4447_ (.Y(_0702_),
    .A(_0060_),
    .B(_0700_));
 sg13g2_nand2b_2 _4448_ (.Y(_0703_),
    .B(net1056),
    .A_N(net1058));
 sg13g2_nor2b_2 _4449_ (.A(_3279_),
    .B_N(_0703_),
    .Y(_0704_));
 sg13g2_nand2_1 _4450_ (.Y(_0705_),
    .A(_3280_),
    .B(_0703_));
 sg13g2_a221oi_1 _4451_ (.B2(net1049),
    .C1(net947),
    .B1(_0705_),
    .A1(_3250_),
    .Y(_0706_),
    .A2(_3257_));
 sg13g2_nand4_1 _4452_ (.B(net947),
    .C(_3250_),
    .A(net1049),
    .Y(_0707_),
    .D(_0690_));
 sg13g2_o21ai_1 _4453_ (.B1(_3244_),
    .Y(_0708_),
    .A1(net1052),
    .A2(_0704_));
 sg13g2_nand3b_1 _4454_ (.B(_0707_),
    .C(_0708_),
    .Y(_0709_),
    .A_N(_0706_));
 sg13g2_nand2_2 _4455_ (.Y(_0710_),
    .A(net1049),
    .B(net948));
 sg13g2_nor2_1 _4456_ (.A(_3279_),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_and2_1 _4457_ (.A(net1058),
    .B(_0642_),
    .X(_0712_));
 sg13g2_a21oi_2 _4458_ (.B1(net947),
    .Y(_0713_),
    .A2(_0712_),
    .A1(_3257_));
 sg13g2_or2_1 _4459_ (.X(_0714_),
    .B(_0640_),
    .A(_3279_));
 sg13g2_or2_1 _4460_ (.X(_0715_),
    .B(_0710_),
    .A(_0703_));
 sg13g2_o21ai_1 _4461_ (.B1(_0715_),
    .Y(_0716_),
    .A1(net1049),
    .A2(_3279_));
 sg13g2_nor2_1 _4462_ (.A(net1045),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_a21oi_2 _4463_ (.B1(_0717_),
    .Y(_0718_),
    .A2(_0714_),
    .A1(_0713_));
 sg13g2_a21o_2 _4464_ (.A2(_0714_),
    .A1(_0713_),
    .B1(_0717_),
    .X(_0719_));
 sg13g2_a22oi_1 _4465_ (.Y(_0720_),
    .B1(_0718_),
    .B2(_3244_),
    .A2(_0711_),
    .A1(net1045));
 sg13g2_a21oi_1 _4466_ (.A1(net889),
    .A2(_0720_),
    .Y(_0721_),
    .B1(net943));
 sg13g2_nor2_1 _4467_ (.A(net945),
    .B(net943),
    .Y(_0722_));
 sg13g2_nand2b_1 _4468_ (.Y(_0723_),
    .B(\vgademo.soundtrack.tri_osc_i[3] ),
    .A_N(\vgademo.soundtrack.tri_osc_i[0] ));
 sg13g2_xor2_1 _4469_ (.B(\vgademo.soundtrack.tri_osc_i[3] ),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(_0724_));
 sg13g2_o21ai_1 _4470_ (.B1(_0629_),
    .Y(_0725_),
    .A1(net944),
    .A2(_0724_));
 sg13g2_nor3_1 _4471_ (.A(net847),
    .B(_0721_),
    .C(_0725_),
    .Y(_0726_));
 sg13g2_a21o_1 _4472_ (.A2(net847),
    .A1(net467),
    .B1(_0726_),
    .X(_0151_));
 sg13g2_nor2b_1 _4473_ (.A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B_N(\vgademo.soundtrack.tri_osc_i[1] ),
    .Y(_0727_));
 sg13g2_xnor2_1 _4474_ (.Y(_0728_),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .B(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_xnor2_1 _4475_ (.Y(_0729_),
    .A(_0723_),
    .B(_0728_));
 sg13g2_nand2b_1 _4476_ (.Y(_0730_),
    .B(_0720_),
    .A_N(net889));
 sg13g2_nor2_1 _4477_ (.A(net1051),
    .B(_3097_),
    .Y(_0731_));
 sg13g2_nand2_1 _4478_ (.Y(_0732_),
    .A(net948),
    .B(net1055));
 sg13g2_a21oi_2 _4479_ (.B1(_3095_),
    .Y(_0733_),
    .A2(_3256_),
    .A1(_3246_));
 sg13g2_nor3_1 _4480_ (.A(net1045),
    .B(_0711_),
    .C(_0733_),
    .Y(_0734_));
 sg13g2_a21oi_2 _4481_ (.B1(_0734_),
    .Y(_0735_),
    .A2(_0711_),
    .A1(net1045));
 sg13g2_nand2_1 _4482_ (.Y(_0736_),
    .A(_0718_),
    .B(_0735_));
 sg13g2_a21oi_1 _4483_ (.A1(net889),
    .A2(_0736_),
    .Y(_0737_),
    .B1(net943));
 sg13g2_a221oi_1 _4484_ (.B2(_0737_),
    .C1(_0678_),
    .B1(_0730_),
    .A1(net943),
    .Y(_0738_),
    .A2(_0729_));
 sg13g2_a21o_1 _4485_ (.A2(net847),
    .A1(net481),
    .B1(_0738_),
    .X(_0152_));
 sg13g2_nand2_1 _4486_ (.Y(_0739_),
    .A(_0710_),
    .B(_0719_));
 sg13g2_nand3_1 _4487_ (.B(_0713_),
    .C(_0719_),
    .A(_0710_),
    .Y(_0740_));
 sg13g2_a21oi_1 _4488_ (.A1(_0718_),
    .A2(_0735_),
    .Y(_0741_),
    .B1(net889));
 sg13g2_nor2_1 _4489_ (.A(net943),
    .B(_0741_),
    .Y(_0742_));
 sg13g2_a21oi_1 _4490_ (.A1(_0723_),
    .A2(_0728_),
    .Y(_0743_),
    .B1(_0727_));
 sg13g2_nand2_1 _4491_ (.Y(_0744_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(_3128_));
 sg13g2_xnor2_1 _4492_ (.Y(_0745_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_nand2b_1 _4493_ (.Y(_0746_),
    .B(_0745_),
    .A_N(_0743_));
 sg13g2_xor2_1 _4494_ (.B(_0745_),
    .A(_0743_),
    .X(_0747_));
 sg13g2_a221oi_1 _4495_ (.B2(net943),
    .C1(_0678_),
    .B1(_0747_),
    .A1(_0740_),
    .Y(_0748_),
    .A2(_0742_));
 sg13g2_a21o_1 _4496_ (.A2(net847),
    .A1(net480),
    .B1(_0748_),
    .X(_0153_));
 sg13g2_nand2_1 _4497_ (.Y(_0749_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(_3129_));
 sg13g2_xor2_1 _4498_ (.B(\vgademo.soundtrack.tri_osc_i[6] ),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .X(_0750_));
 sg13g2_nand3_1 _4499_ (.B(_0746_),
    .C(_0750_),
    .A(_0744_),
    .Y(_0751_));
 sg13g2_a21o_1 _4500_ (.A2(_0746_),
    .A1(_0744_),
    .B1(_0750_),
    .X(_0752_));
 sg13g2_a21oi_1 _4501_ (.A1(_0751_),
    .A2(_0752_),
    .Y(_0753_),
    .B1(net944));
 sg13g2_o21ai_1 _4502_ (.B1(_0713_),
    .Y(_0754_),
    .A1(_3280_),
    .A2(_0710_));
 sg13g2_o21ai_1 _4503_ (.B1(_0754_),
    .Y(_0755_),
    .A1(net1045),
    .A2(_0715_));
 sg13g2_inv_1 _4504_ (.Y(_0756_),
    .A(_0755_));
 sg13g2_nand2_1 _4505_ (.Y(_0757_),
    .A(_0735_),
    .B(_0756_));
 sg13g2_mux2_1 _4506_ (.A0(_0719_),
    .A1(_0739_),
    .S(_0757_),
    .X(_0758_));
 sg13g2_o21ai_1 _4507_ (.B1(net944),
    .Y(_0759_),
    .A1(net889),
    .A2(_0740_));
 sg13g2_a21oi_1 _4508_ (.A1(net890),
    .A2(_0758_),
    .Y(_0760_),
    .B1(_0759_));
 sg13g2_nor2_1 _4509_ (.A(_0753_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_a22oi_1 _4510_ (.Y(_0762_),
    .B1(_0761_),
    .B2(_0677_),
    .A2(net847),
    .A1(net558));
 sg13g2_inv_1 _4511_ (.Y(_0154_),
    .A(_0762_));
 sg13g2_nand2_1 _4512_ (.Y(_0763_),
    .A(net524),
    .B(net848));
 sg13g2_o21ai_1 _4513_ (.B1(_0735_),
    .Y(_0764_),
    .A1(_0718_),
    .A2(_0755_));
 sg13g2_mux2_1 _4514_ (.A0(_0758_),
    .A1(_0764_),
    .S(net889),
    .X(_0765_));
 sg13g2_xor2_1 _4515_ (.B(\vgademo.soundtrack.tri_osc_i[7] ),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .X(_0766_));
 sg13g2_nand3_1 _4516_ (.B(_0752_),
    .C(_0766_),
    .A(_0749_),
    .Y(_0767_));
 sg13g2_a21oi_1 _4517_ (.A1(_0749_),
    .A2(_0752_),
    .Y(_0768_),
    .B1(_0766_));
 sg13g2_nor2_1 _4518_ (.A(net944),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_a22oi_1 _4519_ (.Y(_0770_),
    .B1(_0767_),
    .B2(_0769_),
    .A2(_0765_),
    .A1(net944));
 sg13g2_o21ai_1 _4520_ (.B1(_0763_),
    .Y(_0155_),
    .A1(_0678_),
    .A2(_0770_));
 sg13g2_nand2b_1 _4521_ (.Y(_0771_),
    .B(_0764_),
    .A_N(net890));
 sg13g2_nand3_1 _4522_ (.B(_0719_),
    .C(_0757_),
    .A(net890),
    .Y(_0772_));
 sg13g2_nand3_1 _4523_ (.B(_0771_),
    .C(_0772_),
    .A(net944),
    .Y(_0773_));
 sg13g2_a21oi_1 _4524_ (.A1(\vgademo.soundtrack.tri_osc_i[4] ),
    .A2(_3130_),
    .Y(_0774_),
    .B1(_0768_));
 sg13g2_nor2_1 _4525_ (.A(_3128_),
    .B(\vgademo.soundtrack.tri_osc_i[8] ),
    .Y(_0775_));
 sg13g2_xor2_1 _4526_ (.B(\vgademo.soundtrack.tri_osc_i[8] ),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(_0776_));
 sg13g2_xnor2_1 _4527_ (.Y(_0777_),
    .A(_0774_),
    .B(_0776_));
 sg13g2_a21oi_1 _4528_ (.A1(_0702_),
    .A2(_0777_),
    .Y(_0778_),
    .B1(_0678_));
 sg13g2_a22oi_1 _4529_ (.Y(_0779_),
    .B1(_0773_),
    .B2(_0778_),
    .A2(net848),
    .A1(net571));
 sg13g2_inv_1 _4530_ (.Y(_0156_),
    .A(_0779_));
 sg13g2_a21oi_1 _4531_ (.A1(_3128_),
    .A2(\vgademo.soundtrack.tri_osc_i[8] ),
    .Y(_0780_),
    .B1(_0774_));
 sg13g2_nor3_2 _4532_ (.A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(_0775_),
    .C(_0780_),
    .Y(_0781_));
 sg13g2_o21ai_1 _4533_ (.B1(\vgademo.soundtrack.tri_osc_i[6] ),
    .Y(_0782_),
    .A1(_0775_),
    .A2(_0780_));
 sg13g2_nand2_1 _4534_ (.Y(_0783_),
    .A(net943),
    .B(_0782_));
 sg13g2_o21ai_1 _4535_ (.B1(_0719_),
    .Y(_0784_),
    .A1(net890),
    .A2(_0757_));
 sg13g2_nand2_1 _4536_ (.Y(_0785_),
    .A(net944),
    .B(_0784_));
 sg13g2_o21ai_1 _4537_ (.B1(_0785_),
    .Y(_0786_),
    .A1(_0781_),
    .A2(_0783_));
 sg13g2_a22oi_1 _4538_ (.Y(_0157_),
    .B1(_0786_),
    .B2(_0677_),
    .A2(net848),
    .A1(_3129_));
 sg13g2_xnor2_1 _4539_ (.Y(_0787_),
    .A(_3130_),
    .B(_0781_));
 sg13g2_o21ai_1 _4540_ (.B1(net944),
    .Y(_0788_),
    .A1(net889),
    .A2(_0719_));
 sg13g2_a21oi_1 _4541_ (.A1(net889),
    .A2(_0719_),
    .Y(_0789_),
    .B1(_0788_));
 sg13g2_a21oi_1 _4542_ (.A1(net943),
    .A2(_0787_),
    .Y(_0790_),
    .B1(_0789_));
 sg13g2_a22oi_1 _4543_ (.Y(_0158_),
    .B1(_0790_),
    .B2(_0677_),
    .A2(net847),
    .A1(_3130_));
 sg13g2_a21oi_1 _4544_ (.A1(_3130_),
    .A2(_0781_),
    .Y(_0791_),
    .B1(_3131_));
 sg13g2_o21ai_1 _4545_ (.B1(_0788_),
    .Y(_0792_),
    .A1(_0701_),
    .A2(_0791_));
 sg13g2_a22oi_1 _4546_ (.Y(_0159_),
    .B1(_0792_),
    .B2(_0677_),
    .A2(net848),
    .A1(_3131_));
 sg13g2_nor2_1 _4547_ (.A(net1077),
    .B(net261),
    .Y(_0793_));
 sg13g2_a21oi_2 _4548_ (.B1(_0562_),
    .Y(_0794_),
    .A2(_0563_),
    .A1(_0561_));
 sg13g2_a21oi_1 _4549_ (.A1(net1077),
    .A2(_0794_),
    .Y(_0160_),
    .B1(_0793_));
 sg13g2_mux2_1 _4550_ (.A0(\vgademo.soundtrack.tick_div[0] ),
    .A1(net180),
    .S(net872),
    .X(_0161_));
 sg13g2_a21o_1 _4551_ (.A2(net872),
    .A1(\vgademo.soundtrack.tick_div[0] ),
    .B1(net482),
    .X(_0795_));
 sg13g2_and2_1 _4552_ (.A(_0620_),
    .B(net483),
    .X(_0162_));
 sg13g2_xnor2_1 _4553_ (.Y(_0163_),
    .A(net240),
    .B(_0620_));
 sg13g2_xnor2_1 _4554_ (.Y(_0164_),
    .A(net231),
    .B(_0621_));
 sg13g2_xor2_1 _4555_ (.B(_0622_),
    .A(net216),
    .X(_0165_));
 sg13g2_xor2_1 _4556_ (.B(_0623_),
    .A(net263),
    .X(_0166_));
 sg13g2_a21oi_1 _4557_ (.A1(\vgademo.soundtrack.tick_div[5] ),
    .A2(_0623_),
    .Y(_0796_),
    .B1(net198));
 sg13g2_nor2_1 _4558_ (.A(_0624_),
    .B(net199),
    .Y(_0167_));
 sg13g2_xor2_1 _4559_ (.B(_0624_),
    .A(net270),
    .X(_0168_));
 sg13g2_nand2_1 _4560_ (.Y(_0797_),
    .A(_0093_),
    .B(net870));
 sg13g2_o21ai_1 _4561_ (.B1(_0797_),
    .Y(_0169_),
    .A1(net166),
    .A2(net871));
 sg13g2_nand2_1 _4562_ (.Y(_0798_),
    .A(_0094_),
    .B(net870));
 sg13g2_o21ai_1 _4563_ (.B1(_0798_),
    .Y(_0170_),
    .A1(net174),
    .A2(net870));
 sg13g2_nand2_1 _4564_ (.Y(_0799_),
    .A(_0095_),
    .B(net870));
 sg13g2_o21ai_1 _4565_ (.B1(_0799_),
    .Y(_0171_),
    .A1(net168),
    .A2(net870));
 sg13g2_mux2_1 _4566_ (.A0(net222),
    .A1(_0040_),
    .S(net873),
    .X(_0172_));
 sg13g2_mux2_1 _4567_ (.A0(net229),
    .A1(\vgademo.soundtrack.noise_lfsr[5] ),
    .S(net873),
    .X(_0173_));
 sg13g2_mux2_1 _4568_ (.A0(_0097_),
    .A1(net184),
    .S(net872),
    .X(_0174_));
 sg13g2_mux2_1 _4569_ (.A0(\vgademo.soundtrack.noise_lfsr[6] ),
    .A1(net247),
    .S(net873),
    .X(_0175_));
 sg13g2_mux2_1 _4570_ (.A0(_0098_),
    .A1(net178),
    .S(net872),
    .X(_0176_));
 sg13g2_mux2_1 _4571_ (.A0(net300),
    .A1(\vgademo.soundtrack.noise_lfsr[9] ),
    .S(net872),
    .X(_0177_));
 sg13g2_mux2_1 _4572_ (.A0(net170),
    .A1(\vgademo.soundtrack.noise_lfsr[9] ),
    .S(net870),
    .X(_0178_));
 sg13g2_nand2_1 _4573_ (.Y(_0800_),
    .A(net186),
    .B(net871));
 sg13g2_o21ai_1 _4574_ (.B1(_0800_),
    .Y(_0179_),
    .A1(\vgademo.soundtrack.noise_lfsr[11] ),
    .A2(net870));
 sg13g2_nand2_1 _4575_ (.Y(_0801_),
    .A(_0100_),
    .B(net871));
 sg13g2_o21ai_1 _4576_ (.B1(_0801_),
    .Y(_0180_),
    .A1(net176),
    .A2(net871));
 sg13g2_mux2_1 _4577_ (.A0(_0101_),
    .A1(net182),
    .S(net873),
    .X(_0181_));
 sg13g2_xor2_1 _4578_ (.B(\vgademo.soundtrack.noise_lfsr[14] ),
    .A(\vgademo.soundtrack.noise_lfsr[0] ),
    .X(_0802_));
 sg13g2_mux2_1 _4579_ (.A0(net218),
    .A1(_0802_),
    .S(net872),
    .X(_0182_));
 sg13g2_mux2_1 _4580_ (.A0(net291),
    .A1(\vgademo.soundtrack.noise_lfsr[14] ),
    .S(net870),
    .X(_0183_));
 sg13g2_nand2_1 _4581_ (.Y(_0803_),
    .A(net850),
    .B(_0681_));
 sg13g2_nand3_1 _4582_ (.B(_3268_),
    .C(_3280_),
    .A(net1051),
    .Y(_0804_));
 sg13g2_nand3_1 _4583_ (.B(\vgademo.audio_songpos[6] ),
    .C(_0804_),
    .A(net1046),
    .Y(_0805_));
 sg13g2_nand2_1 _4584_ (.Y(_0806_),
    .A(net904),
    .B(_0805_));
 sg13g2_o21ai_1 _4585_ (.B1(_0696_),
    .Y(_0807_),
    .A1(net1062),
    .A2(_0642_));
 sg13g2_o21ai_1 _4586_ (.B1(net947),
    .Y(_0808_),
    .A1(net1056),
    .A2(_3250_));
 sg13g2_nand2_1 _4587_ (.Y(_0809_),
    .A(_0807_),
    .B(_0808_));
 sg13g2_a22oi_1 _4588_ (.Y(_0810_),
    .B1(_0809_),
    .B2(net904),
    .A2(_0806_),
    .A1(_0703_));
 sg13g2_nor2_1 _4589_ (.A(_3270_),
    .B(_0810_),
    .Y(_0811_));
 sg13g2_nor3_1 _4590_ (.A(_0641_),
    .B(_0643_),
    .C(_0805_),
    .Y(_0812_));
 sg13g2_a21oi_1 _4591_ (.A1(net1052),
    .A2(_0812_),
    .Y(_0813_),
    .B1(_0811_));
 sg13g2_o21ai_1 _4592_ (.B1(_0803_),
    .Y(_0814_),
    .A1(_0629_),
    .A2(_0813_));
 sg13g2_nand3_1 _4593_ (.B(net1028),
    .C(net1019),
    .A(net1024),
    .Y(_0815_));
 sg13g2_or2_1 _4594_ (.X(_0816_),
    .B(_0815_),
    .A(_3134_));
 sg13g2_a21oi_1 _4595_ (.A1(net1028),
    .A2(_0816_),
    .Y(_0817_),
    .B1(net945));
 sg13g2_nand2_1 _4596_ (.Y(_0818_),
    .A(net188),
    .B(_0814_));
 sg13g2_o21ai_1 _4597_ (.B1(_0818_),
    .Y(_0184_),
    .A1(_0814_),
    .A2(_0817_));
 sg13g2_xnor2_1 _4598_ (.Y(_0819_),
    .A(net1024),
    .B(net1028));
 sg13g2_a21oi_1 _4599_ (.A1(_0816_),
    .A2(_0819_),
    .Y(_0820_),
    .B1(net945));
 sg13g2_nand2_1 _4600_ (.Y(_0821_),
    .A(net194),
    .B(_0814_));
 sg13g2_o21ai_1 _4601_ (.B1(_0821_),
    .Y(_0185_),
    .A1(_0814_),
    .A2(_0820_));
 sg13g2_nor2_1 _4602_ (.A(net1014),
    .B(_0815_),
    .Y(_0822_));
 sg13g2_a21oi_1 _4603_ (.A1(net1024),
    .A2(net1028),
    .Y(_0823_),
    .B1(net1019));
 sg13g2_nor4_1 _4604_ (.A(_0628_),
    .B(_0681_),
    .C(_0822_),
    .D(_0823_),
    .Y(_0824_));
 sg13g2_a21oi_1 _4605_ (.A1(_3080_),
    .A2(_0814_),
    .Y(_0186_),
    .B1(_0824_));
 sg13g2_a21oi_1 _4606_ (.A1(_3134_),
    .A2(_0815_),
    .Y(_0825_),
    .B1(net945));
 sg13g2_nand2_1 _4607_ (.Y(_0826_),
    .A(net197),
    .B(_0814_));
 sg13g2_o21ai_1 _4608_ (.B1(_0826_),
    .Y(_0187_),
    .A1(_0814_),
    .A2(_0825_));
 sg13g2_and2_1 _4609_ (.A(net1072),
    .B(net873),
    .X(_0827_));
 sg13g2_nand2_2 _4610_ (.Y(_0828_),
    .A(net1075),
    .B(net873));
 sg13g2_nor3_1 _4611_ (.A(net946),
    .B(\vgademo.audio_songpos[6] ),
    .C(_0710_),
    .Y(_0829_));
 sg13g2_nor2_1 _4612_ (.A(net1029),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_a22oi_1 _4613_ (.Y(_0831_),
    .B1(_0704_),
    .B2(_3264_),
    .A2(_3268_),
    .A1(_3255_));
 sg13g2_a21oi_1 _4614_ (.A1(net1053),
    .A2(_0634_),
    .Y(_0832_),
    .B1(_3095_));
 sg13g2_nor2_1 _4615_ (.A(net946),
    .B(_0832_),
    .Y(_0833_));
 sg13g2_o21ai_1 _4616_ (.B1(_0833_),
    .Y(_0834_),
    .A1(net1047),
    .A2(_0831_));
 sg13g2_nand2_1 _4617_ (.Y(_0835_),
    .A(_3250_),
    .B(_3283_));
 sg13g2_a221oi_1 _4618_ (.B2(_3097_),
    .C1(_3248_),
    .B1(_0835_),
    .A1(net1062),
    .Y(_0836_),
    .A2(_0731_));
 sg13g2_a21oi_1 _4619_ (.A1(\vgademo.audio_songpos[0] ),
    .A2(net1055),
    .Y(_0837_),
    .B1(net1059));
 sg13g2_nand2_1 _4620_ (.Y(_0838_),
    .A(net948),
    .B(_0837_));
 sg13g2_o21ai_1 _4621_ (.B1(_0838_),
    .Y(_0839_),
    .A1(_3246_),
    .A2(_3267_));
 sg13g2_o21ai_1 _4622_ (.B1(_0834_),
    .Y(_0840_),
    .A1(_3245_),
    .A2(_0839_));
 sg13g2_o21ai_1 _4623_ (.B1(net1041),
    .Y(_0841_),
    .A1(_0836_),
    .A2(_0840_));
 sg13g2_nand3b_1 _4624_ (.B(net1045),
    .C(_0640_),
    .Y(_0842_),
    .A_N(_0643_));
 sg13g2_nor2b_1 _4625_ (.A(net1041),
    .B_N(_0842_),
    .Y(_0843_));
 sg13g2_nand4_1 _4626_ (.B(net946),
    .C(_3246_),
    .A(net1048),
    .Y(_0844_),
    .D(_3256_));
 sg13g2_o21ai_1 _4627_ (.B1(_3244_),
    .Y(_0845_),
    .A1(net948),
    .A2(_0704_));
 sg13g2_nand3_1 _4628_ (.B(_0844_),
    .C(_0845_),
    .A(_0843_),
    .Y(_0846_));
 sg13g2_nand3_1 _4629_ (.B(_0841_),
    .C(_0846_),
    .A(net1042),
    .Y(_0847_));
 sg13g2_a21oi_1 _4630_ (.A1(_3265_),
    .A2(_3275_),
    .Y(_0848_),
    .B1(_0635_));
 sg13g2_or2_1 _4631_ (.X(_0849_),
    .B(_0848_),
    .A(net1047));
 sg13g2_a21o_1 _4632_ (.A2(_0835_),
    .A1(_0636_),
    .B1(_3095_),
    .X(_0850_));
 sg13g2_nand2_1 _4633_ (.Y(_0851_),
    .A(_0849_),
    .B(_0850_));
 sg13g2_nor2_1 _4634_ (.A(_3245_),
    .B(_0703_),
    .Y(_0852_));
 sg13g2_a22oi_1 _4635_ (.Y(_0853_),
    .B1(_0852_),
    .B2(_0638_),
    .A2(_0851_),
    .A1(net1043));
 sg13g2_nand2_1 _4636_ (.Y(_0854_),
    .A(_3254_),
    .B(_0732_));
 sg13g2_a21o_1 _4637_ (.A2(_0854_),
    .A1(net1047),
    .B1(_0643_),
    .X(_0855_));
 sg13g2_a21oi_1 _4638_ (.A1(net1043),
    .A2(_0855_),
    .Y(_0856_),
    .B1(_3243_));
 sg13g2_nor2_1 _4639_ (.A(net1043),
    .B(net1042),
    .Y(_0857_));
 sg13g2_a221oi_1 _4640_ (.B2(_0844_),
    .C1(_0857_),
    .B1(_0856_),
    .A1(_3288_),
    .Y(_0858_),
    .A2(_0853_));
 sg13g2_a22oi_1 _4641_ (.Y(_0859_),
    .B1(_0858_),
    .B2(net1029),
    .A2(_0847_),
    .A1(_0830_));
 sg13g2_a21oi_1 _4642_ (.A1(_3266_),
    .A2(_0732_),
    .Y(_0860_),
    .B1(_3095_));
 sg13g2_o21ai_1 _4643_ (.B1(_0856_),
    .Y(_0861_),
    .A1(net1043),
    .A2(_0860_));
 sg13g2_nand3_1 _4644_ (.B(_3250_),
    .C(_3256_),
    .A(net1049),
    .Y(_0862_));
 sg13g2_a221oi_1 _4645_ (.B2(net1051),
    .C1(net1044),
    .B1(_0633_),
    .A1(net1060),
    .Y(_0863_),
    .A2(_3097_));
 sg13g2_a21oi_1 _4646_ (.A1(_3275_),
    .A2(_0863_),
    .Y(_0864_),
    .B1(_3244_));
 sg13g2_nand3_1 _4647_ (.B(_0848_),
    .C(_0862_),
    .A(net1043),
    .Y(_0865_));
 sg13g2_o21ai_1 _4648_ (.B1(_0865_),
    .Y(_0866_),
    .A1(_0643_),
    .A2(_0864_));
 sg13g2_nand2_1 _4649_ (.Y(_0867_),
    .A(_3288_),
    .B(_0866_));
 sg13g2_nand2_1 _4650_ (.Y(_0868_),
    .A(_0861_),
    .B(_0867_));
 sg13g2_nor2_1 _4651_ (.A(_0839_),
    .B(_0864_),
    .Y(_0869_));
 sg13g2_a21oi_1 _4652_ (.A1(net949),
    .A2(_3261_),
    .Y(_0870_),
    .B1(_0710_));
 sg13g2_a21oi_1 _4653_ (.A1(net1043),
    .A2(_0870_),
    .Y(_0871_),
    .B1(_0869_));
 sg13g2_nand3_1 _4654_ (.B(_3244_),
    .C(_0705_),
    .A(net1052),
    .Y(_0872_));
 sg13g2_a221oi_1 _4655_ (.B2(_0843_),
    .C1(_3099_),
    .B1(_0872_),
    .A1(net1041),
    .Y(_0873_),
    .A2(_0871_));
 sg13g2_nor2_1 _4656_ (.A(net1047),
    .B(net1042),
    .Y(_0874_));
 sg13g2_nor2_2 _4657_ (.A(net1042),
    .B(_3245_),
    .Y(_0875_));
 sg13g2_nor4_1 _4658_ (.A(net1029),
    .B(_0829_),
    .C(_0873_),
    .D(_0875_),
    .Y(_0876_));
 sg13g2_a21oi_2 _4659_ (.B1(_0876_),
    .Y(_0877_),
    .A2(_0868_),
    .A1(net1029));
 sg13g2_o21ai_1 _4660_ (.B1(_0646_),
    .Y(_0878_),
    .A1(_3099_),
    .A2(_0844_));
 sg13g2_nand2b_1 _4661_ (.Y(_0879_),
    .B(_0878_),
    .A_N(_3288_));
 sg13g2_nand3_1 _4662_ (.B(_3288_),
    .C(_0849_),
    .A(net1043),
    .Y(_0880_));
 sg13g2_o21ai_1 _4663_ (.B1(_0879_),
    .Y(_0881_),
    .A1(_0870_),
    .A2(_0880_));
 sg13g2_nor3_1 _4664_ (.A(net1047),
    .B(net946),
    .C(_0831_),
    .Y(_0882_));
 sg13g2_o21ai_1 _4665_ (.B1(_3288_),
    .Y(_0883_),
    .A1(_3095_),
    .A2(_0691_));
 sg13g2_nor3_1 _4666_ (.A(_0836_),
    .B(_0882_),
    .C(_0883_),
    .Y(_0884_));
 sg13g2_nor3_2 _4667_ (.A(net946),
    .B(_0641_),
    .C(_0643_),
    .Y(_0885_));
 sg13g2_nor3_1 _4668_ (.A(_3243_),
    .B(_0733_),
    .C(_0885_),
    .Y(_0886_));
 sg13g2_nor4_1 _4669_ (.A(net1029),
    .B(_0874_),
    .C(_0884_),
    .D(_0886_),
    .Y(_0887_));
 sg13g2_a21oi_2 _4670_ (.B1(_0887_),
    .Y(_0888_),
    .A2(_0881_),
    .A1(net1029));
 sg13g2_a21o_2 _4671_ (.A2(_0888_),
    .A1(_0877_),
    .B1(net864),
    .X(_0889_));
 sg13g2_nand2b_1 _4672_ (.Y(_0890_),
    .B(_0877_),
    .A_N(_0888_));
 sg13g2_nand2_1 _4673_ (.Y(_0891_),
    .A(net864),
    .B(_0890_));
 sg13g2_nand2_1 _4674_ (.Y(_0892_),
    .A(_0889_),
    .B(_0891_));
 sg13g2_nand2_1 _4675_ (.Y(_0893_),
    .A(net866),
    .B(_0892_));
 sg13g2_xnor2_1 _4676_ (.Y(_0188_),
    .A(net271),
    .B(_0893_));
 sg13g2_nor2b_1 _4677_ (.A(_0042_),
    .B_N(_0889_),
    .Y(_0894_));
 sg13g2_inv_1 _4678_ (.Y(_0895_),
    .A(_0894_));
 sg13g2_xnor2_1 _4679_ (.Y(_0896_),
    .A(_0042_),
    .B(_0889_));
 sg13g2_nand3_1 _4680_ (.B(_0892_),
    .C(_0896_),
    .A(net271),
    .Y(_0897_));
 sg13g2_a21o_1 _4681_ (.A2(_0892_),
    .A1(\vgademo.soundtrack.pulse_osc_p[0] ),
    .B1(_0896_),
    .X(_0898_));
 sg13g2_nand3_1 _4682_ (.B(_0897_),
    .C(_0898_),
    .A(net866),
    .Y(_0899_));
 sg13g2_o21ai_1 _4683_ (.B1(_0899_),
    .Y(_0189_),
    .A1(_3184_),
    .A2(net866));
 sg13g2_nand2b_1 _4684_ (.Y(_0900_),
    .B(_0890_),
    .A_N(net864));
 sg13g2_or2_1 _4685_ (.X(_0901_),
    .B(_0888_),
    .A(_0877_));
 sg13g2_nand2_1 _4686_ (.Y(_0902_),
    .A(net864),
    .B(_0901_));
 sg13g2_nand2_1 _4687_ (.Y(_0903_),
    .A(_0900_),
    .B(_0902_));
 sg13g2_nor2_1 _4688_ (.A(_3185_),
    .B(_0903_),
    .Y(_0904_));
 sg13g2_xnor2_1 _4689_ (.Y(_0905_),
    .A(_3185_),
    .B(_0903_));
 sg13g2_a21oi_1 _4690_ (.A1(_0895_),
    .A2(_0897_),
    .Y(_0906_),
    .B1(_0905_));
 sg13g2_nand3_1 _4691_ (.B(_0897_),
    .C(_0905_),
    .A(_0895_),
    .Y(_0907_));
 sg13g2_nand3b_1 _4692_ (.B(_0907_),
    .C(net866),
    .Y(_0908_),
    .A_N(_0906_));
 sg13g2_o21ai_1 _4693_ (.B1(_0908_),
    .Y(_0190_),
    .A1(_3185_),
    .A2(net866));
 sg13g2_nand2b_1 _4694_ (.Y(_0909_),
    .B(_0888_),
    .A_N(_0877_));
 sg13g2_mux2_1 _4695_ (.A0(net864),
    .A1(_0891_),
    .S(_0909_),
    .X(_0910_));
 sg13g2_nand2_1 _4696_ (.Y(_0911_),
    .A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .B(_0910_));
 sg13g2_xnor2_1 _4697_ (.Y(_0912_),
    .A(_3186_),
    .B(_0910_));
 sg13g2_o21ai_1 _4698_ (.B1(_0912_),
    .Y(_0913_),
    .A1(_0904_),
    .A2(_0906_));
 sg13g2_or3_1 _4699_ (.A(_0904_),
    .B(_0906_),
    .C(_0912_),
    .X(_0914_));
 sg13g2_a21oi_1 _4700_ (.A1(_0913_),
    .A2(_0914_),
    .Y(_0915_),
    .B1(net865));
 sg13g2_a21oi_1 _4701_ (.A1(_3186_),
    .A2(net865),
    .Y(_0191_),
    .B1(_0915_));
 sg13g2_nand2_1 _4702_ (.Y(_0916_),
    .A(net254),
    .B(net865));
 sg13g2_and3_1 _4703_ (.X(_0917_),
    .A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .B(_0889_),
    .C(_0901_));
 sg13g2_a21oi_1 _4704_ (.A1(_0889_),
    .A2(_0901_),
    .Y(_0918_),
    .B1(\vgademo.soundtrack.pulse_osc_p[4] ));
 sg13g2_or2_1 _4705_ (.X(_0919_),
    .B(_0918_),
    .A(_0917_));
 sg13g2_a21oi_1 _4706_ (.A1(_0911_),
    .A2(_0913_),
    .Y(_0920_),
    .B1(_0919_));
 sg13g2_nand3_1 _4707_ (.B(_0913_),
    .C(_0919_),
    .A(_0911_),
    .Y(_0921_));
 sg13g2_nand2_1 _4708_ (.Y(_0922_),
    .A(net866),
    .B(_0921_));
 sg13g2_o21ai_1 _4709_ (.B1(_0916_),
    .Y(_0192_),
    .A1(_0920_),
    .A2(_0922_));
 sg13g2_nand2_1 _4710_ (.Y(_0923_),
    .A(net297),
    .B(net865));
 sg13g2_nand2_1 _4711_ (.Y(_0924_),
    .A(_0900_),
    .B(_0909_));
 sg13g2_nand3_1 _4712_ (.B(_0900_),
    .C(_0909_),
    .A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .Y(_0925_));
 sg13g2_xnor2_1 _4713_ (.Y(_0926_),
    .A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .B(_0924_));
 sg13g2_nor3_1 _4714_ (.A(_0917_),
    .B(_0920_),
    .C(_0926_),
    .Y(_0927_));
 sg13g2_o21ai_1 _4715_ (.B1(_0926_),
    .Y(_0928_),
    .A1(_0917_),
    .A2(_0920_));
 sg13g2_nand2_1 _4716_ (.Y(_0929_),
    .A(net866),
    .B(_0928_));
 sg13g2_o21ai_1 _4717_ (.B1(_0923_),
    .Y(_0193_),
    .A1(_0927_),
    .A2(_0929_));
 sg13g2_xnor2_1 _4718_ (.Y(_0930_),
    .A(\vgademo.soundtrack.pulse_osc_p[6] ),
    .B(net864));
 sg13g2_a21oi_1 _4719_ (.A1(_0925_),
    .A2(_0928_),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_and3_1 _4720_ (.X(_0932_),
    .A(_0925_),
    .B(_0928_),
    .C(_0930_));
 sg13g2_nor3_1 _4721_ (.A(net865),
    .B(_0931_),
    .C(_0932_),
    .Y(_0933_));
 sg13g2_a21o_1 _4722_ (.A2(net865),
    .A1(net352),
    .B1(_0933_),
    .X(_0194_));
 sg13g2_nor2_1 _4723_ (.A(net320),
    .B(net867),
    .Y(_0934_));
 sg13g2_a21o_1 _4724_ (.A2(_0859_),
    .A1(\vgademo.soundtrack.pulse_osc_p[6] ),
    .B1(_0931_),
    .X(_0935_));
 sg13g2_nor2_1 _4725_ (.A(_3187_),
    .B(_0859_),
    .Y(_0936_));
 sg13g2_xnor2_1 _4726_ (.Y(_0937_),
    .A(net320),
    .B(net864));
 sg13g2_xnor2_1 _4727_ (.Y(_0938_),
    .A(_0935_),
    .B(_0937_));
 sg13g2_a21oi_1 _4728_ (.A1(net867),
    .A2(_0938_),
    .Y(_0195_),
    .B1(_0934_));
 sg13g2_o21ai_1 _4729_ (.B1(net866),
    .Y(_0939_),
    .A1(_0935_),
    .A2(_0936_));
 sg13g2_a21oi_2 _4730_ (.B1(_0939_),
    .Y(_0940_),
    .A2(net864),
    .A1(_3187_));
 sg13g2_xor2_1 _4731_ (.B(_0940_),
    .A(net251),
    .X(_0196_));
 sg13g2_a21oi_1 _4732_ (.A1(\vgademo.soundtrack.pulse_osc_p[8] ),
    .A2(_0940_),
    .Y(_0941_),
    .B1(net233));
 sg13g2_and3_1 _4733_ (.X(_0942_),
    .A(\vgademo.soundtrack.pulse_osc_p[8] ),
    .B(net233),
    .C(_0940_));
 sg13g2_nor2_1 _4734_ (.A(net234),
    .B(_0942_),
    .Y(_0197_));
 sg13g2_and2_1 _4735_ (.A(net224),
    .B(_0942_),
    .X(_0943_));
 sg13g2_xor2_1 _4736_ (.B(_0942_),
    .A(net224),
    .X(_0198_));
 sg13g2_xor2_1 _4737_ (.B(_0943_),
    .A(net267),
    .X(_0199_));
 sg13g2_nand3_1 _4738_ (.B(net267),
    .C(_0943_),
    .A(net543),
    .Y(_0944_));
 sg13g2_a21o_1 _4739_ (.A2(_0943_),
    .A1(net267),
    .B1(net543),
    .X(_0945_));
 sg13g2_and2_1 _4740_ (.A(_0944_),
    .B(_0945_),
    .X(_0200_));
 sg13g2_xnor2_1 _4741_ (.Y(_0201_),
    .A(net243),
    .B(_0944_));
 sg13g2_nor3_1 _4742_ (.A(\vgademo.audio_kick_frames[0] ),
    .B(net847),
    .C(_0722_),
    .Y(_0946_));
 sg13g2_a21o_1 _4743_ (.A2(_0678_),
    .A1(net583),
    .B1(_0946_),
    .X(_0202_));
 sg13g2_nand2b_1 _4744_ (.Y(_0947_),
    .B(_0946_),
    .A_N(net368));
 sg13g2_o21ai_1 _4745_ (.B1(net368),
    .Y(_0948_),
    .A1(\vgademo.audio_kick_frames[0] ),
    .A2(net847));
 sg13g2_nand3_1 _4746_ (.B(net945),
    .C(_0698_),
    .A(net851),
    .Y(_0949_));
 sg13g2_nand3_1 _4747_ (.B(_0948_),
    .C(_0949_),
    .A(_0947_),
    .Y(_0203_));
 sg13g2_xor2_1 _4748_ (.B(_0947_),
    .A(net378),
    .X(_0950_));
 sg13g2_nand2_1 _4749_ (.Y(_0204_),
    .A(_0949_),
    .B(_0950_));
 sg13g2_nand2_1 _4750_ (.Y(_0951_),
    .A(_3268_),
    .B(_0690_));
 sg13g2_nor2_1 _4751_ (.A(_3268_),
    .B(_0731_),
    .Y(_0952_));
 sg13g2_a22oi_1 _4752_ (.Y(_0953_),
    .B1(_0952_),
    .B2(_3265_),
    .A2(_0951_),
    .A1(_0644_));
 sg13g2_o21ai_1 _4753_ (.B1(_0953_),
    .Y(_0954_),
    .A1(_0644_),
    .A2(_0804_));
 sg13g2_nor2_1 _4754_ (.A(_3274_),
    .B(_0639_),
    .Y(_0955_));
 sg13g2_a21oi_1 _4755_ (.A1(_3270_),
    .A2(_0731_),
    .Y(_0956_),
    .B1(_0955_));
 sg13g2_nand2b_1 _4756_ (.Y(_0957_),
    .B(_0837_),
    .A_N(_3282_));
 sg13g2_nor3_1 _4757_ (.A(_3251_),
    .B(_3283_),
    .C(net904),
    .Y(_0958_));
 sg13g2_nand3b_1 _4758_ (.B(net904),
    .C(_0854_),
    .Y(_0959_),
    .A_N(_0639_));
 sg13g2_a21oi_1 _4759_ (.A1(net1051),
    .A2(_3279_),
    .Y(_0960_),
    .B1(_0693_));
 sg13g2_o21ai_1 _4760_ (.B1(_0960_),
    .Y(_0961_),
    .A1(_3274_),
    .A2(_0639_));
 sg13g2_a21oi_1 _4761_ (.A1(net948),
    .A2(_3280_),
    .Y(_0962_),
    .B1(_3281_));
 sg13g2_a21oi_1 _4762_ (.A1(net904),
    .A2(_0961_),
    .Y(_0963_),
    .B1(_0647_));
 sg13g2_o21ai_1 _4763_ (.B1(_0963_),
    .Y(_0964_),
    .A1(net904),
    .A2(_0962_));
 sg13g2_a21oi_1 _4764_ (.A1(_0647_),
    .A2(_0954_),
    .Y(_0965_),
    .B1(_0652_));
 sg13g2_mux2_1 _4765_ (.A0(_0956_),
    .A1(_0957_),
    .S(net904),
    .X(_0966_));
 sg13g2_nor2_1 _4766_ (.A(_0647_),
    .B(_0958_),
    .Y(_0967_));
 sg13g2_a22oi_1 _4767_ (.Y(_0968_),
    .B1(_0967_),
    .B2(_0959_),
    .A2(_0966_),
    .A1(_0647_));
 sg13g2_a221oi_1 _4768_ (.B2(_0652_),
    .C1(_0651_),
    .B1(_0968_),
    .A1(_0964_),
    .Y(_0969_),
    .A2(_0965_));
 sg13g2_nor3_1 _4769_ (.A(_3095_),
    .B(net946),
    .C(_3267_),
    .Y(_0970_));
 sg13g2_o21ai_1 _4770_ (.B1(_0651_),
    .Y(_0971_),
    .A1(_0885_),
    .A2(_0962_));
 sg13g2_nor2_1 _4771_ (.A(_0629_),
    .B(_0969_),
    .Y(_0972_));
 sg13g2_o21ai_1 _4772_ (.B1(_0972_),
    .Y(_0973_),
    .A1(_0970_),
    .A2(_0971_));
 sg13g2_and2_2 _4773_ (.A(_0684_),
    .B(_0973_),
    .X(_0974_));
 sg13g2_o21ai_1 _4774_ (.B1(_0629_),
    .Y(_0975_),
    .A1(_3132_),
    .A2(_3330_));
 sg13g2_mux2_1 _4775_ (.A0(net226),
    .A1(_0975_),
    .S(_0974_),
    .X(_0205_));
 sg13g2_o21ai_1 _4776_ (.B1(_0629_),
    .Y(_0976_),
    .A1(_3330_),
    .A2(_3337_));
 sg13g2_mux2_1 _4777_ (.A0(net227),
    .A1(_0976_),
    .S(_0974_),
    .X(_0206_));
 sg13g2_xor2_1 _4778_ (.B(_3335_),
    .A(\vgademo.soundtrack.pulse_vol[2] ),
    .X(_0977_));
 sg13g2_o21ai_1 _4779_ (.B1(_0629_),
    .Y(_0978_),
    .A1(_3330_),
    .A2(_0977_));
 sg13g2_mux2_1 _4780_ (.A0(net242),
    .A1(_0978_),
    .S(_0974_),
    .X(_0207_));
 sg13g2_a21oi_1 _4781_ (.A1(net1010),
    .A2(_3335_),
    .Y(_0979_),
    .B1(net1009));
 sg13g2_o21ai_1 _4782_ (.B1(_0974_),
    .Y(_0980_),
    .A1(_0628_),
    .A2(_0979_));
 sg13g2_o21ai_1 _4783_ (.B1(_0980_),
    .Y(_0208_),
    .A1(_3079_),
    .A2(_0974_));
 sg13g2_nand2_1 _4784_ (.Y(_0981_),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B(net868));
 sg13g2_xnor2_1 _4785_ (.Y(_0209_),
    .A(net236),
    .B(_0981_));
 sg13g2_nand2_1 _4786_ (.Y(_0982_),
    .A(\vgademo.soundtrack.tri_osc_i[0] ),
    .B(net236));
 sg13g2_xor2_1 _4787_ (.B(\vgademo.soundtrack.tri_osc_p[1] ),
    .A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(_0983_));
 sg13g2_nor2b_1 _4788_ (.A(_0982_),
    .B_N(_0983_),
    .Y(_0984_));
 sg13g2_xor2_1 _4789_ (.B(_0983_),
    .A(_0982_),
    .X(_0985_));
 sg13g2_nand2_1 _4790_ (.Y(_0986_),
    .A(net330),
    .B(net865));
 sg13g2_o21ai_1 _4791_ (.B1(_0986_),
    .Y(_0210_),
    .A1(_0828_),
    .A2(_0985_));
 sg13g2_nor2_1 _4792_ (.A(net411),
    .B(net868),
    .Y(_0987_));
 sg13g2_a21oi_1 _4793_ (.A1(\vgademo.soundtrack.tri_osc_i[1] ),
    .A2(\vgademo.soundtrack.tri_osc_p[1] ),
    .Y(_0988_),
    .B1(_0984_));
 sg13g2_nand2_1 _4794_ (.Y(_0989_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_xnor2_1 _4795_ (.Y(_0990_),
    .A(\vgademo.soundtrack.tri_osc_i[2] ),
    .B(net411));
 sg13g2_or2_1 _4796_ (.X(_0991_),
    .B(_0990_),
    .A(_0988_));
 sg13g2_xnor2_1 _4797_ (.Y(_0992_),
    .A(_0988_),
    .B(_0990_));
 sg13g2_a21oi_1 _4798_ (.A1(net869),
    .A2(_0992_),
    .Y(_0211_),
    .B1(_0987_));
 sg13g2_nor2_1 _4799_ (.A(net400),
    .B(net868),
    .Y(_0993_));
 sg13g2_xnor2_1 _4800_ (.Y(_0994_),
    .A(\vgademo.soundtrack.tri_osc_i[3] ),
    .B(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_a21oi_1 _4801_ (.A1(_0989_),
    .A2(_0991_),
    .Y(_0995_),
    .B1(_0994_));
 sg13g2_nand3_1 _4802_ (.B(_0991_),
    .C(_0994_),
    .A(_0989_),
    .Y(_0996_));
 sg13g2_nand2b_1 _4803_ (.Y(_0997_),
    .B(_0996_),
    .A_N(_0995_));
 sg13g2_a21oi_1 _4804_ (.A1(net868),
    .A2(_0997_),
    .Y(_0212_),
    .B1(_0993_));
 sg13g2_nor2_1 _4805_ (.A(net380),
    .B(net868),
    .Y(_0998_));
 sg13g2_a21oi_1 _4806_ (.A1(\vgademo.soundtrack.tri_osc_i[3] ),
    .A2(\vgademo.soundtrack.tri_osc_p[3] ),
    .Y(_0999_),
    .B1(_0995_));
 sg13g2_nand2_1 _4807_ (.Y(_1000_),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_xnor2_1 _4808_ (.Y(_1001_),
    .A(\vgademo.soundtrack.tri_osc_i[4] ),
    .B(net380));
 sg13g2_xnor2_1 _4809_ (.Y(_1002_),
    .A(_0999_),
    .B(_1001_));
 sg13g2_a21oi_1 _4810_ (.A1(net868),
    .A2(_1002_),
    .Y(_0213_),
    .B1(_0998_));
 sg13g2_o21ai_1 _4811_ (.B1(_1000_),
    .Y(_1003_),
    .A1(_0999_),
    .A2(_1001_));
 sg13g2_nand2_1 _4812_ (.Y(_1004_),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .B(net422));
 sg13g2_xor2_1 _4813_ (.B(net422),
    .A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(_1005_));
 sg13g2_xnor2_1 _4814_ (.Y(_1006_),
    .A(_1003_),
    .B(_1005_));
 sg13g2_nor2_1 _4815_ (.A(net422),
    .B(net868),
    .Y(_1007_));
 sg13g2_a21oi_1 _4816_ (.A1(net868),
    .A2(_1006_),
    .Y(_0214_),
    .B1(_1007_));
 sg13g2_nor2_1 _4817_ (.A(_3129_),
    .B(_3181_),
    .Y(_1008_));
 sg13g2_xnor2_1 _4818_ (.Y(_1009_),
    .A(\vgademo.soundtrack.tri_osc_i[6] ),
    .B(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_o21ai_1 _4819_ (.B1(_1003_),
    .Y(_1010_),
    .A1(\vgademo.soundtrack.tri_osc_i[5] ),
    .A2(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_nand3_1 _4820_ (.B(_1009_),
    .C(_1010_),
    .A(_1004_),
    .Y(_1011_));
 sg13g2_a21oi_1 _4821_ (.A1(_1004_),
    .A2(_1010_),
    .Y(_1012_),
    .B1(_1009_));
 sg13g2_nand3b_1 _4822_ (.B(net869),
    .C(_1011_),
    .Y(_1013_),
    .A_N(_1012_));
 sg13g2_o21ai_1 _4823_ (.B1(_1013_),
    .Y(_0215_),
    .A1(_3181_),
    .A2(net869));
 sg13g2_nand2_1 _4824_ (.Y(_1014_),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .B(net424));
 sg13g2_xor2_1 _4825_ (.B(\vgademo.soundtrack.tri_osc_p[7] ),
    .A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(_1015_));
 sg13g2_or3_1 _4826_ (.A(_1008_),
    .B(_1012_),
    .C(_1015_),
    .X(_1016_));
 sg13g2_o21ai_1 _4827_ (.B1(_1015_),
    .Y(_1017_),
    .A1(_1008_),
    .A2(_1012_));
 sg13g2_nand3_1 _4828_ (.B(_1016_),
    .C(_1017_),
    .A(net869),
    .Y(_1018_));
 sg13g2_o21ai_1 _4829_ (.B1(_1018_),
    .Y(_0216_),
    .A1(_3180_),
    .A2(net869));
 sg13g2_xnor2_1 _4830_ (.Y(_1019_),
    .A(\vgademo.soundtrack.tri_osc_i[8] ),
    .B(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_and3_1 _4831_ (.X(_1020_),
    .A(_1014_),
    .B(_1017_),
    .C(_1019_));
 sg13g2_a21oi_1 _4832_ (.A1(_1014_),
    .A2(_1017_),
    .Y(_1021_),
    .B1(_1019_));
 sg13g2_nor3_1 _4833_ (.A(_0828_),
    .B(_1020_),
    .C(_1021_),
    .Y(_1022_));
 sg13g2_a21o_1 _4834_ (.A2(_0828_),
    .A1(net442),
    .B1(_1022_),
    .X(_0217_));
 sg13g2_a21oi_2 _4835_ (.B1(_1021_),
    .Y(_1023_),
    .A2(\vgademo.soundtrack.tri_osc_p[8] ),
    .A1(\vgademo.soundtrack.tri_osc_i[8] ));
 sg13g2_nand3_1 _4836_ (.B(net867),
    .C(_1023_),
    .A(net393),
    .Y(_1024_));
 sg13g2_nor3_2 _4837_ (.A(net393),
    .B(net865),
    .C(_1023_),
    .Y(_1025_));
 sg13g2_o21ai_1 _4838_ (.B1(_1024_),
    .Y(_1026_),
    .A1(\vgademo.soundtrack.tri_osc_p[9] ),
    .A2(net867));
 sg13g2_nor2_1 _4839_ (.A(net394),
    .B(_1026_),
    .Y(_0218_));
 sg13g2_and2_1 _4840_ (.A(net286),
    .B(_1025_),
    .X(_1027_));
 sg13g2_xor2_1 _4841_ (.B(_1025_),
    .A(net286),
    .X(_0219_));
 sg13g2_xor2_1 _4842_ (.B(_1027_),
    .A(net397),
    .X(_0220_));
 sg13g2_nand3_1 _4843_ (.B(net397),
    .C(_1027_),
    .A(net431),
    .Y(_1028_));
 sg13g2_a21o_1 _4844_ (.A2(_1027_),
    .A1(net397),
    .B1(net431),
    .X(_1029_));
 sg13g2_and2_1 _4845_ (.A(_1028_),
    .B(_1029_),
    .X(_0221_));
 sg13g2_nand4_1 _4846_ (.B(net431),
    .C(net397),
    .A(net318),
    .Y(_1030_),
    .D(_1027_));
 sg13g2_xnor2_1 _4847_ (.Y(_0222_),
    .A(net318),
    .B(_1028_));
 sg13g2_xnor2_1 _4848_ (.Y(_0223_),
    .A(net369),
    .B(_1030_));
 sg13g2_o21ai_1 _4849_ (.B1(net1006),
    .Y(_1031_),
    .A1(_3179_),
    .A2(_1030_));
 sg13g2_o21ai_1 _4850_ (.B1(_1031_),
    .Y(_0224_),
    .A1(_0546_),
    .A2(_1030_));
 sg13g2_nor2_2 _4851_ (.A(net982),
    .B(net985),
    .Y(_1032_));
 sg13g2_or2_1 _4852_ (.X(_1033_),
    .B(net985),
    .A(net983));
 sg13g2_nor2_2 _4853_ (.A(net985),
    .B(net988),
    .Y(_1034_));
 sg13g2_nor3_2 _4854_ (.A(net982),
    .B(net984),
    .C(net989),
    .Y(_1035_));
 sg13g2_or3_1 _4855_ (.A(net982),
    .B(net985),
    .C(net988),
    .X(_1036_));
 sg13g2_nor2_2 _4856_ (.A(net976),
    .B(net979),
    .Y(_1037_));
 sg13g2_nor2_1 _4857_ (.A(net979),
    .B(net982),
    .Y(_1038_));
 sg13g2_nand2_1 _4858_ (.Y(_1039_),
    .A(_1032_),
    .B(_1037_));
 sg13g2_nand3_1 _4859_ (.B(_1035_),
    .C(_1037_),
    .A(net974),
    .Y(_1040_));
 sg13g2_nand2_1 _4860_ (.Y(_1041_),
    .A(\vgademo.a_scrolly[11] ),
    .B(net971));
 sg13g2_nor2_1 _4861_ (.A(_0065_),
    .B(_1041_),
    .Y(_1042_));
 sg13g2_nor2_2 _4862_ (.A(\vgademo.a_scrolly[12] ),
    .B(\vgademo.a_scrolly[13] ),
    .Y(_1043_));
 sg13g2_inv_1 _4863_ (.Y(_1044_),
    .A(_1043_));
 sg13g2_and2_1 _4864_ (.A(net992),
    .B(_1035_),
    .X(_1045_));
 sg13g2_nand2_1 _4865_ (.Y(_1046_),
    .A(net992),
    .B(_1035_));
 sg13g2_and2_1 _4866_ (.A(\vgademo.a_scrolly[10] ),
    .B(net974),
    .X(_1047_));
 sg13g2_nand2_2 _4867_ (.Y(_1048_),
    .A(net971),
    .B(net972));
 sg13g2_nor2b_1 _4868_ (.A(\vgademo.a_scrolly[12] ),
    .B_N(\vgademo.a_scrolly[11] ),
    .Y(_1049_));
 sg13g2_and4_1 _4869_ (.A(_0066_),
    .B(_1037_),
    .C(_1047_),
    .D(_1049_),
    .X(_1050_));
 sg13g2_a22oi_1 _4870_ (.Y(_1051_),
    .B1(_1045_),
    .B2(_1050_),
    .A2(_1042_),
    .A1(_1040_));
 sg13g2_a221oi_1 _4871_ (.B2(_1050_),
    .C1(_1044_),
    .B1(_1045_),
    .A1(_1040_),
    .Y(_1052_),
    .A2(_1042_));
 sg13g2_nand2_2 _4872_ (.Y(_1053_),
    .A(_1043_),
    .B(_1051_));
 sg13g2_nand2_2 _4873_ (.Y(_1054_),
    .A(net993),
    .B(net576));
 sg13g2_and3_1 _4874_ (.X(_1055_),
    .A(net992),
    .B(net984),
    .C(net988));
 sg13g2_nand3_1 _4875_ (.B(net984),
    .C(net988),
    .A(net992),
    .Y(_1056_));
 sg13g2_nor2_1 _4876_ (.A(net981),
    .B(_1055_),
    .Y(_1057_));
 sg13g2_nand2_1 _4877_ (.Y(_1058_),
    .A(_3118_),
    .B(_1056_));
 sg13g2_nor2b_1 _4878_ (.A(net973),
    .B_N(net970),
    .Y(_1059_));
 sg13g2_nand2b_1 _4879_ (.Y(_1060_),
    .B(net970),
    .A_N(net972));
 sg13g2_nand2b_1 _4880_ (.Y(_1061_),
    .B(net979),
    .A_N(net976));
 sg13g2_or2_1 _4881_ (.X(_1062_),
    .B(_1061_),
    .A(_1060_));
 sg13g2_o21ai_1 _4882_ (.B1(net971),
    .Y(_1063_),
    .A1(net972),
    .A2(net977));
 sg13g2_o21ai_1 _4883_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_1057_),
    .A2(_1062_));
 sg13g2_a21oi_1 _4884_ (.A1(_1049_),
    .A2(_1064_),
    .Y(_1065_),
    .B1(_3120_));
 sg13g2_a21o_2 _4885_ (.A2(_1064_),
    .A1(_1049_),
    .B1(_3120_),
    .X(_1066_));
 sg13g2_nor2_1 _4886_ (.A(_0066_),
    .B(_1065_),
    .Y(_1067_));
 sg13g2_nand2_1 _4887_ (.Y(_1068_),
    .A(_3119_),
    .B(_1066_));
 sg13g2_nand2_2 _4888_ (.Y(_1069_),
    .A(\vgademo.a_scrolly[12] ),
    .B(\vgademo.a_scrolly[13] ));
 sg13g2_and2_1 _4889_ (.A(_1037_),
    .B(_1059_),
    .X(_1070_));
 sg13g2_nand3_1 _4890_ (.B(_1037_),
    .C(_1059_),
    .A(_3118_),
    .Y(_1071_));
 sg13g2_nand2_1 _4891_ (.Y(_1072_),
    .A(net970),
    .B(_1071_));
 sg13g2_a221oi_1 _4892_ (.B2(net970),
    .C1(\vgademo.a_scrolly[11] ),
    .B1(_1071_),
    .A1(_1058_),
    .Y(_1073_),
    .A2(_1070_));
 sg13g2_or2_1 _4893_ (.X(_1074_),
    .B(_1073_),
    .A(_1069_));
 sg13g2_and3_1 _4894_ (.X(_1075_),
    .A(_3119_),
    .B(_1066_),
    .C(_1074_));
 sg13g2_nand3_1 _4895_ (.B(_1066_),
    .C(_1074_),
    .A(_3119_),
    .Y(_1076_));
 sg13g2_nor2_1 _4896_ (.A(_3117_),
    .B(_1035_),
    .Y(_1077_));
 sg13g2_a21oi_2 _4897_ (.B1(net977),
    .Y(_1078_),
    .A2(_1036_),
    .A1(net980));
 sg13g2_nor2b_1 _4898_ (.A(_1078_),
    .B_N(net975),
    .Y(_1079_));
 sg13g2_nor2_1 _4899_ (.A(_1048_),
    .B(_1078_),
    .Y(_1080_));
 sg13g2_nand2_2 _4900_ (.Y(_1081_),
    .A(_3113_),
    .B(_1043_));
 sg13g2_nand3b_1 _4901_ (.B(_3113_),
    .C(_0066_),
    .Y(_1082_),
    .A_N(\vgademo.a_scrolly[12] ));
 sg13g2_inv_1 _4902_ (.Y(_1083_),
    .A(_1082_));
 sg13g2_nor4_1 _4903_ (.A(_1046_),
    .B(_1048_),
    .C(_1061_),
    .D(_1082_),
    .Y(_1084_));
 sg13g2_nor3_2 _4904_ (.A(_1080_),
    .B(_1081_),
    .C(_1084_),
    .Y(_1085_));
 sg13g2_nor2b_1 _4905_ (.A(_1085_),
    .B_N(_0064_),
    .Y(_1086_));
 sg13g2_o21ai_1 _4906_ (.B1(_1086_),
    .Y(_1087_),
    .A1(net934),
    .A2(_1075_));
 sg13g2_nand2_1 _4907_ (.Y(_1088_),
    .A(\vgademo.bayer_j[0] ),
    .B(_1087_));
 sg13g2_xnor2_1 _4908_ (.Y(_1089_),
    .A(_3101_),
    .B(_1087_));
 sg13g2_nand2b_1 _4909_ (.Y(_1090_),
    .B(_1089_),
    .A_N(\vgademo.audio_kick_frames[0] ));
 sg13g2_xor2_1 _4910_ (.B(_1089_),
    .A(\vgademo.audio_kick_frames[0] ),
    .X(_1091_));
 sg13g2_nor2_1 _4911_ (.A(net937),
    .B(_1091_),
    .Y(_1092_));
 sg13g2_a21o_1 _4912_ (.A2(_0660_),
    .A1(net465),
    .B1(_1092_),
    .X(_0225_));
 sg13g2_nand2_1 _4913_ (.Y(_1093_),
    .A(_1088_),
    .B(_1090_));
 sg13g2_mux2_1 _4914_ (.A0(net990),
    .A1(_0069_),
    .S(net934),
    .X(_1094_));
 sg13g2_nor2_1 _4915_ (.A(_1085_),
    .B(_1094_),
    .Y(_1095_));
 sg13g2_o21ai_1 _4916_ (.B1(_1095_),
    .Y(_1096_),
    .A1(net934),
    .A2(_1075_));
 sg13g2_xnor2_1 _4917_ (.Y(_1097_),
    .A(_3100_),
    .B(_1096_));
 sg13g2_xor2_1 _4918_ (.B(_1097_),
    .A(_0068_),
    .X(_1098_));
 sg13g2_nand2_1 _4919_ (.Y(_1099_),
    .A(_1093_),
    .B(_1098_));
 sg13g2_xnor2_1 _4920_ (.Y(_1100_),
    .A(_1093_),
    .B(_1098_));
 sg13g2_nor2_1 _4921_ (.A(net937),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_a21o_1 _4922_ (.A2(_0660_),
    .A1(net405),
    .B1(_1101_),
    .X(_0226_));
 sg13g2_a22oi_1 _4923_ (.Y(_1102_),
    .B1(_1097_),
    .B2(_0068_),
    .A2(_1096_),
    .A1(_3121_));
 sg13g2_nand2b_1 _4924_ (.Y(_1103_),
    .B(net934),
    .A_N(net988));
 sg13g2_a221oi_1 _4925_ (.B2(net985),
    .C1(_1085_),
    .B1(_1103_),
    .A1(_1034_),
    .Y(_1104_),
    .A2(net933));
 sg13g2_o21ai_1 _4926_ (.B1(_1104_),
    .Y(_1105_),
    .A1(net933),
    .A2(_1075_));
 sg13g2_xor2_1 _4927_ (.B(_1105_),
    .A(_0071_),
    .X(_1106_));
 sg13g2_nor2b_1 _4928_ (.A(_1102_),
    .B_N(_1106_),
    .Y(_1107_));
 sg13g2_xnor2_1 _4929_ (.Y(_1108_),
    .A(_1102_),
    .B(_1106_));
 sg13g2_xnor2_1 _4930_ (.Y(_1109_),
    .A(_0060_),
    .B(_1108_));
 sg13g2_nor2_1 _4931_ (.A(_1099_),
    .B(_1109_),
    .Y(_1110_));
 sg13g2_xor2_1 _4932_ (.B(_1109_),
    .A(_1099_),
    .X(_1111_));
 sg13g2_mux2_1 _4933_ (.A0(_1111_),
    .A1(net364),
    .S(net937),
    .X(_0227_));
 sg13g2_nor2_1 _4934_ (.A(net361),
    .B(net935),
    .Y(_1112_));
 sg13g2_a21o_1 _4935_ (.A2(_1108_),
    .A1(_0060_),
    .B1(_1107_),
    .X(_1113_));
 sg13g2_nand2b_1 _4936_ (.Y(_1114_),
    .B(_0075_),
    .A_N(net933));
 sg13g2_o21ai_1 _4937_ (.B1(net981),
    .Y(_1115_),
    .A1(net984),
    .A2(net988));
 sg13g2_inv_1 _4938_ (.Y(_1116_),
    .A(_1115_));
 sg13g2_o21ai_1 _4939_ (.B1(net933),
    .Y(_1117_),
    .A1(_1035_),
    .A2(_1116_));
 sg13g2_nand3b_1 _4940_ (.B(_1114_),
    .C(_1117_),
    .Y(_1118_),
    .A_N(_1085_));
 sg13g2_a21oi_2 _4941_ (.B1(_1118_),
    .Y(_1119_),
    .A2(_1076_),
    .A1(_1053_));
 sg13g2_nand2_1 _4942_ (.Y(_1120_),
    .A(_0074_),
    .B(_1119_));
 sg13g2_xor2_1 _4943_ (.B(_1119_),
    .A(_0074_),
    .X(_1121_));
 sg13g2_nor2_1 _4944_ (.A(net968),
    .B(_1105_),
    .Y(_1122_));
 sg13g2_nor2_1 _4945_ (.A(_1121_),
    .B(_1122_),
    .Y(_1123_));
 sg13g2_xor2_1 _4946_ (.B(_1122_),
    .A(_1121_),
    .X(_1124_));
 sg13g2_xnor2_1 _4947_ (.Y(_1125_),
    .A(_1113_),
    .B(_1124_));
 sg13g2_nor3_1 _4948_ (.A(_1099_),
    .B(_1109_),
    .C(_1125_),
    .Y(_1126_));
 sg13g2_xor2_1 _4949_ (.B(_1125_),
    .A(_1110_),
    .X(_1127_));
 sg13g2_a21oi_1 _4950_ (.A1(net935),
    .A2(_1127_),
    .Y(_0228_),
    .B1(_1112_));
 sg13g2_a21oi_1 _4951_ (.A1(_1113_),
    .A2(_1124_),
    .Y(_1128_),
    .B1(_1126_));
 sg13g2_nor3_1 _4952_ (.A(_0066_),
    .B(net933),
    .C(_1065_),
    .Y(_1129_));
 sg13g2_nand2_1 _4953_ (.Y(_1130_),
    .A(net979),
    .B(net981));
 sg13g2_nand3b_1 _4954_ (.B(_1074_),
    .C(_1130_),
    .Y(_1131_),
    .A_N(_1038_));
 sg13g2_nand2_1 _4955_ (.Y(_1132_),
    .A(_0069_),
    .B(_1032_));
 sg13g2_xnor2_1 _4956_ (.Y(_1133_),
    .A(_0078_),
    .B(_1132_));
 sg13g2_a221oi_1 _4957_ (.B2(net934),
    .C1(_1085_),
    .B1(_1133_),
    .A1(_1129_),
    .Y(_1134_),
    .A2(_1131_));
 sg13g2_nand2_1 _4958_ (.Y(_1135_),
    .A(_0077_),
    .B(_1134_));
 sg13g2_xnor2_1 _4959_ (.Y(_1136_),
    .A(_0077_),
    .B(_1134_));
 sg13g2_nand2_1 _4960_ (.Y(_1137_),
    .A(_1120_),
    .B(_1136_));
 sg13g2_xor2_1 _4961_ (.B(_1136_),
    .A(_1120_),
    .X(_1138_));
 sg13g2_xnor2_1 _4962_ (.Y(_1139_),
    .A(_1123_),
    .B(_1138_));
 sg13g2_nor2_1 _4963_ (.A(_1128_),
    .B(_1139_),
    .Y(_1140_));
 sg13g2_xor2_1 _4964_ (.B(_1139_),
    .A(_1128_),
    .X(_1141_));
 sg13g2_mux2_1 _4965_ (.A0(_1141_),
    .A1(net347),
    .S(net937),
    .X(_0229_));
 sg13g2_a21oi_1 _4966_ (.A1(_1123_),
    .A2(_1138_),
    .Y(_1142_),
    .B1(_1140_));
 sg13g2_xor2_1 _4967_ (.B(_1038_),
    .A(_0080_),
    .X(_1143_));
 sg13g2_o21ai_1 _4968_ (.B1(_1143_),
    .Y(_1144_),
    .A1(_1069_),
    .A2(_1073_));
 sg13g2_nand4_1 _4969_ (.B(_1053_),
    .C(_1066_),
    .A(_3119_),
    .Y(_1145_),
    .D(_1144_));
 sg13g2_a21oi_2 _4970_ (.B1(_3117_),
    .Y(_1146_),
    .A2(_1032_),
    .A1(_0069_));
 sg13g2_xnor2_1 _4971_ (.Y(_1147_),
    .A(_0080_),
    .B(_1146_));
 sg13g2_nand2_1 _4972_ (.Y(_1148_),
    .A(net934),
    .B(_1147_));
 sg13g2_a21oi_2 _4973_ (.B1(_1085_),
    .Y(_1149_),
    .A2(_1148_),
    .A1(_1145_));
 sg13g2_and2_1 _4974_ (.A(net965),
    .B(_1149_),
    .X(_1150_));
 sg13g2_or2_1 _4975_ (.X(_1151_),
    .B(_1149_),
    .A(net966));
 sg13g2_xnor2_1 _4976_ (.Y(_1152_),
    .A(net966),
    .B(_1149_));
 sg13g2_or2_1 _4977_ (.X(_1153_),
    .B(_1152_),
    .A(_1135_));
 sg13g2_xnor2_1 _4978_ (.Y(_1154_),
    .A(_1135_),
    .B(_1152_));
 sg13g2_nand2b_1 _4979_ (.Y(_1155_),
    .B(_1154_),
    .A_N(_1137_));
 sg13g2_xor2_1 _4980_ (.B(_1154_),
    .A(_1137_),
    .X(_1156_));
 sg13g2_xor2_1 _4981_ (.B(_1156_),
    .A(_1142_),
    .X(_1157_));
 sg13g2_mux2_1 _4982_ (.A0(_1157_),
    .A1(net464),
    .S(_0658_),
    .X(_0230_));
 sg13g2_nor2_1 _4983_ (.A(net342),
    .B(net935),
    .Y(_1158_));
 sg13g2_o21ai_1 _4984_ (.B1(_1155_),
    .Y(_1159_),
    .A1(_1142_),
    .A2(_1156_));
 sg13g2_nand2b_1 _4985_ (.Y(_1160_),
    .B(_0063_),
    .A_N(_1149_));
 sg13g2_nand2_1 _4986_ (.Y(_1161_),
    .A(_0075_),
    .B(_1037_));
 sg13g2_nand3b_1 _4987_ (.B(_0075_),
    .C(_1037_),
    .Y(_1162_),
    .A_N(net972));
 sg13g2_xor2_1 _4988_ (.B(_1161_),
    .A(net972),
    .X(_1163_));
 sg13g2_o21ai_1 _4989_ (.B1(_1163_),
    .Y(_1164_),
    .A1(_1069_),
    .A2(_1073_));
 sg13g2_nand4_1 _4990_ (.B(_1053_),
    .C(_1066_),
    .A(_3119_),
    .Y(_1165_),
    .D(_1164_));
 sg13g2_a21oi_1 _4991_ (.A1(net976),
    .A2(_1146_),
    .Y(_1166_),
    .B1(net974));
 sg13g2_and3_1 _4992_ (.X(_1167_),
    .A(net974),
    .B(net976),
    .C(_1146_));
 sg13g2_o21ai_1 _4993_ (.B1(net933),
    .Y(_1168_),
    .A1(_1166_),
    .A2(_1167_));
 sg13g2_a21oi_2 _4994_ (.B1(_1085_),
    .Y(_1169_),
    .A2(_1168_),
    .A1(_1165_));
 sg13g2_xnor2_1 _4995_ (.Y(_1170_),
    .A(net964),
    .B(_1169_));
 sg13g2_nand2_1 _4996_ (.Y(_1171_),
    .A(_1160_),
    .B(_1170_));
 sg13g2_xor2_1 _4997_ (.B(_1170_),
    .A(_1160_),
    .X(_1172_));
 sg13g2_xnor2_1 _4998_ (.Y(_1173_),
    .A(_1153_),
    .B(_1172_));
 sg13g2_nor2b_1 _4999_ (.A(_1173_),
    .B_N(_1159_),
    .Y(_1174_));
 sg13g2_xor2_1 _5000_ (.B(_1173_),
    .A(_1159_),
    .X(_1175_));
 sg13g2_a21oi_1 _5001_ (.A1(net935),
    .A2(_1175_),
    .Y(_0231_),
    .B1(_1158_));
 sg13g2_a21o_1 _5002_ (.A2(_1172_),
    .A1(_1153_),
    .B1(_1174_),
    .X(_1176_));
 sg13g2_xor2_1 _5003_ (.B(_1162_),
    .A(_0016_),
    .X(_1177_));
 sg13g2_o21ai_1 _5004_ (.B1(_1177_),
    .Y(_1178_),
    .A1(_1069_),
    .A2(_1073_));
 sg13g2_nand3_1 _5005_ (.B(_1066_),
    .C(_1178_),
    .A(_3119_),
    .Y(_1179_));
 sg13g2_a21oi_1 _5006_ (.A1(net977),
    .A2(_1146_),
    .Y(_1180_),
    .B1(_3115_));
 sg13g2_xnor2_1 _5007_ (.Y(_1181_),
    .A(_3114_),
    .B(_1180_));
 sg13g2_a21o_1 _5008_ (.A2(_1181_),
    .A1(net933),
    .B1(_1085_),
    .X(_1182_));
 sg13g2_a21o_2 _5009_ (.A2(_1179_),
    .A1(_1053_),
    .B1(_1182_),
    .X(_1183_));
 sg13g2_nand2_1 _5010_ (.Y(_1184_),
    .A(_0015_),
    .B(_1183_));
 sg13g2_xor2_1 _5011_ (.B(_1183_),
    .A(_0015_),
    .X(_1185_));
 sg13g2_nor2_2 _5012_ (.A(_3123_),
    .B(_1169_),
    .Y(_1186_));
 sg13g2_nor2_1 _5013_ (.A(_1185_),
    .B(_1186_),
    .Y(_1187_));
 sg13g2_xnor2_1 _5014_ (.Y(_1188_),
    .A(_1185_),
    .B(_1186_));
 sg13g2_nor2_1 _5015_ (.A(_1171_),
    .B(_1188_),
    .Y(_1189_));
 sg13g2_xor2_1 _5016_ (.B(_1188_),
    .A(_1171_),
    .X(_1190_));
 sg13g2_xor2_1 _5017_ (.B(_1190_),
    .A(_1176_),
    .X(_1191_));
 sg13g2_mux2_1 _5018_ (.A0(_1191_),
    .A1(net339),
    .S(net937),
    .X(_0232_));
 sg13g2_a21oi_1 _5019_ (.A1(_1176_),
    .A2(_1190_),
    .Y(_1192_),
    .B1(_1189_));
 sg13g2_xor2_1 _5020_ (.B(_1072_),
    .A(_0020_),
    .X(_1193_));
 sg13g2_nand2_1 _5021_ (.Y(_1194_),
    .A(_1053_),
    .B(_1193_));
 sg13g2_o21ai_1 _5022_ (.B1(net933),
    .Y(_1195_),
    .A1(_1041_),
    .A2(_1166_));
 sg13g2_o21ai_1 _5023_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_1076_),
    .A2(_1194_));
 sg13g2_xnor2_1 _5024_ (.Y(_1197_),
    .A(_0019_),
    .B(_1196_));
 sg13g2_xnor2_1 _5025_ (.Y(_1198_),
    .A(_1184_),
    .B(_1197_));
 sg13g2_xnor2_1 _5026_ (.Y(_1199_),
    .A(_1187_),
    .B(_1198_));
 sg13g2_xnor2_1 _5027_ (.Y(_1200_),
    .A(_1192_),
    .B(_1199_));
 sg13g2_and2_1 _5028_ (.A(net935),
    .B(_1200_),
    .X(_1201_));
 sg13g2_a21o_1 _5029_ (.A2(net937),
    .A1(net307),
    .B1(_1201_),
    .X(_0233_));
 sg13g2_nor2_2 _5030_ (.A(\vgademo.a_scrolly[10] ),
    .B(net974),
    .Y(_1202_));
 sg13g2_nor2_1 _5031_ (.A(net992),
    .B(net988),
    .Y(_1203_));
 sg13g2_or2_2 _5032_ (.X(_1204_),
    .B(net988),
    .A(net991));
 sg13g2_o21ai_1 _5033_ (.B1(net982),
    .Y(_1205_),
    .A1(net985),
    .A2(_1204_));
 sg13g2_nand4_1 _5034_ (.B(_1083_),
    .C(_1202_),
    .A(_1037_),
    .Y(_1206_),
    .D(_1205_));
 sg13g2_nand4_1 _5035_ (.B(_3255_),
    .C(_0875_),
    .A(_3253_),
    .Y(_1207_),
    .D(_1206_));
 sg13g2_o21ai_1 _5036_ (.B1(net912),
    .Y(_1208_),
    .A1(\vgademo.audio_songpos[7] ),
    .A2(_1207_));
 sg13g2_nor2b_1 _5037_ (.A(net994),
    .B_N(_1208_),
    .Y(_1209_));
 sg13g2_a21oi_1 _5038_ (.A1(net994),
    .A2(net912),
    .Y(_0234_),
    .B1(_1209_));
 sg13g2_nand2_1 _5039_ (.Y(_1210_),
    .A(net990),
    .B(net908));
 sg13g2_nand2_1 _5040_ (.Y(_1211_),
    .A(_1054_),
    .B(_1204_));
 sg13g2_o21ai_1 _5041_ (.B1(_1210_),
    .Y(_0235_),
    .A1(_1208_),
    .A2(_1211_));
 sg13g2_nand2_1 _5042_ (.Y(_1212_),
    .A(net986),
    .B(net908));
 sg13g2_xor2_1 _5043_ (.B(_1054_),
    .A(net986),
    .X(_1213_));
 sg13g2_o21ai_1 _5044_ (.B1(_1212_),
    .Y(_0236_),
    .A1(net881),
    .A2(_1213_));
 sg13g2_nand2_1 _5045_ (.Y(_1214_),
    .A(net981),
    .B(net905));
 sg13g2_xnor2_1 _5046_ (.Y(_1215_),
    .A(net595),
    .B(_1056_));
 sg13g2_o21ai_1 _5047_ (.B1(_1214_),
    .Y(_0237_),
    .A1(net881),
    .A2(_1215_));
 sg13g2_nand2_1 _5048_ (.Y(_1216_),
    .A(net980),
    .B(net905));
 sg13g2_nand2_2 _5049_ (.Y(_1217_),
    .A(net983),
    .B(net986));
 sg13g2_xor2_1 _5050_ (.B(_1217_),
    .A(_0078_),
    .X(_1218_));
 sg13g2_nand2_1 _5051_ (.Y(_1219_),
    .A(_0078_),
    .B(_1054_));
 sg13g2_o21ai_1 _5052_ (.B1(_1219_),
    .Y(_1220_),
    .A1(_1054_),
    .A2(_1218_));
 sg13g2_o21ai_1 _5053_ (.B1(_1216_),
    .Y(_0238_),
    .A1(_1208_),
    .A2(_1220_));
 sg13g2_nand2_1 _5054_ (.Y(_1221_),
    .A(net977),
    .B(net905));
 sg13g2_nor3_1 _5055_ (.A(_0078_),
    .B(_1054_),
    .C(_1217_),
    .Y(_1222_));
 sg13g2_xor2_1 _5056_ (.B(_1222_),
    .A(net585),
    .X(_1223_));
 sg13g2_o21ai_1 _5057_ (.B1(_1221_),
    .Y(_0239_),
    .A1(net881),
    .A2(net586));
 sg13g2_nand2_1 _5058_ (.Y(_1224_),
    .A(net972),
    .B(net905));
 sg13g2_nand4_1 _5059_ (.B(net979),
    .C(net981),
    .A(net976),
    .Y(_1225_),
    .D(_1055_));
 sg13g2_nor2_1 _5060_ (.A(_0065_),
    .B(_1225_),
    .Y(_1226_));
 sg13g2_xnor2_1 _5061_ (.Y(_1227_),
    .A(net476),
    .B(_1225_));
 sg13g2_o21ai_1 _5062_ (.B1(_1224_),
    .Y(_0240_),
    .A1(net881),
    .A2(_1227_));
 sg13g2_nand2_1 _5063_ (.Y(_1228_),
    .A(net970),
    .B(net905));
 sg13g2_xor2_1 _5064_ (.B(_1226_),
    .A(net453),
    .X(_1229_));
 sg13g2_o21ai_1 _5065_ (.B1(_1228_),
    .Y(_0241_),
    .A1(net881),
    .A2(net454));
 sg13g2_nand2_1 _5066_ (.Y(_1230_),
    .A(net527),
    .B(net905));
 sg13g2_nor2_1 _5067_ (.A(_1048_),
    .B(_1225_),
    .Y(_1231_));
 sg13g2_nor3_1 _5068_ (.A(_0020_),
    .B(_1048_),
    .C(_1225_),
    .Y(_1232_));
 sg13g2_xor2_1 _5069_ (.B(_1231_),
    .A(_0020_),
    .X(_1233_));
 sg13g2_o21ai_1 _5070_ (.B1(_1230_),
    .Y(_0242_),
    .A1(net881),
    .A2(_1233_));
 sg13g2_nand2_1 _5071_ (.Y(_1234_),
    .A(\vgademo.a_scrolly[12] ),
    .B(net905));
 sg13g2_xnor2_1 _5072_ (.Y(_1235_),
    .A(_3120_),
    .B(_1232_));
 sg13g2_o21ai_1 _5073_ (.B1(_1234_),
    .Y(_0243_),
    .A1(net881),
    .A2(net518));
 sg13g2_nand2_1 _5074_ (.Y(_1236_),
    .A(net441),
    .B(net905));
 sg13g2_and3_1 _5075_ (.X(_1237_),
    .A(\vgademo.a_scrolly[12] ),
    .B(\vgademo.a_scrolly[11] ),
    .C(_1231_));
 sg13g2_xnor2_1 _5076_ (.Y(_1238_),
    .A(_3119_),
    .B(_1237_));
 sg13g2_o21ai_1 _5077_ (.B1(_1236_),
    .Y(_0244_),
    .A1(net881),
    .A2(_1238_));
 sg13g2_nand2_2 _5078_ (.Y(_1239_),
    .A(net941),
    .B(_0585_));
 sg13g2_a21oi_1 _5079_ (.A1(_3198_),
    .A2(_0585_),
    .Y(_1240_),
    .B1(net969));
 sg13g2_nand2_1 _5080_ (.Y(_1241_),
    .A(net969),
    .B(_3198_));
 sg13g2_nor2b_1 _5081_ (.A(_1240_),
    .B_N(_1241_),
    .Y(_0245_));
 sg13g2_xnor2_1 _5082_ (.Y(_0246_),
    .A(net415),
    .B(_1241_));
 sg13g2_nand2_1 _5083_ (.Y(_1242_),
    .A(net968),
    .B(net938));
 sg13g2_nand2_2 _5084_ (.Y(_1243_),
    .A(net415),
    .B(net969));
 sg13g2_nor2_1 _5085_ (.A(_0071_),
    .B(_1243_),
    .Y(_1244_));
 sg13g2_xnor2_1 _5086_ (.Y(_1245_),
    .A(_0071_),
    .B(_1243_));
 sg13g2_o21ai_1 _5087_ (.B1(_1242_),
    .Y(_0247_),
    .A1(_1239_),
    .A2(net416));
 sg13g2_nand2_1 _5088_ (.Y(_1246_),
    .A(net460),
    .B(net938));
 sg13g2_xor2_1 _5089_ (.B(_1244_),
    .A(_0074_),
    .X(_1247_));
 sg13g2_o21ai_1 _5090_ (.B1(_1246_),
    .Y(_0248_),
    .A1(_1239_),
    .A2(_1247_));
 sg13g2_nand2_1 _5091_ (.Y(_1248_),
    .A(net967),
    .B(net938));
 sg13g2_nor2_1 _5092_ (.A(_0582_),
    .B(_1243_),
    .Y(_1249_));
 sg13g2_nor3_1 _5093_ (.A(_0077_),
    .B(_0582_),
    .C(_1243_),
    .Y(_1250_));
 sg13g2_xor2_1 _5094_ (.B(_1249_),
    .A(net563),
    .X(_1251_));
 sg13g2_o21ai_1 _5095_ (.B1(_1248_),
    .Y(_0249_),
    .A1(_1239_),
    .A2(_1251_));
 sg13g2_nand2_1 _5096_ (.Y(_1252_),
    .A(net965),
    .B(net938));
 sg13g2_xor2_1 _5097_ (.B(_1250_),
    .A(net494),
    .X(_1253_));
 sg13g2_o21ai_1 _5098_ (.B1(_1252_),
    .Y(_0250_),
    .A1(_1239_),
    .A2(net495));
 sg13g2_nand2_1 _5099_ (.Y(_1254_),
    .A(net964),
    .B(net939));
 sg13g2_nand3_1 _5100_ (.B(\vgademo.v_count[4] ),
    .C(_1249_),
    .A(net965),
    .Y(_1255_));
 sg13g2_nor2_1 _5101_ (.A(_0017_),
    .B(_1255_),
    .Y(_1256_));
 sg13g2_xnor2_1 _5102_ (.Y(_1257_),
    .A(net534),
    .B(_1255_));
 sg13g2_o21ai_1 _5103_ (.B1(_1254_),
    .Y(_0251_),
    .A1(_1239_),
    .A2(net535));
 sg13g2_nand2_1 _5104_ (.Y(_1258_),
    .A(net963),
    .B(net939));
 sg13g2_xor2_1 _5105_ (.B(_1256_),
    .A(net496),
    .X(_1259_));
 sg13g2_o21ai_1 _5106_ (.B1(_1258_),
    .Y(_0252_),
    .A1(_1239_),
    .A2(net497));
 sg13g2_nand2_1 _5107_ (.Y(_1260_),
    .A(net499),
    .B(net939));
 sg13g2_nor3_1 _5108_ (.A(_0019_),
    .B(_3221_),
    .C(_1255_),
    .Y(_1261_));
 sg13g2_o21ai_1 _5109_ (.B1(_0019_),
    .Y(_1262_),
    .A1(_3221_),
    .A2(_1255_));
 sg13g2_nand2b_1 _5110_ (.Y(_1263_),
    .B(_1262_),
    .A_N(_1239_));
 sg13g2_o21ai_1 _5111_ (.B1(_1260_),
    .Y(_0253_),
    .A1(_1261_),
    .A2(_1263_));
 sg13g2_nand2_1 _5112_ (.Y(_1264_),
    .A(net962),
    .B(net938));
 sg13g2_xor2_1 _5113_ (.B(_1261_),
    .A(net389),
    .X(_1265_));
 sg13g2_o21ai_1 _5114_ (.B1(_1264_),
    .Y(_0254_),
    .A1(_1239_),
    .A2(net390));
 sg13g2_nand2_1 _5115_ (.Y(_1266_),
    .A(net997),
    .B(_3188_));
 sg13g2_xnor2_1 _5116_ (.Y(_1267_),
    .A(net996),
    .B(\vgademo.scanline_audio_sample[6] ));
 sg13g2_nand3_1 _5117_ (.B(_1266_),
    .C(_1267_),
    .A(_0037_),
    .Y(_1268_));
 sg13g2_nor2b_1 _5118_ (.A(\vgademo.scanline_audio_sample[4] ),
    .B_N(net998),
    .Y(_1269_));
 sg13g2_nand2b_1 _5119_ (.Y(_1270_),
    .B(\vgademo.scanline_audio_sample[4] ),
    .A_N(net998));
 sg13g2_o21ai_1 _5120_ (.B1(_1270_),
    .Y(_1271_),
    .A1(net997),
    .A2(_3188_));
 sg13g2_nor3_1 _5121_ (.A(_1268_),
    .B(_1269_),
    .C(_1271_),
    .Y(_1272_));
 sg13g2_nand2_1 _5122_ (.Y(_1273_),
    .A(_3108_),
    .B(\vgademo.scanline_audio_sample[2] ));
 sg13g2_nand2b_1 _5123_ (.Y(_1274_),
    .B(net1002),
    .A_N(\vgademo.scanline_audio_sample[2] ));
 sg13g2_nand2_1 _5124_ (.Y(_1275_),
    .A(_1273_),
    .B(_1274_));
 sg13g2_nand2_1 _5125_ (.Y(_1276_),
    .A(net1000),
    .B(_3189_));
 sg13g2_xnor2_1 _5126_ (.Y(_1277_),
    .A(net1000),
    .B(\vgademo.scanline_audio_sample[3] ));
 sg13g2_nand4_1 _5127_ (.B(_1273_),
    .C(_1274_),
    .A(_1272_),
    .Y(_1278_),
    .D(_1277_));
 sg13g2_xor2_1 _5128_ (.B(\vgademo.scanline_audio_sample[1] ),
    .A(net1003),
    .X(_1279_));
 sg13g2_a21oi_1 _5129_ (.A1(net1005),
    .A2(_3190_),
    .Y(_1280_),
    .B1(_1279_));
 sg13g2_a21o_1 _5130_ (.A2(\vgademo.scanline_audio_sample[1] ),
    .A1(_3106_),
    .B1(_1280_),
    .X(_1281_));
 sg13g2_nand2b_1 _5131_ (.Y(_1282_),
    .B(_1281_),
    .A_N(_1278_));
 sg13g2_nor2_1 _5132_ (.A(\vgademo.h_count[7] ),
    .B(\vgademo.h_count[6] ),
    .Y(_1283_));
 sg13g2_nor2b_1 _5133_ (.A(_1268_),
    .B_N(_1271_),
    .Y(_1284_));
 sg13g2_a21oi_1 _5134_ (.A1(\vgademo.scanline_audio_sample[6] ),
    .A2(_1283_),
    .Y(_1285_),
    .B1(_1284_));
 sg13g2_o21ai_1 _5135_ (.B1(_1273_),
    .Y(_1286_),
    .A1(net1000),
    .A2(_3189_));
 sg13g2_nand3_1 _5136_ (.B(_1276_),
    .C(_1286_),
    .A(_1272_),
    .Y(_1287_));
 sg13g2_nand3_1 _5137_ (.B(_1285_),
    .C(_1287_),
    .A(_1282_),
    .Y(_1288_));
 sg13g2_inv_1 _5138_ (.Y(_1289_),
    .A(_1288_));
 sg13g2_o21ai_1 _5139_ (.B1(_1280_),
    .Y(_1290_),
    .A1(net1005),
    .A2(_3190_));
 sg13g2_nor2_1 _5140_ (.A(_1278_),
    .B(_1290_),
    .Y(_1291_));
 sg13g2_nand2_1 _5141_ (.Y(_1292_),
    .A(net995),
    .B(_3227_));
 sg13g2_nor3_2 _5142_ (.A(_1289_),
    .B(_1291_),
    .C(_1292_),
    .Y(_1293_));
 sg13g2_inv_1 _5143_ (.Y(_1294_),
    .A(net863));
 sg13g2_xor2_1 _5144_ (.B(_1105_),
    .A(\vgademo.v_count[2] ),
    .X(_1295_));
 sg13g2_nand4_1 _5145_ (.B(_1097_),
    .C(_1121_),
    .A(_1088_),
    .Y(_1296_),
    .D(_1295_));
 sg13g2_nor2_1 _5146_ (.A(_3121_),
    .B(_1096_),
    .Y(_1297_));
 sg13g2_nand3_1 _5147_ (.B(_1295_),
    .C(_1297_),
    .A(_1121_),
    .Y(_1298_));
 sg13g2_a22oi_1 _5148_ (.Y(_1299_),
    .B1(_1121_),
    .B2(_1122_),
    .A2(_1119_),
    .A1(_3102_));
 sg13g2_nand3_1 _5149_ (.B(_1298_),
    .C(_1299_),
    .A(_1296_),
    .Y(_1300_));
 sg13g2_nand2b_1 _5150_ (.Y(_1301_),
    .B(_1185_),
    .A_N(_1170_));
 sg13g2_nor2_1 _5151_ (.A(net962),
    .B(_1197_),
    .Y(_1302_));
 sg13g2_nor4_1 _5152_ (.A(net962),
    .B(_1136_),
    .C(_1152_),
    .D(_1197_),
    .Y(_1303_));
 sg13g2_nor2b_1 _5153_ (.A(_1301_),
    .B_N(_1303_),
    .Y(_1304_));
 sg13g2_and2_1 _5154_ (.A(_3222_),
    .B(_1196_),
    .X(_1305_));
 sg13g2_nand2_1 _5155_ (.Y(_1306_),
    .A(_3104_),
    .B(_1134_));
 sg13g2_a21o_1 _5156_ (.A2(_1306_),
    .A1(_1151_),
    .B1(_1150_),
    .X(_1307_));
 sg13g2_a22oi_1 _5157_ (.Y(_1308_),
    .B1(_1185_),
    .B2(_1186_),
    .A2(_1183_),
    .A1(_3105_));
 sg13g2_o21ai_1 _5158_ (.B1(_1308_),
    .Y(_1309_),
    .A1(_1301_),
    .A2(_1307_));
 sg13g2_a221oi_1 _5159_ (.B2(_1302_),
    .C1(_1305_),
    .B1(_1309_),
    .A1(_1300_),
    .Y(_1310_),
    .A2(_1304_));
 sg13g2_and4_1 _5160_ (.A(_1089_),
    .B(_1097_),
    .C(_1121_),
    .D(_1295_),
    .X(_1311_));
 sg13g2_and2_1 _5161_ (.A(_1304_),
    .B(_1311_),
    .X(_1312_));
 sg13g2_nand2_2 _5162_ (.Y(_1313_),
    .A(_1304_),
    .B(_1311_));
 sg13g2_nor2_1 _5163_ (.A(_1310_),
    .B(_1312_),
    .Y(_1314_));
 sg13g2_nand2b_1 _5164_ (.Y(_1315_),
    .B(_1313_),
    .A_N(_1310_));
 sg13g2_mux2_1 _5165_ (.A0(_0077_),
    .A1(_0052_),
    .S(net857),
    .X(_1316_));
 sg13g2_nor2_1 _5166_ (.A(\vgademo.b_cos[9] ),
    .B(_1316_),
    .Y(_1317_));
 sg13g2_mux2_1 _5167_ (.A0(_0074_),
    .A1(_0051_),
    .S(net857),
    .X(_1318_));
 sg13g2_nor2_1 _5168_ (.A(\vgademo.b_cos[8] ),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_mux2_1 _5169_ (.A0(_0071_),
    .A1(_0049_),
    .S(net857),
    .X(_1320_));
 sg13g2_nand2b_1 _5170_ (.Y(_1321_),
    .B(_3145_),
    .A_N(_1320_));
 sg13g2_xnor2_1 _5171_ (.Y(_1322_),
    .A(\vgademo.b_cos[7] ),
    .B(_1320_));
 sg13g2_nor2_1 _5172_ (.A(_3144_),
    .B(\vgademo.plane_du[2] ),
    .Y(_1323_));
 sg13g2_nand2_1 _5173_ (.Y(_1324_),
    .A(\vgademo.b_cos[6] ),
    .B(_1323_));
 sg13g2_nor2_1 _5174_ (.A(net959),
    .B(_1323_),
    .Y(_1325_));
 sg13g2_o21ai_1 _5175_ (.B1(_1324_),
    .Y(_1326_),
    .A1(_3192_),
    .A2(_1325_));
 sg13g2_nand2_1 _5176_ (.Y(_1327_),
    .A(net857),
    .B(_1326_));
 sg13g2_nor2_1 _5177_ (.A(net969),
    .B(_3144_),
    .Y(_1328_));
 sg13g2_nor2_1 _5178_ (.A(net959),
    .B(_1328_),
    .Y(_1329_));
 sg13g2_nand2_1 _5179_ (.Y(_1330_),
    .A(net959),
    .B(_1328_));
 sg13g2_a21o_1 _5180_ (.A2(_1330_),
    .A1(_3121_),
    .B1(_1329_),
    .X(_1331_));
 sg13g2_o21ai_1 _5181_ (.B1(_1327_),
    .Y(_1332_),
    .A1(net857),
    .A2(_1331_));
 sg13g2_o21ai_1 _5182_ (.B1(_1321_),
    .Y(_1333_),
    .A1(_1322_),
    .A2(_1332_));
 sg13g2_xor2_1 _5183_ (.B(_1318_),
    .A(net958),
    .X(_1334_));
 sg13g2_a21oi_1 _5184_ (.A1(_1333_),
    .A2(_1334_),
    .Y(_1335_),
    .B1(_1319_));
 sg13g2_xnor2_1 _5185_ (.Y(_1336_),
    .A(_3147_),
    .B(_1316_));
 sg13g2_nor2b_1 _5186_ (.A(_1335_),
    .B_N(_1336_),
    .Y(_1337_));
 sg13g2_nor2_1 _5187_ (.A(_1317_),
    .B(_1337_),
    .Y(_1338_));
 sg13g2_mux2_1 _5188_ (.A0(_0063_),
    .A1(_0053_),
    .S(net857),
    .X(_1339_));
 sg13g2_xnor2_1 _5189_ (.Y(_1340_),
    .A(net956),
    .B(_1339_));
 sg13g2_o21ai_1 _5190_ (.B1(_1340_),
    .Y(_1341_),
    .A1(_1317_),
    .A2(_1337_));
 sg13g2_xnor2_1 _5191_ (.Y(_1342_),
    .A(_1338_),
    .B(_1340_));
 sg13g2_inv_1 _5192_ (.Y(_1343_),
    .A(_1342_));
 sg13g2_xor2_1 _5193_ (.B(_1336_),
    .A(_1335_),
    .X(_1344_));
 sg13g2_inv_1 _5194_ (.Y(_1345_),
    .A(_1344_));
 sg13g2_xor2_1 _5195_ (.B(_1332_),
    .A(_1322_),
    .X(_1346_));
 sg13g2_xnor2_1 _5196_ (.Y(_1347_),
    .A(_1322_),
    .B(_1332_));
 sg13g2_xor2_1 _5197_ (.B(_1334_),
    .A(_1333_),
    .X(_1348_));
 sg13g2_inv_2 _5198_ (.Y(_1349_),
    .A(net845));
 sg13g2_nor2_2 _5199_ (.A(net846),
    .B(_1349_),
    .Y(_1350_));
 sg13g2_nand2_1 _5200_ (.Y(_1351_),
    .A(_1346_),
    .B(net845));
 sg13g2_nand2_1 _5201_ (.Y(_1352_),
    .A(net985),
    .B(_1204_));
 sg13g2_nand2_1 _5202_ (.Y(_1353_),
    .A(net977),
    .B(_3117_));
 sg13g2_nor2_1 _5203_ (.A(net982),
    .B(_1353_),
    .Y(_1354_));
 sg13g2_a21oi_1 _5204_ (.A1(_1352_),
    .A2(_1354_),
    .Y(_1355_),
    .B1(_0080_));
 sg13g2_and4_1 _5205_ (.A(net985),
    .B(_1083_),
    .C(_1203_),
    .D(_1354_),
    .X(_1356_));
 sg13g2_o21ai_1 _5206_ (.B1(net974),
    .Y(_1357_),
    .A1(_1355_),
    .A2(_1356_));
 sg13g2_nand4_1 _5207_ (.B(_3114_),
    .C(_1043_),
    .A(_3113_),
    .Y(_1358_),
    .D(_1357_));
 sg13g2_inv_1 _5208_ (.Y(_1359_),
    .A(_1358_));
 sg13g2_nor2_1 _5209_ (.A(net971),
    .B(_1079_),
    .Y(_1360_));
 sg13g2_nand2_1 _5210_ (.Y(_1361_),
    .A(\vgademo.a_scrolly[13] ),
    .B(\vgademo.a_scrolly[11] ));
 sg13g2_o21ai_1 _5211_ (.B1(_1069_),
    .Y(_1362_),
    .A1(_1360_),
    .A2(_1361_));
 sg13g2_a21oi_2 _5212_ (.B1(_1359_),
    .Y(_1363_),
    .A2(net888),
    .A1(_1067_));
 sg13g2_a21o_2 _5213_ (.A2(_1362_),
    .A1(_1067_),
    .B1(_1359_),
    .X(_1364_));
 sg13g2_nor2_1 _5214_ (.A(_1060_),
    .B(_1353_),
    .Y(_1365_));
 sg13g2_a21oi_1 _5215_ (.A1(_1115_),
    .A2(_1365_),
    .Y(_1366_),
    .B1(_1063_));
 sg13g2_and4_1 _5216_ (.A(net991),
    .B(net982),
    .C(_1034_),
    .D(_1365_),
    .X(_1367_));
 sg13g2_nor3_2 _5217_ (.A(_1081_),
    .B(_1366_),
    .C(_1367_),
    .Y(_1368_));
 sg13g2_inv_1 _5218_ (.Y(_1369_),
    .A(_1368_));
 sg13g2_xnor2_1 _5219_ (.Y(_1370_),
    .A(net986),
    .B(_1204_));
 sg13g2_a221oi_1 _5220_ (.B2(net888),
    .C1(_1364_),
    .B1(_1370_),
    .A1(net986),
    .Y(_1371_),
    .A2(_1368_));
 sg13g2_nor2_1 _5221_ (.A(_0030_),
    .B(net858),
    .Y(_1372_));
 sg13g2_nor3_1 _5222_ (.A(net1003),
    .B(net1000),
    .C(net1002),
    .Y(_1373_));
 sg13g2_nor2b_1 _5223_ (.A(net998),
    .B_N(_1373_),
    .Y(_1374_));
 sg13g2_nor2_1 _5224_ (.A(_3109_),
    .B(_1374_),
    .Y(_1375_));
 sg13g2_xnor2_1 _5225_ (.Y(_1376_),
    .A(_0036_),
    .B(_1375_));
 sg13g2_a21oi_2 _5226_ (.B1(_1372_),
    .Y(_1377_),
    .A2(_1376_),
    .A1(net858));
 sg13g2_nor2b_2 _5227_ (.A(_1377_),
    .B_N(_1371_),
    .Y(_1378_));
 sg13g2_nand2b_1 _5228_ (.Y(_1379_),
    .B(_1371_),
    .A_N(_1377_));
 sg13g2_nand2_1 _5229_ (.Y(_1380_),
    .A(_1068_),
    .B(net888));
 sg13g2_nand3_1 _5230_ (.B(_1211_),
    .C(net888),
    .A(_1068_),
    .Y(_1381_));
 sg13g2_o21ai_1 _5231_ (.B1(_1381_),
    .Y(_1382_),
    .A1(_0069_),
    .A2(_1369_));
 sg13g2_nand2_2 _5232_ (.Y(_1383_),
    .A(_1358_),
    .B(_1382_));
 sg13g2_xnor2_1 _5233_ (.Y(_1384_),
    .A(_3109_),
    .B(_1374_));
 sg13g2_mux2_2 _5234_ (.A0(_0047_),
    .A1(_1384_),
    .S(net858),
    .X(_1385_));
 sg13g2_nor2_2 _5235_ (.A(_1383_),
    .B(_1385_),
    .Y(_1386_));
 sg13g2_or2_1 _5236_ (.X(_1387_),
    .B(_1385_),
    .A(_1383_));
 sg13g2_a221oi_1 _5237_ (.B2(_0064_),
    .C1(_1364_),
    .B1(_1368_),
    .A1(net993),
    .Y(_1388_),
    .A2(net888));
 sg13g2_xor2_1 _5238_ (.B(_1373_),
    .A(_0044_),
    .X(_1389_));
 sg13g2_o21ai_1 _5239_ (.B1(_0029_),
    .Y(_1390_),
    .A1(_1310_),
    .A2(_1312_));
 sg13g2_nand3b_1 _5240_ (.B(_1313_),
    .C(_1389_),
    .Y(_1391_),
    .A_N(_1310_));
 sg13g2_and3_1 _5241_ (.X(_1392_),
    .A(_1388_),
    .B(_1390_),
    .C(_1391_));
 sg13g2_nand3_1 _5242_ (.B(_1390_),
    .C(_1391_),
    .A(_1388_),
    .Y(_1393_));
 sg13g2_o21ai_1 _5243_ (.B1(_3191_),
    .Y(_1394_),
    .A1(_1310_),
    .A2(_1312_));
 sg13g2_xnor2_1 _5244_ (.Y(_1395_),
    .A(_0034_),
    .B(_3232_));
 sg13g2_nand3b_1 _5245_ (.B(_1313_),
    .C(_1395_),
    .Y(_1396_),
    .A_N(_1310_));
 sg13g2_and2_1 _5246_ (.A(_1394_),
    .B(_1396_),
    .X(_1397_));
 sg13g2_xnor2_1 _5247_ (.Y(_1398_),
    .A(net1004),
    .B(\vgademo.h_count[2] ));
 sg13g2_o21ai_1 _5248_ (.B1(_3169_),
    .Y(_1399_),
    .A1(_1310_),
    .A2(_1312_));
 sg13g2_nand3b_1 _5249_ (.B(_1313_),
    .C(_1398_),
    .Y(_1400_),
    .A_N(_1310_));
 sg13g2_nand4_1 _5250_ (.B(_1396_),
    .C(_1399_),
    .A(_1394_),
    .Y(_1401_),
    .D(_1400_));
 sg13g2_a21o_1 _5251_ (.A2(_1391_),
    .A1(_1390_),
    .B1(_1388_),
    .X(_1402_));
 sg13g2_and4_2 _5252_ (.A(_1363_),
    .B(_1393_),
    .C(_1401_),
    .D(_1402_),
    .X(_1403_));
 sg13g2_nand4_1 _5253_ (.B(_1393_),
    .C(_1401_),
    .A(_1363_),
    .Y(_1404_),
    .D(_1402_));
 sg13g2_xor2_1 _5254_ (.B(_1385_),
    .A(_1383_),
    .X(_1405_));
 sg13g2_xnor2_1 _5255_ (.Y(_1406_),
    .A(_1383_),
    .B(_1385_));
 sg13g2_a21oi_2 _5256_ (.B1(_1406_),
    .Y(_1407_),
    .A2(_1404_),
    .A1(_1393_));
 sg13g2_o21ai_1 _5257_ (.B1(_1405_),
    .Y(_1408_),
    .A1(_1392_),
    .A2(_1403_));
 sg13g2_xnor2_1 _5258_ (.Y(_1409_),
    .A(_1371_),
    .B(_1377_));
 sg13g2_xor2_1 _5259_ (.B(_1377_),
    .A(_1371_),
    .X(_1410_));
 sg13g2_a21oi_2 _5260_ (.B1(_1410_),
    .Y(_1411_),
    .A2(_1408_),
    .A1(_1387_));
 sg13g2_o21ai_1 _5261_ (.B1(_1409_),
    .Y(_1412_),
    .A1(_1386_),
    .A2(_1407_));
 sg13g2_nand2_1 _5262_ (.Y(_1413_),
    .A(_1033_),
    .B(_1217_));
 sg13g2_nand2_1 _5263_ (.Y(_1414_),
    .A(_0075_),
    .B(_1352_));
 sg13g2_xor2_1 _5264_ (.B(_1352_),
    .A(_0075_),
    .X(_1415_));
 sg13g2_a221oi_1 _5265_ (.B2(net888),
    .C1(_1364_),
    .B1(_1415_),
    .A1(_1368_),
    .Y(_1416_),
    .A2(_1413_));
 sg13g2_nand2_1 _5266_ (.Y(_1417_),
    .A(net996),
    .B(_1375_));
 sg13g2_inv_1 _5267_ (.Y(_1418_),
    .A(_1417_));
 sg13g2_xnor2_1 _5268_ (.Y(_1419_),
    .A(_3110_),
    .B(_1417_));
 sg13g2_nor2_1 _5269_ (.A(_0046_),
    .B(net858),
    .Y(_1420_));
 sg13g2_a21oi_2 _5270_ (.B1(_1420_),
    .Y(_1421_),
    .A2(_1419_),
    .A1(net858));
 sg13g2_inv_1 _5271_ (.Y(_1422_),
    .A(_1421_));
 sg13g2_nand2_2 _5272_ (.Y(_1423_),
    .A(_1416_),
    .B(_1422_));
 sg13g2_inv_1 _5273_ (.Y(_1424_),
    .A(_1423_));
 sg13g2_xnor2_1 _5274_ (.Y(_1425_),
    .A(_1416_),
    .B(_1421_));
 sg13g2_xor2_1 _5275_ (.B(_1421_),
    .A(_1416_),
    .X(_1426_));
 sg13g2_a21oi_2 _5276_ (.B1(_1426_),
    .Y(_1427_),
    .A2(_1412_),
    .A1(_1379_));
 sg13g2_o21ai_1 _5277_ (.B1(_1425_),
    .Y(_1428_),
    .A1(_1378_),
    .A2(_1411_));
 sg13g2_nor3_2 _5278_ (.A(_1378_),
    .B(_1411_),
    .C(_1425_),
    .Y(_1429_));
 sg13g2_nand3_1 _5279_ (.B(_1412_),
    .C(_1426_),
    .A(_1379_),
    .Y(_1430_));
 sg13g2_o21ai_1 _5280_ (.B1(_1426_),
    .Y(_1431_),
    .A1(_1378_),
    .A2(_1411_));
 sg13g2_nand3_1 _5281_ (.B(_1412_),
    .C(_1425_),
    .A(_1379_),
    .Y(_1432_));
 sg13g2_nor2_2 _5282_ (.A(_1427_),
    .B(_1429_),
    .Y(_1433_));
 sg13g2_nand2_1 _5283_ (.Y(_1434_),
    .A(net842),
    .B(net840));
 sg13g2_nor3_2 _5284_ (.A(_1386_),
    .B(_1407_),
    .C(_1409_),
    .Y(_1435_));
 sg13g2_nand3_1 _5285_ (.B(_1408_),
    .C(_1410_),
    .A(_1387_),
    .Y(_1436_));
 sg13g2_nand3_1 _5286_ (.B(_1408_),
    .C(_1409_),
    .A(_1387_),
    .Y(_1437_));
 sg13g2_o21ai_1 _5287_ (.B1(_1410_),
    .Y(_1438_),
    .A1(_1386_),
    .A2(_1407_));
 sg13g2_nor2_2 _5288_ (.A(_1411_),
    .B(_1435_),
    .Y(_1439_));
 sg13g2_nand2_2 _5289_ (.Y(_1440_),
    .A(_1412_),
    .B(_1436_));
 sg13g2_a21oi_2 _5290_ (.B1(_1439_),
    .Y(_1441_),
    .A2(net840),
    .A1(net842));
 sg13g2_nor3_2 _5291_ (.A(_1392_),
    .B(_1403_),
    .C(_1405_),
    .Y(_1442_));
 sg13g2_nand3_1 _5292_ (.B(_1404_),
    .C(_1406_),
    .A(_1393_),
    .Y(_1443_));
 sg13g2_nor2_2 _5293_ (.A(_1407_),
    .B(_1442_),
    .Y(_1444_));
 sg13g2_nand2_2 _5294_ (.Y(_1445_),
    .A(_1408_),
    .B(_1443_));
 sg13g2_a22oi_1 _5295_ (.Y(_1446_),
    .B1(_1402_),
    .B2(_1393_),
    .A2(_1401_),
    .A1(_1363_));
 sg13g2_nor2_1 _5296_ (.A(_1403_),
    .B(_1446_),
    .Y(_1447_));
 sg13g2_or2_2 _5297_ (.X(_1448_),
    .B(_1446_),
    .A(_1403_));
 sg13g2_o21ai_1 _5298_ (.B1(_1448_),
    .Y(_1449_),
    .A1(_1407_),
    .A2(_1442_));
 sg13g2_a22oi_1 _5299_ (.Y(_1450_),
    .B1(_1445_),
    .B2(_1448_),
    .A2(_1438_),
    .A1(_1437_));
 sg13g2_a21oi_1 _5300_ (.A1(net841),
    .A2(net839),
    .Y(_1451_),
    .B1(_1450_));
 sg13g2_nand3_1 _5301_ (.B(_1399_),
    .C(_1400_),
    .A(_1363_),
    .Y(_1452_));
 sg13g2_xnor2_1 _5302_ (.Y(_1453_),
    .A(_1397_),
    .B(_1452_));
 sg13g2_nand2_2 _5303_ (.Y(_1454_),
    .A(_1448_),
    .B(_1453_));
 sg13g2_nand2_1 _5304_ (.Y(_1455_),
    .A(_1444_),
    .B(_1454_));
 sg13g2_a22oi_1 _5305_ (.Y(_1456_),
    .B1(_1444_),
    .B2(_1454_),
    .A2(_1436_),
    .A1(_1412_));
 sg13g2_nor3_1 _5306_ (.A(_1427_),
    .B(_1429_),
    .C(_1456_),
    .Y(_1457_));
 sg13g2_nor2_1 _5307_ (.A(_1451_),
    .B(_1457_),
    .Y(_1458_));
 sg13g2_o21ai_1 _5308_ (.B1(_1036_),
    .Y(_1459_),
    .A1(_1034_),
    .A2(_1414_));
 sg13g2_nor3_1 _5309_ (.A(_3117_),
    .B(_1034_),
    .C(_1414_),
    .Y(_1460_));
 sg13g2_xnor2_1 _5310_ (.Y(_1461_),
    .A(_3117_),
    .B(_1459_));
 sg13g2_a221oi_1 _5311_ (.B2(net888),
    .C1(_1364_),
    .B1(_1461_),
    .A1(_1218_),
    .Y(_1462_),
    .A2(_1368_));
 sg13g2_nor2_1 _5312_ (.A(_0031_),
    .B(net858),
    .Y(_1463_));
 sg13g2_nand2_1 _5313_ (.Y(_1464_),
    .A(_0037_),
    .B(_1417_));
 sg13g2_xor2_1 _5314_ (.B(_1464_),
    .A(_0038_),
    .X(_1465_));
 sg13g2_a21oi_2 _5315_ (.B1(_1463_),
    .Y(_1466_),
    .A2(_1465_),
    .A1(net858));
 sg13g2_nand2b_1 _5316_ (.Y(_1467_),
    .B(_1462_),
    .A_N(_1466_));
 sg13g2_xor2_1 _5317_ (.B(_1466_),
    .A(_1462_),
    .X(_1468_));
 sg13g2_a21o_2 _5318_ (.A2(net843),
    .A1(_1423_),
    .B1(_1468_),
    .X(_1469_));
 sg13g2_xnor2_1 _5319_ (.Y(_1470_),
    .A(_0080_),
    .B(_1077_));
 sg13g2_and2_1 _5320_ (.A(_1460_),
    .B(_1470_),
    .X(_1471_));
 sg13g2_or2_1 _5321_ (.X(_1472_),
    .B(_1470_),
    .A(_1460_));
 sg13g2_inv_1 _5322_ (.Y(_1473_),
    .A(_1472_));
 sg13g2_or3_1 _5323_ (.A(_1380_),
    .B(_1471_),
    .C(_1473_),
    .X(_1474_));
 sg13g2_o21ai_1 _5324_ (.B1(net978),
    .Y(_1475_),
    .A1(net980),
    .A2(_1033_));
 sg13g2_nand3_1 _5325_ (.B(_1033_),
    .C(_1217_),
    .A(_0078_),
    .Y(_1476_));
 sg13g2_nand3_1 _5326_ (.B(_1475_),
    .C(_1476_),
    .A(_1039_),
    .Y(_1477_));
 sg13g2_or2_1 _5327_ (.X(_1478_),
    .B(_1476_),
    .A(_3116_));
 sg13g2_nand3_1 _5328_ (.B(_1477_),
    .C(_1478_),
    .A(_1368_),
    .Y(_1479_));
 sg13g2_a21o_1 _5329_ (.A2(_1479_),
    .A1(_1474_),
    .B1(_1359_),
    .X(_1480_));
 sg13g2_nor2_1 _5330_ (.A(_0045_),
    .B(net858),
    .Y(_1481_));
 sg13g2_nor3_2 _5331_ (.A(\vgademo.h_count[7] ),
    .B(\vgademo.h_count[8] ),
    .C(_1418_),
    .Y(_1482_));
 sg13g2_xnor2_1 _5332_ (.Y(_1483_),
    .A(\vgademo.h_count[9] ),
    .B(_1482_));
 sg13g2_a21oi_2 _5333_ (.B1(_1481_),
    .Y(_1484_),
    .A2(_1483_),
    .A1(net859));
 sg13g2_or2_1 _5334_ (.X(_1485_),
    .B(_1484_),
    .A(_1480_));
 sg13g2_xnor2_1 _5335_ (.Y(_1486_),
    .A(_1480_),
    .B(_1484_));
 sg13g2_inv_1 _5336_ (.Y(_1487_),
    .A(_1486_));
 sg13g2_a21o_1 _5337_ (.A2(_1469_),
    .A1(_1467_),
    .B1(_1486_),
    .X(_1488_));
 sg13g2_nand3_1 _5338_ (.B(_1469_),
    .C(_1487_),
    .A(_1467_),
    .Y(_1489_));
 sg13g2_a21o_1 _5339_ (.A2(_1469_),
    .A1(_1467_),
    .B1(_1487_),
    .X(_1490_));
 sg13g2_nand2_2 _5340_ (.Y(_1491_),
    .A(_1489_),
    .B(_1490_));
 sg13g2_and2_1 _5341_ (.A(_1489_),
    .B(_1490_),
    .X(_1492_));
 sg13g2_nand2b_1 _5342_ (.Y(_1493_),
    .B(_1453_),
    .A_N(_1449_));
 sg13g2_xnor2_1 _5343_ (.Y(_1494_),
    .A(_1444_),
    .B(_1454_));
 sg13g2_nor2_1 _5344_ (.A(_1439_),
    .B(_1494_),
    .Y(_1495_));
 sg13g2_nand3_1 _5345_ (.B(_1443_),
    .C(_1447_),
    .A(_1408_),
    .Y(_1496_));
 sg13g2_nand2_1 _5346_ (.Y(_1497_),
    .A(_1449_),
    .B(_1496_));
 sg13g2_nor2_1 _5347_ (.A(_1440_),
    .B(_1497_),
    .Y(_1498_));
 sg13g2_nand4_1 _5348_ (.B(_1436_),
    .C(_1449_),
    .A(_1412_),
    .Y(_1499_),
    .D(_1496_));
 sg13g2_mux2_1 _5349_ (.A0(_1495_),
    .A1(_1498_),
    .S(_1434_),
    .X(_1500_));
 sg13g2_nor2_1 _5350_ (.A(_1351_),
    .B(_1500_),
    .Y(_1501_));
 sg13g2_nor2_1 _5351_ (.A(_1491_),
    .B(_1501_),
    .Y(_1502_));
 sg13g2_o21ai_1 _5352_ (.B1(_1502_),
    .Y(_1503_),
    .A1(_1350_),
    .A2(_1458_));
 sg13g2_nand3_1 _5353_ (.B(net843),
    .C(_1468_),
    .A(_1423_),
    .Y(_1504_));
 sg13g2_nand3b_1 _5354_ (.B(net843),
    .C(_1423_),
    .Y(_1505_),
    .A_N(_1468_));
 sg13g2_o21ai_1 _5355_ (.B1(_1468_),
    .Y(_1506_),
    .A1(_1424_),
    .A2(_1427_));
 sg13g2_nand2_1 _5356_ (.Y(_1507_),
    .A(_1505_),
    .B(_1506_));
 sg13g2_nand2_2 _5357_ (.Y(_1508_),
    .A(_1469_),
    .B(_1504_));
 sg13g2_mux2_1 _5358_ (.A0(_1448_),
    .A1(_1454_),
    .S(_1445_),
    .X(_1509_));
 sg13g2_a221oi_1 _5359_ (.B2(_1509_),
    .C1(_1450_),
    .B1(_1440_),
    .A1(net842),
    .Y(_1510_),
    .A2(net840));
 sg13g2_a221oi_1 _5360_ (.B2(_1509_),
    .C1(_1456_),
    .B1(_1439_),
    .A1(_1431_),
    .Y(_1511_),
    .A2(_1432_));
 sg13g2_o21ai_1 _5361_ (.B1(net846),
    .Y(_1512_),
    .A1(_1510_),
    .A2(_1511_));
 sg13g2_nor3_1 _5362_ (.A(_1427_),
    .B(_1429_),
    .C(_1440_),
    .Y(_1513_));
 sg13g2_nand3_1 _5363_ (.B(net840),
    .C(_1439_),
    .A(net841),
    .Y(_1514_));
 sg13g2_nand4_1 _5364_ (.B(net840),
    .C(_1439_),
    .A(net842),
    .Y(_1515_),
    .D(_1455_));
 sg13g2_or3_1 _5365_ (.A(_1403_),
    .B(_1446_),
    .C(_1453_),
    .X(_1516_));
 sg13g2_nand3b_1 _5366_ (.B(_1443_),
    .C(_1408_),
    .Y(_1517_),
    .A_N(_1516_));
 sg13g2_o21ai_1 _5367_ (.B1(_1517_),
    .Y(_1518_),
    .A1(_1411_),
    .A2(_1435_));
 sg13g2_a221oi_1 _5368_ (.B2(_1448_),
    .C1(_1518_),
    .B1(_1445_),
    .A1(net841),
    .Y(_1519_),
    .A2(net839));
 sg13g2_nand3b_1 _5369_ (.B(_1346_),
    .C(_1515_),
    .Y(_1520_),
    .A_N(_1519_));
 sg13g2_a21oi_1 _5370_ (.A1(_1512_),
    .A2(_1520_),
    .Y(_1521_),
    .B1(net845));
 sg13g2_nor3_1 _5371_ (.A(_1433_),
    .B(_1450_),
    .C(_1495_),
    .Y(_1522_));
 sg13g2_a21o_1 _5372_ (.A2(_1499_),
    .A1(_1457_),
    .B1(_1522_),
    .X(_1523_));
 sg13g2_nor2_2 _5373_ (.A(_1346_),
    .B(_1349_),
    .Y(_1524_));
 sg13g2_nand4_1 _5374_ (.B(net839),
    .C(_1439_),
    .A(net841),
    .Y(_1525_),
    .D(_1509_));
 sg13g2_nand4_1 _5375_ (.B(_1432_),
    .C(_1440_),
    .A(_1431_),
    .Y(_1526_),
    .D(_1509_));
 sg13g2_and2_1 _5376_ (.A(_1525_),
    .B(_1526_),
    .X(_1527_));
 sg13g2_a221oi_1 _5377_ (.B2(_1527_),
    .C1(_1521_),
    .B1(_1524_),
    .A1(_1350_),
    .Y(_1528_),
    .A2(_1523_));
 sg13g2_and2_1 _5378_ (.A(_1445_),
    .B(_1516_),
    .X(_1529_));
 sg13g2_o21ai_1 _5379_ (.B1(_1516_),
    .Y(_1530_),
    .A1(_1407_),
    .A2(_1442_));
 sg13g2_nand4_1 _5380_ (.B(_1438_),
    .C(_1517_),
    .A(_1437_),
    .Y(_1531_),
    .D(_1530_));
 sg13g2_nand4_1 _5381_ (.B(net839),
    .C(_1499_),
    .A(net843),
    .Y(_1532_),
    .D(_1531_));
 sg13g2_nand4_1 _5382_ (.B(_1432_),
    .C(_1440_),
    .A(_1431_),
    .Y(_1533_),
    .D(_1494_));
 sg13g2_nor3_2 _5383_ (.A(_1411_),
    .B(_1435_),
    .C(_1445_),
    .Y(_1534_));
 sg13g2_nand3_1 _5384_ (.B(_1436_),
    .C(_1444_),
    .A(_1412_),
    .Y(_1535_));
 sg13g2_o21ai_1 _5385_ (.B1(_1534_),
    .Y(_1536_),
    .A1(_1427_),
    .A2(_1429_));
 sg13g2_nand3_1 _5386_ (.B(_1533_),
    .C(_1536_),
    .A(_1532_),
    .Y(_1537_));
 sg13g2_a21oi_1 _5387_ (.A1(_1508_),
    .A2(_1537_),
    .Y(_1538_),
    .B1(net834));
 sg13g2_o21ai_1 _5388_ (.B1(_1538_),
    .Y(_1539_),
    .A1(_1508_),
    .A2(_1528_));
 sg13g2_a21o_1 _5389_ (.A2(_1539_),
    .A1(_1503_),
    .B1(_1344_),
    .X(_1540_));
 sg13g2_nor2_1 _5390_ (.A(_1514_),
    .B(_1517_),
    .Y(_1541_));
 sg13g2_nand2_1 _5391_ (.Y(_1542_),
    .A(net833),
    .B(_1541_));
 sg13g2_o21ai_1 _5392_ (.B1(_1445_),
    .Y(_1543_),
    .A1(_1411_),
    .A2(_1435_));
 sg13g2_nand4_1 _5393_ (.B(net839),
    .C(_1497_),
    .A(net841),
    .Y(_1544_),
    .D(_1543_));
 sg13g2_nand4_1 _5394_ (.B(_1432_),
    .C(_1494_),
    .A(_1431_),
    .Y(_1545_),
    .D(_1535_));
 sg13g2_and2_1 _5395_ (.A(_1544_),
    .B(_1545_),
    .X(_1546_));
 sg13g2_a22oi_1 _5396_ (.Y(_1547_),
    .B1(_1544_),
    .B2(_1545_),
    .A2(_1506_),
    .A1(_1505_));
 sg13g2_nand4_1 _5397_ (.B(net839),
    .C(_1497_),
    .A(net841),
    .Y(_1548_),
    .D(_1518_));
 sg13g2_nand2_1 _5398_ (.Y(_1549_),
    .A(_1533_),
    .B(_1548_));
 sg13g2_a21oi_2 _5399_ (.B1(_1547_),
    .Y(_1550_),
    .A2(_1549_),
    .A1(_1508_));
 sg13g2_o21ai_1 _5400_ (.B1(_1346_),
    .Y(_1551_),
    .A1(net833),
    .A2(_1550_));
 sg13g2_o21ai_1 _5401_ (.B1(net846),
    .Y(_1552_),
    .A1(net834),
    .A2(_1546_));
 sg13g2_a22oi_1 _5402_ (.Y(_1553_),
    .B1(_1551_),
    .B2(_1552_),
    .A2(_1541_),
    .A1(net833));
 sg13g2_a21oi_1 _5403_ (.A1(_1508_),
    .A2(_1537_),
    .Y(_1554_),
    .B1(_1547_));
 sg13g2_nand3b_1 _5404_ (.B(_1489_),
    .C(_1490_),
    .Y(_1555_),
    .A_N(_1458_));
 sg13g2_o21ai_1 _5405_ (.B1(_1555_),
    .Y(_1556_),
    .A1(net833),
    .A2(_1554_));
 sg13g2_nand2_1 _5406_ (.Y(_1557_),
    .A(_1491_),
    .B(_1550_));
 sg13g2_a221oi_1 _5407_ (.B2(_1524_),
    .C1(_1345_),
    .B1(_1557_),
    .A1(_1350_),
    .Y(_1558_),
    .A2(_1556_));
 sg13g2_o21ai_1 _5408_ (.B1(_1558_),
    .Y(_1559_),
    .A1(net845),
    .A2(_1553_));
 sg13g2_a21o_1 _5409_ (.A2(_1559_),
    .A1(_1540_),
    .B1(_1343_),
    .X(_1560_));
 sg13g2_mux2_1 _5410_ (.A0(_1495_),
    .A1(_1498_),
    .S(_1433_),
    .X(_1561_));
 sg13g2_nand2b_1 _5411_ (.Y(_1562_),
    .B(_1507_),
    .A_N(_1561_));
 sg13g2_nand2_1 _5412_ (.Y(_1563_),
    .A(_1508_),
    .B(_1527_));
 sg13g2_a21oi_1 _5413_ (.A1(_1562_),
    .A2(_1563_),
    .Y(_1564_),
    .B1(net835));
 sg13g2_a21o_1 _5414_ (.A2(_1563_),
    .A1(_1562_),
    .B1(net835),
    .X(_1565_));
 sg13g2_o21ai_1 _5415_ (.B1(_1526_),
    .Y(_1566_),
    .A1(_1494_),
    .A2(_1514_));
 sg13g2_mux2_1 _5416_ (.A0(_1561_),
    .A1(_1566_),
    .S(_1508_),
    .X(_1567_));
 sg13g2_nor2_1 _5417_ (.A(net835),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_nand3b_1 _5418_ (.B(_1491_),
    .C(_1346_),
    .Y(_1569_),
    .A_N(_1567_));
 sg13g2_nand4_1 _5419_ (.B(_1432_),
    .C(_1440_),
    .A(_1431_),
    .Y(_1570_),
    .D(_1493_));
 sg13g2_nand4_1 _5420_ (.B(_1436_),
    .C(_1444_),
    .A(_1412_),
    .Y(_1571_),
    .D(_1454_));
 sg13g2_nand4_1 _5421_ (.B(net839),
    .C(_1518_),
    .A(net841),
    .Y(_1572_),
    .D(_1571_));
 sg13g2_nand4_1 _5422_ (.B(_1506_),
    .C(_1570_),
    .A(_1505_),
    .Y(_1573_),
    .D(_1572_));
 sg13g2_nand4_1 _5423_ (.B(_1504_),
    .C(_1525_),
    .A(_1469_),
    .Y(_1574_),
    .D(_1526_));
 sg13g2_a21oi_1 _5424_ (.A1(_1573_),
    .A2(_1574_),
    .Y(_1575_),
    .B1(net834));
 sg13g2_a221oi_1 _5425_ (.B2(_1574_),
    .C1(_1346_),
    .B1(_1573_),
    .A1(_1489_),
    .Y(_1576_),
    .A2(_1490_));
 sg13g2_nor2_1 _5426_ (.A(net845),
    .B(_1576_),
    .Y(_1577_));
 sg13g2_a22oi_1 _5427_ (.Y(_1578_),
    .B1(_1569_),
    .B2(_1577_),
    .A2(_1565_),
    .A1(_1524_));
 sg13g2_a21oi_1 _5428_ (.A1(net841),
    .A2(net839),
    .Y(_1579_),
    .B1(_1543_));
 sg13g2_nor2_1 _5429_ (.A(_1514_),
    .B(_1529_),
    .Y(_1580_));
 sg13g2_a221oi_1 _5430_ (.B2(_1580_),
    .C1(_1491_),
    .B1(_1517_),
    .A1(_1441_),
    .Y(_1581_),
    .A2(_1445_));
 sg13g2_and2_1 _5431_ (.A(_1491_),
    .B(_1523_),
    .X(_1582_));
 sg13g2_a21oi_1 _5432_ (.A1(_1491_),
    .A2(_1523_),
    .Y(_1583_),
    .B1(_1351_));
 sg13g2_a21oi_1 _5433_ (.A1(_1542_),
    .A2(_1583_),
    .Y(_1584_),
    .B1(_1344_));
 sg13g2_o21ai_1 _5434_ (.B1(_1584_),
    .Y(_1585_),
    .A1(_1578_),
    .A2(_1581_));
 sg13g2_a22oi_1 _5435_ (.Y(_1586_),
    .B1(_1513_),
    .B2(_1449_),
    .A2(_1456_),
    .A1(_1434_));
 sg13g2_a221oi_1 _5436_ (.B2(_1433_),
    .C1(net846),
    .B1(_1534_),
    .A1(_1441_),
    .Y(_1587_),
    .A2(_1529_));
 sg13g2_a21oi_1 _5437_ (.A1(net846),
    .A2(_1586_),
    .Y(_1588_),
    .B1(_1587_));
 sg13g2_a22oi_1 _5438_ (.Y(_1589_),
    .B1(_1579_),
    .B2(_1448_),
    .A2(_1534_),
    .A1(_1433_));
 sg13g2_nor2_1 _5439_ (.A(_1454_),
    .B(_1579_),
    .Y(_1590_));
 sg13g2_nor3_1 _5440_ (.A(_1351_),
    .B(_1589_),
    .C(_1590_),
    .Y(_1591_));
 sg13g2_a21oi_1 _5441_ (.A1(_1507_),
    .A2(_1590_),
    .Y(_1592_),
    .B1(_1589_));
 sg13g2_a221oi_1 _5442_ (.B2(_1524_),
    .C1(_1591_),
    .B1(_1592_),
    .A1(_1349_),
    .Y(_1593_),
    .A2(_1588_));
 sg13g2_o21ai_1 _5443_ (.B1(_1542_),
    .Y(_1594_),
    .A1(net833),
    .A2(_1593_));
 sg13g2_a21oi_1 _5444_ (.A1(_1344_),
    .A2(_1594_),
    .Y(_1595_),
    .B1(_1342_));
 sg13g2_o21ai_1 _5445_ (.B1(_1341_),
    .Y(_1596_),
    .A1(_3148_),
    .A2(_1339_));
 sg13g2_nand2_2 _5446_ (.Y(_1597_),
    .A(net956),
    .B(_3149_));
 sg13g2_xnor2_1 _5447_ (.Y(_1598_),
    .A(net956),
    .B(\vgademo.b_cos[11] ));
 sg13g2_xor2_1 _5448_ (.B(\vgademo.b_cos[11] ),
    .A(\vgademo.b_cos[10] ),
    .X(_1599_));
 sg13g2_mux2_1 _5449_ (.A0(net964),
    .A1(\vgademo.plane_du[8] ),
    .S(net857),
    .X(_1600_));
 sg13g2_xnor2_1 _5450_ (.Y(_1601_),
    .A(_1599_),
    .B(_1600_));
 sg13g2_xnor2_1 _5451_ (.Y(_1602_),
    .A(_1596_),
    .B(_1601_));
 sg13g2_a21oi_1 _5452_ (.A1(_1585_),
    .A2(_1595_),
    .Y(_1603_),
    .B1(_1602_));
 sg13g2_o21ai_1 _5453_ (.B1(net846),
    .Y(_1604_),
    .A1(net833),
    .A2(_1554_));
 sg13g2_a21o_1 _5454_ (.A2(_1604_),
    .A1(_1551_),
    .B1(net845),
    .X(_1605_));
 sg13g2_o21ai_1 _5455_ (.B1(_1524_),
    .Y(_1606_),
    .A1(net833),
    .A2(_1550_));
 sg13g2_o21ai_1 _5456_ (.B1(_1350_),
    .Y(_1607_),
    .A1(net833),
    .A2(_1546_));
 sg13g2_and3_1 _5457_ (.X(_1608_),
    .A(_1344_),
    .B(_1606_),
    .C(_1607_));
 sg13g2_mux4_1 _5458_ (.S0(_1348_),
    .A0(_1564_),
    .A1(_1575_),
    .A2(_1582_),
    .A3(_1568_),
    .S1(_1347_),
    .X(_1609_));
 sg13g2_o21ai_1 _5459_ (.B1(_1343_),
    .Y(_1610_),
    .A1(_1491_),
    .A2(_1500_));
 sg13g2_a221oi_1 _5460_ (.B2(_1345_),
    .C1(_1610_),
    .B1(_1609_),
    .A1(_1605_),
    .Y(_1611_),
    .A2(_1608_));
 sg13g2_nand3_1 _5461_ (.B(_1441_),
    .C(_1529_),
    .A(net846),
    .Y(_1612_));
 sg13g2_a22oi_1 _5462_ (.Y(_1613_),
    .B1(_1513_),
    .B2(_1454_),
    .A2(_1496_),
    .A1(_1441_));
 sg13g2_o21ai_1 _5463_ (.B1(_1612_),
    .Y(_1614_),
    .A1(net846),
    .A2(_1613_));
 sg13g2_o21ai_1 _5464_ (.B1(_1508_),
    .Y(_1615_),
    .A1(_1580_),
    .A2(_1614_));
 sg13g2_a221oi_1 _5465_ (.B2(_1433_),
    .C1(_1346_),
    .B1(_1534_),
    .A1(_1441_),
    .Y(_1616_),
    .A2(_1529_));
 sg13g2_a21oi_1 _5466_ (.A1(_1346_),
    .A2(_1586_),
    .Y(_1617_),
    .B1(_1616_));
 sg13g2_a21oi_1 _5467_ (.A1(_1507_),
    .A2(_1617_),
    .Y(_1618_),
    .B1(_1349_));
 sg13g2_nand2_1 _5468_ (.Y(_1619_),
    .A(_1347_),
    .B(_1590_));
 sg13g2_nand2_1 _5469_ (.Y(_1620_),
    .A(_1592_),
    .B(_1619_));
 sg13g2_a221oi_1 _5470_ (.B2(_1349_),
    .C1(net835),
    .B1(_1620_),
    .A1(_1615_),
    .Y(_1621_),
    .A2(_1618_));
 sg13g2_nand2_1 _5471_ (.Y(_1622_),
    .A(_1342_),
    .B(_1555_));
 sg13g2_o21ai_1 _5472_ (.B1(_1602_),
    .Y(_1623_),
    .A1(_1621_),
    .A2(_1622_));
 sg13g2_nand2_1 _5473_ (.Y(_1624_),
    .A(_1485_),
    .B(_1488_));
 sg13g2_xnor2_1 _5474_ (.Y(_1625_),
    .A(net974),
    .B(_1078_));
 sg13g2_nor2_1 _5475_ (.A(_1473_),
    .B(_1625_),
    .Y(_1626_));
 sg13g2_nor2_1 _5476_ (.A(_1080_),
    .B(_1360_),
    .Y(_1627_));
 sg13g2_xnor2_1 _5477_ (.Y(_1628_),
    .A(_1626_),
    .B(_1627_));
 sg13g2_o21ai_1 _5478_ (.B1(_1369_),
    .Y(_1629_),
    .A1(_1380_),
    .A2(_1628_));
 sg13g2_and2_1 _5479_ (.A(_1475_),
    .B(_1477_),
    .X(_1630_));
 sg13g2_nor3_1 _5480_ (.A(_1047_),
    .B(_1202_),
    .C(_1630_),
    .Y(_1631_));
 sg13g2_a21oi_1 _5481_ (.A1(net971),
    .A2(_1475_),
    .Y(_1632_),
    .B1(_1631_));
 sg13g2_o21ai_1 _5482_ (.B1(_1358_),
    .Y(_1633_),
    .A1(_1369_),
    .A2(_1632_));
 sg13g2_nand2b_1 _5483_ (.Y(_1634_),
    .B(_1629_),
    .A_N(_1633_));
 sg13g2_or3_1 _5484_ (.A(\vgademo.h_count[10] ),
    .B(_3111_),
    .C(_1482_),
    .X(_1635_));
 sg13g2_nand3_1 _5485_ (.B(net859),
    .C(_1635_),
    .A(_0061_),
    .Y(_1636_));
 sg13g2_o21ai_1 _5486_ (.B1(_1636_),
    .Y(_1637_),
    .A1(_3174_),
    .A2(net859));
 sg13g2_xor2_1 _5487_ (.B(_1637_),
    .A(_1634_),
    .X(_1638_));
 sg13g2_xor2_1 _5488_ (.B(_1630_),
    .A(net975),
    .X(_1639_));
 sg13g2_xnor2_1 _5489_ (.Y(_1640_),
    .A(_1472_),
    .B(_1625_));
 sg13g2_a221oi_1 _5490_ (.B2(net888),
    .C1(_1364_),
    .B1(_1640_),
    .A1(_1368_),
    .Y(_1641_),
    .A2(_1639_));
 sg13g2_o21ai_1 _5491_ (.B1(\vgademo.h_count[10] ),
    .Y(_1642_),
    .A1(_3111_),
    .A2(_1482_));
 sg13g2_nand3_1 _5492_ (.B(_1635_),
    .C(_1642_),
    .A(net859),
    .Y(_1643_));
 sg13g2_o21ai_1 _5493_ (.B1(_1643_),
    .Y(_1644_),
    .A1(_0032_),
    .A2(net859));
 sg13g2_a22oi_1 _5494_ (.Y(_1645_),
    .B1(_1641_),
    .B2(_1644_),
    .A2(_1638_),
    .A1(_1624_));
 sg13g2_or2_1 _5495_ (.X(_1646_),
    .B(_1644_),
    .A(_1641_));
 sg13g2_and2_1 _5496_ (.A(_1638_),
    .B(_1646_),
    .X(_1647_));
 sg13g2_a21oi_1 _5497_ (.A1(_1485_),
    .A2(_1488_),
    .Y(_1648_),
    .B1(_1647_));
 sg13g2_mux2_1 _5498_ (.A0(_1648_),
    .A1(_1647_),
    .S(_1645_),
    .X(_1649_));
 sg13g2_o21ai_1 _5499_ (.B1(_1649_),
    .Y(_1650_),
    .A1(_1611_),
    .A2(_1623_));
 sg13g2_a21oi_1 _5500_ (.A1(_1560_),
    .A2(_1603_),
    .Y(_1651_),
    .B1(_1650_));
 sg13g2_a21o_1 _5501_ (.A2(_1603_),
    .A1(_1560_),
    .B1(_1650_),
    .X(_1652_));
 sg13g2_xnor2_1 _5502_ (.Y(_1653_),
    .A(net957),
    .B(\vgademo.b_cos[10] ));
 sg13g2_nand2b_1 _5503_ (.Y(_1654_),
    .B(\vgademo.v_count[3] ),
    .A_N(net958));
 sg13g2_nand2_1 _5504_ (.Y(_1655_),
    .A(_3102_),
    .B(net958));
 sg13g2_o21ai_1 _5505_ (.B1(_3100_),
    .Y(_1656_),
    .A1(net959),
    .A2(_1328_));
 sg13g2_a22oi_1 _5506_ (.Y(_1657_),
    .B1(_1330_),
    .B2(_1656_),
    .A2(_3145_),
    .A1(net968));
 sg13g2_o21ai_1 _5507_ (.B1(_1655_),
    .Y(_1658_),
    .A1(net968),
    .A2(_3145_));
 sg13g2_o21ai_1 _5508_ (.B1(_1654_),
    .Y(_1659_),
    .A1(_1657_),
    .A2(_1658_));
 sg13g2_xnor2_1 _5509_ (.Y(_1660_),
    .A(_0063_),
    .B(_1653_));
 sg13g2_o21ai_1 _5510_ (.B1(_1659_),
    .Y(_1661_),
    .A1(net967),
    .A2(net957));
 sg13g2_o21ai_1 _5511_ (.B1(_1661_),
    .Y(_1662_),
    .A1(_3104_),
    .A2(_3147_));
 sg13g2_a22oi_1 _5512_ (.Y(_1663_),
    .B1(_1660_),
    .B2(_1662_),
    .A2(_1653_),
    .A1(net965));
 sg13g2_nor2_1 _5513_ (.A(net957),
    .B(\vgademo.b_cos[11] ),
    .Y(_1664_));
 sg13g2_a21oi_2 _5514_ (.B1(_1664_),
    .Y(_1665_),
    .A2(_1598_),
    .A1(net957));
 sg13g2_xnor2_1 _5515_ (.Y(_1666_),
    .A(_3123_),
    .B(_1665_));
 sg13g2_a22oi_1 _5516_ (.Y(_1667_),
    .B1(_1665_),
    .B2(net964),
    .A2(_3124_),
    .A1(net963));
 sg13g2_o21ai_1 _5517_ (.B1(_1667_),
    .Y(_1668_),
    .A1(_1663_),
    .A2(_1666_));
 sg13g2_or2_1 _5518_ (.X(_1669_),
    .B(_1597_),
    .A(_3147_));
 sg13g2_nand3_1 _5519_ (.B(_0019_),
    .C(_1669_),
    .A(net963),
    .Y(_1670_));
 sg13g2_o21ai_1 _5520_ (.B1(_1670_),
    .Y(_1671_),
    .A1(_0019_),
    .A2(_1669_));
 sg13g2_nor2_1 _5521_ (.A(_3224_),
    .B(_1669_),
    .Y(_1672_));
 sg13g2_o21ai_1 _5522_ (.B1(_3147_),
    .Y(_1673_),
    .A1(net967),
    .A2(_1659_));
 sg13g2_a22oi_1 _5523_ (.Y(_1674_),
    .B1(_1659_),
    .B2(net967),
    .A2(net956),
    .A1(net965));
 sg13g2_xnor2_1 _5524_ (.Y(_1675_),
    .A(_0017_),
    .B(_1598_));
 sg13g2_a221oi_1 _5525_ (.B2(_1674_),
    .C1(_1675_),
    .B1(_1673_),
    .A1(_3103_),
    .Y(_1676_),
    .A2(_3148_));
 sg13g2_a221oi_1 _5526_ (.B2(net964),
    .C1(_1676_),
    .B1(_1599_),
    .A1(net963),
    .Y(_1677_),
    .A2(_1597_));
 sg13g2_o21ai_1 _5527_ (.B1(_0019_),
    .Y(_1678_),
    .A1(net963),
    .A2(_1597_));
 sg13g2_o21ai_1 _5528_ (.B1(_0022_),
    .Y(_1679_),
    .A1(_1677_),
    .A2(_1678_));
 sg13g2_a21oi_1 _5529_ (.A1(_3222_),
    .A2(_1679_),
    .Y(_1680_),
    .B1(_1672_));
 sg13g2_a21oi_2 _5530_ (.B1(_1680_),
    .Y(_1681_),
    .A2(_1671_),
    .A1(_1668_));
 sg13g2_inv_1 _5531_ (.Y(_1682_),
    .A(_1681_));
 sg13g2_nor2_1 _5532_ (.A(net829),
    .B(_1682_),
    .Y(_1683_));
 sg13g2_nand2_1 _5533_ (.Y(_1684_),
    .A(net832),
    .B(_1681_));
 sg13g2_nand2_1 _5534_ (.Y(_1685_),
    .A(_1345_),
    .B(_1444_));
 sg13g2_nand2_1 _5535_ (.Y(_1686_),
    .A(net845),
    .B(_1447_));
 sg13g2_xnor2_1 _5536_ (.Y(_1687_),
    .A(_1344_),
    .B(_1445_));
 sg13g2_o21ai_1 _5537_ (.B1(_1685_),
    .Y(_1688_),
    .A1(_1686_),
    .A2(_1687_));
 sg13g2_xnor2_1 _5538_ (.Y(_1689_),
    .A(_1342_),
    .B(_1440_));
 sg13g2_xnor2_1 _5539_ (.Y(_1690_),
    .A(_1688_),
    .B(_1689_));
 sg13g2_inv_1 _5540_ (.Y(_1691_),
    .A(_1690_));
 sg13g2_nand3_1 _5541_ (.B(_1681_),
    .C(_1690_),
    .A(net832),
    .Y(_1692_));
 sg13g2_and2_1 _5542_ (.A(net861),
    .B(_1692_),
    .X(_1693_));
 sg13g2_nand2_2 _5543_ (.Y(_1694_),
    .A(_1294_),
    .B(_1692_));
 sg13g2_nand2_1 _5544_ (.Y(_1695_),
    .A(\vgademo.plane_du[8] ),
    .B(_1665_));
 sg13g2_xnor2_1 _5545_ (.Y(_1696_),
    .A(_0053_),
    .B(_1653_));
 sg13g2_nand2b_1 _5546_ (.Y(_1697_),
    .B(net958),
    .A_N(\vgademo.plane_du[5] ));
 sg13g2_nand2b_1 _5547_ (.Y(_1698_),
    .B(\vgademo.plane_du[5] ),
    .A_N(net958));
 sg13g2_a221oi_1 _5548_ (.B2(\vgademo.plane_du[3] ),
    .C1(_1325_),
    .B1(_1324_),
    .A1(_3145_),
    .Y(_1699_),
    .A2(\vgademo.plane_du[4] ));
 sg13g2_o21ai_1 _5549_ (.B1(_1697_),
    .Y(_1700_),
    .A1(_3145_),
    .A2(\vgademo.plane_du[4] ));
 sg13g2_o21ai_1 _5550_ (.B1(_1698_),
    .Y(_1701_),
    .A1(_1699_),
    .A2(_1700_));
 sg13g2_and2_1 _5551_ (.A(\vgademo.plane_du[6] ),
    .B(_1701_),
    .X(_1702_));
 sg13g2_or2_1 _5552_ (.X(_1703_),
    .B(_1701_),
    .A(\vgademo.plane_du[6] ));
 sg13g2_a21o_1 _5553_ (.A2(_1703_),
    .A1(net957),
    .B1(_1702_),
    .X(_1704_));
 sg13g2_a22oi_1 _5554_ (.Y(_1705_),
    .B1(_1696_),
    .B2(_1704_),
    .A2(_1653_),
    .A1(\vgademo.plane_du[7] ));
 sg13g2_xor2_1 _5555_ (.B(_1665_),
    .A(_0054_),
    .X(_1706_));
 sg13g2_o21ai_1 _5556_ (.B1(_1695_),
    .Y(_1707_),
    .A1(_1705_),
    .A2(_1706_));
 sg13g2_nand3_1 _5557_ (.B(_1669_),
    .C(_1707_),
    .A(net950),
    .Y(_1708_));
 sg13g2_a221oi_1 _5558_ (.B2(_3147_),
    .C1(_1702_),
    .B1(_1703_),
    .A1(net956),
    .Y(_1709_),
    .A2(\vgademo.plane_du[7] ));
 sg13g2_xnor2_1 _5559_ (.Y(_1710_),
    .A(_0054_),
    .B(_1599_));
 sg13g2_o21ai_1 _5560_ (.B1(_1710_),
    .Y(_1711_),
    .A1(net956),
    .A2(\vgademo.plane_du[7] ));
 sg13g2_a22oi_1 _5561_ (.Y(_1712_),
    .B1(_1599_),
    .B2(\vgademo.plane_du[8] ),
    .A2(_1597_),
    .A1(net950));
 sg13g2_o21ai_1 _5562_ (.B1(_1712_),
    .Y(_1713_),
    .A1(_1709_),
    .A2(_1711_));
 sg13g2_or2_1 _5563_ (.X(_1714_),
    .B(_1597_),
    .A(net950));
 sg13g2_and3_2 _5564_ (.X(_1715_),
    .A(_1708_),
    .B(_1713_),
    .C(_1714_));
 sg13g2_nand3_1 _5565_ (.B(_1713_),
    .C(_1714_),
    .A(_1708_),
    .Y(_1716_));
 sg13g2_nand2_1 _5566_ (.Y(_1717_),
    .A(net831),
    .B(net853));
 sg13g2_and2_1 _5567_ (.A(net980),
    .B(\vgademo.plane_du[8] ),
    .X(_1718_));
 sg13g2_and2_1 _5568_ (.A(net990),
    .B(\vgademo.plane_du[5] ),
    .X(_1719_));
 sg13g2_nand2_1 _5569_ (.Y(_1720_),
    .A(net990),
    .B(\vgademo.plane_du[5] ));
 sg13g2_nand2_1 _5570_ (.Y(_1721_),
    .A(net994),
    .B(\vgademo.plane_du[4] ));
 sg13g2_nor2_1 _5571_ (.A(net990),
    .B(\vgademo.plane_du[5] ),
    .Y(_1722_));
 sg13g2_or3_1 _5572_ (.A(_1719_),
    .B(_1721_),
    .C(_1722_),
    .X(_1723_));
 sg13g2_xnor2_1 _5573_ (.Y(_1724_),
    .A(net986),
    .B(\vgademo.plane_du[6] ));
 sg13g2_a21oi_1 _5574_ (.A1(_1720_),
    .A2(_1723_),
    .Y(_1725_),
    .B1(_1724_));
 sg13g2_a21oi_1 _5575_ (.A1(net986),
    .A2(\vgademo.plane_du[6] ),
    .Y(_1726_),
    .B1(_1725_));
 sg13g2_xor2_1 _5576_ (.B(\vgademo.plane_du[7] ),
    .A(net983),
    .X(_1727_));
 sg13g2_nand2b_1 _5577_ (.Y(_1728_),
    .B(_1727_),
    .A_N(_1726_));
 sg13g2_o21ai_1 _5578_ (.B1(_1728_),
    .Y(_1729_),
    .A1(_3118_),
    .A2(_3163_));
 sg13g2_xor2_1 _5579_ (.B(\vgademo.plane_du[8] ),
    .A(net980),
    .X(_1730_));
 sg13g2_a21o_1 _5580_ (.A2(_1730_),
    .A1(_1729_),
    .B1(_1718_),
    .X(_1731_));
 sg13g2_and2_1 _5581_ (.A(net978),
    .B(net950),
    .X(_1732_));
 sg13g2_xor2_1 _5582_ (.B(net950),
    .A(net978),
    .X(_1733_));
 sg13g2_xnor2_1 _5583_ (.Y(_1734_),
    .A(_1731_),
    .B(_1733_));
 sg13g2_and2_1 _5584_ (.A(\vgademo.a_cos[12] ),
    .B(\vgademo.plane_u[17] ),
    .X(_1735_));
 sg13g2_and2_1 _5585_ (.A(\vgademo.a_cos[11] ),
    .B(\vgademo.plane_u[16] ),
    .X(_1736_));
 sg13g2_nand2_1 _5586_ (.Y(_1737_),
    .A(\vgademo.a_cos[10] ),
    .B(\vgademo.plane_u[15] ));
 sg13g2_nor2_1 _5587_ (.A(\vgademo.a_cos[10] ),
    .B(\vgademo.plane_u[15] ),
    .Y(_1738_));
 sg13g2_xor2_1 _5588_ (.B(\vgademo.plane_u[15] ),
    .A(\vgademo.a_cos[10] ),
    .X(_1739_));
 sg13g2_nand2_1 _5589_ (.Y(_1740_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.plane_u[12] ));
 sg13g2_xnor2_1 _5590_ (.Y(_1741_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.plane_u[12] ));
 sg13g2_or2_1 _5591_ (.X(_1742_),
    .B(\vgademo.plane_u[10] ),
    .A(\vgademo.a_cos[5] ));
 sg13g2_nand3_1 _5592_ (.B(\vgademo.plane_u[9] ),
    .C(_1742_),
    .A(\vgademo.a_cos[4] ),
    .Y(_1743_));
 sg13g2_a22oi_1 _5593_ (.Y(_1744_),
    .B1(\vgademo.plane_u[11] ),
    .B2(\vgademo.a_cos[6] ),
    .A2(\vgademo.plane_u[10] ),
    .A1(\vgademo.a_cos[5] ));
 sg13g2_a22oi_1 _5594_ (.Y(_1745_),
    .B1(_1743_),
    .B2(_1744_),
    .A2(_3167_),
    .A1(_3141_));
 sg13g2_nand2b_1 _5595_ (.Y(_1746_),
    .B(_1745_),
    .A_N(_1741_));
 sg13g2_xnor2_1 _5596_ (.Y(_1747_),
    .A(\vgademo.a_cos[8] ),
    .B(\vgademo.plane_u[13] ));
 sg13g2_a21oi_2 _5597_ (.B1(_1747_),
    .Y(_1748_),
    .A2(_1746_),
    .A1(_1740_));
 sg13g2_a21o_1 _5598_ (.A2(\vgademo.plane_u[13] ),
    .A1(\vgademo.a_cos[8] ),
    .B1(_1748_),
    .X(_1749_));
 sg13g2_a21o_1 _5599_ (.A2(\vgademo.plane_u[14] ),
    .A1(\vgademo.a_cos[9] ),
    .B1(_1749_),
    .X(_1750_));
 sg13g2_o21ai_1 _5600_ (.B1(_1750_),
    .Y(_1751_),
    .A1(\vgademo.a_cos[9] ),
    .A2(\vgademo.plane_u[14] ));
 sg13g2_o21ai_1 _5601_ (.B1(_1737_),
    .Y(_1752_),
    .A1(_1738_),
    .A2(_1751_));
 sg13g2_xor2_1 _5602_ (.B(\vgademo.plane_u[16] ),
    .A(\vgademo.a_cos[11] ),
    .X(_1753_));
 sg13g2_a21o_1 _5603_ (.A2(_1753_),
    .A1(_1752_),
    .B1(_1736_),
    .X(_1754_));
 sg13g2_xor2_1 _5604_ (.B(\vgademo.plane_u[17] ),
    .A(\vgademo.a_cos[12] ),
    .X(_1755_));
 sg13g2_a21o_1 _5605_ (.A2(_1755_),
    .A1(_1754_),
    .B1(_1735_),
    .X(_1756_));
 sg13g2_xor2_1 _5606_ (.B(\vgademo.plane_u[18] ),
    .A(\vgademo.a_cos[13] ),
    .X(_1757_));
 sg13g2_xnor2_1 _5607_ (.Y(_1758_),
    .A(_1756_),
    .B(_1757_));
 sg13g2_nor2_1 _5608_ (.A(_1734_),
    .B(_1758_),
    .Y(_1759_));
 sg13g2_xor2_1 _5609_ (.B(_1758_),
    .A(_1734_),
    .X(_1760_));
 sg13g2_xnor2_1 _5610_ (.Y(_1761_),
    .A(_1729_),
    .B(_1730_));
 sg13g2_xnor2_1 _5611_ (.Y(_1762_),
    .A(_1754_),
    .B(_1755_));
 sg13g2_xor2_1 _5612_ (.B(_1762_),
    .A(_1761_),
    .X(_1763_));
 sg13g2_xnor2_1 _5613_ (.Y(_1764_),
    .A(_1752_),
    .B(_1753_));
 sg13g2_inv_1 _5614_ (.Y(_1765_),
    .A(_1764_));
 sg13g2_xnor2_1 _5615_ (.Y(_1766_),
    .A(_1726_),
    .B(_1727_));
 sg13g2_xnor2_1 _5616_ (.Y(_1767_),
    .A(net1054),
    .B(_1766_));
 sg13g2_xor2_1 _5617_ (.B(_1764_),
    .A(net1061),
    .X(_1768_));
 sg13g2_nand3_1 _5618_ (.B(_1767_),
    .C(_1768_),
    .A(net1041),
    .Y(_1769_));
 sg13g2_xnor2_1 _5619_ (.Y(_1770_),
    .A(_3097_),
    .B(_1763_));
 sg13g2_xnor2_1 _5620_ (.Y(_1771_),
    .A(net949),
    .B(_1760_));
 sg13g2_nor3_1 _5621_ (.A(_1769_),
    .B(_1770_),
    .C(_1771_),
    .Y(_1772_));
 sg13g2_inv_1 _5622_ (.Y(_1773_),
    .A(_1772_));
 sg13g2_xor2_1 _5623_ (.B(_1766_),
    .A(_1764_),
    .X(_1774_));
 sg13g2_nand3_1 _5624_ (.B(_1766_),
    .C(_1773_),
    .A(_1764_),
    .Y(_1775_));
 sg13g2_nor3_1 _5625_ (.A(_1764_),
    .B(_1766_),
    .C(net844),
    .Y(_1776_));
 sg13g2_nor2_2 _5626_ (.A(net844),
    .B(_1774_),
    .Y(_1777_));
 sg13g2_inv_1 _5627_ (.Y(_1778_),
    .A(_1777_));
 sg13g2_o21ai_1 _5628_ (.B1(_1721_),
    .Y(_1779_),
    .A1(_1719_),
    .A2(_1722_));
 sg13g2_nand3_1 _5629_ (.B(_1777_),
    .C(_1779_),
    .A(_1723_),
    .Y(_1780_));
 sg13g2_nand2_1 _5630_ (.Y(_1781_),
    .A(_1765_),
    .B(_1766_));
 sg13g2_nand3_1 _5631_ (.B(_1765_),
    .C(_1766_),
    .A(_1763_),
    .Y(_1782_));
 sg13g2_o21ai_1 _5632_ (.B1(_1782_),
    .Y(_1783_),
    .A1(_1761_),
    .A2(_1762_));
 sg13g2_a21oi_1 _5633_ (.A1(_1760_),
    .A2(_1783_),
    .Y(_1784_),
    .B1(_1759_));
 sg13g2_a21o_1 _5634_ (.A2(\vgademo.plane_u[18] ),
    .A1(\vgademo.a_cos[13] ),
    .B1(_1756_),
    .X(_1785_));
 sg13g2_o21ai_1 _5635_ (.B1(_1785_),
    .Y(_1786_),
    .A1(\vgademo.a_cos[13] ),
    .A2(\vgademo.plane_u[18] ));
 sg13g2_a21oi_1 _5636_ (.A1(_1731_),
    .A2(_1733_),
    .Y(_1787_),
    .B1(_1732_));
 sg13g2_xor2_1 _5637_ (.B(\vgademo.a_cos[14] ),
    .A(net975),
    .X(_1788_));
 sg13g2_xor2_1 _5638_ (.B(\vgademo.plane_u[19] ),
    .A(\vgademo.plane_du[10] ),
    .X(_1789_));
 sg13g2_xnor2_1 _5639_ (.Y(_1790_),
    .A(_1788_),
    .B(_1789_));
 sg13g2_xnor2_1 _5640_ (.Y(_1791_),
    .A(_1787_),
    .B(_1790_));
 sg13g2_xnor2_1 _5641_ (.Y(_1792_),
    .A(_1786_),
    .B(_1791_));
 sg13g2_xnor2_1 _5642_ (.Y(_1793_),
    .A(_1784_),
    .B(_1792_));
 sg13g2_xnor2_1 _5643_ (.Y(_1794_),
    .A(_1760_),
    .B(_1783_));
 sg13g2_xor2_1 _5644_ (.B(_1781_),
    .A(_1763_),
    .X(_1795_));
 sg13g2_o21ai_1 _5645_ (.B1(_1795_),
    .Y(_1796_),
    .A1(_3256_),
    .A2(_1774_));
 sg13g2_o21ai_1 _5646_ (.B1(net1054),
    .Y(_1797_),
    .A1(net1057),
    .A2(_1774_));
 sg13g2_nor2_1 _5647_ (.A(\vgademo.audio_songpos[4] ),
    .B(_1794_),
    .Y(_1798_));
 sg13g2_a21oi_1 _5648_ (.A1(_1796_),
    .A2(_1797_),
    .Y(_1799_),
    .B1(_1798_));
 sg13g2_a221oi_1 _5649_ (.B2(\vgademo.audio_songpos[4] ),
    .C1(_1799_),
    .B1(_1794_),
    .A1(\vgademo.audio_songpos[5] ),
    .Y(_1800_),
    .A2(_1793_));
 sg13g2_o21ai_1 _5650_ (.B1(_3288_),
    .Y(_1801_),
    .A1(\vgademo.audio_songpos[5] ),
    .A2(_1793_));
 sg13g2_nor2_2 _5651_ (.A(_1800_),
    .B(_1801_),
    .Y(_1802_));
 sg13g2_nor2_2 _5652_ (.A(net844),
    .B(_1802_),
    .Y(_1803_));
 sg13g2_inv_1 _5653_ (.Y(_1804_),
    .A(_1803_));
 sg13g2_a21oi_2 _5654_ (.B1(_1802_),
    .Y(_1805_),
    .A2(net844),
    .A1(_0062_));
 sg13g2_nand2_1 _5655_ (.Y(_1806_),
    .A(_1780_),
    .B(_1805_));
 sg13g2_o21ai_1 _5656_ (.B1(_1806_),
    .Y(_1807_),
    .A1(net828),
    .A2(net852));
 sg13g2_a21oi_2 _5657_ (.B1(_1802_),
    .Y(_1808_),
    .A2(net844),
    .A1(_0055_));
 sg13g2_nand2_2 _5658_ (.Y(_1809_),
    .A(_1775_),
    .B(_1808_));
 sg13g2_nand3_1 _5659_ (.B(net853),
    .C(_1809_),
    .A(net830),
    .Y(_1810_));
 sg13g2_nand3_1 _5660_ (.B(_1807_),
    .C(_1810_),
    .A(net854),
    .Y(_1811_));
 sg13g2_nand2_1 _5661_ (.Y(_1812_),
    .A(net1066),
    .B(net979));
 sg13g2_nand2_1 _5662_ (.Y(_1813_),
    .A(net981),
    .B(net1065));
 sg13g2_nand2_1 _5663_ (.Y(_1814_),
    .A(net979),
    .B(net1065));
 sg13g2_nand2_1 _5664_ (.Y(_1815_),
    .A(net1066),
    .B(net981));
 sg13g2_xor2_1 _5665_ (.B(_1815_),
    .A(_1814_),
    .X(_1816_));
 sg13g2_nand2_1 _5666_ (.Y(_1817_),
    .A(\vgademo.linelfsr[8] ),
    .B(_1816_));
 sg13g2_o21ai_1 _5667_ (.B1(_1817_),
    .Y(_1818_),
    .A1(_1814_),
    .A2(_1815_));
 sg13g2_nand2_1 _5668_ (.Y(_1819_),
    .A(net1066),
    .B(net976));
 sg13g2_nand2_1 _5669_ (.Y(_1820_),
    .A(net976),
    .B(net1065));
 sg13g2_xor2_1 _5670_ (.B(_1820_),
    .A(_1812_),
    .X(_1821_));
 sg13g2_nand2_1 _5671_ (.Y(_1822_),
    .A(\vgademo.linelfsr[9] ),
    .B(_1821_));
 sg13g2_xnor2_1 _5672_ (.Y(_1823_),
    .A(\vgademo.linelfsr[9] ),
    .B(_1821_));
 sg13g2_nor2b_1 _5673_ (.A(_1823_),
    .B_N(_1818_),
    .Y(_1824_));
 sg13g2_nand2b_1 _5674_ (.Y(_1825_),
    .B(_1823_),
    .A_N(_1818_));
 sg13g2_nand2b_1 _5675_ (.Y(_1826_),
    .B(_1825_),
    .A_N(_1824_));
 sg13g2_a21o_1 _5676_ (.A2(_1825_),
    .A1(net973),
    .B1(_1824_),
    .X(_1827_));
 sg13g2_o21ai_1 _5677_ (.B1(_1822_),
    .Y(_1828_),
    .A1(_1812_),
    .A2(_1820_));
 sg13g2_nand2_1 _5678_ (.Y(_1829_),
    .A(net972),
    .B(net1065));
 sg13g2_xor2_1 _5679_ (.B(_1829_),
    .A(_1819_),
    .X(_1830_));
 sg13g2_nand2_1 _5680_ (.Y(_1831_),
    .A(\vgademo.linelfsr[10] ),
    .B(_1830_));
 sg13g2_xnor2_1 _5681_ (.Y(_1832_),
    .A(\vgademo.linelfsr[10] ),
    .B(_1830_));
 sg13g2_nand2b_1 _5682_ (.Y(_1833_),
    .B(_1828_),
    .A_N(_1832_));
 sg13g2_xor2_1 _5683_ (.B(_1832_),
    .A(_1828_),
    .X(_1834_));
 sg13g2_xnor2_1 _5684_ (.Y(_1835_),
    .A(_3114_),
    .B(_1834_));
 sg13g2_nor2b_1 _5685_ (.A(_1835_),
    .B_N(_1827_),
    .Y(_1836_));
 sg13g2_xor2_1 _5686_ (.B(_1835_),
    .A(_1827_),
    .X(_1837_));
 sg13g2_nand2_1 _5687_ (.Y(_1838_),
    .A(net984),
    .B(net1064));
 sg13g2_nand2_1 _5688_ (.Y(_1839_),
    .A(net1067),
    .B(net984));
 sg13g2_xor2_1 _5689_ (.B(_1839_),
    .A(_1813_),
    .X(_1840_));
 sg13g2_nand2_1 _5690_ (.Y(_1841_),
    .A(\vgademo.linelfsr[7] ),
    .B(_1840_));
 sg13g2_o21ai_1 _5691_ (.B1(_1841_),
    .Y(_1842_),
    .A1(_1813_),
    .A2(_1839_));
 sg13g2_xnor2_1 _5692_ (.Y(_1843_),
    .A(\vgademo.linelfsr[8] ),
    .B(_1816_));
 sg13g2_nand2b_1 _5693_ (.Y(_1844_),
    .B(_1842_),
    .A_N(_1843_));
 sg13g2_xor2_1 _5694_ (.B(_1843_),
    .A(_1842_),
    .X(_1845_));
 sg13g2_o21ai_1 _5695_ (.B1(_1844_),
    .Y(_1846_),
    .A1(_3116_),
    .A2(_1845_));
 sg13g2_xor2_1 _5696_ (.B(_1826_),
    .A(net973),
    .X(_1847_));
 sg13g2_nand2b_1 _5697_ (.Y(_1848_),
    .B(_1846_),
    .A_N(_1847_));
 sg13g2_nor2b_1 _5698_ (.A(_1846_),
    .B_N(_1847_),
    .Y(_1849_));
 sg13g2_nand2_1 _5699_ (.Y(_1850_),
    .A(net1067),
    .B(net989));
 sg13g2_xor2_1 _5700_ (.B(_1850_),
    .A(_1838_),
    .X(_1851_));
 sg13g2_nand2_1 _5701_ (.Y(_1852_),
    .A(\vgademo.linelfsr[6] ),
    .B(_1851_));
 sg13g2_o21ai_1 _5702_ (.B1(_1852_),
    .Y(_1853_),
    .A1(_1838_),
    .A2(_1850_));
 sg13g2_xnor2_1 _5703_ (.Y(_1854_),
    .A(\vgademo.linelfsr[7] ),
    .B(_1840_));
 sg13g2_nand2b_1 _5704_ (.Y(_1855_),
    .B(_1853_),
    .A_N(_1854_));
 sg13g2_xor2_1 _5705_ (.B(_1854_),
    .A(_1853_),
    .X(_1856_));
 sg13g2_o21ai_1 _5706_ (.B1(_1855_),
    .Y(_1857_),
    .A1(_3117_),
    .A2(_1856_));
 sg13g2_xnor2_1 _5707_ (.Y(_1858_),
    .A(_3116_),
    .B(_1845_));
 sg13g2_nor2b_1 _5708_ (.A(_1858_),
    .B_N(_1857_),
    .Y(_1859_));
 sg13g2_xnor2_1 _5709_ (.Y(_1860_),
    .A(_1857_),
    .B(_1858_));
 sg13g2_and4_1 _5710_ (.A(net1067),
    .B(net991),
    .C(net989),
    .D(net1064),
    .X(_1861_));
 sg13g2_a22oi_1 _5711_ (.Y(_1862_),
    .B1(net989),
    .B2(net1064),
    .A2(net991),
    .A1(net1067));
 sg13g2_nor3_1 _5712_ (.A(_3177_),
    .B(_1861_),
    .C(_1862_),
    .Y(_1863_));
 sg13g2_or2_1 _5713_ (.X(_1864_),
    .B(_1863_),
    .A(_1861_));
 sg13g2_xnor2_1 _5714_ (.Y(_1865_),
    .A(\vgademo.linelfsr[6] ),
    .B(_1851_));
 sg13g2_nand2b_1 _5715_ (.Y(_1866_),
    .B(_1864_),
    .A_N(_1865_));
 sg13g2_xor2_1 _5716_ (.B(_1865_),
    .A(_1864_),
    .X(_1867_));
 sg13g2_o21ai_1 _5717_ (.B1(_1866_),
    .Y(_1868_),
    .A1(_3118_),
    .A2(_1867_));
 sg13g2_xnor2_1 _5718_ (.Y(_1869_),
    .A(_3117_),
    .B(_1856_));
 sg13g2_nand2b_1 _5719_ (.Y(_1870_),
    .B(_1868_),
    .A_N(_1869_));
 sg13g2_nand2b_1 _5720_ (.Y(_1871_),
    .B(_1869_),
    .A_N(_1868_));
 sg13g2_inv_1 _5721_ (.Y(_1872_),
    .A(_1871_));
 sg13g2_and3_1 _5722_ (.X(_1873_),
    .A(net991),
    .B(net1064),
    .C(\vgademo.linelfsr[4] ));
 sg13g2_a21oi_1 _5723_ (.A1(net991),
    .A2(net1064),
    .Y(_1874_),
    .B1(\vgademo.linelfsr[4] ));
 sg13g2_nor2_1 _5724_ (.A(_1873_),
    .B(_1874_),
    .Y(_1875_));
 sg13g2_a21o_1 _5725_ (.A2(_1875_),
    .A1(net989),
    .B1(_1873_),
    .X(_1876_));
 sg13g2_o21ai_1 _5726_ (.B1(_3177_),
    .Y(_1877_),
    .A1(_1861_),
    .A2(_1862_));
 sg13g2_nand2b_1 _5727_ (.Y(_1878_),
    .B(_1877_),
    .A_N(_1863_));
 sg13g2_nor2b_1 _5728_ (.A(_1878_),
    .B_N(_1876_),
    .Y(_1879_));
 sg13g2_xnor2_1 _5729_ (.Y(_1880_),
    .A(_1876_),
    .B(_1878_));
 sg13g2_a21o_1 _5730_ (.A2(_1880_),
    .A1(net984),
    .B1(_1879_),
    .X(_1881_));
 sg13g2_xnor2_1 _5731_ (.Y(_1882_),
    .A(_3118_),
    .B(_1867_));
 sg13g2_nor2b_1 _5732_ (.A(_1882_),
    .B_N(_1881_),
    .Y(_1883_));
 sg13g2_xnor2_1 _5733_ (.Y(_1884_),
    .A(net984),
    .B(_1880_));
 sg13g2_xnor2_1 _5734_ (.Y(_1885_),
    .A(net989),
    .B(_1875_));
 sg13g2_nand2_1 _5735_ (.Y(_1886_),
    .A(\vgademo.linelfsr[3] ),
    .B(net991));
 sg13g2_nor2_1 _5736_ (.A(_1885_),
    .B(_1886_),
    .Y(_1887_));
 sg13g2_nor2b_1 _5737_ (.A(_1884_),
    .B_N(_1887_),
    .Y(_1888_));
 sg13g2_xor2_1 _5738_ (.B(_1882_),
    .A(_1881_),
    .X(_1889_));
 sg13g2_inv_1 _5739_ (.Y(_1890_),
    .A(_1889_));
 sg13g2_a21oi_1 _5740_ (.A1(_1888_),
    .A2(_1890_),
    .Y(_1891_),
    .B1(_1883_));
 sg13g2_a21oi_1 _5741_ (.A1(_1870_),
    .A2(_1891_),
    .Y(_1892_),
    .B1(_1872_));
 sg13g2_a21oi_1 _5742_ (.A1(_1860_),
    .A2(_1892_),
    .Y(_1893_),
    .B1(_1859_));
 sg13g2_a21oi_1 _5743_ (.A1(_1848_),
    .A2(_1893_),
    .Y(_1894_),
    .B1(_1849_));
 sg13g2_nor2b_1 _5744_ (.A(_1837_),
    .B_N(_1894_),
    .Y(_1895_));
 sg13g2_nor2_1 _5745_ (.A(_1836_),
    .B(_1895_),
    .Y(_1896_));
 sg13g2_o21ai_1 _5746_ (.B1(_1833_),
    .Y(_1897_),
    .A1(_3114_),
    .A2(_1834_));
 sg13g2_o21ai_1 _5747_ (.B1(_1831_),
    .Y(_1898_),
    .A1(_1819_),
    .A2(_1829_));
 sg13g2_nand2_1 _5748_ (.Y(_1899_),
    .A(net1066),
    .B(net970));
 sg13g2_nor2_1 _5749_ (.A(_1829_),
    .B(_1899_),
    .Y(_1900_));
 sg13g2_a22oi_1 _5750_ (.Y(_1901_),
    .B1(net1065),
    .B2(net970),
    .A2(net972),
    .A1(net1066));
 sg13g2_nor2_1 _5751_ (.A(_1900_),
    .B(_1901_),
    .Y(_1902_));
 sg13g2_xnor2_1 _5752_ (.Y(_1903_),
    .A(\vgademo.linelfsr[11] ),
    .B(_1902_));
 sg13g2_nand2b_1 _5753_ (.Y(_1904_),
    .B(_1898_),
    .A_N(_1903_));
 sg13g2_xor2_1 _5754_ (.B(_1903_),
    .A(_1898_),
    .X(_1905_));
 sg13g2_xnor2_1 _5755_ (.Y(_1906_),
    .A(_3113_),
    .B(_1905_));
 sg13g2_nand2b_1 _5756_ (.Y(_1907_),
    .B(_1897_),
    .A_N(_1906_));
 sg13g2_xor2_1 _5757_ (.B(_1906_),
    .A(_1897_),
    .X(_1908_));
 sg13g2_xor2_1 _5758_ (.B(_1908_),
    .A(_1896_),
    .X(_1909_));
 sg13g2_xnor2_1 _5759_ (.Y(_1910_),
    .A(\vgademo.linelfsr[3] ),
    .B(net991));
 sg13g2_inv_1 _5760_ (.Y(_1911_),
    .A(_1910_));
 sg13g2_nand2b_1 _5761_ (.Y(_1912_),
    .B(_1911_),
    .A_N(_1885_));
 sg13g2_nor2_1 _5762_ (.A(_1884_),
    .B(_1912_),
    .Y(_1913_));
 sg13g2_xor2_1 _5763_ (.B(_1887_),
    .A(_1884_),
    .X(_1914_));
 sg13g2_a21o_1 _5764_ (.A2(_1914_),
    .A1(_1912_),
    .B1(_1913_),
    .X(_1915_));
 sg13g2_xor2_1 _5765_ (.B(_1886_),
    .A(_1885_),
    .X(_1916_));
 sg13g2_mux2_1 _5766_ (.A0(_1885_),
    .A1(_1916_),
    .S(_1910_),
    .X(_1917_));
 sg13g2_and2_1 _5767_ (.A(_3134_),
    .B(_1917_),
    .X(_1918_));
 sg13g2_inv_1 _5768_ (.Y(_1919_),
    .A(_1918_));
 sg13g2_xnor2_1 _5769_ (.Y(_1920_),
    .A(net1015),
    .B(_1917_));
 sg13g2_nand2b_1 _5770_ (.Y(_1921_),
    .B(\vgademo.linelfsr[2] ),
    .A_N(\vgademo.audio_snare_frames[1] ));
 sg13g2_xor2_1 _5771_ (.B(_1910_),
    .A(net1019),
    .X(_1922_));
 sg13g2_or2_1 _5772_ (.X(_1923_),
    .B(_1922_),
    .A(_1921_));
 sg13g2_o21ai_1 _5773_ (.B1(_1923_),
    .Y(_1924_),
    .A1(net1019),
    .A2(_1911_));
 sg13g2_nand2_1 _5774_ (.Y(_1925_),
    .A(_1920_),
    .B(_1924_));
 sg13g2_a21oi_1 _5775_ (.A1(_1919_),
    .A2(_1925_),
    .Y(_1926_),
    .B1(_1915_));
 sg13g2_inv_1 _5776_ (.Y(_1927_),
    .A(_1926_));
 sg13g2_nand2_1 _5777_ (.Y(_1928_),
    .A(_1870_),
    .B(_1871_));
 sg13g2_nor3_2 _5778_ (.A(_1889_),
    .B(_1927_),
    .C(_1928_),
    .Y(_1929_));
 sg13g2_xnor2_1 _5779_ (.Y(_1930_),
    .A(_1846_),
    .B(_1847_));
 sg13g2_xor2_1 _5780_ (.B(_1892_),
    .A(_1860_),
    .X(_1931_));
 sg13g2_inv_1 _5781_ (.Y(_1932_),
    .A(_1931_));
 sg13g2_xor2_1 _5782_ (.B(_1928_),
    .A(_1891_),
    .X(_1933_));
 sg13g2_inv_1 _5783_ (.Y(_1934_),
    .A(_1933_));
 sg13g2_xnor2_1 _5784_ (.Y(_1935_),
    .A(_1888_),
    .B(_1889_));
 sg13g2_nand3_1 _5785_ (.B(_1933_),
    .C(_1935_),
    .A(_1913_),
    .Y(_1936_));
 sg13g2_or2_1 _5786_ (.X(_1937_),
    .B(_1936_),
    .A(_1932_));
 sg13g2_xnor2_1 _5787_ (.Y(_1938_),
    .A(_1931_),
    .B(_1936_));
 sg13g2_nand2_1 _5788_ (.Y(_1939_),
    .A(_1860_),
    .B(_1929_));
 sg13g2_nand3_1 _5789_ (.B(_1929_),
    .C(_1930_),
    .A(_1860_),
    .Y(_1940_));
 sg13g2_xnor2_1 _5790_ (.Y(_1941_),
    .A(_1837_),
    .B(_1894_));
 sg13g2_xnor2_1 _5791_ (.Y(_1942_),
    .A(_1893_),
    .B(_1930_));
 sg13g2_nor2b_1 _5792_ (.A(_1937_),
    .B_N(_1942_),
    .Y(_1943_));
 sg13g2_and2_1 _5793_ (.A(_1941_),
    .B(_1943_),
    .X(_1944_));
 sg13g2_xnor2_1 _5794_ (.Y(_1945_),
    .A(_1941_),
    .B(_1943_));
 sg13g2_nor2_1 _5795_ (.A(_1940_),
    .B(_1945_),
    .Y(_1946_));
 sg13g2_nand2_1 _5796_ (.Y(_1947_),
    .A(_1909_),
    .B(_1946_));
 sg13g2_o21ai_1 _5797_ (.B1(_1907_),
    .Y(_1948_),
    .A1(_1896_),
    .A2(_1908_));
 sg13g2_o21ai_1 _5798_ (.B1(_1904_),
    .Y(_1949_),
    .A1(_3113_),
    .A2(_1905_));
 sg13g2_a21oi_1 _5799_ (.A1(\vgademo.linelfsr[11] ),
    .A2(_1902_),
    .Y(_1950_),
    .B1(_1900_));
 sg13g2_xnor2_1 _5800_ (.Y(_1951_),
    .A(_3087_),
    .B(_1899_));
 sg13g2_nand2_1 _5801_ (.Y(_1952_),
    .A(\vgademo.a_scrolly[11] ),
    .B(net1065));
 sg13g2_xor2_1 _5802_ (.B(_1952_),
    .A(\vgademo.a_scrolly[12] ),
    .X(_1953_));
 sg13g2_xnor2_1 _5803_ (.Y(_1954_),
    .A(_1951_),
    .B(_1953_));
 sg13g2_xnor2_1 _5804_ (.Y(_1955_),
    .A(_1950_),
    .B(_1954_));
 sg13g2_xnor2_1 _5805_ (.Y(_1956_),
    .A(_1949_),
    .B(_1955_));
 sg13g2_xor2_1 _5806_ (.B(_1956_),
    .A(_1948_),
    .X(_1957_));
 sg13g2_and2_1 _5807_ (.A(_1909_),
    .B(_1944_),
    .X(_1958_));
 sg13g2_nor2_1 _5808_ (.A(_1957_),
    .B(_1958_),
    .Y(_1959_));
 sg13g2_and2_1 _5809_ (.A(_1957_),
    .B(_1958_),
    .X(_1960_));
 sg13g2_nand2_1 _5810_ (.Y(_1961_),
    .A(_1957_),
    .B(_1958_));
 sg13g2_o21ai_1 _5811_ (.B1(_1947_),
    .Y(_1962_),
    .A1(_1959_),
    .A2(_1960_));
 sg13g2_inv_1 _5812_ (.Y(_1963_),
    .A(_1962_));
 sg13g2_nor2_1 _5813_ (.A(_1944_),
    .B(_1946_),
    .Y(_1964_));
 sg13g2_xor2_1 _5814_ (.B(_1964_),
    .A(_1909_),
    .X(_1965_));
 sg13g2_nand2_1 _5815_ (.Y(_1966_),
    .A(\vgademo.h_count[9] ),
    .B(_1965_));
 sg13g2_xor2_1 _5816_ (.B(_1945_),
    .A(_1940_),
    .X(_1967_));
 sg13g2_nor2_1 _5817_ (.A(_0038_),
    .B(_1967_),
    .Y(_1968_));
 sg13g2_or2_1 _5818_ (.X(_1969_),
    .B(_1926_),
    .A(_1913_));
 sg13g2_nand2_1 _5819_ (.Y(_1970_),
    .A(_1935_),
    .B(_1969_));
 sg13g2_xor2_1 _5820_ (.B(_1969_),
    .A(_1935_),
    .X(_1971_));
 sg13g2_nand3_1 _5821_ (.B(_1919_),
    .C(_1925_),
    .A(_1915_),
    .Y(_1972_));
 sg13g2_nand2_1 _5822_ (.Y(_1973_),
    .A(_1927_),
    .B(_1972_));
 sg13g2_xnor2_1 _5823_ (.Y(_1974_),
    .A(_1920_),
    .B(_1924_));
 sg13g2_nor2b_1 _5824_ (.A(\vgademo.linelfsr[2] ),
    .B_N(\vgademo.audio_snare_frames[1] ),
    .Y(_1975_));
 sg13g2_a21o_1 _5825_ (.A2(_1921_),
    .A1(net1005),
    .B1(_1975_),
    .X(_1976_));
 sg13g2_o21ai_1 _5826_ (.B1(_1976_),
    .Y(_1977_),
    .A1(net1003),
    .A2(_1922_));
 sg13g2_nand2_1 _5827_ (.Y(_1978_),
    .A(net1003),
    .B(_1922_));
 sg13g2_nand3_1 _5828_ (.B(_1977_),
    .C(_1978_),
    .A(_1923_),
    .Y(_1979_));
 sg13g2_a21oi_1 _5829_ (.A1(_3175_),
    .A2(_1979_),
    .Y(_1980_),
    .B1(_1974_));
 sg13g2_a21oi_1 _5830_ (.A1(_0033_),
    .A2(_1979_),
    .Y(_1981_),
    .B1(net1002));
 sg13g2_a21oi_1 _5831_ (.A1(_1974_),
    .A2(_1981_),
    .Y(_1982_),
    .B1(_1980_));
 sg13g2_a21o_1 _5832_ (.A2(_1982_),
    .A1(_1973_),
    .B1(net1000),
    .X(_1983_));
 sg13g2_o21ai_1 _5833_ (.B1(_1983_),
    .Y(_1984_),
    .A1(_1973_),
    .A2(_1982_));
 sg13g2_o21ai_1 _5834_ (.B1(_1984_),
    .Y(_1985_),
    .A1(_0044_),
    .A2(_1971_));
 sg13g2_xor2_1 _5835_ (.B(_1933_),
    .A(_0035_),
    .X(_1986_));
 sg13g2_xor2_1 _5836_ (.B(_1986_),
    .A(_1970_),
    .X(_1987_));
 sg13g2_a21oi_1 _5837_ (.A1(_0044_),
    .A2(_1971_),
    .Y(_1988_),
    .B1(_1987_));
 sg13g2_xnor2_1 _5838_ (.Y(_1989_),
    .A(_1934_),
    .B(_1970_));
 sg13g2_a22oi_1 _5839_ (.Y(_1990_),
    .B1(_1989_),
    .B2(net997),
    .A2(_1988_),
    .A1(_1985_));
 sg13g2_xnor2_1 _5840_ (.Y(_1991_),
    .A(_1929_),
    .B(_1938_));
 sg13g2_xor2_1 _5841_ (.B(_1991_),
    .A(_0036_),
    .X(_1992_));
 sg13g2_nor2_1 _5842_ (.A(_1990_),
    .B(_1992_),
    .Y(_1993_));
 sg13g2_nand2_1 _5843_ (.Y(_1994_),
    .A(_1937_),
    .B(_1939_));
 sg13g2_xor2_1 _5844_ (.B(_1994_),
    .A(_1942_),
    .X(_1995_));
 sg13g2_a21oi_1 _5845_ (.A1(net996),
    .A2(_1991_),
    .Y(_1996_),
    .B1(_1993_));
 sg13g2_o21ai_1 _5846_ (.B1(_1996_),
    .Y(_1997_),
    .A1(_3110_),
    .A2(_1995_));
 sg13g2_a22oi_1 _5847_ (.Y(_1998_),
    .B1(_1995_),
    .B2(_3110_),
    .A2(_1967_),
    .A1(_0038_));
 sg13g2_a21oi_1 _5848_ (.A1(_1997_),
    .A2(_1998_),
    .Y(_1999_),
    .B1(_1968_));
 sg13g2_xnor2_1 _5849_ (.Y(_2000_),
    .A(_3176_),
    .B(_1965_));
 sg13g2_o21ai_1 _5850_ (.B1(_1966_),
    .Y(_2001_),
    .A1(_1999_),
    .A2(_2000_));
 sg13g2_xor2_1 _5851_ (.B(_1962_),
    .A(net995),
    .X(_2002_));
 sg13g2_a22oi_1 _5852_ (.Y(_2003_),
    .B1(_2001_),
    .B2(_2002_),
    .A2(_1963_),
    .A1(\vgademo.h_count[10] ));
 sg13g2_a21oi_1 _5853_ (.A1(_1947_),
    .A2(_1961_),
    .Y(_2004_),
    .B1(_1959_));
 sg13g2_nand2b_1 _5854_ (.Y(_2005_),
    .B(\vgademo.h_count[8] ),
    .A_N(_1941_));
 sg13g2_nor2_1 _5855_ (.A(_0044_),
    .B(_1935_),
    .Y(_2006_));
 sg13g2_nand2b_1 _5856_ (.Y(_2007_),
    .B(\vgademo.linelfsr[2] ),
    .A_N(net1005));
 sg13g2_o21ai_1 _5857_ (.B1(_2007_),
    .Y(_2008_),
    .A1(net1003),
    .A2(_1910_));
 sg13g2_o21ai_1 _5858_ (.B1(_2008_),
    .Y(_2009_),
    .A1(_3106_),
    .A2(_1911_));
 sg13g2_nand3_1 _5859_ (.B(_1916_),
    .C(_2009_),
    .A(_3175_),
    .Y(_2010_));
 sg13g2_a21oi_1 _5860_ (.A1(_0033_),
    .A2(_2009_),
    .Y(_2011_),
    .B1(net1002));
 sg13g2_o21ai_1 _5861_ (.B1(_2010_),
    .Y(_2012_),
    .A1(_1916_),
    .A2(_2011_));
 sg13g2_o21ai_1 _5862_ (.B1(_2012_),
    .Y(_2013_),
    .A1(net1000),
    .A2(_1914_));
 sg13g2_a21oi_1 _5863_ (.A1(net1000),
    .A2(_1914_),
    .Y(_2014_),
    .B1(_2006_));
 sg13g2_a22oi_1 _5864_ (.Y(_2015_),
    .B1(_2013_),
    .B2(_2014_),
    .A2(_1935_),
    .A1(_0044_));
 sg13g2_a22oi_1 _5865_ (.Y(_2016_),
    .B1(_1986_),
    .B2(_2015_),
    .A2(_1934_),
    .A1(net997));
 sg13g2_xnor2_1 _5866_ (.Y(_2017_),
    .A(_0036_),
    .B(_1931_));
 sg13g2_nor2_1 _5867_ (.A(_2016_),
    .B(_2017_),
    .Y(_2018_));
 sg13g2_nor2_1 _5868_ (.A(_3110_),
    .B(_1942_),
    .Y(_2019_));
 sg13g2_a21oi_1 _5869_ (.A1(net996),
    .A2(_1932_),
    .Y(_2020_),
    .B1(_2018_));
 sg13g2_a21oi_1 _5870_ (.A1(_3110_),
    .A2(_1942_),
    .Y(_2021_),
    .B1(_2020_));
 sg13g2_xor2_1 _5871_ (.B(_1941_),
    .A(_0038_),
    .X(_2022_));
 sg13g2_o21ai_1 _5872_ (.B1(_2022_),
    .Y(_2023_),
    .A1(_2019_),
    .A2(_2021_));
 sg13g2_a22oi_1 _5873_ (.Y(_2024_),
    .B1(_2005_),
    .B2(_2023_),
    .A2(_1909_),
    .A1(_3111_));
 sg13g2_nor2_1 _5874_ (.A(net995),
    .B(_1957_),
    .Y(_2025_));
 sg13g2_nor2_1 _5875_ (.A(_3111_),
    .B(_1909_),
    .Y(_2026_));
 sg13g2_nor3_1 _5876_ (.A(_2024_),
    .B(_2025_),
    .C(_2026_),
    .Y(_2027_));
 sg13g2_nor2_2 _5877_ (.A(\vgademo.v_count[8] ),
    .B(net975),
    .Y(_2028_));
 sg13g2_nor2_1 _5878_ (.A(net962),
    .B(net971),
    .Y(_2029_));
 sg13g2_xnor2_1 _5879_ (.Y(_2030_),
    .A(net962),
    .B(net971));
 sg13g2_nand2b_1 _5880_ (.Y(_2031_),
    .B(_2030_),
    .A_N(_2028_));
 sg13g2_nand2_1 _5881_ (.Y(_2032_),
    .A(net963),
    .B(net978));
 sg13g2_xor2_1 _5882_ (.B(net975),
    .A(\vgademo.v_count[8] ),
    .X(_2033_));
 sg13g2_or2_1 _5883_ (.X(_2034_),
    .B(_2033_),
    .A(_2032_));
 sg13g2_nor2_1 _5884_ (.A(net964),
    .B(net980),
    .Y(_2035_));
 sg13g2_xnor2_1 _5885_ (.Y(_2036_),
    .A(net963),
    .B(net978));
 sg13g2_nor2_1 _5886_ (.A(_2035_),
    .B(_2036_),
    .Y(_2037_));
 sg13g2_nor2_1 _5887_ (.A(net966),
    .B(net983),
    .Y(_2038_));
 sg13g2_xor2_1 _5888_ (.B(net980),
    .A(net964),
    .X(_2039_));
 sg13g2_nor2_1 _5889_ (.A(_2038_),
    .B(_2039_),
    .Y(_2040_));
 sg13g2_or2_1 _5890_ (.X(_2041_),
    .B(net987),
    .A(net967));
 sg13g2_xnor2_1 _5891_ (.Y(_2042_),
    .A(net966),
    .B(net983));
 sg13g2_or2_1 _5892_ (.X(_2043_),
    .B(_2042_),
    .A(_2041_));
 sg13g2_nor2_1 _5893_ (.A(net968),
    .B(net993),
    .Y(_2044_));
 sg13g2_xnor2_1 _5894_ (.Y(_2045_),
    .A(net967),
    .B(net986));
 sg13g2_o21ai_1 _5895_ (.B1(_2045_),
    .Y(_2046_),
    .A1(\vgademo.v_count[3] ),
    .A2(net990));
 sg13g2_a21oi_1 _5896_ (.A1(\vgademo.v_count[3] ),
    .A2(net990),
    .Y(_2047_),
    .B1(_2045_));
 sg13g2_or2_1 _5897_ (.X(_2048_),
    .B(_2047_),
    .A(_2044_));
 sg13g2_nand2_1 _5898_ (.Y(_2049_),
    .A(_2043_),
    .B(_2046_));
 sg13g2_nor2b_1 _5899_ (.A(_2046_),
    .B_N(_2043_),
    .Y(_2050_));
 sg13g2_a21oi_1 _5900_ (.A1(_2041_),
    .A2(_2042_),
    .Y(_2051_),
    .B1(_2050_));
 sg13g2_o21ai_1 _5901_ (.B1(_2051_),
    .Y(_2052_),
    .A1(_2048_),
    .A2(_2049_));
 sg13g2_xnor2_1 _5902_ (.Y(_2053_),
    .A(_2038_),
    .B(_2039_));
 sg13g2_inv_1 _5903_ (.Y(_2054_),
    .A(_2053_));
 sg13g2_a21oi_1 _5904_ (.A1(_2052_),
    .A2(_2054_),
    .Y(_2055_),
    .B1(_2040_));
 sg13g2_inv_1 _5905_ (.Y(_2056_),
    .A(_2055_));
 sg13g2_xor2_1 _5906_ (.B(_2036_),
    .A(_2035_),
    .X(_2057_));
 sg13g2_a21oi_1 _5907_ (.A1(_2056_),
    .A2(_2057_),
    .Y(_2058_),
    .B1(_2037_));
 sg13g2_xnor2_1 _5908_ (.Y(_2059_),
    .A(_2032_),
    .B(_2033_));
 sg13g2_o21ai_1 _5909_ (.B1(_2034_),
    .Y(_2060_),
    .A1(_2058_),
    .A2(_2059_));
 sg13g2_xor2_1 _5910_ (.B(_2030_),
    .A(_2028_),
    .X(_2061_));
 sg13g2_nand2b_1 _5911_ (.Y(_2062_),
    .B(_2060_),
    .A_N(_2061_));
 sg13g2_xnor2_1 _5912_ (.Y(_2063_),
    .A(_3113_),
    .B(_2029_));
 sg13g2_a21oi_1 _5913_ (.A1(_2031_),
    .A2(_2062_),
    .Y(_2064_),
    .B1(_2063_));
 sg13g2_nor2_1 _5914_ (.A(_0020_),
    .B(_2029_),
    .Y(_2065_));
 sg13g2_nor2_1 _5915_ (.A(_2064_),
    .B(_2065_),
    .Y(_2066_));
 sg13g2_nor3_1 _5916_ (.A(\vgademo.a_scrolly[12] ),
    .B(_2064_),
    .C(_2065_),
    .Y(_2067_));
 sg13g2_nand2_1 _5917_ (.Y(_2068_),
    .A(_1043_),
    .B(_2066_));
 sg13g2_o21ai_1 _5918_ (.B1(_2068_),
    .Y(_2069_),
    .A1(_3112_),
    .A2(_2067_));
 sg13g2_xnor2_1 _5919_ (.Y(_2070_),
    .A(_0067_),
    .B(_2066_));
 sg13g2_nor2_1 _5920_ (.A(_2069_),
    .B(_2070_),
    .Y(_2071_));
 sg13g2_nand2b_1 _5921_ (.Y(_2072_),
    .B(_2061_),
    .A_N(_2060_));
 sg13g2_a21oi_1 _5922_ (.A1(_2062_),
    .A2(_2072_),
    .Y(_2073_),
    .B1(_2069_));
 sg13g2_nor2_1 _5923_ (.A(\vgademo.a_scrolly[13] ),
    .B(_2067_),
    .Y(_2074_));
 sg13g2_xnor2_1 _5924_ (.Y(_2075_),
    .A(_3119_),
    .B(_2074_));
 sg13g2_nand3_1 _5925_ (.B(_2062_),
    .C(_2063_),
    .A(_2031_),
    .Y(_2076_));
 sg13g2_nor2b_1 _5926_ (.A(_2064_),
    .B_N(_2076_),
    .Y(_2077_));
 sg13g2_xor2_1 _5927_ (.B(_2059_),
    .A(_2058_),
    .X(_2078_));
 sg13g2_xnor2_1 _5928_ (.Y(_2079_),
    .A(_2052_),
    .B(_2053_));
 sg13g2_xnor2_1 _5929_ (.Y(_2080_),
    .A(_2055_),
    .B(_2057_));
 sg13g2_nand4_1 _5930_ (.B(_2078_),
    .C(_2079_),
    .A(_2077_),
    .Y(_2081_),
    .D(_2080_));
 sg13g2_nor2b_1 _5931_ (.A(_2069_),
    .B_N(_2081_),
    .Y(_2082_));
 sg13g2_nor2_1 _5932_ (.A(_2069_),
    .B(_2077_),
    .Y(_2083_));
 sg13g2_nor4_2 _5933_ (.A(_2071_),
    .B(_2073_),
    .C(_2075_),
    .Y(_2084_),
    .D(_2082_));
 sg13g2_nor2_1 _5934_ (.A(_2027_),
    .B(_2084_),
    .Y(_2085_));
 sg13g2_o21ai_1 _5935_ (.B1(_2085_),
    .Y(_2086_),
    .A1(_2003_),
    .A2(_2004_));
 sg13g2_a21oi_2 _5936_ (.B1(_2086_),
    .Y(_2087_),
    .A2(_1957_),
    .A1(net995));
 sg13g2_nor2_2 _5937_ (.A(net855),
    .B(_2087_),
    .Y(_2088_));
 sg13g2_inv_1 _5938_ (.Y(_2089_),
    .A(_2088_));
 sg13g2_nor4_2 _5939_ (.A(net992),
    .B(\vgademo.a_scrolly[10] ),
    .C(net974),
    .Y(_2090_),
    .D(_1353_));
 sg13g2_a22oi_1 _5940_ (.Y(_2091_),
    .B1(_2090_),
    .B2(_1035_),
    .A2(_1202_),
    .A1(_3116_));
 sg13g2_and3_1 _5941_ (.X(_2092_),
    .A(_1035_),
    .B(_1083_),
    .C(_2090_));
 sg13g2_nor3_2 _5942_ (.A(_1081_),
    .B(_2091_),
    .C(_2092_),
    .Y(_2093_));
 sg13g2_a21oi_2 _5943_ (.B1(_2089_),
    .Y(_2094_),
    .A2(_2093_),
    .A1(_0069_));
 sg13g2_nor2_1 _5944_ (.A(_1683_),
    .B(_2088_),
    .Y(_2095_));
 sg13g2_nor2_1 _5945_ (.A(_1683_),
    .B(_2094_),
    .Y(_2096_));
 sg13g2_nor2_2 _5946_ (.A(_2075_),
    .B(_2093_),
    .Y(_2097_));
 sg13g2_o21ai_1 _5947_ (.B1(_2097_),
    .Y(_2098_),
    .A1(_2069_),
    .A2(_2078_));
 sg13g2_a21oi_1 _5948_ (.A1(_2094_),
    .A2(_2098_),
    .Y(_2099_),
    .B1(net827));
 sg13g2_a21o_2 _5949_ (.A2(_2099_),
    .A1(_1811_),
    .B1(_1694_),
    .X(_2100_));
 sg13g2_xnor2_1 _5950_ (.Y(_2101_),
    .A(net1004),
    .B(net993));
 sg13g2_xnor2_1 _5951_ (.Y(_2102_),
    .A(_3100_),
    .B(_2101_));
 sg13g2_inv_1 _5952_ (.Y(_2103_),
    .A(_2102_));
 sg13g2_and2_1 _5953_ (.A(_2100_),
    .B(_2103_),
    .X(_2104_));
 sg13g2_xnor2_1 _5954_ (.Y(_2105_),
    .A(net845),
    .B(_1447_));
 sg13g2_inv_1 _5955_ (.Y(_2106_),
    .A(_2105_));
 sg13g2_nand2_1 _5956_ (.Y(_2107_),
    .A(_1294_),
    .B(_2106_));
 sg13g2_xnor2_1 _5957_ (.Y(_2108_),
    .A(_1686_),
    .B(_1687_));
 sg13g2_inv_1 _5958_ (.Y(_2109_),
    .A(_2108_));
 sg13g2_nor2_2 _5959_ (.A(_1684_),
    .B(_2109_),
    .Y(_2110_));
 sg13g2_nand3_1 _5960_ (.B(_1681_),
    .C(_2108_),
    .A(net832),
    .Y(_2111_));
 sg13g2_nand3_1 _5961_ (.B(_1692_),
    .C(_2111_),
    .A(net861),
    .Y(_2112_));
 sg13g2_nand3_1 _5962_ (.B(_1690_),
    .C(_2108_),
    .A(net861),
    .Y(_2113_));
 sg13g2_and2_1 _5963_ (.A(_2112_),
    .B(_2113_),
    .X(_2114_));
 sg13g2_nand3_1 _5964_ (.B(_2112_),
    .C(_2113_),
    .A(_2107_),
    .Y(_2115_));
 sg13g2_nand3_1 _5965_ (.B(_1723_),
    .C(_1724_),
    .A(_1720_),
    .Y(_2116_));
 sg13g2_nand3b_1 _5966_ (.B(_1777_),
    .C(_2116_),
    .Y(_2117_),
    .A_N(_1725_));
 sg13g2_nor2_1 _5967_ (.A(_0057_),
    .B(_1802_),
    .Y(_2118_));
 sg13g2_nor2_1 _5968_ (.A(_1803_),
    .B(_2118_),
    .Y(_2119_));
 sg13g2_o21ai_1 _5969_ (.B1(_2117_),
    .Y(_2120_),
    .A1(_1803_),
    .A2(_2118_));
 sg13g2_inv_1 _5970_ (.Y(_2121_),
    .A(_2120_));
 sg13g2_or2_1 _5971_ (.X(_2122_),
    .B(_1774_),
    .A(_1761_));
 sg13g2_and2_2 _5972_ (.A(_1803_),
    .B(_2122_),
    .X(_2123_));
 sg13g2_o21ai_1 _5973_ (.B1(_2121_),
    .Y(_2124_),
    .A1(net828),
    .A2(net852));
 sg13g2_nand3_1 _5974_ (.B(net853),
    .C(_2123_),
    .A(net830),
    .Y(_2125_));
 sg13g2_nand3_1 _5975_ (.B(_2124_),
    .C(_2125_),
    .A(net854),
    .Y(_2126_));
 sg13g2_and2_1 _5976_ (.A(_0056_),
    .B(_2093_),
    .X(_2127_));
 sg13g2_o21ai_1 _5977_ (.B1(net860),
    .Y(_2128_),
    .A1(_2087_),
    .A2(_2127_));
 sg13g2_nand2_1 _5978_ (.Y(_2129_),
    .A(net860),
    .B(_2097_));
 sg13g2_o21ai_1 _5979_ (.B1(_2128_),
    .Y(_2130_),
    .A1(_2073_),
    .A2(_2129_));
 sg13g2_inv_1 _5980_ (.Y(_2131_),
    .A(_2130_));
 sg13g2_a21o_1 _5981_ (.A2(_2131_),
    .A1(_2126_),
    .B1(net827),
    .X(_2132_));
 sg13g2_nand2_1 _5982_ (.Y(_2133_),
    .A(_2115_),
    .B(_2132_));
 sg13g2_xnor2_1 _5983_ (.Y(_2134_),
    .A(_2100_),
    .B(_2102_));
 sg13g2_a21oi_1 _5984_ (.A1(_2133_),
    .A2(_2134_),
    .Y(_2135_),
    .B1(_2104_));
 sg13g2_nand3_1 _5985_ (.B(net826),
    .C(_1809_),
    .A(net854),
    .Y(_2136_));
 sg13g2_a21oi_1 _5986_ (.A1(_0075_),
    .A2(_2093_),
    .Y(_2137_),
    .B1(_2087_));
 sg13g2_nor2_1 _5987_ (.A(net855),
    .B(_2137_),
    .Y(_2138_));
 sg13g2_nor2_1 _5988_ (.A(_2083_),
    .B(_2129_),
    .Y(_2139_));
 sg13g2_nor2_1 _5989_ (.A(_2138_),
    .B(_2139_),
    .Y(_2140_));
 sg13g2_a21oi_1 _5990_ (.A1(_2136_),
    .A2(_2140_),
    .Y(_2141_),
    .B1(net827));
 sg13g2_nor2_1 _5991_ (.A(_1687_),
    .B(_2105_),
    .Y(_2142_));
 sg13g2_nand4_1 _5992_ (.B(_1681_),
    .C(_1690_),
    .A(net832),
    .Y(_2143_),
    .D(_2142_));
 sg13g2_nand2_2 _5993_ (.Y(_2144_),
    .A(net861),
    .B(_2143_));
 sg13g2_nor2_1 _5994_ (.A(_2141_),
    .B(_2144_),
    .Y(_2145_));
 sg13g2_or2_1 _5995_ (.X(_2146_),
    .B(_2144_),
    .A(_2141_));
 sg13g2_xor2_1 _5996_ (.B(net993),
    .A(\vgademo.h_count[0] ),
    .X(_2147_));
 sg13g2_xnor2_1 _5997_ (.Y(_2148_),
    .A(\vgademo.h_count[0] ),
    .B(net993));
 sg13g2_a21o_1 _5998_ (.A2(_2132_),
    .A1(_2115_),
    .B1(_2148_),
    .X(_2149_));
 sg13g2_nor2_1 _5999_ (.A(_2133_),
    .B(_2147_),
    .Y(_2150_));
 sg13g2_nand3_1 _6000_ (.B(_2132_),
    .C(_2148_),
    .A(_2115_),
    .Y(_2151_));
 sg13g2_and3_1 _6001_ (.X(_2152_),
    .A(_2146_),
    .B(_2149_),
    .C(_2151_));
 sg13g2_a21oi_1 _6002_ (.A1(_2149_),
    .A2(_2151_),
    .Y(_2153_),
    .B1(_2146_));
 sg13g2_o21ai_1 _6003_ (.B1(_2135_),
    .Y(_2154_),
    .A1(_2152_),
    .A2(_2153_));
 sg13g2_a21oi_2 _6004_ (.B1(_1802_),
    .Y(_2155_),
    .A2(net844),
    .A1(_0058_));
 sg13g2_o21ai_1 _6005_ (.B1(_2155_),
    .Y(_2156_),
    .A1(_3158_),
    .A2(_1778_));
 sg13g2_o21ai_1 _6006_ (.B1(_2156_),
    .Y(_2157_),
    .A1(net828),
    .A2(net852));
 sg13g2_nand3_1 _6007_ (.B(net853),
    .C(_1806_),
    .A(net831),
    .Y(_2158_));
 sg13g2_nand3_1 _6008_ (.B(_2157_),
    .C(_2158_),
    .A(net856),
    .Y(_2159_));
 sg13g2_o21ai_1 _6009_ (.B1(_2097_),
    .Y(_2160_),
    .A1(_2069_),
    .A2(_2079_));
 sg13g2_a21oi_1 _6010_ (.A1(_2088_),
    .A2(_2160_),
    .Y(_2161_),
    .B1(net827));
 sg13g2_a21oi_2 _6011_ (.B1(net863),
    .Y(_2162_),
    .A2(_2161_),
    .A1(_2159_));
 sg13g2_nor2_1 _6012_ (.A(_2101_),
    .B(_2162_),
    .Y(_2163_));
 sg13g2_nand2_1 _6013_ (.Y(_2164_),
    .A(_0064_),
    .B(_2093_));
 sg13g2_a22oi_1 _6014_ (.Y(_2165_),
    .B1(_2088_),
    .B2(_2164_),
    .A2(_1681_),
    .A1(net830));
 sg13g2_o21ai_1 _6015_ (.B1(_2097_),
    .Y(_2166_),
    .A1(_2069_),
    .A2(_2080_));
 sg13g2_a21oi_1 _6016_ (.A1(net830),
    .A2(_1681_),
    .Y(_2167_),
    .B1(_2166_));
 sg13g2_or2_1 _6017_ (.X(_2168_),
    .B(_2167_),
    .A(_2165_));
 sg13g2_or2_1 _6018_ (.X(_2169_),
    .B(\vgademo.plane_du[4] ),
    .A(net993));
 sg13g2_nand3_1 _6019_ (.B(_1777_),
    .C(_2169_),
    .A(_1721_),
    .Y(_2170_));
 sg13g2_a21oi_2 _6020_ (.B1(_1802_),
    .Y(_2171_),
    .A2(net844),
    .A1(_0059_));
 sg13g2_nand2_1 _6021_ (.Y(_2172_),
    .A(_2170_),
    .B(_2171_));
 sg13g2_o21ai_1 _6022_ (.B1(_2172_),
    .Y(_2173_),
    .A1(net828),
    .A2(net852));
 sg13g2_o21ai_1 _6023_ (.B1(_2173_),
    .Y(_2174_),
    .A1(net826),
    .A2(_2121_));
 sg13g2_o21ai_1 _6024_ (.B1(_2168_),
    .Y(_2175_),
    .A1(net860),
    .A2(_2174_));
 sg13g2_nand2_1 _6025_ (.Y(_2176_),
    .A(net861),
    .B(_2175_));
 sg13g2_xor2_1 _6026_ (.B(_2162_),
    .A(_2101_),
    .X(_2177_));
 sg13g2_a21oi_1 _6027_ (.A1(_2176_),
    .A2(_2177_),
    .Y(_2178_),
    .B1(_2163_));
 sg13g2_xnor2_1 _6028_ (.Y(_2179_),
    .A(_2133_),
    .B(_2134_));
 sg13g2_nor2_1 _6029_ (.A(_2178_),
    .B(_2179_),
    .Y(_2180_));
 sg13g2_xor2_1 _6030_ (.B(_2179_),
    .A(_2178_),
    .X(_2181_));
 sg13g2_nor3_1 _6031_ (.A(_2135_),
    .B(_2152_),
    .C(_2153_),
    .Y(_2182_));
 sg13g2_or3_1 _6032_ (.A(_2135_),
    .B(_2152_),
    .C(_2153_),
    .X(_2183_));
 sg13g2_nor2_1 _6033_ (.A(\vgademo.scanline_audio_sample[4] ),
    .B(\vgademo.scanline_audio_sample[3] ),
    .Y(_2184_));
 sg13g2_nand2_1 _6034_ (.Y(_2185_),
    .A(_0043_),
    .B(_2184_));
 sg13g2_xor2_1 _6035_ (.B(_2185_),
    .A(\vgademo.scanline_audio_sample[6] ),
    .X(_2186_));
 sg13g2_xnor2_1 _6036_ (.Y(_2187_),
    .A(_0036_),
    .B(_2186_));
 sg13g2_xnor2_1 _6037_ (.Y(_2188_),
    .A(_0043_),
    .B(_2184_));
 sg13g2_xor2_1 _6038_ (.B(_2188_),
    .A(_0035_),
    .X(_2189_));
 sg13g2_xor2_1 _6039_ (.B(\vgademo.scanline_audio_sample[3] ),
    .A(\vgademo.scanline_audio_sample[4] ),
    .X(_2190_));
 sg13g2_nor2b_1 _6040_ (.A(_2190_),
    .B_N(_0044_),
    .Y(_2191_));
 sg13g2_xnor2_1 _6041_ (.Y(_2192_),
    .A(_0044_),
    .B(_2190_));
 sg13g2_nand4_1 _6042_ (.B(_2187_),
    .C(_2189_),
    .A(_0037_),
    .Y(_2193_),
    .D(_2192_));
 sg13g2_nor2_1 _6043_ (.A(_1275_),
    .B(_1277_),
    .Y(_2194_));
 sg13g2_nor2_1 _6044_ (.A(_1273_),
    .B(_1277_),
    .Y(_2195_));
 sg13g2_a221oi_1 _6045_ (.B2(_2194_),
    .C1(_2195_),
    .B1(_1281_),
    .A1(_3107_),
    .Y(_2196_),
    .A2(_3189_));
 sg13g2_nor2b_1 _6046_ (.A(_2186_),
    .B_N(_1283_),
    .Y(_2197_));
 sg13g2_a22oi_1 _6047_ (.Y(_2198_),
    .B1(_2189_),
    .B2(_2191_),
    .A2(_2188_),
    .A1(_3109_));
 sg13g2_nand3b_1 _6048_ (.B(_2187_),
    .C(_0037_),
    .Y(_2199_),
    .A_N(_2198_));
 sg13g2_o21ai_1 _6049_ (.B1(_2199_),
    .Y(_2200_),
    .A1(_2193_),
    .A2(_2196_));
 sg13g2_nor2_1 _6050_ (.A(_1290_),
    .B(_2193_),
    .Y(_2201_));
 sg13g2_a21oi_1 _6051_ (.A1(_2194_),
    .A2(_2201_),
    .Y(_2202_),
    .B1(_1292_));
 sg13g2_o21ai_1 _6052_ (.B1(_2202_),
    .Y(_2203_),
    .A1(_2197_),
    .A2(_2200_));
 sg13g2_nor2_1 _6053_ (.A(net861),
    .B(_2203_),
    .Y(_2204_));
 sg13g2_inv_1 _6054_ (.Y(_2205_),
    .A(_2204_));
 sg13g2_nor2_1 _6055_ (.A(net860),
    .B(_2123_),
    .Y(_2206_));
 sg13g2_o21ai_1 _6056_ (.B1(_2206_),
    .Y(_2207_),
    .A1(net828),
    .A2(net852));
 sg13g2_a21oi_1 _6057_ (.A1(_0078_),
    .A2(_2093_),
    .Y(_2208_),
    .B1(_2087_));
 sg13g2_nor2_2 _6058_ (.A(net855),
    .B(_2208_),
    .Y(_2209_));
 sg13g2_nor2_1 _6059_ (.A(_2071_),
    .B(_2129_),
    .Y(_2210_));
 sg13g2_nor2_1 _6060_ (.A(_2209_),
    .B(_2210_),
    .Y(_2211_));
 sg13g2_a21oi_1 _6061_ (.A1(_2207_),
    .A2(_2211_),
    .Y(_2212_),
    .B1(net827));
 sg13g2_o21ai_1 _6062_ (.B1(_2205_),
    .Y(_2213_),
    .A1(_2144_),
    .A2(_2212_));
 sg13g2_xnor2_1 _6063_ (.Y(_2214_),
    .A(\vgademo.h_count[2] ),
    .B(net993));
 sg13g2_nor2_1 _6064_ (.A(_2213_),
    .B(_2214_),
    .Y(_2215_));
 sg13g2_a22oi_1 _6065_ (.Y(_2216_),
    .B1(_2213_),
    .B2(_2214_),
    .A2(_2175_),
    .A1(net861));
 sg13g2_o21ai_1 _6066_ (.B1(_2100_),
    .Y(_2217_),
    .A1(_2215_),
    .A2(_2216_));
 sg13g2_nor3_1 _6067_ (.A(_2100_),
    .B(_2215_),
    .C(_2216_),
    .Y(_2218_));
 sg13g2_xnor2_1 _6068_ (.Y(_2219_),
    .A(_2176_),
    .B(_2177_));
 sg13g2_o21ai_1 _6069_ (.B1(_2217_),
    .Y(_2220_),
    .A1(_2218_),
    .A2(_2219_));
 sg13g2_nand4_1 _6070_ (.B(_2181_),
    .C(_2183_),
    .A(_2154_),
    .Y(_2221_),
    .D(_2220_));
 sg13g2_o21ai_1 _6071_ (.B1(_2149_),
    .Y(_2222_),
    .A1(_2145_),
    .A2(_2150_));
 sg13g2_xnor2_1 _6072_ (.Y(_2223_),
    .A(net969),
    .B(_2147_));
 sg13g2_xnor2_1 _6073_ (.Y(_2224_),
    .A(_2146_),
    .B(net942));
 sg13g2_xnor2_1 _6074_ (.Y(_2225_),
    .A(_2213_),
    .B(_2224_));
 sg13g2_a221oi_1 _6075_ (.B2(_2225_),
    .C1(_2182_),
    .B1(_2222_),
    .A1(_2154_),
    .Y(_2226_),
    .A2(_2180_));
 sg13g2_nor2_1 _6076_ (.A(_2222_),
    .B(_2225_),
    .Y(_2227_));
 sg13g2_a21oi_1 _6077_ (.A1(_2221_),
    .A2(_2226_),
    .Y(_2228_),
    .B1(_2227_));
 sg13g2_a21o_1 _6078_ (.A2(net942),
    .A1(_2145_),
    .B1(_2213_),
    .X(_2229_));
 sg13g2_o21ai_1 _6079_ (.B1(_2213_),
    .Y(_2230_),
    .A1(_2145_),
    .A2(net942));
 sg13g2_and2_1 _6080_ (.A(_2229_),
    .B(_2230_),
    .X(_2231_));
 sg13g2_nand2_1 _6081_ (.Y(_2232_),
    .A(_2228_),
    .B(_2231_));
 sg13g2_nor4_1 _6082_ (.A(net1000),
    .B(net1002),
    .C(net997),
    .D(net998),
    .Y(_2233_));
 sg13g2_o21ai_1 _6083_ (.B1(_3227_),
    .Y(_2234_),
    .A1(_3193_),
    .A2(_2233_));
 sg13g2_nor2b_2 _6084_ (.A(net995),
    .B_N(_2234_),
    .Y(_2235_));
 sg13g2_nor4_1 _6085_ (.A(net539),
    .B(net969),
    .C(\vgademo.v_count[3] ),
    .D(net968),
    .Y(_2236_));
 sg13g2_and2_1 _6086_ (.A(_3225_),
    .B(_2236_),
    .X(_2237_));
 sg13g2_or4_2 _6087_ (.A(net962),
    .B(_3223_),
    .C(_2235_),
    .D(_2237_),
    .X(_2238_));
 sg13g2_inv_1 _6088_ (.Y(_2239_),
    .A(_2238_));
 sg13g2_o21ai_1 _6089_ (.B1(_2239_),
    .Y(_2240_),
    .A1(_2228_),
    .A2(_2231_));
 sg13g2_nor2b_1 _6090_ (.A(_2240_),
    .B_N(_2232_),
    .Y(_0255_));
 sg13g2_a21oi_1 _6091_ (.A1(_2229_),
    .A2(_2232_),
    .Y(_0256_),
    .B1(_2238_));
 sg13g2_nand2_1 _6092_ (.Y(_2241_),
    .A(\vgademo.a_sin[6] ),
    .B(net909));
 sg13g2_xnor2_1 _6093_ (.Y(_0257_),
    .A(net249),
    .B(_2241_));
 sg13g2_nor2_1 _6094_ (.A(net324),
    .B(net910),
    .Y(_2242_));
 sg13g2_nand2b_1 _6095_ (.Y(_2243_),
    .B(\vgademo.a_sin[6] ),
    .A_N(net249));
 sg13g2_nor2b_1 _6096_ (.A(\vgademo.a_sin[7] ),
    .B_N(\vgademo.a_cos[1] ),
    .Y(_2244_));
 sg13g2_xnor2_1 _6097_ (.Y(_2245_),
    .A(\vgademo.a_sin[7] ),
    .B(net324));
 sg13g2_xnor2_1 _6098_ (.Y(_2246_),
    .A(_2243_),
    .B(_2245_));
 sg13g2_a21oi_1 _6099_ (.A1(net910),
    .A2(_2246_),
    .Y(_0258_),
    .B1(_2242_));
 sg13g2_nor2_1 _6100_ (.A(net306),
    .B(net910),
    .Y(_2247_));
 sg13g2_a21o_1 _6101_ (.A2(_2245_),
    .A1(_2243_),
    .B1(_2244_),
    .X(_2248_));
 sg13g2_nand2b_1 _6102_ (.Y(_2249_),
    .B(net306),
    .A_N(\vgademo.a_sin[8] ));
 sg13g2_xnor2_1 _6103_ (.Y(_2250_),
    .A(\vgademo.a_sin[8] ),
    .B(net306));
 sg13g2_nand2_1 _6104_ (.Y(_2251_),
    .A(_2248_),
    .B(_2250_));
 sg13g2_xnor2_1 _6105_ (.Y(_2252_),
    .A(_2248_),
    .B(_2250_));
 sg13g2_a21oi_1 _6106_ (.A1(net910),
    .A2(_2252_),
    .Y(_0259_),
    .B1(_2247_));
 sg13g2_nor2_1 _6107_ (.A(_3136_),
    .B(\vgademo.a_sin[9] ),
    .Y(_2253_));
 sg13g2_xor2_1 _6108_ (.B(\vgademo.a_sin[9] ),
    .A(\vgademo.a_cos[3] ),
    .X(_2254_));
 sg13g2_nand3_1 _6109_ (.B(_2251_),
    .C(_2254_),
    .A(_2249_),
    .Y(_2255_));
 sg13g2_a21oi_1 _6110_ (.A1(_2249_),
    .A2(_2251_),
    .Y(_2256_),
    .B1(_2254_));
 sg13g2_nand3b_1 _6111_ (.B(net914),
    .C(_2255_),
    .Y(_2257_),
    .A_N(_2256_));
 sg13g2_o21ai_1 _6112_ (.B1(_2257_),
    .Y(_0260_),
    .A1(_3136_),
    .A2(net914));
 sg13g2_xnor2_1 _6113_ (.Y(_2258_),
    .A(\vgademo.a_cos[4] ),
    .B(\vgademo.a_sin[10] ));
 sg13g2_or3_1 _6114_ (.A(_2253_),
    .B(_2256_),
    .C(_2258_),
    .X(_2259_));
 sg13g2_o21ai_1 _6115_ (.B1(_2258_),
    .Y(_2260_),
    .A1(_2253_),
    .A2(_2256_));
 sg13g2_a21oi_1 _6116_ (.A1(_2259_),
    .A2(_2260_),
    .Y(_2261_),
    .B1(net907));
 sg13g2_a21oi_1 _6117_ (.A1(_3138_),
    .A2(net906),
    .Y(_0261_),
    .B1(_2261_));
 sg13g2_o21ai_1 _6118_ (.B1(_2260_),
    .Y(_2262_),
    .A1(_3138_),
    .A2(\vgademo.a_sin[10] ));
 sg13g2_nor2b_1 _6119_ (.A(\vgademo.a_sin[11] ),
    .B_N(\vgademo.a_cos[5] ),
    .Y(_2263_));
 sg13g2_nand2b_1 _6120_ (.Y(_2264_),
    .B(\vgademo.a_sin[11] ),
    .A_N(\vgademo.a_cos[5] ));
 sg13g2_nor2b_1 _6121_ (.A(_2263_),
    .B_N(_2264_),
    .Y(_2265_));
 sg13g2_nor2_1 _6122_ (.A(net437),
    .B(net915),
    .Y(_2266_));
 sg13g2_xnor2_1 _6123_ (.Y(_2267_),
    .A(_2262_),
    .B(_2265_));
 sg13g2_a21oi_1 _6124_ (.A1(net911),
    .A2(_2267_),
    .Y(_0262_),
    .B1(net438));
 sg13g2_nor2_1 _6125_ (.A(_3141_),
    .B(\vgademo.a_sin[12] ),
    .Y(_2268_));
 sg13g2_xor2_1 _6126_ (.B(\vgademo.a_sin[12] ),
    .A(\vgademo.a_cos[6] ),
    .X(_2269_));
 sg13g2_a21oi_1 _6127_ (.A1(_2262_),
    .A2(_2264_),
    .Y(_2270_),
    .B1(_2263_));
 sg13g2_nor2_1 _6128_ (.A(_2269_),
    .B(_2270_),
    .Y(_2271_));
 sg13g2_xor2_1 _6129_ (.B(_2270_),
    .A(_2269_),
    .X(_2272_));
 sg13g2_nand2_1 _6130_ (.Y(_2273_),
    .A(net915),
    .B(_2272_));
 sg13g2_o21ai_1 _6131_ (.B1(_2273_),
    .Y(_0263_),
    .A1(_3141_),
    .A2(net911));
 sg13g2_xnor2_1 _6132_ (.Y(_2274_),
    .A(\vgademo.a_cos[7] ),
    .B(\vgademo.a_sin[13] ));
 sg13g2_o21ai_1 _6133_ (.B1(_2274_),
    .Y(_2275_),
    .A1(_2268_),
    .A2(_2271_));
 sg13g2_or3_1 _6134_ (.A(_2268_),
    .B(_2271_),
    .C(_2274_),
    .X(_2276_));
 sg13g2_and2_1 _6135_ (.A(_2275_),
    .B(_2276_),
    .X(_2277_));
 sg13g2_nand2_1 _6136_ (.Y(_2278_),
    .A(net911),
    .B(_2277_));
 sg13g2_o21ai_1 _6137_ (.B1(_2278_),
    .Y(_0264_),
    .A1(_3143_),
    .A2(net911));
 sg13g2_o21ai_1 _6138_ (.B1(_2275_),
    .Y(_2279_),
    .A1(_3143_),
    .A2(\vgademo.a_sin[13] ));
 sg13g2_xnor2_1 _6139_ (.Y(_2280_),
    .A(\vgademo.a_cos[8] ),
    .B(net961));
 sg13g2_and2_1 _6140_ (.A(_2279_),
    .B(_2280_),
    .X(_2281_));
 sg13g2_xor2_1 _6141_ (.B(_2280_),
    .A(_2279_),
    .X(_2282_));
 sg13g2_mux2_1 _6142_ (.A0(net570),
    .A1(_2282_),
    .S(net909),
    .X(_0265_));
 sg13g2_nor2_1 _6143_ (.A(net568),
    .B(net915),
    .Y(_2283_));
 sg13g2_xnor2_1 _6144_ (.Y(_2284_),
    .A(\vgademo.a_cos[9] ),
    .B(net960));
 sg13g2_a21oi_1 _6145_ (.A1(\vgademo.a_cos[8] ),
    .A2(_3155_),
    .Y(_2285_),
    .B1(_2281_));
 sg13g2_xor2_1 _6146_ (.B(_2285_),
    .A(_2284_),
    .X(_2286_));
 sg13g2_a21oi_1 _6147_ (.A1(net915),
    .A2(_2286_),
    .Y(_0266_),
    .B1(_2283_));
 sg13g2_xnor2_1 _6148_ (.Y(_2287_),
    .A(\vgademo.a_cos[10] ),
    .B(net961));
 sg13g2_o21ai_1 _6149_ (.B1(_3155_),
    .Y(_2288_),
    .A1(\vgademo.a_cos[8] ),
    .A2(\vgademo.a_cos[9] ));
 sg13g2_inv_1 _6150_ (.Y(_2289_),
    .A(_2288_));
 sg13g2_a21oi_1 _6151_ (.A1(_2281_),
    .A2(_2284_),
    .Y(_2290_),
    .B1(_2289_));
 sg13g2_nand2b_1 _6152_ (.Y(_2291_),
    .B(_2287_),
    .A_N(_2290_));
 sg13g2_xnor2_1 _6153_ (.Y(_2292_),
    .A(_2287_),
    .B(_2290_));
 sg13g2_nand2_1 _6154_ (.Y(_2293_),
    .A(net912),
    .B(_2292_));
 sg13g2_o21ai_1 _6155_ (.B1(_2293_),
    .Y(_0267_),
    .A1(_3146_),
    .A2(net912));
 sg13g2_nor2_1 _6156_ (.A(net532),
    .B(net913),
    .Y(_2294_));
 sg13g2_xnor2_1 _6157_ (.Y(_2295_),
    .A(\vgademo.a_cos[11] ),
    .B(net960));
 sg13g2_o21ai_1 _6158_ (.B1(_2291_),
    .Y(_2296_),
    .A1(_3146_),
    .A2(net960));
 sg13g2_xnor2_1 _6159_ (.Y(_2297_),
    .A(_2295_),
    .B(_2296_));
 sg13g2_a21oi_1 _6160_ (.A1(net913),
    .A2(_2297_),
    .Y(_0268_),
    .B1(_2294_));
 sg13g2_nor2_1 _6161_ (.A(net515),
    .B(net913),
    .Y(_2298_));
 sg13g2_nand4_1 _6162_ (.B(_2284_),
    .C(_2287_),
    .A(_2281_),
    .Y(_2299_),
    .D(_2295_));
 sg13g2_o21ai_1 _6163_ (.B1(_3155_),
    .Y(_2300_),
    .A1(\vgademo.a_cos[10] ),
    .A2(\vgademo.a_cos[11] ));
 sg13g2_nand3_1 _6164_ (.B(_2299_),
    .C(_2300_),
    .A(_2288_),
    .Y(_2301_));
 sg13g2_nor2b_1 _6165_ (.A(net960),
    .B_N(\vgademo.a_cos[12] ),
    .Y(_2302_));
 sg13g2_xnor2_1 _6166_ (.Y(_2303_),
    .A(\vgademo.a_cos[12] ),
    .B(net960));
 sg13g2_xnor2_1 _6167_ (.Y(_2304_),
    .A(_2301_),
    .B(_2303_));
 sg13g2_a21oi_1 _6168_ (.A1(net913),
    .A2(_2304_),
    .Y(_0269_),
    .B1(_2298_));
 sg13g2_nor2_1 _6169_ (.A(net215),
    .B(net913),
    .Y(_2305_));
 sg13g2_a21oi_1 _6170_ (.A1(_2301_),
    .A2(_2303_),
    .Y(_2306_),
    .B1(_2302_));
 sg13g2_nand2_1 _6171_ (.Y(_2307_),
    .A(\vgademo.a_cos[13] ),
    .B(_3155_));
 sg13g2_nor2_1 _6172_ (.A(\vgademo.a_cos[13] ),
    .B(_3155_),
    .Y(_2308_));
 sg13g2_xnor2_1 _6173_ (.Y(_2309_),
    .A(\vgademo.a_cos[13] ),
    .B(net960));
 sg13g2_xnor2_1 _6174_ (.Y(_2310_),
    .A(_2306_),
    .B(_2309_));
 sg13g2_a21oi_1 _6175_ (.A1(net913),
    .A2(_2310_),
    .Y(_0270_),
    .B1(_2305_));
 sg13g2_nor2_1 _6176_ (.A(net459),
    .B(net913),
    .Y(_2311_));
 sg13g2_o21ai_1 _6177_ (.B1(_2307_),
    .Y(_2312_),
    .A1(_2306_),
    .A2(_2308_));
 sg13g2_xnor2_1 _6178_ (.Y(_2313_),
    .A(\vgademo.a_cos[14] ),
    .B(net960));
 sg13g2_xnor2_1 _6179_ (.Y(_2314_),
    .A(_2312_),
    .B(_2313_));
 sg13g2_inv_2 _6180_ (.Y(_2315_),
    .A(net838));
 sg13g2_a21oi_1 _6181_ (.A1(net913),
    .A2(net838),
    .Y(_0271_),
    .B1(_2311_));
 sg13g2_xnor2_1 _6182_ (.Y(_0272_),
    .A(net253),
    .B(_2273_));
 sg13g2_nand2_1 _6183_ (.Y(_2316_),
    .A(net253),
    .B(_2272_));
 sg13g2_xnor2_1 _6184_ (.Y(_2317_),
    .A(net299),
    .B(_2277_));
 sg13g2_nor2_1 _6185_ (.A(_2316_),
    .B(_2317_),
    .Y(_2318_));
 sg13g2_nand2_1 _6186_ (.Y(_2319_),
    .A(net299),
    .B(net906));
 sg13g2_a21o_1 _6187_ (.A2(_2317_),
    .A1(_2316_),
    .B1(net906),
    .X(_2320_));
 sg13g2_o21ai_1 _6188_ (.B1(_2319_),
    .Y(_0273_),
    .A1(_2318_),
    .A2(_2320_));
 sg13g2_a21oi_1 _6189_ (.A1(net600),
    .A2(_2277_),
    .Y(_2321_),
    .B1(_2318_));
 sg13g2_and2_1 _6190_ (.A(\vgademo.a_sin[2] ),
    .B(_2282_),
    .X(_2322_));
 sg13g2_xnor2_1 _6191_ (.Y(_2323_),
    .A(\vgademo.a_sin[2] ),
    .B(_2282_));
 sg13g2_nor2_1 _6192_ (.A(_2321_),
    .B(_2323_),
    .Y(_2324_));
 sg13g2_nand2_1 _6193_ (.Y(_2325_),
    .A(net288),
    .B(net906));
 sg13g2_a21o_1 _6194_ (.A2(_2323_),
    .A1(_2321_),
    .B1(net906),
    .X(_2326_));
 sg13g2_o21ai_1 _6195_ (.B1(_2325_),
    .Y(_0274_),
    .A1(_2324_),
    .A2(_2326_));
 sg13g2_or2_1 _6196_ (.X(_2327_),
    .B(_2286_),
    .A(_3150_));
 sg13g2_xnor2_1 _6197_ (.Y(_2328_),
    .A(\vgademo.a_sin[3] ),
    .B(_2286_));
 sg13g2_o21ai_1 _6198_ (.B1(_2328_),
    .Y(_2329_),
    .A1(_2322_),
    .A2(_2324_));
 sg13g2_or3_1 _6199_ (.A(_2322_),
    .B(_2324_),
    .C(_2328_),
    .X(_2330_));
 sg13g2_nand3_1 _6200_ (.B(_2329_),
    .C(_2330_),
    .A(net909),
    .Y(_2331_));
 sg13g2_o21ai_1 _6201_ (.B1(_2331_),
    .Y(_0275_),
    .A1(_3150_),
    .A2(net909));
 sg13g2_and2_1 _6202_ (.A(\vgademo.a_sin[4] ),
    .B(_2292_),
    .X(_2332_));
 sg13g2_xnor2_1 _6203_ (.Y(_2333_),
    .A(\vgademo.a_sin[4] ),
    .B(_2292_));
 sg13g2_a21oi_1 _6204_ (.A1(_2327_),
    .A2(_2329_),
    .Y(_2334_),
    .B1(_2333_));
 sg13g2_nand3_1 _6205_ (.B(_2329_),
    .C(_2333_),
    .A(_2327_),
    .Y(_2335_));
 sg13g2_nand2_1 _6206_ (.Y(_2336_),
    .A(net312),
    .B(net907));
 sg13g2_nand2_1 _6207_ (.Y(_2337_),
    .A(net909),
    .B(_2335_));
 sg13g2_o21ai_1 _6208_ (.B1(_2336_),
    .Y(_0276_),
    .A1(_2334_),
    .A2(_2337_));
 sg13g2_nand2b_1 _6209_ (.Y(_2338_),
    .B(net349),
    .A_N(_2297_));
 sg13g2_xnor2_1 _6210_ (.Y(_2339_),
    .A(\vgademo.a_sin[5] ),
    .B(_2297_));
 sg13g2_o21ai_1 _6211_ (.B1(_2339_),
    .Y(_2340_),
    .A1(_2332_),
    .A2(_2334_));
 sg13g2_or3_1 _6212_ (.A(_2332_),
    .B(_2334_),
    .C(_2339_),
    .X(_2341_));
 sg13g2_nand3_1 _6213_ (.B(_2340_),
    .C(_2341_),
    .A(net912),
    .Y(_2342_));
 sg13g2_o21ai_1 _6214_ (.B1(_2342_),
    .Y(_0277_),
    .A1(_3151_),
    .A2(net909));
 sg13g2_nor2_1 _6215_ (.A(_3091_),
    .B(_2304_),
    .Y(_2343_));
 sg13g2_xnor2_1 _6216_ (.Y(_2344_),
    .A(_3091_),
    .B(_2304_));
 sg13g2_a21oi_1 _6217_ (.A1(_2338_),
    .A2(_2340_),
    .Y(_2345_),
    .B1(_2344_));
 sg13g2_nand3_1 _6218_ (.B(_2340_),
    .C(_2344_),
    .A(_2338_),
    .Y(_2346_));
 sg13g2_nand3b_1 _6219_ (.B(_2346_),
    .C(net909),
    .Y(_2347_),
    .A_N(_2345_));
 sg13g2_o21ai_1 _6220_ (.B1(_2347_),
    .Y(_0278_),
    .A1(_3091_),
    .A2(net909));
 sg13g2_nand2_1 _6221_ (.Y(_2348_),
    .A(\vgademo.a_sin[7] ),
    .B(_2310_));
 sg13g2_xnor2_1 _6222_ (.Y(_2349_),
    .A(_3152_),
    .B(_2310_));
 sg13g2_o21ai_1 _6223_ (.B1(_2349_),
    .Y(_2350_),
    .A1(_2343_),
    .A2(_2345_));
 sg13g2_or3_1 _6224_ (.A(_2343_),
    .B(_2345_),
    .C(_2349_),
    .X(_2351_));
 sg13g2_nand3_1 _6225_ (.B(_2350_),
    .C(_2351_),
    .A(net910),
    .Y(_2352_));
 sg13g2_o21ai_1 _6226_ (.B1(_2352_),
    .Y(_0279_),
    .A1(_3152_),
    .A2(net910));
 sg13g2_xor2_1 _6227_ (.B(net838),
    .A(\vgademo.a_sin[8] ),
    .X(_2353_));
 sg13g2_a21oi_1 _6228_ (.A1(_2348_),
    .A2(_2350_),
    .Y(_2354_),
    .B1(_2353_));
 sg13g2_nand3_1 _6229_ (.B(_2350_),
    .C(_2353_),
    .A(_2348_),
    .Y(_2355_));
 sg13g2_nand2_1 _6230_ (.Y(_2356_),
    .A(net469),
    .B(net906));
 sg13g2_nand2_1 _6231_ (.Y(_2357_),
    .A(net910),
    .B(_2355_));
 sg13g2_o21ai_1 _6232_ (.B1(_2356_),
    .Y(_0280_),
    .A1(_2354_),
    .A2(_2357_));
 sg13g2_nor2_1 _6233_ (.A(net501),
    .B(net914),
    .Y(_2358_));
 sg13g2_a21oi_1 _6234_ (.A1(\vgademo.a_sin[8] ),
    .A2(_2315_),
    .Y(_2359_),
    .B1(_2354_));
 sg13g2_xnor2_1 _6235_ (.Y(_2360_),
    .A(\vgademo.a_sin[9] ),
    .B(net838));
 sg13g2_xor2_1 _6236_ (.B(_2360_),
    .A(_2359_),
    .X(_2361_));
 sg13g2_a21oi_1 _6237_ (.A1(net910),
    .A2(_2361_),
    .Y(_0281_),
    .B1(_2358_));
 sg13g2_nor2_1 _6238_ (.A(net521),
    .B(net914),
    .Y(_2362_));
 sg13g2_o21ai_1 _6239_ (.B1(_2315_),
    .Y(_2363_),
    .A1(\vgademo.a_sin[8] ),
    .A2(\vgademo.a_sin[9] ));
 sg13g2_and2_1 _6240_ (.A(_2354_),
    .B(_2360_),
    .X(_2364_));
 sg13g2_nor2b_1 _6241_ (.A(_2364_),
    .B_N(_2363_),
    .Y(_2365_));
 sg13g2_nand2_1 _6242_ (.Y(_2366_),
    .A(\vgademo.a_sin[10] ),
    .B(_2315_));
 sg13g2_xor2_1 _6243_ (.B(net838),
    .A(\vgademo.a_sin[10] ),
    .X(_2367_));
 sg13g2_xnor2_1 _6244_ (.Y(_2368_),
    .A(_2365_),
    .B(_2367_));
 sg13g2_a21oi_1 _6245_ (.A1(net914),
    .A2(_2368_),
    .Y(_0282_),
    .B1(_2362_));
 sg13g2_nor2_1 _6246_ (.A(net531),
    .B(net914),
    .Y(_2369_));
 sg13g2_o21ai_1 _6247_ (.B1(_2366_),
    .Y(_2370_),
    .A1(_2365_),
    .A2(_2367_));
 sg13g2_xnor2_1 _6248_ (.Y(_2371_),
    .A(\vgademo.a_sin[11] ),
    .B(net838));
 sg13g2_xnor2_1 _6249_ (.Y(_2372_),
    .A(_2370_),
    .B(_2371_));
 sg13g2_a21oi_1 _6250_ (.A1(net914),
    .A2(_2372_),
    .Y(_0283_),
    .B1(_2369_));
 sg13g2_a21oi_1 _6251_ (.A1(_3153_),
    .A2(net838),
    .Y(_2373_),
    .B1(_2367_));
 sg13g2_o21ai_1 _6252_ (.B1(_2315_),
    .Y(_2374_),
    .A1(\vgademo.a_sin[10] ),
    .A2(\vgademo.a_sin[11] ));
 sg13g2_nand2_1 _6253_ (.Y(_2375_),
    .A(_2363_),
    .B(_2374_));
 sg13g2_a21oi_1 _6254_ (.A1(_2364_),
    .A2(_2373_),
    .Y(_2376_),
    .B1(_2375_));
 sg13g2_xnor2_1 _6255_ (.Y(_2377_),
    .A(\vgademo.a_sin[12] ),
    .B(net838));
 sg13g2_nor2b_1 _6256_ (.A(_2376_),
    .B_N(_2377_),
    .Y(_2378_));
 sg13g2_nor2b_1 _6257_ (.A(_2377_),
    .B_N(_2376_),
    .Y(_2379_));
 sg13g2_nor3_1 _6258_ (.A(net906),
    .B(_2378_),
    .C(_2379_),
    .Y(_2380_));
 sg13g2_a21o_1 _6259_ (.A2(net906),
    .A1(net544),
    .B1(_2380_),
    .X(_0284_));
 sg13g2_a21oi_1 _6260_ (.A1(\vgademo.a_sin[12] ),
    .A2(_2315_),
    .Y(_2381_),
    .B1(_2378_));
 sg13g2_xnor2_1 _6261_ (.Y(_2382_),
    .A(_2315_),
    .B(_2381_));
 sg13g2_nand2_1 _6262_ (.Y(_2383_),
    .A(net914),
    .B(_2382_));
 sg13g2_xnor2_1 _6263_ (.Y(_0285_),
    .A(net561),
    .B(_2383_));
 sg13g2_a21oi_1 _6264_ (.A1(_2314_),
    .A2(_2378_),
    .Y(_2384_),
    .B1(_3154_));
 sg13g2_a21oi_1 _6265_ (.A1(_2315_),
    .A2(_2381_),
    .Y(_2385_),
    .B1(\vgademo.a_sin[13] ));
 sg13g2_nor3_2 _6266_ (.A(net907),
    .B(_2384_),
    .C(_2385_),
    .Y(_2386_));
 sg13g2_xnor2_1 _6267_ (.Y(_0286_),
    .A(_3155_),
    .B(_2386_));
 sg13g2_and4_1 _6268_ (.A(\vgademo.h_count[10] ),
    .B(net1078),
    .C(_3227_),
    .D(_0575_),
    .X(_2387_));
 sg13g2_nand2_1 _6269_ (.Y(_2388_),
    .A(_0494_),
    .B(net899));
 sg13g2_o21ai_1 _6270_ (.B1(_2388_),
    .Y(_0287_),
    .A1(_3190_),
    .A2(net895));
 sg13g2_mux2_1 _6271_ (.A0(net379),
    .A1(_0508_),
    .S(net895),
    .X(_0288_));
 sg13g2_mux2_1 _6272_ (.A0(net362),
    .A1(_0522_),
    .S(net899),
    .X(_0289_));
 sg13g2_nand2_1 _6273_ (.Y(_2389_),
    .A(_0538_),
    .B(net895));
 sg13g2_o21ai_1 _6274_ (.B1(_2389_),
    .Y(_0290_),
    .A1(_3189_),
    .A2(net895));
 sg13g2_mux2_1 _6275_ (.A0(net485),
    .A1(_0552_),
    .S(net895),
    .X(_0291_));
 sg13g2_nand2_1 _6276_ (.Y(_2390_),
    .A(_0558_),
    .B(net895));
 sg13g2_o21ai_1 _6277_ (.B1(_2390_),
    .Y(_0292_),
    .A1(_3188_),
    .A2(net895));
 sg13g2_mux2_1 _6278_ (.A0(net468),
    .A1(_0557_),
    .S(net895),
    .X(_0293_));
 sg13g2_o21ai_1 _6279_ (.B1(net308),
    .Y(_2391_),
    .A1(_3135_),
    .A2(net918));
 sg13g2_nor2_2 _6280_ (.A(net308),
    .B(_3135_),
    .Y(_2392_));
 sg13g2_nor2_1 _6281_ (.A(net929),
    .B(net917),
    .Y(_2393_));
 sg13g2_nand2_2 _6282_ (.Y(_2394_),
    .A(net927),
    .B(net919));
 sg13g2_a22oi_1 _6283_ (.Y(_2395_),
    .B1(_2392_),
    .B2(_2393_),
    .A2(net892),
    .A1(\vgademo.a_cos[3] ));
 sg13g2_o21ai_1 _6284_ (.B1(_2395_),
    .Y(_0294_),
    .A1(net892),
    .A2(_2391_));
 sg13g2_nor2_1 _6285_ (.A(net343),
    .B(net920),
    .Y(_2396_));
 sg13g2_xnor2_1 _6286_ (.Y(_2397_),
    .A(\vgademo.b_cos[1] ),
    .B(\vgademo.b_sin[8] ));
 sg13g2_nor2b_1 _6287_ (.A(_2392_),
    .B_N(_2397_),
    .Y(_2398_));
 sg13g2_xor2_1 _6288_ (.B(_2397_),
    .A(_2392_),
    .X(_2399_));
 sg13g2_a221oi_1 _6289_ (.B2(_2399_),
    .C1(_2396_),
    .B1(net887),
    .A1(_3138_),
    .Y(_0295_),
    .A2(net892));
 sg13g2_a21oi_1 _6290_ (.A1(net343),
    .A2(_3137_),
    .Y(_2400_),
    .B1(_2398_));
 sg13g2_xnor2_1 _6291_ (.Y(_2401_),
    .A(net429),
    .B(\vgademo.b_sin[9] ));
 sg13g2_nor2b_1 _6292_ (.A(_2400_),
    .B_N(_2401_),
    .Y(_2402_));
 sg13g2_xor2_1 _6293_ (.B(_2401_),
    .A(_2400_),
    .X(_2403_));
 sg13g2_nand2b_1 _6294_ (.Y(_2404_),
    .B(net892),
    .A_N(\vgademo.a_cos[5] ));
 sg13g2_o21ai_1 _6295_ (.B1(_2404_),
    .Y(_2405_),
    .A1(net429),
    .A2(net920));
 sg13g2_a21oi_1 _6296_ (.A1(net887),
    .A2(_2403_),
    .Y(_0296_),
    .B1(net430));
 sg13g2_a21oi_1 _6297_ (.A1(\vgademo.b_cos[2] ),
    .A2(_3139_),
    .Y(_2406_),
    .B1(_2402_));
 sg13g2_xnor2_1 _6298_ (.Y(_2407_),
    .A(\vgademo.b_cos[3] ),
    .B(\vgademo.b_sin[10] ));
 sg13g2_nor2b_1 _6299_ (.A(_2406_),
    .B_N(_2407_),
    .Y(_2408_));
 sg13g2_xor2_1 _6300_ (.B(_2407_),
    .A(_2406_),
    .X(_2409_));
 sg13g2_nor2_1 _6301_ (.A(net385),
    .B(net920),
    .Y(_2410_));
 sg13g2_a221oi_1 _6302_ (.B2(_2409_),
    .C1(_2410_),
    .B1(net887),
    .A1(_3141_),
    .Y(_0297_),
    .A2(net892));
 sg13g2_a21oi_2 _6303_ (.B1(_2408_),
    .Y(_2411_),
    .A2(_3140_),
    .A1(net385));
 sg13g2_xnor2_1 _6304_ (.Y(_2412_),
    .A(\vgademo.b_cos[4] ),
    .B(net952));
 sg13g2_nor2b_1 _6305_ (.A(_2411_),
    .B_N(_2412_),
    .Y(_2413_));
 sg13g2_xor2_1 _6306_ (.B(_2412_),
    .A(_2411_),
    .X(_2414_));
 sg13g2_nor2_1 _6307_ (.A(net407),
    .B(net919),
    .Y(_2415_));
 sg13g2_a221oi_1 _6308_ (.B2(_2414_),
    .C1(_2415_),
    .B1(net887),
    .A1(_3143_),
    .Y(_0298_),
    .A2(net893));
 sg13g2_xnor2_1 _6309_ (.Y(_2416_),
    .A(net952),
    .B(\vgademo.b_cos[5] ));
 sg13g2_a21oi_1 _6310_ (.A1(\vgademo.b_cos[4] ),
    .A2(_3142_),
    .Y(_2417_),
    .B1(_2413_));
 sg13g2_a21o_1 _6311_ (.A2(net919),
    .A1(\vgademo.a_cos[8] ),
    .B1(net887),
    .X(_2418_));
 sg13g2_xnor2_1 _6312_ (.Y(_2419_),
    .A(_2416_),
    .B(_2417_));
 sg13g2_o21ai_1 _6313_ (.B1(_2418_),
    .Y(_2420_),
    .A1(net931),
    .A2(_2419_));
 sg13g2_o21ai_1 _6314_ (.B1(_2420_),
    .Y(_0299_),
    .A1(_3144_),
    .A2(net919));
 sg13g2_o21ai_1 _6315_ (.B1(_3142_),
    .Y(_2421_),
    .A1(\vgademo.b_cos[4] ),
    .A2(\vgademo.b_cos[5] ));
 sg13g2_nand2_1 _6316_ (.Y(_2422_),
    .A(_2413_),
    .B(_2416_));
 sg13g2_xor2_1 _6317_ (.B(net959),
    .A(net952),
    .X(_2423_));
 sg13g2_a21oi_1 _6318_ (.A1(_2421_),
    .A2(_2422_),
    .Y(_2424_),
    .B1(_2423_));
 sg13g2_nand3_1 _6319_ (.B(_2422_),
    .C(_2423_),
    .A(_2421_),
    .Y(_2425_));
 sg13g2_nand2_1 _6320_ (.Y(_2426_),
    .A(net886),
    .B(_2425_));
 sg13g2_a22oi_1 _6321_ (.Y(_2427_),
    .B1(net891),
    .B2(net568),
    .A2(net916),
    .A1(net959));
 sg13g2_o21ai_1 _6322_ (.B1(net569),
    .Y(_0300_),
    .A1(_2424_),
    .A2(_2426_));
 sg13g2_xnor2_1 _6323_ (.Y(_2428_),
    .A(net951),
    .B(\vgademo.b_cos[7] ));
 sg13g2_a21oi_1 _6324_ (.A1(_3142_),
    .A2(net959),
    .Y(_2429_),
    .B1(_2424_));
 sg13g2_xnor2_1 _6325_ (.Y(_2430_),
    .A(_2428_),
    .B(_2429_));
 sg13g2_nand2_1 _6326_ (.Y(_2431_),
    .A(net488),
    .B(net891));
 sg13g2_a22oi_1 _6327_ (.Y(_2432_),
    .B1(net886),
    .B2(_2430_),
    .A2(net916),
    .A1(\vgademo.b_cos[7] ));
 sg13g2_nand2_1 _6328_ (.Y(_0301_),
    .A(_2431_),
    .B(_2432_));
 sg13g2_nor2_1 _6329_ (.A(_2422_),
    .B(_2423_),
    .Y(_2433_));
 sg13g2_o21ai_1 _6330_ (.B1(_3142_),
    .Y(_2434_),
    .A1(net959),
    .A2(\vgademo.b_cos[7] ));
 sg13g2_nand2_1 _6331_ (.Y(_2435_),
    .A(_2421_),
    .B(_2434_));
 sg13g2_a21oi_2 _6332_ (.B1(_2435_),
    .Y(_2436_),
    .A2(_2433_),
    .A1(_2428_));
 sg13g2_inv_1 _6333_ (.Y(_2437_),
    .A(_2436_));
 sg13g2_nor2b_1 _6334_ (.A(net951),
    .B_N(net958),
    .Y(_2438_));
 sg13g2_xnor2_1 _6335_ (.Y(_2439_),
    .A(net951),
    .B(net958));
 sg13g2_inv_1 _6336_ (.Y(_2440_),
    .A(_2439_));
 sg13g2_xnor2_1 _6337_ (.Y(_2441_),
    .A(_2436_),
    .B(_2439_));
 sg13g2_nand2_1 _6338_ (.Y(_2442_),
    .A(net532),
    .B(net891));
 sg13g2_a22oi_1 _6339_ (.Y(_2443_),
    .B1(net886),
    .B2(_2441_),
    .A2(net916),
    .A1(net958));
 sg13g2_nand2_1 _6340_ (.Y(_0302_),
    .A(_2442_),
    .B(_2443_));
 sg13g2_nor2_1 _6341_ (.A(net951),
    .B(_3147_),
    .Y(_2444_));
 sg13g2_xor2_1 _6342_ (.B(net957),
    .A(net951),
    .X(_2445_));
 sg13g2_a21oi_1 _6343_ (.A1(_2437_),
    .A2(_2439_),
    .Y(_2446_),
    .B1(_2438_));
 sg13g2_xor2_1 _6344_ (.B(_2446_),
    .A(_2445_),
    .X(_2447_));
 sg13g2_nand2_1 _6345_ (.Y(_2448_),
    .A(net515),
    .B(net891));
 sg13g2_a22oi_1 _6346_ (.Y(_2449_),
    .B1(net886),
    .B2(_2447_),
    .A2(net916),
    .A1(net957));
 sg13g2_nand2_1 _6347_ (.Y(_0303_),
    .A(_2448_),
    .B(_2449_));
 sg13g2_nor3_1 _6348_ (.A(_2436_),
    .B(_2440_),
    .C(_2445_),
    .Y(_2450_));
 sg13g2_nor3_1 _6349_ (.A(_2438_),
    .B(_2444_),
    .C(_2450_),
    .Y(_2451_));
 sg13g2_xnor2_1 _6350_ (.Y(_2452_),
    .A(net951),
    .B(net956));
 sg13g2_nand2b_1 _6351_ (.Y(_2453_),
    .B(_2452_),
    .A_N(_2451_));
 sg13g2_xnor2_1 _6352_ (.Y(_2454_),
    .A(_2451_),
    .B(_2452_));
 sg13g2_a22oi_1 _6353_ (.Y(_2455_),
    .B1(net886),
    .B2(_2454_),
    .A2(net891),
    .A1(net580));
 sg13g2_o21ai_1 _6354_ (.B1(_2455_),
    .Y(_0304_),
    .A1(_3148_),
    .A2(net919));
 sg13g2_o21ai_1 _6355_ (.B1(_2453_),
    .Y(_2456_),
    .A1(net951),
    .A2(_3148_));
 sg13g2_xor2_1 _6356_ (.B(\vgademo.b_cos[11] ),
    .A(net951),
    .X(_2457_));
 sg13g2_xnor2_1 _6357_ (.Y(_2458_),
    .A(_2456_),
    .B(_2457_));
 sg13g2_a22oi_1 _6358_ (.Y(_2459_),
    .B1(net886),
    .B2(_2458_),
    .A2(net891),
    .A1(net459));
 sg13g2_o21ai_1 _6359_ (.B1(_2459_),
    .Y(_0305_),
    .A1(_3149_),
    .A2(net919));
 sg13g2_mux2_1 _6360_ (.A0(net340),
    .A1(_0225_),
    .S(_0663_),
    .X(_0306_));
 sg13g2_nand2b_1 _6361_ (.Y(_2460_),
    .B(net900),
    .A_N(net508));
 sg13g2_xor2_1 _6362_ (.B(\vgademo.plane_dx_div.d[17] ),
    .A(\vgademo.plane_dx_div.d[16] ),
    .X(_2461_));
 sg13g2_nor2_1 _6363_ (.A(net953),
    .B(_2461_),
    .Y(_2462_));
 sg13g2_a21oi_1 _6364_ (.A1(net953),
    .A2(_0070_),
    .Y(_2463_),
    .B1(_2462_));
 sg13g2_nand2_1 _6365_ (.Y(_2464_),
    .A(net340),
    .B(_2463_));
 sg13g2_xnor2_1 _6366_ (.Y(_2465_),
    .A(net340),
    .B(_2463_));
 sg13g2_a21oi_1 _6367_ (.A1(net902),
    .A2(_2465_),
    .Y(_2466_),
    .B1(_1092_));
 sg13g2_o21ai_1 _6368_ (.B1(_2460_),
    .Y(_2467_),
    .A1(_1101_),
    .A2(_2466_));
 sg13g2_a21oi_1 _6369_ (.A1(_1091_),
    .A2(_1101_),
    .Y(_0307_),
    .B1(_2467_));
 sg13g2_nor2_1 _6370_ (.A(_1091_),
    .B(_1100_),
    .Y(_2468_));
 sg13g2_nor2_1 _6371_ (.A(_1111_),
    .B(_2468_),
    .Y(_2469_));
 sg13g2_xnor2_1 _6372_ (.Y(_2470_),
    .A(_1111_),
    .B(_2468_));
 sg13g2_nor2_1 _6373_ (.A(net358),
    .B(_0663_),
    .Y(_2471_));
 sg13g2_o21ai_1 _6374_ (.B1(\vgademo.plane_dx_div.d[18] ),
    .Y(_2472_),
    .A1(\vgademo.plane_dx_div.d[16] ),
    .A2(\vgademo.plane_dx_div.d[17] ));
 sg13g2_or3_2 _6375_ (.A(\vgademo.plane_dx_div.d[16] ),
    .B(\vgademo.plane_dx_div.d[17] ),
    .C(\vgademo.plane_dx_div.d[18] ),
    .X(_2473_));
 sg13g2_a21oi_1 _6376_ (.A1(_2472_),
    .A2(_2473_),
    .Y(_2474_),
    .B1(net953));
 sg13g2_a21oi_1 _6377_ (.A1(net953),
    .A2(_0073_),
    .Y(_2475_),
    .B1(_2474_));
 sg13g2_nand2_1 _6378_ (.Y(_2476_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_2475_));
 sg13g2_xnor2_1 _6379_ (.Y(_2477_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_2475_));
 sg13g2_xnor2_1 _6380_ (.Y(_2478_),
    .A(_2464_),
    .B(_2477_));
 sg13g2_a221oi_1 _6381_ (.B2(net902),
    .C1(_2471_),
    .B1(_2478_),
    .A1(net935),
    .Y(_0308_),
    .A2(_2470_));
 sg13g2_nand2_1 _6382_ (.Y(_2479_),
    .A(_1127_),
    .B(_2469_));
 sg13g2_xnor2_1 _6383_ (.Y(_2480_),
    .A(_1127_),
    .B(_2469_));
 sg13g2_nor2_1 _6384_ (.A(net365),
    .B(_0663_),
    .Y(_2481_));
 sg13g2_o21ai_1 _6385_ (.B1(_2476_),
    .Y(_2482_),
    .A1(_2464_),
    .A2(_2477_));
 sg13g2_xor2_1 _6386_ (.B(_2473_),
    .A(\vgademo.plane_dx_div.d[19] ),
    .X(_2483_));
 sg13g2_nor2_1 _6387_ (.A(net953),
    .B(_2483_),
    .Y(_2484_));
 sg13g2_a21oi_1 _6388_ (.A1(net953),
    .A2(_0076_),
    .Y(_2485_),
    .B1(_2484_));
 sg13g2_and2_1 _6389_ (.A(\vgademo.plane_dx_div.r[18] ),
    .B(_2485_),
    .X(_2486_));
 sg13g2_xor2_1 _6390_ (.B(_2485_),
    .A(net358),
    .X(_2487_));
 sg13g2_xnor2_1 _6391_ (.Y(_2488_),
    .A(_2482_),
    .B(_2487_));
 sg13g2_a221oi_1 _6392_ (.B2(net902),
    .C1(_2481_),
    .B1(_2488_),
    .A1(net935),
    .Y(_0309_),
    .A2(_2480_));
 sg13g2_nor2_1 _6393_ (.A(_1141_),
    .B(_2479_),
    .Y(_2489_));
 sg13g2_xnor2_1 _6394_ (.Y(_2490_),
    .A(_1141_),
    .B(_2479_));
 sg13g2_nor2_1 _6395_ (.A(net278),
    .B(_0663_),
    .Y(_2491_));
 sg13g2_a21oi_1 _6396_ (.A1(_2482_),
    .A2(_2487_),
    .Y(_2492_),
    .B1(_2486_));
 sg13g2_o21ai_1 _6397_ (.B1(\vgademo.plane_dx_div.d[20] ),
    .Y(_2493_),
    .A1(\vgademo.plane_dx_div.d[19] ),
    .A2(_2473_));
 sg13g2_or3_2 _6398_ (.A(\vgademo.plane_dx_div.d[19] ),
    .B(\vgademo.plane_dx_div.d[20] ),
    .C(_2473_),
    .X(_2494_));
 sg13g2_a21oi_1 _6399_ (.A1(_2493_),
    .A2(_2494_),
    .Y(_2495_),
    .B1(net953));
 sg13g2_a21oi_1 _6400_ (.A1(net953),
    .A2(_0079_),
    .Y(_2496_),
    .B1(_2495_));
 sg13g2_nand2_1 _6401_ (.Y(_2497_),
    .A(\vgademo.plane_dx_div.r[19] ),
    .B(_2496_));
 sg13g2_xnor2_1 _6402_ (.Y(_2498_),
    .A(\vgademo.plane_dx_div.r[19] ),
    .B(_2496_));
 sg13g2_xnor2_1 _6403_ (.Y(_2499_),
    .A(_2492_),
    .B(_2498_));
 sg13g2_a221oi_1 _6404_ (.B2(net902),
    .C1(_2491_),
    .B1(_2499_),
    .A1(net935),
    .Y(_0310_),
    .A2(_2490_));
 sg13g2_nand2b_1 _6405_ (.Y(_2500_),
    .B(_2489_),
    .A_N(_1157_));
 sg13g2_xor2_1 _6406_ (.B(_2489_),
    .A(_1157_),
    .X(_2501_));
 sg13g2_nor2_1 _6407_ (.A(net363),
    .B(_0663_),
    .Y(_2502_));
 sg13g2_o21ai_1 _6408_ (.B1(_2497_),
    .Y(_2503_),
    .A1(_2492_),
    .A2(_2498_));
 sg13g2_xor2_1 _6409_ (.B(_2494_),
    .A(\vgademo.plane_dx_div.d[21] ),
    .X(_2504_));
 sg13g2_nor2_1 _6410_ (.A(net954),
    .B(_2504_),
    .Y(_2505_));
 sg13g2_and2_1 _6411_ (.A(net954),
    .B(_0013_),
    .X(_2506_));
 sg13g2_nor3_1 _6412_ (.A(_3122_),
    .B(_2505_),
    .C(_2506_),
    .Y(_2507_));
 sg13g2_o21ai_1 _6413_ (.B1(_3122_),
    .Y(_2508_),
    .A1(_2505_),
    .A2(_2506_));
 sg13g2_nor2b_1 _6414_ (.A(_2507_),
    .B_N(_2508_),
    .Y(_2509_));
 sg13g2_xnor2_1 _6415_ (.Y(_2510_),
    .A(_2503_),
    .B(_2509_));
 sg13g2_a221oi_1 _6416_ (.B2(net903),
    .C1(_2502_),
    .B1(_2510_),
    .A1(net936),
    .Y(_0311_),
    .A2(_2501_));
 sg13g2_nand2b_1 _6417_ (.Y(_2511_),
    .B(_1175_),
    .A_N(_2500_));
 sg13g2_xor2_1 _6418_ (.B(_2500_),
    .A(_1175_),
    .X(_2512_));
 sg13g2_nor2_1 _6419_ (.A(net360),
    .B(_0663_),
    .Y(_2513_));
 sg13g2_a21oi_1 _6420_ (.A1(_2503_),
    .A2(_2508_),
    .Y(_2514_),
    .B1(_2507_));
 sg13g2_nand2b_1 _6421_ (.Y(_2515_),
    .B(net954),
    .A_N(_0014_));
 sg13g2_o21ai_1 _6422_ (.B1(\vgademo.plane_dx_div.d[22] ),
    .Y(_2516_),
    .A1(\vgademo.plane_dx_div.d[21] ),
    .A2(_2494_));
 sg13g2_nor3_2 _6423_ (.A(\vgademo.plane_dx_div.d[21] ),
    .B(\vgademo.plane_dx_div.d[22] ),
    .C(_2494_),
    .Y(_2517_));
 sg13g2_nand2b_1 _6424_ (.Y(_2518_),
    .B(_2516_),
    .A_N(net954));
 sg13g2_o21ai_1 _6425_ (.B1(_2515_),
    .Y(_2519_),
    .A1(_2517_),
    .A2(_2518_));
 sg13g2_nor2_1 _6426_ (.A(\vgademo.plane_dx_div.r[21] ),
    .B(_2519_),
    .Y(_2520_));
 sg13g2_and2_1 _6427_ (.A(\vgademo.plane_dx_div.r[21] ),
    .B(_2519_),
    .X(_2521_));
 sg13g2_nor2_1 _6428_ (.A(_2520_),
    .B(_2521_),
    .Y(_2522_));
 sg13g2_xor2_1 _6429_ (.B(_2522_),
    .A(_2514_),
    .X(_2523_));
 sg13g2_a221oi_1 _6430_ (.B2(net903),
    .C1(_2513_),
    .B1(_2523_),
    .A1(net936),
    .Y(_0312_),
    .A2(_2512_));
 sg13g2_nand2_1 _6431_ (.Y(_2524_),
    .A(_1191_),
    .B(_2511_));
 sg13g2_nor2_1 _6432_ (.A(_1191_),
    .B(_2511_),
    .Y(_2525_));
 sg13g2_nand2b_1 _6433_ (.Y(_2526_),
    .B(\vgademo.plane_dx_div.d[23] ),
    .A_N(_2517_));
 sg13g2_nand2b_1 _6434_ (.Y(_2527_),
    .B(_2517_),
    .A_N(\vgademo.plane_dx_div.d[23] ));
 sg13g2_a21oi_1 _6435_ (.A1(_2526_),
    .A2(_2527_),
    .Y(_2528_),
    .B1(net954));
 sg13g2_a21oi_1 _6436_ (.A1(net954),
    .A2(_0018_),
    .Y(_2529_),
    .B1(_2528_));
 sg13g2_and2_1 _6437_ (.A(\vgademo.plane_dx_div.r[22] ),
    .B(_2529_),
    .X(_2530_));
 sg13g2_xor2_1 _6438_ (.B(_2529_),
    .A(\vgademo.plane_dx_div.r[22] ),
    .X(_2531_));
 sg13g2_nor2b_1 _6439_ (.A(_2521_),
    .B_N(_2514_),
    .Y(_2532_));
 sg13g2_nor2_1 _6440_ (.A(_2520_),
    .B(_2532_),
    .Y(_2533_));
 sg13g2_and2_1 _6441_ (.A(_2531_),
    .B(_2533_),
    .X(_2534_));
 sg13g2_xor2_1 _6442_ (.B(_2533_),
    .A(_2531_),
    .X(_2535_));
 sg13g2_nor2_1 _6443_ (.A(_0660_),
    .B(_2525_),
    .Y(_2536_));
 sg13g2_a221oi_1 _6444_ (.B2(_2524_),
    .C1(net900),
    .B1(_2536_),
    .A1(_0660_),
    .Y(_2537_),
    .A2(_2535_));
 sg13g2_a21oi_1 _6445_ (.A1(_3126_),
    .A2(net901),
    .Y(_0313_),
    .B1(_2537_));
 sg13g2_o21ai_1 _6446_ (.B1(_1200_),
    .Y(_2538_),
    .A1(_1191_),
    .A2(_2511_));
 sg13g2_nand2_1 _6447_ (.Y(_2539_),
    .A(\vgademo.plane_dx_div.d[24] ),
    .B(_2527_));
 sg13g2_nor2_1 _6448_ (.A(\vgademo.plane_dx_div.d[24] ),
    .B(_2527_),
    .Y(_2540_));
 sg13g2_nor2_1 _6449_ (.A(\vgademo.plane_dx_div.r[25] ),
    .B(_2540_),
    .Y(_2541_));
 sg13g2_a22oi_1 _6450_ (.Y(_2542_),
    .B1(_2539_),
    .B2(_2541_),
    .A2(_3125_),
    .A1(net955));
 sg13g2_xnor2_1 _6451_ (.Y(_2543_),
    .A(\vgademo.plane_dx_div.r[23] ),
    .B(_2542_));
 sg13g2_nor3_1 _6452_ (.A(_2530_),
    .B(_2534_),
    .C(_2543_),
    .Y(_2544_));
 sg13g2_o21ai_1 _6453_ (.B1(_2543_),
    .Y(_2545_),
    .A1(_2530_),
    .A2(_2534_));
 sg13g2_nor2b_1 _6454_ (.A(_2544_),
    .B_N(_2545_),
    .Y(_2546_));
 sg13g2_or2_1 _6455_ (.X(_2547_),
    .B(_2536_),
    .A(_1201_));
 sg13g2_a221oi_1 _6456_ (.B2(_2538_),
    .C1(net901),
    .B1(_2547_),
    .A1(_0660_),
    .Y(_2548_),
    .A2(_2546_));
 sg13g2_a21oi_1 _6457_ (.A1(_3127_),
    .A2(net900),
    .Y(_0314_),
    .B1(_2548_));
 sg13g2_nor2_1 _6458_ (.A(net345),
    .B(_0663_),
    .Y(_2549_));
 sg13g2_o21ai_1 _6459_ (.B1(_2545_),
    .Y(_2550_),
    .A1(_3126_),
    .A2(_2542_));
 sg13g2_xnor2_1 _6460_ (.Y(_2551_),
    .A(\vgademo.plane_dx_div.r[24] ),
    .B(_2541_));
 sg13g2_xnor2_1 _6461_ (.Y(_2552_),
    .A(_2550_),
    .B(_2551_));
 sg13g2_a21oi_1 _6462_ (.A1(_0660_),
    .A2(_2552_),
    .Y(_2553_),
    .B1(_2547_));
 sg13g2_a21oi_1 _6463_ (.A1(_0663_),
    .A2(_2553_),
    .Y(_0315_),
    .B1(_2549_));
 sg13g2_and2_1 _6464_ (.A(net863),
    .B(_2203_),
    .X(_2554_));
 sg13g2_nor2_1 _6465_ (.A(_1734_),
    .B(_1774_),
    .Y(_2555_));
 sg13g2_nor2_2 _6466_ (.A(_1804_),
    .B(_2555_),
    .Y(_2556_));
 sg13g2_nor2_1 _6467_ (.A(net860),
    .B(_2556_),
    .Y(_2557_));
 sg13g2_nand2_1 _6468_ (.Y(_2558_),
    .A(net826),
    .B(_2557_));
 sg13g2_nand2_1 _6469_ (.Y(_2559_),
    .A(_1691_),
    .B(_2106_));
 sg13g2_a21oi_1 _6470_ (.A1(_2105_),
    .A2(_2108_),
    .Y(_2560_),
    .B1(_1690_));
 sg13g2_nor2_1 _6471_ (.A(_1683_),
    .B(_2209_),
    .Y(_2561_));
 sg13g2_a221oi_1 _6472_ (.B2(_2558_),
    .C1(net862),
    .B1(_2561_),
    .A1(net827),
    .Y(_2562_),
    .A2(_2560_));
 sg13g2_nor2_2 _6473_ (.A(_2554_),
    .B(_2562_),
    .Y(_2563_));
 sg13g2_nor2_1 _6474_ (.A(net827),
    .B(_2138_),
    .Y(_2564_));
 sg13g2_o21ai_1 _6475_ (.B1(_1808_),
    .Y(_2565_),
    .A1(net844),
    .A2(_2122_));
 sg13g2_nand3_1 _6476_ (.B(net826),
    .C(_2565_),
    .A(net854),
    .Y(_2566_));
 sg13g2_a22oi_1 _6477_ (.Y(_2567_),
    .B1(_2564_),
    .B2(_2566_),
    .A2(_2559_),
    .A1(_2110_));
 sg13g2_nor2_1 _6478_ (.A(net863),
    .B(_2567_),
    .Y(_2568_));
 sg13g2_or2_1 _6479_ (.X(_2569_),
    .B(_2567_),
    .A(net862));
 sg13g2_a21oi_1 _6480_ (.A1(_2223_),
    .A2(_2568_),
    .Y(_2570_),
    .B1(_2563_));
 sg13g2_inv_1 _6481_ (.Y(_2571_),
    .A(_2570_));
 sg13g2_o21ai_1 _6482_ (.B1(_2563_),
    .Y(_2572_),
    .A1(net942),
    .A2(_2568_));
 sg13g2_nor2b_1 _6483_ (.A(_2570_),
    .B_N(_2572_),
    .Y(_2573_));
 sg13g2_inv_1 _6484_ (.Y(_2574_),
    .A(_2573_));
 sg13g2_nor2b_2 _6485_ (.A(_2119_),
    .B_N(_1775_),
    .Y(_2575_));
 sg13g2_o21ai_1 _6486_ (.B1(_2575_),
    .Y(_2576_),
    .A1(net828),
    .A2(net852));
 sg13g2_nand3_1 _6487_ (.B(net853),
    .C(_2556_),
    .A(net830),
    .Y(_2577_));
 sg13g2_nand3_1 _6488_ (.B(_2576_),
    .C(_2577_),
    .A(net854),
    .Y(_2578_));
 sg13g2_a21oi_2 _6489_ (.B1(net827),
    .Y(_2579_),
    .A2(_2578_),
    .A1(_2128_));
 sg13g2_nor2_1 _6490_ (.A(_2114_),
    .B(_2579_),
    .Y(_2580_));
 sg13g2_o21ai_1 _6491_ (.B1(_2147_),
    .Y(_2581_),
    .A1(_2114_),
    .A2(_2579_));
 sg13g2_or3_1 _6492_ (.A(_2114_),
    .B(_2147_),
    .C(_2579_),
    .X(_2582_));
 sg13g2_nand3_1 _6493_ (.B(_2581_),
    .C(_2582_),
    .A(_2569_),
    .Y(_2583_));
 sg13g2_nand2_1 _6494_ (.Y(_2584_),
    .A(_2581_),
    .B(_2583_));
 sg13g2_xnor2_1 _6495_ (.Y(_2585_),
    .A(net942),
    .B(_2569_));
 sg13g2_xnor2_1 _6496_ (.Y(_2586_),
    .A(_2563_),
    .B(_2585_));
 sg13g2_or2_1 _6497_ (.X(_2587_),
    .B(_2586_),
    .A(_2584_));
 sg13g2_inv_1 _6498_ (.Y(_2588_),
    .A(_2587_));
 sg13g2_nand2_1 _6499_ (.Y(_2589_),
    .A(_2155_),
    .B(_2170_));
 sg13g2_o21ai_1 _6500_ (.B1(_2589_),
    .Y(_2590_),
    .A1(net829),
    .A2(_1716_));
 sg13g2_nand2_1 _6501_ (.Y(_2591_),
    .A(_1805_),
    .B(_2117_));
 sg13g2_nand3_1 _6502_ (.B(net853),
    .C(_2591_),
    .A(net831),
    .Y(_2592_));
 sg13g2_nand3_1 _6503_ (.B(_2590_),
    .C(_2592_),
    .A(net856),
    .Y(_2593_));
 sg13g2_a21oi_1 _6504_ (.A1(_2095_),
    .A2(_2593_),
    .Y(_2594_),
    .B1(net862));
 sg13g2_nor2_1 _6505_ (.A(_2101_),
    .B(_2594_),
    .Y(_2595_));
 sg13g2_nand2_1 _6506_ (.Y(_2596_),
    .A(_1780_),
    .B(_2171_));
 sg13g2_a21oi_1 _6507_ (.A1(_1717_),
    .A2(_2596_),
    .Y(_2597_),
    .B1(net860));
 sg13g2_o21ai_1 _6508_ (.B1(_2597_),
    .Y(_2598_),
    .A1(net826),
    .A2(_2575_));
 sg13g2_a21oi_2 _6509_ (.B1(net862),
    .Y(_2599_),
    .A2(_2598_),
    .A1(_2165_));
 sg13g2_xnor2_1 _6510_ (.Y(_2600_),
    .A(_2101_),
    .B(_2594_));
 sg13g2_nor2_1 _6511_ (.A(_2599_),
    .B(_2600_),
    .Y(_2601_));
 sg13g2_nand3_1 _6512_ (.B(_1715_),
    .C(_2565_),
    .A(net830),
    .Y(_2602_));
 sg13g2_o21ai_1 _6513_ (.B1(_2591_),
    .Y(_2603_),
    .A1(net829),
    .A2(_1716_));
 sg13g2_nand3_1 _6514_ (.B(_2602_),
    .C(_2603_),
    .A(net854),
    .Y(_2604_));
 sg13g2_nand2_1 _6515_ (.Y(_2605_),
    .A(_1691_),
    .B(_2105_));
 sg13g2_or4_1 _6516_ (.A(net829),
    .B(_1682_),
    .C(_2109_),
    .D(_2605_),
    .X(_2606_));
 sg13g2_nand3_1 _6517_ (.B(_2143_),
    .C(_2606_),
    .A(net861),
    .Y(_2607_));
 sg13g2_a21oi_1 _6518_ (.A1(_2096_),
    .A2(_2604_),
    .Y(_2608_),
    .B1(_2607_));
 sg13g2_or2_1 _6519_ (.X(_2609_),
    .B(_2608_),
    .A(_2102_));
 sg13g2_xnor2_1 _6520_ (.Y(_2610_),
    .A(_2102_),
    .B(_2608_));
 sg13g2_xor2_1 _6521_ (.B(_2610_),
    .A(_2580_),
    .X(_2611_));
 sg13g2_or3_1 _6522_ (.A(_2595_),
    .B(_2601_),
    .C(_2611_),
    .X(_2612_));
 sg13g2_xor2_1 _6523_ (.B(_2600_),
    .A(_2599_),
    .X(_2613_));
 sg13g2_nand2b_1 _6524_ (.Y(_2614_),
    .B(_2562_),
    .A_N(_2214_));
 sg13g2_a22oi_1 _6525_ (.Y(_2615_),
    .B1(_2599_),
    .B2(_2614_),
    .A2(_2563_),
    .A1(_2214_));
 sg13g2_or2_1 _6526_ (.X(_2616_),
    .B(_2615_),
    .A(_2613_));
 sg13g2_o21ai_1 _6527_ (.B1(_2611_),
    .Y(_2617_),
    .A1(_2595_),
    .A2(_2601_));
 sg13g2_and3_1 _6528_ (.X(_2618_),
    .A(_2612_),
    .B(_2616_),
    .C(_2617_));
 sg13g2_a221oi_1 _6529_ (.B2(_2615_),
    .C1(_2607_),
    .B1(_2613_),
    .A1(_2096_),
    .Y(_2619_),
    .A2(_2604_));
 sg13g2_o21ai_1 _6530_ (.B1(_2609_),
    .Y(_2620_),
    .A1(_2580_),
    .A2(_2610_));
 sg13g2_a21o_1 _6531_ (.A2(_2582_),
    .A1(_2581_),
    .B1(_2569_),
    .X(_2621_));
 sg13g2_and3_1 _6532_ (.X(_2622_),
    .A(_2583_),
    .B(_2620_),
    .C(_2621_));
 sg13g2_nand3_1 _6533_ (.B(_2620_),
    .C(_2621_),
    .A(_2583_),
    .Y(_2623_));
 sg13g2_a21oi_1 _6534_ (.A1(_2583_),
    .A2(_2621_),
    .Y(_2624_),
    .B1(_2620_));
 sg13g2_nor3_1 _6535_ (.A(_2619_),
    .B(_2622_),
    .C(_2624_),
    .Y(_2625_));
 sg13g2_o21ai_1 _6536_ (.B1(_2623_),
    .Y(_2626_),
    .A1(_2617_),
    .A2(_2624_));
 sg13g2_a221oi_1 _6537_ (.B2(_2625_),
    .C1(_2626_),
    .B1(_2618_),
    .A1(_2584_),
    .Y(_2627_),
    .A2(_2586_));
 sg13g2_o21ai_1 _6538_ (.B1(_2574_),
    .Y(_2628_),
    .A1(_2588_),
    .A2(_2627_));
 sg13g2_nand3b_1 _6539_ (.B(_2573_),
    .C(_2587_),
    .Y(_2629_),
    .A_N(_2627_));
 sg13g2_and3_1 _6540_ (.X(_0316_),
    .A(_2239_),
    .B(_2628_),
    .C(_2629_));
 sg13g2_a21oi_1 _6541_ (.A1(_2571_),
    .A2(_2629_),
    .Y(_0317_),
    .B1(_2238_));
 sg13g2_nand2_1 _6542_ (.Y(_2630_),
    .A(\vgademo.b_sin[0] ),
    .B(_2430_));
 sg13g2_xnor2_1 _6543_ (.Y(_2631_),
    .A(\vgademo.b_sin[0] ),
    .B(_2430_));
 sg13g2_a22oi_1 _6544_ (.Y(_2632_),
    .B1(net891),
    .B2(net382),
    .A2(net916),
    .A1(\vgademo.b_sin[0] ));
 sg13g2_o21ai_1 _6545_ (.B1(net383),
    .Y(_0318_),
    .A1(_2394_),
    .A2(_2631_));
 sg13g2_nand2_1 _6546_ (.Y(_2633_),
    .A(\vgademo.b_sin[1] ),
    .B(_2441_));
 sg13g2_xnor2_1 _6547_ (.Y(_2634_),
    .A(\vgademo.b_sin[1] ),
    .B(_2441_));
 sg13g2_xnor2_1 _6548_ (.Y(_2635_),
    .A(_2630_),
    .B(_2634_));
 sg13g2_a22oi_1 _6549_ (.Y(_2636_),
    .B1(net894),
    .B2(net312),
    .A2(net916),
    .A1(\vgademo.b_sin[1] ));
 sg13g2_o21ai_1 _6550_ (.B1(net313),
    .Y(_0319_),
    .A1(_2394_),
    .A2(_2635_));
 sg13g2_o21ai_1 _6551_ (.B1(_2633_),
    .Y(_2637_),
    .A1(_2630_),
    .A2(_2634_));
 sg13g2_xor2_1 _6552_ (.B(_2447_),
    .A(\vgademo.b_sin[2] ),
    .X(_2638_));
 sg13g2_and2_1 _6553_ (.A(_2637_),
    .B(_2638_),
    .X(_2639_));
 sg13g2_o21ai_1 _6554_ (.B1(net886),
    .Y(_2640_),
    .A1(_2637_),
    .A2(_2638_));
 sg13g2_a22oi_1 _6555_ (.Y(_2641_),
    .B1(net894),
    .B2(net349),
    .A2(net916),
    .A1(\vgademo.b_sin[2] ));
 sg13g2_o21ai_1 _6556_ (.B1(net350),
    .Y(_0320_),
    .A1(_2639_),
    .A2(_2640_));
 sg13g2_a21oi_1 _6557_ (.A1(\vgademo.b_sin[2] ),
    .A2(_2447_),
    .Y(_2642_),
    .B1(_2639_));
 sg13g2_nand2_1 _6558_ (.Y(_2643_),
    .A(\vgademo.b_sin[3] ),
    .B(_2454_));
 sg13g2_xnor2_1 _6559_ (.Y(_2644_),
    .A(\vgademo.b_sin[3] ),
    .B(_2454_));
 sg13g2_or2_1 _6560_ (.X(_2645_),
    .B(_2644_),
    .A(_2642_));
 sg13g2_a21oi_1 _6561_ (.A1(_2642_),
    .A2(_2644_),
    .Y(_2646_),
    .B1(_2394_));
 sg13g2_nand2_1 _6562_ (.Y(_2647_),
    .A(_2645_),
    .B(_2646_));
 sg13g2_a22oi_1 _6563_ (.Y(_2648_),
    .B1(net893),
    .B2(net433),
    .A2(net918),
    .A1(\vgademo.b_sin[3] ));
 sg13g2_nand2_1 _6564_ (.Y(_0321_),
    .A(_2647_),
    .B(net434));
 sg13g2_xnor2_1 _6565_ (.Y(_2649_),
    .A(\vgademo.b_sin[4] ),
    .B(_2458_));
 sg13g2_nand3_1 _6566_ (.B(_2645_),
    .C(_2649_),
    .A(_2643_),
    .Y(_2650_));
 sg13g2_a21oi_2 _6567_ (.B1(_2649_),
    .Y(_2651_),
    .A2(_2645_),
    .A1(_2643_));
 sg13g2_nand2_1 _6568_ (.Y(_2652_),
    .A(net886),
    .B(_2650_));
 sg13g2_a22oi_1 _6569_ (.Y(_2653_),
    .B1(net893),
    .B2(\vgademo.a_sin[7] ),
    .A2(net918),
    .A1(net443));
 sg13g2_o21ai_1 _6570_ (.B1(net444),
    .Y(_0322_),
    .A1(_2651_),
    .A2(_2652_));
 sg13g2_nand2_1 _6571_ (.Y(_2654_),
    .A(net284),
    .B(net917));
 sg13g2_xor2_1 _6572_ (.B(net837),
    .A(net284),
    .X(_2655_));
 sg13g2_a21oi_1 _6573_ (.A1(\vgademo.b_sin[4] ),
    .A2(net837),
    .Y(_2656_),
    .B1(_2651_));
 sg13g2_o21ai_1 _6574_ (.B1(net926),
    .Y(_2657_),
    .A1(_2655_),
    .A2(_2656_));
 sg13g2_a21oi_1 _6575_ (.A1(_2655_),
    .A2(_2656_),
    .Y(_2658_),
    .B1(_2657_));
 sg13g2_o21ai_1 _6576_ (.B1(net920),
    .Y(_2659_),
    .A1(\vgademo.a_sin[8] ),
    .A2(net926));
 sg13g2_o21ai_1 _6577_ (.B1(_2654_),
    .Y(_0323_),
    .A1(_2658_),
    .A2(_2659_));
 sg13g2_o21ai_1 _6578_ (.B1(net837),
    .Y(_2660_),
    .A1(\vgademo.b_sin[4] ),
    .A2(\vgademo.b_sin[5] ));
 sg13g2_nand2_1 _6579_ (.Y(_2661_),
    .A(_2651_),
    .B(_2655_));
 sg13g2_nand2_1 _6580_ (.Y(_2662_),
    .A(_2660_),
    .B(_2661_));
 sg13g2_xnor2_1 _6581_ (.Y(_2663_),
    .A(\vgademo.b_sin[6] ),
    .B(net836));
 sg13g2_inv_1 _6582_ (.Y(_2664_),
    .A(_2663_));
 sg13g2_a21oi_1 _6583_ (.A1(_2660_),
    .A2(_2661_),
    .Y(_2665_),
    .B1(_2663_));
 sg13g2_o21ai_1 _6584_ (.B1(net887),
    .Y(_2666_),
    .A1(_2662_),
    .A2(_2664_));
 sg13g2_a22oi_1 _6585_ (.Y(_2667_),
    .B1(net892),
    .B2(\vgademo.a_sin[9] ),
    .A2(net917),
    .A1(net455));
 sg13g2_o21ai_1 _6586_ (.B1(net456),
    .Y(_0324_),
    .A1(_2665_),
    .A2(_2666_));
 sg13g2_nand2_1 _6587_ (.Y(_2668_),
    .A(net304),
    .B(net917));
 sg13g2_a21oi_1 _6588_ (.A1(\vgademo.b_sin[6] ),
    .A2(net836),
    .Y(_2669_),
    .B1(_2665_));
 sg13g2_xnor2_1 _6589_ (.Y(_2670_),
    .A(_3135_),
    .B(net836));
 sg13g2_o21ai_1 _6590_ (.B1(net926),
    .Y(_2671_),
    .A1(_2669_),
    .A2(_2670_));
 sg13g2_a21oi_1 _6591_ (.A1(_2669_),
    .A2(_2670_),
    .Y(_2672_),
    .B1(_2671_));
 sg13g2_o21ai_1 _6592_ (.B1(net919),
    .Y(_2673_),
    .A1(\vgademo.a_sin[10] ),
    .A2(net926));
 sg13g2_o21ai_1 _6593_ (.B1(_2668_),
    .Y(_0325_),
    .A1(_2672_),
    .A2(_2673_));
 sg13g2_nor2_1 _6594_ (.A(_2661_),
    .B(_2663_),
    .Y(_2674_));
 sg13g2_o21ai_1 _6595_ (.B1(_2674_),
    .Y(_2675_),
    .A1(\vgademo.b_sin[7] ),
    .A2(net836));
 sg13g2_o21ai_1 _6596_ (.B1(net836),
    .Y(_2676_),
    .A1(\vgademo.b_sin[7] ),
    .A2(\vgademo.b_sin[6] ));
 sg13g2_nand3_1 _6597_ (.B(_2675_),
    .C(_2676_),
    .A(_2660_),
    .Y(_2677_));
 sg13g2_xnor2_1 _6598_ (.Y(_2678_),
    .A(\vgademo.b_sin[8] ),
    .B(net836));
 sg13g2_inv_1 _6599_ (.Y(_2679_),
    .A(_2678_));
 sg13g2_and2_1 _6600_ (.A(_2677_),
    .B(_2679_),
    .X(_2680_));
 sg13g2_o21ai_1 _6601_ (.B1(net887),
    .Y(_2681_),
    .A1(_2677_),
    .A2(_2679_));
 sg13g2_a22oi_1 _6602_ (.Y(_2682_),
    .B1(net892),
    .B2(\vgademo.a_sin[11] ),
    .A2(net917),
    .A1(net474));
 sg13g2_o21ai_1 _6603_ (.B1(net475),
    .Y(_0326_),
    .A1(_2680_),
    .A2(_2681_));
 sg13g2_a21oi_1 _6604_ (.A1(\vgademo.b_sin[8] ),
    .A2(net836),
    .Y(_2683_),
    .B1(_2680_));
 sg13g2_nor2_1 _6605_ (.A(\vgademo.b_sin[9] ),
    .B(net837),
    .Y(_2684_));
 sg13g2_xnor2_1 _6606_ (.Y(_2685_),
    .A(\vgademo.b_sin[9] ),
    .B(net837));
 sg13g2_nor2_1 _6607_ (.A(_2683_),
    .B(_2684_),
    .Y(_2686_));
 sg13g2_xnor2_1 _6608_ (.Y(_2687_),
    .A(_2683_),
    .B(_2685_));
 sg13g2_a22oi_1 _6609_ (.Y(_2688_),
    .B1(net892),
    .B2(\vgademo.a_sin[12] ),
    .A2(net917),
    .A1(net537));
 sg13g2_o21ai_1 _6610_ (.B1(net538),
    .Y(_0327_),
    .A1(_2394_),
    .A2(_2687_));
 sg13g2_xnor2_1 _6611_ (.Y(_2689_),
    .A(\vgademo.b_sin[10] ),
    .B(net836));
 sg13g2_a21oi_1 _6612_ (.A1(\vgademo.b_sin[9] ),
    .A2(net837),
    .Y(_2690_),
    .B1(_2686_));
 sg13g2_nor2_1 _6613_ (.A(_2689_),
    .B(_2690_),
    .Y(_2691_));
 sg13g2_a21o_1 _6614_ (.A2(_2690_),
    .A1(_2689_),
    .B1(_2394_),
    .X(_2692_));
 sg13g2_a22oi_1 _6615_ (.Y(_2693_),
    .B1(net893),
    .B2(\vgademo.a_sin[13] ),
    .A2(net917),
    .A1(net462));
 sg13g2_o21ai_1 _6616_ (.B1(net463),
    .Y(_0328_),
    .A1(_2691_),
    .A2(_2692_));
 sg13g2_nand2_1 _6617_ (.Y(_2694_),
    .A(net952),
    .B(net916));
 sg13g2_a21o_1 _6618_ (.A2(net837),
    .A1(\vgademo.b_sin[10] ),
    .B1(_2691_),
    .X(_2695_));
 sg13g2_xor2_1 _6619_ (.B(_2456_),
    .A(\vgademo.b_cos[11] ),
    .X(_2696_));
 sg13g2_o21ai_1 _6620_ (.B1(net927),
    .Y(_2697_),
    .A1(_2695_),
    .A2(_2696_));
 sg13g2_a21oi_1 _6621_ (.A1(_2695_),
    .A2(_2696_),
    .Y(_2698_),
    .B1(_2697_));
 sg13g2_o21ai_1 _6622_ (.B1(net919),
    .Y(_2699_),
    .A1(net961),
    .A2(net927));
 sg13g2_o21ai_1 _6623_ (.B1(_2694_),
    .Y(_0329_),
    .A1(_2698_),
    .A2(_2699_));
 sg13g2_nand2_1 _6624_ (.Y(_2700_),
    .A(net922),
    .B(_2235_));
 sg13g2_nand2_2 _6625_ (.Y(_2701_),
    .A(net1079),
    .B(_2700_));
 sg13g2_inv_2 _6626_ (.Y(_2702_),
    .A(net880));
 sg13g2_nand2_1 _6627_ (.Y(_2703_),
    .A(net258),
    .B(\vgademo.plane_du[0] ));
 sg13g2_nand2_1 _6628_ (.Y(_2704_),
    .A(net295),
    .B(net337));
 sg13g2_xor2_1 _6629_ (.B(\vgademo.plane_du[1] ),
    .A(\vgademo.plane_u[1] ),
    .X(_2705_));
 sg13g2_nand2b_1 _6630_ (.Y(_2706_),
    .B(_2705_),
    .A_N(_2703_));
 sg13g2_xor2_1 _6631_ (.B(_2705_),
    .A(_2703_),
    .X(_2707_));
 sg13g2_nor2_1 _6632_ (.A(net930),
    .B(_2707_),
    .Y(_2708_));
 sg13g2_a21oi_1 _6633_ (.A1(\vgademo.plane_dx[0] ),
    .A2(net930),
    .Y(_2709_),
    .B1(_2708_));
 sg13g2_nand2_1 _6634_ (.Y(_2710_),
    .A(net295),
    .B(net877));
 sg13g2_o21ai_1 _6635_ (.B1(_2710_),
    .Y(_0330_),
    .A1(net877),
    .A2(_2709_));
 sg13g2_nand2_1 _6636_ (.Y(_2711_),
    .A(net376),
    .B(\vgademo.plane_du[2] ));
 sg13g2_xnor2_1 _6637_ (.Y(_2712_),
    .A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ));
 sg13g2_nand3_1 _6638_ (.B(_2706_),
    .C(_2712_),
    .A(_2704_),
    .Y(_2713_));
 sg13g2_a21o_1 _6639_ (.A2(_2706_),
    .A1(_2704_),
    .B1(_2712_),
    .X(_2714_));
 sg13g2_nand3_1 _6640_ (.B(_2713_),
    .C(_2714_),
    .A(net925),
    .Y(_2715_));
 sg13g2_nor2b_1 _6641_ (.A(net1040),
    .B_N(net955),
    .Y(_2716_));
 sg13g2_xnor2_1 _6642_ (.Y(_2717_),
    .A(net1040),
    .B(net955));
 sg13g2_a21oi_1 _6643_ (.A1(net929),
    .A2(_2717_),
    .Y(_2718_),
    .B1(net878));
 sg13g2_a22oi_1 _6644_ (.Y(_0331_),
    .B1(_2715_),
    .B2(_2718_),
    .A2(net877),
    .A1(_3156_));
 sg13g2_nand2_1 _6645_ (.Y(_2719_),
    .A(\vgademo.plane_u[3] ),
    .B(\vgademo.plane_du[3] ));
 sg13g2_xnor2_1 _6646_ (.Y(_2720_),
    .A(\vgademo.plane_u[3] ),
    .B(\vgademo.plane_du[3] ));
 sg13g2_nand3_1 _6647_ (.B(_2714_),
    .C(_2720_),
    .A(_2711_),
    .Y(_2721_));
 sg13g2_a21o_1 _6648_ (.A2(_2714_),
    .A1(_2711_),
    .B1(_2720_),
    .X(_2722_));
 sg13g2_nand3_1 _6649_ (.B(_2721_),
    .C(_2722_),
    .A(net925),
    .Y(_2723_));
 sg13g2_and2_1 _6650_ (.A(_3084_),
    .B(_2716_),
    .X(_2724_));
 sg13g2_xnor2_1 _6651_ (.Y(_2725_),
    .A(\vgademo.plane_dx[2] ),
    .B(_2716_));
 sg13g2_a21oi_1 _6652_ (.A1(net929),
    .A2(_2725_),
    .Y(_2726_),
    .B1(net878));
 sg13g2_a22oi_1 _6653_ (.Y(_0332_),
    .B1(_2723_),
    .B2(_2726_),
    .A2(net878),
    .A1(_3157_));
 sg13g2_xnor2_1 _6654_ (.Y(_2727_),
    .A(\vgademo.plane_u[4] ),
    .B(\vgademo.plane_du[4] ));
 sg13g2_a21oi_1 _6655_ (.A1(_2719_),
    .A2(_2722_),
    .Y(_2728_),
    .B1(_2727_));
 sg13g2_and3_1 _6656_ (.X(_2729_),
    .A(_2719_),
    .B(_2722_),
    .C(_2727_));
 sg13g2_o21ai_1 _6657_ (.B1(net925),
    .Y(_2730_),
    .A1(_2728_),
    .A2(_2729_));
 sg13g2_nor2_1 _6658_ (.A(\vgademo.plane_dx[3] ),
    .B(_2724_),
    .Y(_2731_));
 sg13g2_xnor2_1 _6659_ (.Y(_2732_),
    .A(\vgademo.plane_dx[3] ),
    .B(_2724_));
 sg13g2_o21ai_1 _6660_ (.B1(_2730_),
    .Y(_2733_),
    .A1(net927),
    .A2(_2732_));
 sg13g2_nand2_1 _6661_ (.Y(_2734_),
    .A(net272),
    .B(net878));
 sg13g2_o21ai_1 _6662_ (.B1(_2734_),
    .Y(_0333_),
    .A1(net880),
    .A2(_2733_));
 sg13g2_a21o_1 _6663_ (.A2(\vgademo.plane_du[4] ),
    .A1(\vgademo.plane_u[4] ),
    .B1(_2728_),
    .X(_2735_));
 sg13g2_nand2_1 _6664_ (.Y(_2736_),
    .A(net290),
    .B(\vgademo.plane_du[5] ));
 sg13g2_or2_1 _6665_ (.X(_2737_),
    .B(\vgademo.plane_du[5] ),
    .A(\vgademo.plane_u[5] ));
 sg13g2_nand2_1 _6666_ (.Y(_2738_),
    .A(_2736_),
    .B(_2737_));
 sg13g2_xnor2_1 _6667_ (.Y(_2739_),
    .A(_2735_),
    .B(_2738_));
 sg13g2_nand2b_1 _6668_ (.Y(_2740_),
    .B(\vgademo.plane_dx[0] ),
    .A_N(_0024_));
 sg13g2_xnor2_1 _6669_ (.Y(_2741_),
    .A(\vgademo.plane_dx[0] ),
    .B(net1039));
 sg13g2_nand2_1 _6670_ (.Y(_2742_),
    .A(_0023_),
    .B(_2741_));
 sg13g2_xnor2_1 _6671_ (.Y(_2743_),
    .A(_0023_),
    .B(_2741_));
 sg13g2_xnor2_1 _6672_ (.Y(_2744_),
    .A(_2731_),
    .B(_2743_));
 sg13g2_a21oi_1 _6673_ (.A1(net929),
    .A2(_2744_),
    .Y(_2745_),
    .B1(net878));
 sg13g2_o21ai_1 _6674_ (.B1(_2745_),
    .Y(_2746_),
    .A1(net929),
    .A2(_2739_));
 sg13g2_o21ai_1 _6675_ (.B1(_2746_),
    .Y(_0334_),
    .A1(_3159_),
    .A2(_2702_));
 sg13g2_nand2_1 _6676_ (.Y(_2747_),
    .A(net357),
    .B(\vgademo.plane_du[6] ));
 sg13g2_xnor2_1 _6677_ (.Y(_2748_),
    .A(\vgademo.plane_u[6] ),
    .B(\vgademo.plane_du[6] ));
 sg13g2_nand2_1 _6678_ (.Y(_2749_),
    .A(_2735_),
    .B(_2737_));
 sg13g2_nand3_1 _6679_ (.B(_2748_),
    .C(_2749_),
    .A(_2736_),
    .Y(_2750_));
 sg13g2_a21o_1 _6680_ (.A2(_2749_),
    .A1(_2736_),
    .B1(_2748_),
    .X(_2751_));
 sg13g2_nand3_1 _6681_ (.B(_2750_),
    .C(_2751_),
    .A(net925),
    .Y(_2752_));
 sg13g2_o21ai_1 _6682_ (.B1(_2742_),
    .Y(_2753_),
    .A1(_2731_),
    .A2(_2743_));
 sg13g2_nand2_1 _6683_ (.Y(_2754_),
    .A(net1038),
    .B(\vgademo.plane_dx[1] ));
 sg13g2_nor2_1 _6684_ (.A(net1038),
    .B(net1040),
    .Y(_2755_));
 sg13g2_xor2_1 _6685_ (.B(net1040),
    .A(net1038),
    .X(_2756_));
 sg13g2_xnor2_1 _6686_ (.Y(_2757_),
    .A(_2740_),
    .B(_2756_));
 sg13g2_xnor2_1 _6687_ (.Y(_2758_),
    .A(net955),
    .B(_2757_));
 sg13g2_nor2b_1 _6688_ (.A(_2741_),
    .B_N(_2758_),
    .Y(_2759_));
 sg13g2_xnor2_1 _6689_ (.Y(_2760_),
    .A(_2741_),
    .B(_2758_));
 sg13g2_and2_1 _6690_ (.A(_2753_),
    .B(_2760_),
    .X(_2761_));
 sg13g2_o21ai_1 _6691_ (.B1(net929),
    .Y(_2762_),
    .A1(_2753_),
    .A2(_2760_));
 sg13g2_nor2_1 _6692_ (.A(_2761_),
    .B(_2762_),
    .Y(_2763_));
 sg13g2_nor2_1 _6693_ (.A(net877),
    .B(_2763_),
    .Y(_2764_));
 sg13g2_a22oi_1 _6694_ (.Y(_0335_),
    .B1(_2752_),
    .B2(_2764_),
    .A2(net877),
    .A1(_3161_));
 sg13g2_nand2_1 _6695_ (.Y(_2765_),
    .A(\vgademo.plane_u[7] ),
    .B(\vgademo.plane_du[7] ));
 sg13g2_xnor2_1 _6696_ (.Y(_2766_),
    .A(\vgademo.plane_u[7] ),
    .B(\vgademo.plane_du[7] ));
 sg13g2_nand3_1 _6697_ (.B(_2751_),
    .C(_2766_),
    .A(_2747_),
    .Y(_2767_));
 sg13g2_a21o_1 _6698_ (.A2(_2751_),
    .A1(_2747_),
    .B1(_2766_),
    .X(_2768_));
 sg13g2_nand3_1 _6699_ (.B(_2767_),
    .C(_2768_),
    .A(net924),
    .Y(_2769_));
 sg13g2_nor2_1 _6700_ (.A(_2759_),
    .B(_2761_),
    .Y(_2770_));
 sg13g2_nand2_1 _6701_ (.Y(_2771_),
    .A(\vgademo.plane_dx[0] ),
    .B(_2757_));
 sg13g2_o21ai_1 _6702_ (.B1(_2754_),
    .Y(_2772_),
    .A1(_2740_),
    .A2(_2755_));
 sg13g2_inv_1 _6703_ (.Y(_2773_),
    .A(_2772_));
 sg13g2_nand2_1 _6704_ (.Y(_2774_),
    .A(\vgademo.plane_dx_div.q[5] ),
    .B(\vgademo.plane_dx[2] ));
 sg13g2_xnor2_1 _6705_ (.Y(_2775_),
    .A(\vgademo.plane_dx_div.q[5] ),
    .B(\vgademo.plane_dx[2] ));
 sg13g2_xnor2_1 _6706_ (.Y(_2776_),
    .A(_2772_),
    .B(_2775_));
 sg13g2_xnor2_1 _6707_ (.Y(_2777_),
    .A(_0025_),
    .B(_2776_));
 sg13g2_nand2b_1 _6708_ (.Y(_2778_),
    .B(_2771_),
    .A_N(_2777_));
 sg13g2_xor2_1 _6709_ (.B(_2777_),
    .A(_2771_),
    .X(_2779_));
 sg13g2_xor2_1 _6710_ (.B(_2779_),
    .A(_2758_),
    .X(_2780_));
 sg13g2_nor2b_1 _6711_ (.A(_2780_),
    .B_N(_2770_),
    .Y(_2781_));
 sg13g2_nor2b_1 _6712_ (.A(_2770_),
    .B_N(_2780_),
    .Y(_2782_));
 sg13g2_inv_1 _6713_ (.Y(_2783_),
    .A(_2782_));
 sg13g2_nor3_1 _6714_ (.A(net924),
    .B(_2781_),
    .C(_2782_),
    .Y(_2784_));
 sg13g2_nor2_1 _6715_ (.A(net877),
    .B(_2784_),
    .Y(_2785_));
 sg13g2_a22oi_1 _6716_ (.Y(_0336_),
    .B1(_2769_),
    .B2(_2785_),
    .A2(net877),
    .A1(_3162_));
 sg13g2_xnor2_1 _6717_ (.Y(_2786_),
    .A(\vgademo.plane_u[8] ),
    .B(\vgademo.plane_du[8] ));
 sg13g2_a21oi_1 _6718_ (.A1(_2765_),
    .A2(_2768_),
    .Y(_2787_),
    .B1(_2786_));
 sg13g2_nand3_1 _6719_ (.B(_2768_),
    .C(_2786_),
    .A(_2765_),
    .Y(_2788_));
 sg13g2_nor2b_1 _6720_ (.A(_2787_),
    .B_N(_2788_),
    .Y(_2789_));
 sg13g2_o21ai_1 _6721_ (.B1(_2783_),
    .Y(_2790_),
    .A1(_2758_),
    .A2(_2779_));
 sg13g2_nand2_1 _6722_ (.Y(_2791_),
    .A(net1040),
    .B(_2776_));
 sg13g2_o21ai_1 _6723_ (.B1(_2774_),
    .Y(_2792_),
    .A1(_2773_),
    .A2(_2775_));
 sg13g2_xor2_1 _6724_ (.B(\vgademo.plane_dx[3] ),
    .A(net1035),
    .X(_2793_));
 sg13g2_xnor2_1 _6725_ (.Y(_2794_),
    .A(_2792_),
    .B(_2793_));
 sg13g2_xor2_1 _6726_ (.B(_2794_),
    .A(_0026_),
    .X(_2795_));
 sg13g2_nand2b_1 _6727_ (.Y(_2796_),
    .B(_2791_),
    .A_N(_2795_));
 sg13g2_xor2_1 _6728_ (.B(_2795_),
    .A(_2791_),
    .X(_2797_));
 sg13g2_xor2_1 _6729_ (.B(_2797_),
    .A(_2778_),
    .X(_2798_));
 sg13g2_nor2_1 _6730_ (.A(_2790_),
    .B(_2798_),
    .Y(_2799_));
 sg13g2_nand2_1 _6731_ (.Y(_2800_),
    .A(_2790_),
    .B(_2798_));
 sg13g2_nor2_1 _6732_ (.A(net924),
    .B(_2799_),
    .Y(_2801_));
 sg13g2_a221oi_1 _6733_ (.B2(_2801_),
    .C1(net879),
    .B1(_2800_),
    .A1(net924),
    .Y(_2802_),
    .A2(_2789_));
 sg13g2_a21oi_1 _6734_ (.A1(_3164_),
    .A2(net879),
    .Y(_0337_),
    .B1(_2802_));
 sg13g2_a21o_1 _6735_ (.A2(\vgademo.plane_du[8] ),
    .A1(\vgademo.plane_u[8] ),
    .B1(_2787_),
    .X(_2803_));
 sg13g2_or2_1 _6736_ (.X(_2804_),
    .B(\vgademo.plane_du[9] ),
    .A(\vgademo.plane_u[9] ));
 sg13g2_xnor2_1 _6737_ (.Y(_2805_),
    .A(\vgademo.plane_u[9] ),
    .B(net950));
 sg13g2_xnor2_1 _6738_ (.Y(_2806_),
    .A(_2803_),
    .B(_2805_));
 sg13g2_o21ai_1 _6739_ (.B1(_2800_),
    .Y(_2807_),
    .A1(_2778_),
    .A2(_2797_));
 sg13g2_nor2_1 _6740_ (.A(_3084_),
    .B(_2794_),
    .Y(_2808_));
 sg13g2_a22oi_1 _6741_ (.Y(_2809_),
    .B1(_2792_),
    .B2(_2793_),
    .A2(_3160_),
    .A1(net1035));
 sg13g2_xnor2_1 _6742_ (.Y(_2810_),
    .A(\vgademo.plane_dx_div.q[7] ),
    .B(net1039));
 sg13g2_nand2b_1 _6743_ (.Y(_2811_),
    .B(_2810_),
    .A_N(_2809_));
 sg13g2_xnor2_1 _6744_ (.Y(_2812_),
    .A(_2809_),
    .B(_2810_));
 sg13g2_xnor2_1 _6745_ (.Y(_2813_),
    .A(\vgademo.plane_dx[3] ),
    .B(net955));
 sg13g2_nor2b_1 _6746_ (.A(_2812_),
    .B_N(_2813_),
    .Y(_2814_));
 sg13g2_xnor2_1 _6747_ (.Y(_2815_),
    .A(_2812_),
    .B(_2813_));
 sg13g2_nand2b_1 _6748_ (.Y(_2816_),
    .B(_2815_),
    .A_N(_2808_));
 sg13g2_xor2_1 _6749_ (.B(_2815_),
    .A(_2808_),
    .X(_2817_));
 sg13g2_nor2_1 _6750_ (.A(_2796_),
    .B(_2817_),
    .Y(_2818_));
 sg13g2_xor2_1 _6751_ (.B(_2817_),
    .A(_2796_),
    .X(_2819_));
 sg13g2_nor2_1 _6752_ (.A(_2807_),
    .B(_2819_),
    .Y(_2820_));
 sg13g2_nand2_1 _6753_ (.Y(_2821_),
    .A(_2807_),
    .B(_2819_));
 sg13g2_nor2_1 _6754_ (.A(net924),
    .B(_2820_),
    .Y(_2822_));
 sg13g2_a221oi_1 _6755_ (.B2(_2822_),
    .C1(net879),
    .B1(_2821_),
    .A1(net924),
    .Y(_2823_),
    .A2(_2806_));
 sg13g2_a21oi_1 _6756_ (.A1(_3165_),
    .A2(net879),
    .Y(_0338_),
    .B1(_2823_));
 sg13g2_nand2_1 _6757_ (.Y(_2824_),
    .A(\vgademo.plane_u[10] ),
    .B(\vgademo.plane_du[10] ));
 sg13g2_xor2_1 _6758_ (.B(\vgademo.plane_du[10] ),
    .A(\vgademo.plane_u[10] ),
    .X(_2825_));
 sg13g2_a21o_1 _6759_ (.A2(net950),
    .A1(\vgademo.plane_u[9] ),
    .B1(_2803_),
    .X(_2826_));
 sg13g2_a21oi_1 _6760_ (.A1(_2804_),
    .A2(_2826_),
    .Y(_2827_),
    .B1(_2825_));
 sg13g2_nand3_1 _6761_ (.B(_2825_),
    .C(_2826_),
    .A(_2804_),
    .Y(_2828_));
 sg13g2_nor2_1 _6762_ (.A(net929),
    .B(_2827_),
    .Y(_2829_));
 sg13g2_a21oi_1 _6763_ (.A1(_2807_),
    .A2(_2819_),
    .Y(_2830_),
    .B1(_2818_));
 sg13g2_a21oi_1 _6764_ (.A1(_3083_),
    .A2(net955),
    .Y(_2831_),
    .B1(_2814_));
 sg13g2_xor2_1 _6765_ (.B(net1039),
    .A(net1040),
    .X(_2832_));
 sg13g2_inv_1 _6766_ (.Y(_2833_),
    .A(_2832_));
 sg13g2_o21ai_1 _6767_ (.B1(_2811_),
    .Y(_2834_),
    .A1(_3082_),
    .A2(net1039));
 sg13g2_nand2_1 _6768_ (.Y(_2835_),
    .A(net1032),
    .B(net1038));
 sg13g2_xor2_1 _6769_ (.B(net1037),
    .A(net1032),
    .X(_2836_));
 sg13g2_xnor2_1 _6770_ (.Y(_2837_),
    .A(_2834_),
    .B(_2836_));
 sg13g2_xnor2_1 _6771_ (.Y(_2838_),
    .A(_2832_),
    .B(_2837_));
 sg13g2_nand2b_1 _6772_ (.Y(_2839_),
    .B(_2838_),
    .A_N(_2831_));
 sg13g2_xor2_1 _6773_ (.B(_2838_),
    .A(_2831_),
    .X(_2840_));
 sg13g2_nor2_1 _6774_ (.A(_2816_),
    .B(_2840_),
    .Y(_2841_));
 sg13g2_xnor2_1 _6775_ (.Y(_2842_),
    .A(_2816_),
    .B(_2840_));
 sg13g2_or2_1 _6776_ (.X(_2843_),
    .B(_2842_),
    .A(_2830_));
 sg13g2_a21oi_1 _6777_ (.A1(_2830_),
    .A2(_2842_),
    .Y(_2844_),
    .B1(net924));
 sg13g2_a221oi_1 _6778_ (.B2(_2844_),
    .C1(net879),
    .B1(_2843_),
    .A1(_2828_),
    .Y(_2845_),
    .A2(_2829_));
 sg13g2_a21oi_1 _6779_ (.A1(_3166_),
    .A2(net879),
    .Y(_0339_),
    .B1(_2845_));
 sg13g2_a21oi_2 _6780_ (.B1(_0027_),
    .Y(_2846_),
    .A2(_2828_),
    .A1(_2824_));
 sg13g2_nand3_1 _6781_ (.B(_2824_),
    .C(_2828_),
    .A(_0027_),
    .Y(_2847_));
 sg13g2_nor2_1 _6782_ (.A(net929),
    .B(_2846_),
    .Y(_2848_));
 sg13g2_nor2b_1 _6783_ (.A(_2841_),
    .B_N(_2843_),
    .Y(_2849_));
 sg13g2_a22oi_1 _6784_ (.Y(_2850_),
    .B1(_2833_),
    .B2(_2837_),
    .A2(_0025_),
    .A1(net1039));
 sg13g2_xnor2_1 _6785_ (.Y(_2851_),
    .A(\vgademo.plane_dx_div.q[9] ),
    .B(net1036));
 sg13g2_o21ai_1 _6786_ (.B1(_2834_),
    .Y(_2852_),
    .A1(net1032),
    .A2(net1038));
 sg13g2_nand2_1 _6787_ (.Y(_2853_),
    .A(_2835_),
    .B(_2852_));
 sg13g2_a21oi_1 _6788_ (.A1(_2835_),
    .A2(_2852_),
    .Y(_2854_),
    .B1(_2851_));
 sg13g2_xor2_1 _6789_ (.B(_2853_),
    .A(_2851_),
    .X(_2855_));
 sg13g2_xor2_1 _6790_ (.B(\vgademo.plane_dx[2] ),
    .A(net1037),
    .X(_2856_));
 sg13g2_xnor2_1 _6791_ (.Y(_2857_),
    .A(_2855_),
    .B(_2856_));
 sg13g2_nor2_1 _6792_ (.A(_2850_),
    .B(_2857_),
    .Y(_2858_));
 sg13g2_xnor2_1 _6793_ (.Y(_2859_),
    .A(_2850_),
    .B(_2857_));
 sg13g2_xnor2_1 _6794_ (.Y(_2860_),
    .A(_2839_),
    .B(_2859_));
 sg13g2_nor2_1 _6795_ (.A(_2849_),
    .B(_2860_),
    .Y(_2861_));
 sg13g2_inv_1 _6796_ (.Y(_2862_),
    .A(_2861_));
 sg13g2_a21oi_1 _6797_ (.A1(_2849_),
    .A2(_2860_),
    .Y(_2863_),
    .B1(net924));
 sg13g2_a221oi_1 _6798_ (.B2(_2863_),
    .C1(net879),
    .B1(_2862_),
    .A1(_2847_),
    .Y(_2864_),
    .A2(_2848_));
 sg13g2_a21oi_1 _6799_ (.A1(_3167_),
    .A2(net879),
    .Y(_0340_),
    .B1(_2864_));
 sg13g2_xnor2_1 _6800_ (.Y(_2865_),
    .A(_0028_),
    .B(_2846_));
 sg13g2_o21ai_1 _6801_ (.B1(_2862_),
    .Y(_2866_),
    .A1(_2839_),
    .A2(_2859_));
 sg13g2_nor2b_1 _6802_ (.A(net1037),
    .B_N(_0026_),
    .Y(_2867_));
 sg13g2_a21o_1 _6803_ (.A2(_2856_),
    .A1(_2855_),
    .B1(_2867_),
    .X(_2868_));
 sg13g2_a21oi_1 _6804_ (.A1(\vgademo.plane_dx_div.q[9] ),
    .A2(net1036),
    .Y(_2869_),
    .B1(_2854_));
 sg13g2_nor2b_1 _6805_ (.A(_2869_),
    .B_N(net1035),
    .Y(_2870_));
 sg13g2_xnor2_1 _6806_ (.Y(_2871_),
    .A(net1034),
    .B(_2869_));
 sg13g2_xor2_1 _6807_ (.B(\vgademo.plane_dx[3] ),
    .A(net1036),
    .X(_2872_));
 sg13g2_nand2b_1 _6808_ (.Y(_2873_),
    .B(_2872_),
    .A_N(_2871_));
 sg13g2_xnor2_1 _6809_ (.Y(_2874_),
    .A(_2871_),
    .B(_2872_));
 sg13g2_nand2_1 _6810_ (.Y(_2875_),
    .A(_2868_),
    .B(_2874_));
 sg13g2_xor2_1 _6811_ (.B(_2874_),
    .A(_2868_),
    .X(_2876_));
 sg13g2_xnor2_1 _6812_ (.Y(_2877_),
    .A(_2858_),
    .B(_2876_));
 sg13g2_nand2b_1 _6813_ (.Y(_2878_),
    .B(_2877_),
    .A_N(_2866_));
 sg13g2_nor2b_1 _6814_ (.A(_2877_),
    .B_N(_2866_),
    .Y(_2879_));
 sg13g2_nor2_1 _6815_ (.A(net926),
    .B(_2879_),
    .Y(_2880_));
 sg13g2_a221oi_1 _6816_ (.B2(_2880_),
    .C1(net880),
    .B1(_2878_),
    .A1(net926),
    .Y(_2881_),
    .A2(_2865_));
 sg13g2_a21oi_1 _6817_ (.A1(_3168_),
    .A2(net880),
    .Y(_0341_),
    .B1(_2881_));
 sg13g2_a21oi_1 _6818_ (.A1(_2858_),
    .A2(_2876_),
    .Y(_2882_),
    .B1(_2879_));
 sg13g2_o21ai_1 _6819_ (.B1(_2873_),
    .Y(_2883_),
    .A1(net1036),
    .A2(_3160_));
 sg13g2_xnor2_1 _6820_ (.Y(_2884_),
    .A(net1033),
    .B(_2870_));
 sg13g2_nor2b_1 _6821_ (.A(net1035),
    .B_N(net1039),
    .Y(_2885_));
 sg13g2_xnor2_1 _6822_ (.Y(_2886_),
    .A(net1035),
    .B(net1039));
 sg13g2_xnor2_1 _6823_ (.Y(_2887_),
    .A(_2884_),
    .B(_2886_));
 sg13g2_nor2b_1 _6824_ (.A(_2887_),
    .B_N(_2883_),
    .Y(_2888_));
 sg13g2_xor2_1 _6825_ (.B(_2887_),
    .A(_2883_),
    .X(_2889_));
 sg13g2_nor2_1 _6826_ (.A(_2875_),
    .B(_2889_),
    .Y(_2890_));
 sg13g2_xor2_1 _6827_ (.B(_2889_),
    .A(_2875_),
    .X(_2891_));
 sg13g2_nor2b_1 _6828_ (.A(_2882_),
    .B_N(_2891_),
    .Y(_2892_));
 sg13g2_nor2b_1 _6829_ (.A(_2891_),
    .B_N(_2882_),
    .Y(_2893_));
 sg13g2_nor3_1 _6830_ (.A(net926),
    .B(_2892_),
    .C(_2893_),
    .Y(_2894_));
 sg13g2_a21oi_1 _6831_ (.A1(\vgademo.plane_u[12] ),
    .A2(_2846_),
    .Y(_2895_),
    .B1(net406));
 sg13g2_and3_1 _6832_ (.X(_2896_),
    .A(\vgademo.plane_u[12] ),
    .B(\vgademo.plane_u[13] ),
    .C(_2846_));
 sg13g2_nor3_1 _6833_ (.A(net931),
    .B(_2895_),
    .C(_2896_),
    .Y(_2897_));
 sg13g2_nor3_1 _6834_ (.A(net876),
    .B(_2894_),
    .C(_2897_),
    .Y(_2898_));
 sg13g2_a21oi_1 _6835_ (.A1(_3170_),
    .A2(net876),
    .Y(_0342_),
    .B1(_2898_));
 sg13g2_a21oi_2 _6836_ (.B1(_2885_),
    .Y(_2899_),
    .A2(_2886_),
    .A1(_2884_));
 sg13g2_nand3_1 _6837_ (.B(net1033),
    .C(_2870_),
    .A(net1031),
    .Y(_2900_));
 sg13g2_a21o_1 _6838_ (.A2(_2870_),
    .A1(net1033),
    .B1(net1031),
    .X(_2901_));
 sg13g2_nand2_1 _6839_ (.Y(_2902_),
    .A(_2900_),
    .B(_2901_));
 sg13g2_xor2_1 _6840_ (.B(net1037),
    .A(net1033),
    .X(_2903_));
 sg13g2_nand2_1 _6841_ (.Y(_2904_),
    .A(_2902_),
    .B(_2903_));
 sg13g2_xnor2_1 _6842_ (.Y(_2905_),
    .A(_2902_),
    .B(_2903_));
 sg13g2_nor2_1 _6843_ (.A(_2899_),
    .B(_2905_),
    .Y(_2906_));
 sg13g2_xor2_1 _6844_ (.B(_2905_),
    .A(_2899_),
    .X(_2907_));
 sg13g2_nand2_1 _6845_ (.Y(_2908_),
    .A(_2888_),
    .B(_2907_));
 sg13g2_xnor2_1 _6846_ (.Y(_2909_),
    .A(_2888_),
    .B(_2907_));
 sg13g2_inv_1 _6847_ (.Y(_2910_),
    .A(_2909_));
 sg13g2_o21ai_1 _6848_ (.B1(_2910_),
    .Y(_2911_),
    .A1(_2890_),
    .A2(_2892_));
 sg13g2_or3_1 _6849_ (.A(_2890_),
    .B(_2892_),
    .C(_2910_),
    .X(_2912_));
 sg13g2_nand2_1 _6850_ (.Y(_2913_),
    .A(_2911_),
    .B(_2912_));
 sg13g2_xnor2_1 _6851_ (.Y(_2914_),
    .A(net458),
    .B(_2896_));
 sg13g2_nand2_1 _6852_ (.Y(_2915_),
    .A(net927),
    .B(_2914_));
 sg13g2_a21oi_1 _6853_ (.A1(net930),
    .A2(_2913_),
    .Y(_2916_),
    .B1(net880));
 sg13g2_a22oi_1 _6854_ (.Y(_2917_),
    .B1(_2915_),
    .B2(_2916_),
    .A2(net875),
    .A1(net458));
 sg13g2_inv_1 _6855_ (.Y(_0343_),
    .A(_2917_));
 sg13g2_o21ai_1 _6856_ (.B1(_2904_),
    .Y(_2918_),
    .A1(net1033),
    .A2(net1037));
 sg13g2_xor2_1 _6857_ (.B(net1036),
    .A(net1031),
    .X(_2919_));
 sg13g2_xor2_1 _6858_ (.B(_2900_),
    .A(net1030),
    .X(_2920_));
 sg13g2_nand2_1 _6859_ (.Y(_2921_),
    .A(_2919_),
    .B(_2920_));
 sg13g2_xor2_1 _6860_ (.B(_2920_),
    .A(_2919_),
    .X(_2922_));
 sg13g2_nand2_1 _6861_ (.Y(_2923_),
    .A(_2918_),
    .B(_2922_));
 sg13g2_xnor2_1 _6862_ (.Y(_2924_),
    .A(_2918_),
    .B(_2922_));
 sg13g2_or3_1 _6863_ (.A(_2899_),
    .B(_2905_),
    .C(_2924_),
    .X(_2925_));
 sg13g2_xor2_1 _6864_ (.B(_2924_),
    .A(_2906_),
    .X(_2926_));
 sg13g2_a21o_1 _6865_ (.A2(_2911_),
    .A1(_2908_),
    .B1(_2926_),
    .X(_2927_));
 sg13g2_nand3_1 _6866_ (.B(_2911_),
    .C(_2926_),
    .A(_2908_),
    .Y(_2928_));
 sg13g2_nand3_1 _6867_ (.B(_2927_),
    .C(_2928_),
    .A(net931),
    .Y(_2929_));
 sg13g2_nor2b_1 _6868_ (.A(_0029_),
    .B_N(_2896_),
    .Y(_2930_));
 sg13g2_xnor2_1 _6869_ (.Y(_2931_),
    .A(_3171_),
    .B(_2930_));
 sg13g2_a21oi_1 _6870_ (.A1(net927),
    .A2(_2931_),
    .Y(_2932_),
    .B1(net875));
 sg13g2_a22oi_1 _6871_ (.Y(_0344_),
    .B1(_2929_),
    .B2(_2932_),
    .A2(net875),
    .A1(_3171_));
 sg13g2_o21ai_1 _6872_ (.B1(_2921_),
    .Y(_2933_),
    .A1(net1031),
    .A2(net1036));
 sg13g2_nand3_1 _6873_ (.B(net1034),
    .C(_2900_),
    .A(net1030),
    .Y(_2934_));
 sg13g2_o21ai_1 _6874_ (.B1(_2934_),
    .Y(_2935_),
    .A1(net1030),
    .A2(net1034));
 sg13g2_and2_1 _6875_ (.A(_2933_),
    .B(_2935_),
    .X(_2936_));
 sg13g2_xnor2_1 _6876_ (.Y(_2937_),
    .A(_2933_),
    .B(_2935_));
 sg13g2_nor2_1 _6877_ (.A(_2923_),
    .B(_2937_),
    .Y(_2938_));
 sg13g2_xnor2_1 _6878_ (.Y(_2939_),
    .A(_2923_),
    .B(_2937_));
 sg13g2_a21oi_1 _6879_ (.A1(_2925_),
    .A2(_2927_),
    .Y(_2940_),
    .B1(_2939_));
 sg13g2_and3_1 _6880_ (.X(_2941_),
    .A(_2925_),
    .B(_2927_),
    .C(_2939_));
 sg13g2_and3_1 _6881_ (.X(_2942_),
    .A(\vgademo.plane_u[14] ),
    .B(\vgademo.plane_u[15] ),
    .C(_2896_));
 sg13g2_o21ai_1 _6882_ (.B1(net931),
    .Y(_2943_),
    .A1(_2940_),
    .A2(_2941_));
 sg13g2_xor2_1 _6883_ (.B(_2942_),
    .A(_0030_),
    .X(_2944_));
 sg13g2_a21oi_1 _6884_ (.A1(net923),
    .A2(_2944_),
    .Y(_2945_),
    .B1(net874));
 sg13g2_a22oi_1 _6885_ (.Y(_2946_),
    .B1(_2943_),
    .B2(_2945_),
    .A2(net874),
    .A1(net409));
 sg13g2_inv_1 _6886_ (.Y(_0345_),
    .A(net410));
 sg13g2_nand2_1 _6887_ (.Y(_2947_),
    .A(net387),
    .B(net874));
 sg13g2_a21oi_2 _6888_ (.B1(net1033),
    .Y(_2948_),
    .A2(net1034),
    .A1(net1030));
 sg13g2_nand3_1 _6889_ (.B(net1033),
    .C(net1034),
    .A(net1030),
    .Y(_2949_));
 sg13g2_nor2b_1 _6890_ (.A(_2948_),
    .B_N(_2949_),
    .Y(_2950_));
 sg13g2_nand2_1 _6891_ (.Y(_2951_),
    .A(_2936_),
    .B(_2950_));
 sg13g2_xnor2_1 _6892_ (.Y(_2952_),
    .A(_2936_),
    .B(_2950_));
 sg13g2_inv_1 _6893_ (.Y(_2953_),
    .A(_2952_));
 sg13g2_o21ai_1 _6894_ (.B1(_2953_),
    .Y(_2954_),
    .A1(_2938_),
    .A2(_2940_));
 sg13g2_or3_1 _6895_ (.A(_2938_),
    .B(_2940_),
    .C(_2953_),
    .X(_2955_));
 sg13g2_and2_1 _6896_ (.A(_2954_),
    .B(_2955_),
    .X(_2956_));
 sg13g2_nand3_1 _6897_ (.B(\vgademo.plane_u[17] ),
    .C(_2942_),
    .A(\vgademo.plane_u[16] ),
    .Y(_2957_));
 sg13g2_inv_1 _6898_ (.Y(_2958_),
    .A(_2957_));
 sg13g2_a21oi_1 _6899_ (.A1(\vgademo.plane_u[16] ),
    .A2(_2942_),
    .Y(_2959_),
    .B1(net387));
 sg13g2_o21ai_1 _6900_ (.B1(net923),
    .Y(_2960_),
    .A1(_2958_),
    .A2(_2959_));
 sg13g2_o21ai_1 _6901_ (.B1(_2960_),
    .Y(_2961_),
    .A1(net923),
    .A2(_2956_));
 sg13g2_o21ai_1 _6902_ (.B1(_2947_),
    .Y(_0346_),
    .A1(net874),
    .A2(_2961_));
 sg13g2_xnor2_1 _6903_ (.Y(_2962_),
    .A(net1031),
    .B(_2948_));
 sg13g2_and3_1 _6904_ (.X(_2963_),
    .A(_2951_),
    .B(_2954_),
    .C(_2962_));
 sg13g2_a21oi_1 _6905_ (.A1(_2951_),
    .A2(_2954_),
    .Y(_2964_),
    .B1(_2962_));
 sg13g2_o21ai_1 _6906_ (.B1(net931),
    .Y(_2965_),
    .A1(_2963_),
    .A2(_2964_));
 sg13g2_xor2_1 _6907_ (.B(_2957_),
    .A(\vgademo.plane_u[18] ),
    .X(_2966_));
 sg13g2_a21oi_1 _6908_ (.A1(net923),
    .A2(_2966_),
    .Y(_2967_),
    .B1(net874));
 sg13g2_a22oi_1 _6909_ (.Y(_2968_),
    .B1(_2965_),
    .B2(_2967_),
    .A2(net874),
    .A1(net504));
 sg13g2_inv_1 _6910_ (.Y(_0347_),
    .A(_2968_));
 sg13g2_a21o_1 _6911_ (.A2(_2948_),
    .A1(net1031),
    .B1(_2964_),
    .X(_2969_));
 sg13g2_nor2_1 _6912_ (.A(net1030),
    .B(net1031),
    .Y(_2970_));
 sg13g2_nand2_1 _6913_ (.Y(_2971_),
    .A(net1030),
    .B(net1031));
 sg13g2_nor2b_1 _6914_ (.A(_2970_),
    .B_N(_2971_),
    .Y(_2972_));
 sg13g2_xnor2_1 _6915_ (.Y(_2973_),
    .A(_2969_),
    .B(_2972_));
 sg13g2_nor2_1 _6916_ (.A(_0031_),
    .B(_2957_),
    .Y(_2974_));
 sg13g2_xnor2_1 _6917_ (.Y(_2975_),
    .A(\vgademo.plane_u[19] ),
    .B(_2974_));
 sg13g2_a21oi_1 _6918_ (.A1(net922),
    .A2(_2975_),
    .Y(_2976_),
    .B1(net874));
 sg13g2_o21ai_1 _6919_ (.B1(_2976_),
    .Y(_2977_),
    .A1(net922),
    .A2(_2973_));
 sg13g2_o21ai_1 _6920_ (.B1(_2977_),
    .Y(_0348_),
    .A1(_3172_),
    .A2(_2702_));
 sg13g2_a21oi_1 _6921_ (.A1(_2964_),
    .A2(_2970_),
    .Y(_2978_),
    .B1(net927));
 sg13g2_o21ai_1 _6922_ (.B1(_2978_),
    .Y(_2979_),
    .A1(_2969_),
    .A2(_2971_));
 sg13g2_nand3_1 _6923_ (.B(\vgademo.plane_u[19] ),
    .C(_2958_),
    .A(\vgademo.plane_u[18] ),
    .Y(_2980_));
 sg13g2_xnor2_1 _6924_ (.Y(_2981_),
    .A(net335),
    .B(_2980_));
 sg13g2_a21oi_1 _6925_ (.A1(net922),
    .A2(_2981_),
    .Y(_2982_),
    .B1(net874));
 sg13g2_a22oi_1 _6926_ (.Y(_0349_),
    .B1(_2979_),
    .B2(_2982_),
    .A2(net875),
    .A1(_3173_));
 sg13g2_nor2_1 _6927_ (.A(_0032_),
    .B(_2980_),
    .Y(_2983_));
 sg13g2_a21oi_1 _6928_ (.A1(net446),
    .A2(_2983_),
    .Y(_2984_),
    .B1(net932));
 sg13g2_o21ai_1 _6929_ (.B1(_2984_),
    .Y(_2985_),
    .A1(net446),
    .A2(_2983_));
 sg13g2_nor2_1 _6930_ (.A(net876),
    .B(_2978_),
    .Y(_2986_));
 sg13g2_a22oi_1 _6931_ (.Y(_0350_),
    .B1(_2985_),
    .B2(_2986_),
    .A2(net875),
    .A1(_3174_));
 sg13g2_nor2_1 _6932_ (.A(_1762_),
    .B(_1774_),
    .Y(_2987_));
 sg13g2_nor2_2 _6933_ (.A(_1804_),
    .B(_2987_),
    .Y(_2988_));
 sg13g2_nor2_1 _6934_ (.A(net860),
    .B(_2988_),
    .Y(_2989_));
 sg13g2_a21o_1 _6935_ (.A2(_2989_),
    .A1(net826),
    .B1(_2209_),
    .X(_2990_));
 sg13g2_a21oi_1 _6936_ (.A1(_1684_),
    .A2(_2990_),
    .Y(_2991_),
    .B1(_2112_));
 sg13g2_or2_1 _6937_ (.X(_2992_),
    .B(_2991_),
    .A(_2204_));
 sg13g2_nand2b_2 _6938_ (.Y(_2993_),
    .B(_1808_),
    .A_N(_1776_));
 sg13g2_nand3_1 _6939_ (.B(net826),
    .C(_2993_),
    .A(net854),
    .Y(_2994_));
 sg13g2_a221oi_1 _6940_ (.B2(_2564_),
    .C1(net862),
    .B1(_2994_),
    .A1(_2110_),
    .Y(_2995_),
    .A2(_2605_));
 sg13g2_nor2_2 _6941_ (.A(_2554_),
    .B(_2995_),
    .Y(_2996_));
 sg13g2_a21o_1 _6942_ (.A2(_2996_),
    .A1(net942),
    .B1(_2992_),
    .X(_2997_));
 sg13g2_o21ai_1 _6943_ (.B1(_2992_),
    .Y(_2998_),
    .A1(net942),
    .A2(_2996_));
 sg13g2_and2_1 _6944_ (.A(_2997_),
    .B(_2998_),
    .X(_2999_));
 sg13g2_inv_1 _6945_ (.Y(_3000_),
    .A(_2999_));
 sg13g2_xor2_1 _6946_ (.B(\vgademo.plane_u[14] ),
    .A(\vgademo.a_cos[9] ),
    .X(_3001_));
 sg13g2_xnor2_1 _6947_ (.Y(_3002_),
    .A(_1749_),
    .B(_3001_));
 sg13g2_o21ai_1 _6948_ (.B1(_1805_),
    .Y(_3003_),
    .A1(_1778_),
    .A2(_3002_));
 sg13g2_nand3_1 _6949_ (.B(_1715_),
    .C(_3003_),
    .A(net830),
    .Y(_3004_));
 sg13g2_xor2_1 _6950_ (.B(_1745_),
    .A(_1741_),
    .X(_3005_));
 sg13g2_o21ai_1 _6951_ (.B1(_2155_),
    .Y(_3006_),
    .A1(_1778_),
    .A2(_3005_));
 sg13g2_o21ai_1 _6952_ (.B1(_3006_),
    .Y(_3007_),
    .A1(net829),
    .A2(_1716_));
 sg13g2_nand3_1 _6953_ (.B(_3004_),
    .C(_3007_),
    .A(net856),
    .Y(_3008_));
 sg13g2_a21oi_2 _6954_ (.B1(net862),
    .Y(_3009_),
    .A2(_3008_),
    .A1(_2095_));
 sg13g2_nor2_1 _6955_ (.A(_2101_),
    .B(_3009_),
    .Y(_3010_));
 sg13g2_xnor2_1 _6956_ (.Y(_3011_),
    .A(_1739_),
    .B(_1751_));
 sg13g2_a21oi_2 _6957_ (.B1(_2119_),
    .Y(_3012_),
    .A2(_3011_),
    .A1(_1777_));
 sg13g2_nand3_1 _6958_ (.B(_1746_),
    .C(_1747_),
    .A(_1740_),
    .Y(_3013_));
 sg13g2_nand2_1 _6959_ (.Y(_3014_),
    .A(_1777_),
    .B(_3013_));
 sg13g2_o21ai_1 _6960_ (.B1(_2171_),
    .Y(_3015_),
    .A1(_1748_),
    .A2(_3014_));
 sg13g2_a21oi_1 _6961_ (.A1(_1717_),
    .A2(_3015_),
    .Y(_3016_),
    .B1(_1314_));
 sg13g2_o21ai_1 _6962_ (.B1(_3016_),
    .Y(_3017_),
    .A1(net826),
    .A2(_3012_));
 sg13g2_a21oi_1 _6963_ (.A1(_2165_),
    .A2(_3017_),
    .Y(_3018_),
    .B1(net862));
 sg13g2_a21o_1 _6964_ (.A2(_3017_),
    .A1(_2165_),
    .B1(net862),
    .X(_3019_));
 sg13g2_xor2_1 _6965_ (.B(_3009_),
    .A(_2101_),
    .X(_3020_));
 sg13g2_a21oi_1 _6966_ (.A1(_3019_),
    .A2(_3020_),
    .Y(_3021_),
    .B1(_3010_));
 sg13g2_o21ai_1 _6967_ (.B1(_3012_),
    .Y(_3022_),
    .A1(net828),
    .A2(net852));
 sg13g2_nand3_1 _6968_ (.B(net853),
    .C(_2988_),
    .A(net830),
    .Y(_3023_));
 sg13g2_nand3_1 _6969_ (.B(_3022_),
    .C(_3023_),
    .A(net855),
    .Y(_3024_));
 sg13g2_and2_1 _6970_ (.A(_1684_),
    .B(_2128_),
    .X(_3025_));
 sg13g2_a21oi_2 _6971_ (.B1(_2110_),
    .Y(_3026_),
    .A2(_3025_),
    .A1(_3024_));
 sg13g2_a21o_1 _6972_ (.A2(_3025_),
    .A1(_3024_),
    .B1(_2110_),
    .X(_3027_));
 sg13g2_nor2_1 _6973_ (.A(_1694_),
    .B(_3026_),
    .Y(_3028_));
 sg13g2_nand2_1 _6974_ (.Y(_3029_),
    .A(_1693_),
    .B(_3027_));
 sg13g2_o21ai_1 _6975_ (.B1(_3003_),
    .Y(_3030_),
    .A1(net828),
    .A2(net852));
 sg13g2_nand3_1 _6976_ (.B(net853),
    .C(_2993_),
    .A(net831),
    .Y(_3031_));
 sg13g2_nand3_1 _6977_ (.B(_3030_),
    .C(_3031_),
    .A(net854),
    .Y(_3032_));
 sg13g2_a21o_2 _6978_ (.A2(_3032_),
    .A1(_2096_),
    .B1(_2144_),
    .X(_3033_));
 sg13g2_and2_1 _6979_ (.A(_2205_),
    .B(_3033_),
    .X(_3034_));
 sg13g2_and3_1 _6980_ (.X(_3035_),
    .A(_2103_),
    .B(_2205_),
    .C(_3033_));
 sg13g2_nand3_1 _6981_ (.B(_2205_),
    .C(_3033_),
    .A(_2103_),
    .Y(_3036_));
 sg13g2_a21oi_1 _6982_ (.A1(_2205_),
    .A2(_3033_),
    .Y(_3037_),
    .B1(_2103_));
 sg13g2_a21o_1 _6983_ (.A2(_3033_),
    .A1(_2205_),
    .B1(_2103_),
    .X(_3038_));
 sg13g2_nor3_1 _6984_ (.A(_3028_),
    .B(_3035_),
    .C(_3037_),
    .Y(_3039_));
 sg13g2_nand3_1 _6985_ (.B(_3036_),
    .C(_3038_),
    .A(_3029_),
    .Y(_3040_));
 sg13g2_a21oi_1 _6986_ (.A1(_3036_),
    .A2(_3038_),
    .Y(_3041_),
    .B1(_3029_));
 sg13g2_o21ai_1 _6987_ (.B1(_3028_),
    .Y(_3042_),
    .A1(_3035_),
    .A2(_3037_));
 sg13g2_nor3_1 _6988_ (.A(_3021_),
    .B(_3039_),
    .C(_3041_),
    .Y(_3043_));
 sg13g2_a21oi_1 _6989_ (.A1(_3029_),
    .A2(_3038_),
    .Y(_3044_),
    .B1(_3035_));
 sg13g2_a21oi_1 _6990_ (.A1(_1693_),
    .A2(_3027_),
    .Y(_3045_),
    .B1(_2148_));
 sg13g2_o21ai_1 _6991_ (.B1(_2147_),
    .Y(_3046_),
    .A1(_1694_),
    .A2(_3026_));
 sg13g2_nor3_1 _6992_ (.A(_1694_),
    .B(_2147_),
    .C(_3026_),
    .Y(_3047_));
 sg13g2_nand3_1 _6993_ (.B(_2148_),
    .C(_3027_),
    .A(_1693_),
    .Y(_3048_));
 sg13g2_nor3_2 _6994_ (.A(_2996_),
    .B(_3045_),
    .C(_3047_),
    .Y(_3049_));
 sg13g2_a221oi_1 _6995_ (.B2(_3048_),
    .C1(_2995_),
    .B1(_3046_),
    .A1(net863),
    .Y(_3050_),
    .A2(_2203_));
 sg13g2_nor3_1 _6996_ (.A(_3044_),
    .B(_3049_),
    .C(_3050_),
    .Y(_3051_));
 sg13g2_or2_1 _6997_ (.X(_3052_),
    .B(_3051_),
    .A(_3043_));
 sg13g2_o21ai_1 _6998_ (.B1(_3044_),
    .Y(_3053_),
    .A1(_3049_),
    .A2(_3050_));
 sg13g2_xnor2_1 _6999_ (.Y(_3054_),
    .A(_3018_),
    .B(_3020_));
 sg13g2_or2_1 _7000_ (.X(_3055_),
    .B(_3054_),
    .A(_3034_));
 sg13g2_and2_1 _7001_ (.A(_3053_),
    .B(_3055_),
    .X(_3056_));
 sg13g2_a221oi_1 _7002_ (.B2(_3042_),
    .C1(_3010_),
    .B1(_3040_),
    .A1(_3019_),
    .Y(_3057_),
    .A2(_3020_));
 sg13g2_o21ai_1 _7003_ (.B1(_3018_),
    .Y(_3058_),
    .A1(_2214_),
    .A2(_2991_));
 sg13g2_nand2_1 _7004_ (.Y(_3059_),
    .A(_2214_),
    .B(_2992_));
 sg13g2_a22oi_1 _7005_ (.Y(_3060_),
    .B1(_3058_),
    .B2(_3059_),
    .A2(_3054_),
    .A1(_3034_));
 sg13g2_nor4_1 _7006_ (.A(_3043_),
    .B(_3051_),
    .C(_3057_),
    .D(_3060_),
    .Y(_3061_));
 sg13g2_nor2_1 _7007_ (.A(_3045_),
    .B(_3049_),
    .Y(_3062_));
 sg13g2_xnor2_1 _7008_ (.Y(_3063_),
    .A(net942),
    .B(_2996_));
 sg13g2_xnor2_1 _7009_ (.Y(_3064_),
    .A(_2992_),
    .B(_3063_));
 sg13g2_nor2_1 _7010_ (.A(_3062_),
    .B(_3064_),
    .Y(_3065_));
 sg13g2_a221oi_1 _7011_ (.B2(_3061_),
    .C1(_3065_),
    .B1(_3056_),
    .A1(_3052_),
    .Y(_3066_),
    .A2(_3053_));
 sg13g2_nand2_1 _7012_ (.Y(_3067_),
    .A(_3062_),
    .B(_3064_));
 sg13g2_inv_1 _7013_ (.Y(_3068_),
    .A(_3067_));
 sg13g2_o21ai_1 _7014_ (.B1(_3000_),
    .Y(_3069_),
    .A1(_3066_),
    .A2(_3068_));
 sg13g2_nand3b_1 _7015_ (.B(_3067_),
    .C(_2999_),
    .Y(_3070_),
    .A_N(_3066_));
 sg13g2_and3_1 _7016_ (.X(_0351_),
    .A(_2239_),
    .B(_3069_),
    .C(_3070_));
 sg13g2_a21oi_1 _7017_ (.A1(_2997_),
    .A2(_3070_),
    .Y(_0352_),
    .B1(_2238_));
 sg13g2_nor2_1 _7018_ (.A(net280),
    .B(net897),
    .Y(_3071_));
 sg13g2_a21oi_1 _7019_ (.A1(_3086_),
    .A2(net897),
    .Y(_0353_),
    .B1(_3071_));
 sg13g2_nor2_1 _7020_ (.A(net337),
    .B(net897),
    .Y(_3072_));
 sg13g2_a21oi_1 _7021_ (.A1(_3085_),
    .A2(net896),
    .Y(_0354_),
    .B1(_3072_));
 sg13g2_nor2_1 _7022_ (.A(net439),
    .B(net896),
    .Y(_3073_));
 sg13g2_a21oi_1 _7023_ (.A1(_3084_),
    .A2(net896),
    .Y(_0355_),
    .B1(_3073_));
 sg13g2_nor2_1 _7024_ (.A(net486),
    .B(net896),
    .Y(_3074_));
 sg13g2_a21oi_1 _7025_ (.A1(_3083_),
    .A2(net896),
    .Y(_0356_),
    .B1(_3074_));
 sg13g2_nor2_1 _7026_ (.A(\vgademo.plane_du[4] ),
    .B(net896),
    .Y(_3075_));
 sg13g2_a21oi_1 _7027_ (.A1(net1039),
    .A2(net896),
    .Y(_0357_),
    .B1(_3075_));
 sg13g2_mux2_1 _7028_ (.A0(net578),
    .A1(net1037),
    .S(net898),
    .X(_0358_));
 sg13g2_mux2_1 _7029_ (.A0(net597),
    .A1(net1036),
    .S(net898),
    .X(_0359_));
 sg13g2_mux2_1 _7030_ (.A0(net588),
    .A1(net1034),
    .S(net898),
    .X(_0360_));
 sg13g2_nor2_1 _7031_ (.A(net457),
    .B(net898),
    .Y(_3076_));
 sg13g2_a21oi_1 _7032_ (.A1(_3082_),
    .A2(net898),
    .Y(_0361_),
    .B1(_3076_));
 sg13g2_mux2_1 _7033_ (.A0(net950),
    .A1(net1032),
    .S(net897),
    .X(_0362_));
 sg13g2_mux2_1 _7034_ (.A0(\vgademo.plane_du[10] ),
    .A1(net413),
    .S(net896),
    .X(_0363_));
 sg13g2_a21oi_1 _7035_ (.A1(\vgademo.plane_du[0] ),
    .A2(_2702_),
    .Y(_3077_),
    .B1(net258));
 sg13g2_a21oi_1 _7036_ (.A1(net925),
    .A2(_2703_),
    .Y(_3078_),
    .B1(net877));
 sg13g2_nor2_1 _7037_ (.A(net259),
    .B(_3078_),
    .Y(_0364_));
 sg13g2_dfrbp_1 _7038_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net33),
    .D(_0111_),
    .Q_N(_3548_),
    .Q(\vgademo.linelfsr[0] ));
 sg13g2_dfrbp_1 _7039_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net31),
    .D(net507),
    .Q_N(_3547_),
    .Q(\vgademo.linelfsr[1] ));
 sg13g2_dfrbp_1 _7040_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net29),
    .D(net327),
    .Q_N(_3546_),
    .Q(\vgademo.linelfsr[2] ));
 sg13g2_dfrbp_1 _7041_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net27),
    .D(_0114_),
    .Q_N(_3545_),
    .Q(\vgademo.linelfsr[3] ));
 sg13g2_dfrbp_1 _7042_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net25),
    .D(_0115_),
    .Q_N(_3544_),
    .Q(\vgademo.linelfsr[4] ));
 sg13g2_dfrbp_1 _7043_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net23),
    .D(net303),
    .Q_N(_3543_),
    .Q(\vgademo.linelfsr[5] ));
 sg13g2_dfrbp_1 _7044_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net21),
    .D(net375),
    .Q_N(_3542_),
    .Q(\vgademo.linelfsr[6] ));
 sg13g2_dfrbp_1 _7045_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net19),
    .D(net427),
    .Q_N(_3541_),
    .Q(\vgademo.linelfsr[7] ));
 sg13g2_dfrbp_1 _7046_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net17),
    .D(_0119_),
    .Q_N(_3540_),
    .Q(\vgademo.linelfsr[8] ));
 sg13g2_dfrbp_1 _7047_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net15),
    .D(net403),
    .Q_N(_3539_),
    .Q(\vgademo.linelfsr[9] ));
 sg13g2_dfrbp_1 _7048_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net162),
    .D(net311),
    .Q_N(_3538_),
    .Q(\vgademo.linelfsr[10] ));
 sg13g2_dfrbp_1 _7049_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net160),
    .D(_0122_),
    .Q_N(_3537_),
    .Q(\vgademo.linelfsr[11] ));
 sg13g2_dfrbp_1 _7050_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net158),
    .D(_0123_),
    .Q_N(_3536_),
    .Q(\vgademo.linelfsr[12] ));
 sg13g2_dfrbp_1 _7051_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1070),
    .D(net276),
    .Q_N(\vgademo.audio_songpos[0] ),
    .Q(_0085_));
 sg13g2_dfrbp_1 _7052_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1073),
    .D(net204),
    .Q_N(\vgademo.audio_songpos[1] ),
    .Q(_0086_));
 sg13g2_dfrbp_1 _7053_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1073),
    .D(_0126_),
    .Q_N(\vgademo.audio_songpos[2] ),
    .Q(_0087_));
 sg13g2_dfrbp_1 _7054_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1073),
    .D(_0127_),
    .Q_N(\vgademo.audio_songpos[3] ),
    .Q(_0088_));
 sg13g2_dfrbp_1 _7055_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1074),
    .D(_0128_),
    .Q_N(\vgademo.audio_songpos[4] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 _7056_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1073),
    .D(_0129_),
    .Q_N(\vgademo.audio_songpos[5] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 _7057_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1069),
    .D(_0130_),
    .Q_N(\vgademo.audio_songpos[6] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 _7058_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1069),
    .D(net192),
    .Q_N(\vgademo.audio_songpos[7] ),
    .Q(_0092_));
 sg13g2_dfrbp_1 _7059_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net140),
    .D(net565),
    .Q_N(_0025_),
    .Q(\vgademo.plane_dx[1] ));
 sg13g2_dfrbp_1 _7060_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net138),
    .D(_0133_),
    .Q_N(_0026_),
    .Q(\vgademo.plane_dx[2] ));
 sg13g2_dfrbp_1 _7061_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net136),
    .D(_0134_),
    .Q_N(_0023_),
    .Q(\vgademo.plane_dx[3] ));
 sg13g2_dfrbp_1 _7062_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net134),
    .D(_0135_),
    .Q_N(_0024_),
    .Q(\vgademo.plane_dx_div.q[3] ));
 sg13g2_dfrbp_1 _7063_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net132),
    .D(_0136_),
    .Q_N(_3535_),
    .Q(\vgademo.plane_dx_div.q[4] ));
 sg13g2_dfrbp_1 _7064_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net130),
    .D(_0137_),
    .Q_N(_3534_),
    .Q(\vgademo.plane_dx_div.q[5] ));
 sg13g2_dfrbp_1 _7065_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net128),
    .D(_0138_),
    .Q_N(_3533_),
    .Q(\vgademo.plane_dx_div.q[6] ));
 sg13g2_dfrbp_1 _7066_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net126),
    .D(_0139_),
    .Q_N(_3532_),
    .Q(\vgademo.plane_dx_div.q[7] ));
 sg13g2_dfrbp_1 _7067_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net124),
    .D(_0140_),
    .Q_N(_3531_),
    .Q(\vgademo.plane_dx_div.q[8] ));
 sg13g2_dfrbp_1 _7068_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net122),
    .D(_0141_),
    .Q_N(_3530_),
    .Q(\vgademo.plane_dx_div.q[9] ));
 sg13g2_dfrbp_1 _7069_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net120),
    .D(net173),
    .Q_N(_0084_),
    .Q(\vgademo.plane_dx_div.i[0] ));
 sg13g2_dfrbp_1 _7070_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net118),
    .D(net334),
    .Q_N(_3529_),
    .Q(\vgademo.plane_dx_div.i[1] ));
 sg13g2_dfrbp_1 _7071_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net116),
    .D(_0144_),
    .Q_N(_3528_),
    .Q(\vgademo.plane_dx_div.i[2] ));
 sg13g2_dfrbp_1 _7072_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net34),
    .D(_0145_),
    .Q_N(_3549_),
    .Q(\vgademo.plane_dx_div.i[3] ));
 sg13g2_dfrbp_1 _7073_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1072),
    .D(\vgademo.soundtrack.sigma_delta_accum_[0] ),
    .Q_N(_3550_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[0] ));
 sg13g2_dfrbp_1 _7074_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1072),
    .D(\vgademo.soundtrack.sigma_delta_accum_[1] ),
    .Q_N(_3551_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[1] ));
 sg13g2_dfrbp_1 _7075_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net1071),
    .D(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .Q_N(_3552_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[2] ));
 sg13g2_dfrbp_1 _7076_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1068),
    .D(net317),
    .Q_N(_3553_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[3] ));
 sg13g2_dfrbp_1 _7077_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1068),
    .D(net551),
    .Q_N(_3554_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[4] ));
 sg13g2_dfrbp_1 _7078_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1068),
    .D(\vgademo.soundtrack.sigma_delta_accum_[5] ),
    .Q_N(_3555_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[5] ));
 sg13g2_dfrbp_1 _7079_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1068),
    .D(net547),
    .Q_N(_3556_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[6] ));
 sg13g2_dfrbp_1 _7080_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1068),
    .D(net503),
    .Q_N(_3557_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[7] ));
 sg13g2_dfrbp_1 _7081_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1068),
    .D(\vgademo.soundtrack.sigma_delta_accum_[8] ),
    .Q_N(_3558_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[8] ));
 sg13g2_dfrbp_1 _7082_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1070),
    .D(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .Q_N(_3559_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[9] ));
 sg13g2_dfrbp_1 _7083_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1070),
    .D(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .Q_N(_3560_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[10] ));
 sg13g2_dfrbp_1 _7084_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1070),
    .D(net530),
    .Q_N(_3561_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[11] ));
 sg13g2_dfrbp_1 _7085_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1069),
    .D(net523),
    .Q_N(_3562_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[12] ));
 sg13g2_dfrbp_1 _7086_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1069),
    .D(net513),
    .Q_N(_3563_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[13] ));
 sg13g2_dfrbp_1 _7087_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1069),
    .D(\vgademo.soundtrack.sigma_delta_accum_[14] ),
    .Q_N(_3564_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[14] ));
 sg13g2_dfrbp_1 _7088_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1069),
    .D(\vgademo.soundtrack.sigma_delta_accum_[15] ),
    .Q_N(_3527_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[15] ));
 sg13g2_dfrbp_1 _7089_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1074),
    .D(net323),
    .Q_N(_0058_),
    .Q(\vgademo.audio_beat_out[0] ));
 sg13g2_dfrbp_1 _7090_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1074),
    .D(net372),
    .Q_N(_0059_),
    .Q(\vgademo.audio_beat_out[1] ));
 sg13g2_dfrbp_1 _7091_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1073),
    .D(_0148_),
    .Q_N(_0062_),
    .Q(\vgademo.audio_beat_out[2] ));
 sg13g2_dfrbp_1 _7092_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1073),
    .D(net354),
    .Q_N(_0057_),
    .Q(\vgademo.audio_beat_out[3] ));
 sg13g2_dfrbp_1 _7093_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1073),
    .D(net492),
    .Q_N(_0055_),
    .Q(\vgademo.audio_beat_out[4] ));
 sg13g2_dfrbp_1 _7094_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1075),
    .D(_0151_),
    .Q_N(_3526_),
    .Q(\vgademo.soundtrack.tri_osc_i[0] ));
 sg13g2_dfrbp_1 _7095_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1072),
    .D(_0152_),
    .Q_N(_3525_),
    .Q(\vgademo.soundtrack.tri_osc_i[1] ));
 sg13g2_dfrbp_1 _7096_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1072),
    .D(_0153_),
    .Q_N(_3524_),
    .Q(\vgademo.soundtrack.tri_osc_i[2] ));
 sg13g2_dfrbp_1 _7097_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1072),
    .D(_0154_),
    .Q_N(_3523_),
    .Q(\vgademo.soundtrack.tri_osc_i[3] ));
 sg13g2_dfrbp_1 _7098_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1081),
    .D(_0155_),
    .Q_N(_3522_),
    .Q(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_dfrbp_1 _7099_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1085),
    .D(_0156_),
    .Q_N(_3521_),
    .Q(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_dfrbp_1 _7100_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1088),
    .D(_0157_),
    .Q_N(_3520_),
    .Q(\vgademo.soundtrack.tri_osc_i[6] ));
 sg13g2_dfrbp_1 _7101_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1081),
    .D(_0158_),
    .Q_N(_3519_),
    .Q(\vgademo.soundtrack.tri_osc_i[7] ));
 sg13g2_dfrbp_1 _7102_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1081),
    .D(_0159_),
    .Q_N(_3518_),
    .Q(\vgademo.soundtrack.tri_osc_i[8] ));
 sg13g2_dfrbp_1 _7103_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net113),
    .D(net262),
    .Q_N(_3517_),
    .Q(audio));
 sg13g2_dfrbp_1 _7104_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1082),
    .D(net181),
    .Q_N(\vgademo.soundtrack.tick_div_[0] ),
    .Q(\vgademo.soundtrack.tick_div[0] ));
 sg13g2_dfrbp_1 _7105_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1082),
    .D(net484),
    .Q_N(_3516_),
    .Q(\vgademo.soundtrack.tick_div[1] ));
 sg13g2_dfrbp_1 _7106_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1082),
    .D(net241),
    .Q_N(_3515_),
    .Q(\vgademo.soundtrack.tick_div[2] ));
 sg13g2_dfrbp_1 _7107_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1082),
    .D(net232),
    .Q_N(_3514_),
    .Q(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_dfrbp_1 _7108_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1082),
    .D(net217),
    .Q_N(_3513_),
    .Q(\vgademo.soundtrack.tick_div[4] ));
 sg13g2_dfrbp_1 _7109_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1087),
    .D(net264),
    .Q_N(_3512_),
    .Q(\vgademo.soundtrack.tick_div[5] ));
 sg13g2_dfrbp_1 _7110_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1087),
    .D(net200),
    .Q_N(_3511_),
    .Q(\vgademo.soundtrack.tick_div[6] ));
 sg13g2_dfrbp_1 _7111_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1085),
    .D(_0168_),
    .Q_N(_3510_),
    .Q(\vgademo.soundtrack.tick_div[7] ));
 sg13g2_dfrbp_1 _7112_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1080),
    .D(net167),
    .Q_N(\vgademo.soundtrack.noise_lfsr[0] ),
    .Q(_0093_));
 sg13g2_dfrbp_1 _7113_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1080),
    .D(net175),
    .Q_N(\vgademo.soundtrack.noise_lfsr[1] ),
    .Q(_0094_));
 sg13g2_dfrbp_1 _7114_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1080),
    .D(net169),
    .Q_N(\vgademo.soundtrack.noise_lfsr[2] ),
    .Q(_0095_));
 sg13g2_dfrbp_1 _7115_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1072),
    .D(net223),
    .Q_N(\vgademo.soundtrack.noise_lfsr[3] ),
    .Q(_0096_));
 sg13g2_dfrbp_1 _7116_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1080),
    .D(net230),
    .Q_N(_0040_),
    .Q(\vgademo.soundtrack.noise_lfsr[4] ));
 sg13g2_dfrbp_1 _7117_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1081),
    .D(net185),
    .Q_N(\vgademo.soundtrack.noise_lfsr[5] ),
    .Q(_0097_));
 sg13g2_dfrbp_1 _7118_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1081),
    .D(net248),
    .Q_N(_0083_),
    .Q(\vgademo.soundtrack.noise_lfsr[6] ));
 sg13g2_dfrbp_1 _7119_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1081),
    .D(net179),
    .Q_N(\vgademo.soundtrack.noise_lfsr[7] ),
    .Q(_0098_));
 sg13g2_dfrbp_1 _7120_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1080),
    .D(net301),
    .Q_N(_0082_),
    .Q(\vgademo.soundtrack.noise_lfsr[8] ));
 sg13g2_dfrbp_1 _7121_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1080),
    .D(net171),
    .Q_N(_3509_),
    .Q(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_dfrbp_1 _7122_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1080),
    .D(net187),
    .Q_N(\vgademo.soundtrack.noise_lfsr[10] ),
    .Q(_0099_));
 sg13g2_dfrbp_1 _7123_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1080),
    .D(net177),
    .Q_N(\vgademo.soundtrack.noise_lfsr[11] ),
    .Q(_0100_));
 sg13g2_dfrbp_1 _7124_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1084),
    .D(net183),
    .Q_N(\vgademo.soundtrack.noise_lfsr[12] ),
    .Q(_0101_));
 sg13g2_dfrbp_1 _7125_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1084),
    .D(net219),
    .Q_N(_0081_),
    .Q(\vgademo.soundtrack.noise_lfsr[13] ));
 sg13g2_dfrbp_1 _7126_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1081),
    .D(net292),
    .Q_N(_3508_),
    .Q(\vgademo.soundtrack.noise_lfsr[14] ));
 sg13g2_dfrbp_1 _7127_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1085),
    .D(net189),
    .Q_N(\vgademo.audio_snare_frames[0] ),
    .Q(_0102_));
 sg13g2_dfrbp_1 _7128_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1085),
    .D(net195),
    .Q_N(\vgademo.audio_snare_frames[1] ),
    .Q(_0103_));
 sg13g2_dfrbp_1 _7129_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1074),
    .D(net214),
    .Q_N(\vgademo.audio_snare_frames[2] ),
    .Q(_0104_));
 sg13g2_dfrbp_1 _7130_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1074),
    .D(_0187_),
    .Q_N(\vgademo.audio_snare_frames[3] ),
    .Q(_0105_));
 sg13g2_dfrbp_1 _7131_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net86),
    .D(_0188_),
    .Q_N(_3507_),
    .Q(\vgademo.soundtrack.pulse_osc_p[0] ));
 sg13g2_dfrbp_1 _7132_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net85),
    .D(net266),
    .Q_N(_0042_),
    .Q(\vgademo.soundtrack.pulse_osc_p[1] ));
 sg13g2_dfrbp_1 _7133_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net84),
    .D(net329),
    .Q_N(_3506_),
    .Q(\vgademo.soundtrack.pulse_osc_p[2] ));
 sg13g2_dfrbp_1 _7134_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net83),
    .D(_0191_),
    .Q_N(_3505_),
    .Q(\vgademo.soundtrack.pulse_osc_p[3] ));
 sg13g2_dfrbp_1 _7135_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net79),
    .D(net255),
    .Q_N(_3504_),
    .Q(\vgademo.soundtrack.pulse_osc_p[4] ));
 sg13g2_dfrbp_1 _7136_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net78),
    .D(net298),
    .Q_N(_3503_),
    .Q(\vgademo.soundtrack.pulse_osc_p[5] ));
 sg13g2_dfrbp_1 _7137_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net77),
    .D(_0194_),
    .Q_N(_3502_),
    .Q(\vgademo.soundtrack.pulse_osc_p[6] ));
 sg13g2_dfrbp_1 _7138_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net76),
    .D(_0195_),
    .Q_N(_3501_),
    .Q(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_dfrbp_1 _7139_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net75),
    .D(net252),
    .Q_N(_3500_),
    .Q(\vgademo.soundtrack.pulse_osc_p[8] ));
 sg13g2_dfrbp_1 _7140_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net74),
    .D(net235),
    .Q_N(_3499_),
    .Q(\vgademo.soundtrack.pulse_osc_p[9] ));
 sg13g2_dfrbp_1 _7141_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net73),
    .D(net225),
    .Q_N(_3498_),
    .Q(\vgademo.soundtrack.pulse_osc_p[10] ));
 sg13g2_dfrbp_1 _7142_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net72),
    .D(_0199_),
    .Q_N(_3497_),
    .Q(\vgademo.soundtrack.pulse_osc_p[11] ));
 sg13g2_dfrbp_1 _7143_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net71),
    .D(_0200_),
    .Q_N(_3496_),
    .Q(\vgademo.soundtrack.pulse_osc_p[12] ));
 sg13g2_dfrbp_1 _7144_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net70),
    .D(net244),
    .Q_N(_3495_),
    .Q(\vgademo.soundtrack.pulse_osc_p[13] ));
 sg13g2_dfrbp_1 _7145_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1085),
    .D(_0202_),
    .Q_N(_3494_),
    .Q(\vgademo.audio_kick_frames[0] ));
 sg13g2_dfrbp_1 _7146_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1085),
    .D(_0203_),
    .Q_N(_0068_),
    .Q(\vgademo.audio_kick_frames[1] ));
 sg13g2_dfrbp_1 _7147_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1085),
    .D(_0204_),
    .Q_N(_0060_),
    .Q(\vgademo.audio_kick_frames[2] ));
 sg13g2_dfrbp_1 _7148_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1068),
    .D(_0205_),
    .Q_N(\vgademo.soundtrack.pulse_vol[0] ),
    .Q(_0106_));
 sg13g2_dfrbp_1 _7149_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1071),
    .D(_0206_),
    .Q_N(\vgademo.soundtrack.pulse_vol[1] ),
    .Q(_0107_));
 sg13g2_dfrbp_1 _7150_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1068),
    .D(_0207_),
    .Q_N(\vgademo.soundtrack.pulse_vol[2] ),
    .Q(_0108_));
 sg13g2_dfrbp_1 _7151_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1072),
    .D(net212),
    .Q_N(\vgademo.soundtrack.pulse_vol[3] ),
    .Q(_0109_));
 sg13g2_dfrbp_1 _7152_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1082),
    .D(net165),
    .Q_N(\vgademo.soundtrack.sample_div_[0] ),
    .Q(\vgademo.soundtrack.sample_div[0] ));
 sg13g2_dfrbp_1 _7153_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1083),
    .D(net221),
    .Q_N(_3565_),
    .Q(\vgademo.soundtrack.sample_div[1] ));
 sg13g2_dfrbp_1 _7154_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1083),
    .D(net473),
    .Q_N(_3566_),
    .Q(\vgademo.soundtrack.sample_div[2] ));
 sg13g2_dfrbp_1 _7155_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1083),
    .D(net246),
    .Q_N(_3567_),
    .Q(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_dfrbp_1 _7156_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1082),
    .D(net206),
    .Q_N(_3568_),
    .Q(\vgademo.soundtrack.sample_div[4] ));
 sg13g2_dfrbp_1 _7157_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1082),
    .D(\vgademo.soundtrack.sample_div_[5] ),
    .Q_N(_3569_),
    .Q(\vgademo.soundtrack.sample_div[5] ));
 sg13g2_dfrbp_1 _7158_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1083),
    .D(\vgademo.soundtrack.sample_div_[6] ),
    .Q_N(_3570_),
    .Q(\vgademo.soundtrack.sample_div[6] ));
 sg13g2_dfrbp_1 _7159_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1084),
    .D(net239),
    .Q_N(_3571_),
    .Q(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_dfrbp_1 _7160_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1084),
    .D(net208),
    .Q_N(_3572_),
    .Q(\vgademo.soundtrack.sample_div[8] ));
 sg13g2_dfrbp_1 _7161_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1084),
    .D(\vgademo.soundtrack.sample_div_[9] ),
    .Q_N(_3493_),
    .Q(\vgademo.soundtrack.sample_div[9] ));
 sg13g2_dfrbp_1 _7162_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net61),
    .D(net237),
    .Q_N(_3492_),
    .Q(\vgademo.soundtrack.tri_osc_p[0] ));
 sg13g2_dfrbp_1 _7163_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net60),
    .D(net331),
    .Q_N(_3491_),
    .Q(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_dfrbp_1 _7164_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net59),
    .D(net412),
    .Q_N(_3490_),
    .Q(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_dfrbp_1 _7165_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net58),
    .D(net401),
    .Q_N(_3489_),
    .Q(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_dfrbp_1 _7166_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net57),
    .D(_0213_),
    .Q_N(_3488_),
    .Q(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_dfrbp_1 _7167_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net56),
    .D(net423),
    .Q_N(_3487_),
    .Q(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_dfrbp_1 _7168_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net55),
    .D(_0215_),
    .Q_N(_3486_),
    .Q(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_dfrbp_1 _7169_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net54),
    .D(_0216_),
    .Q_N(_3485_),
    .Q(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_dfrbp_1 _7170_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net53),
    .D(_0217_),
    .Q_N(_3484_),
    .Q(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_dfrbp_1 _7171_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net52),
    .D(net395),
    .Q_N(_0041_),
    .Q(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_dfrbp_1 _7172_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net51),
    .D(net287),
    .Q_N(_3483_),
    .Q(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_dfrbp_1 _7173_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net50),
    .D(_0220_),
    .Q_N(_3482_),
    .Q(\vgademo.soundtrack.tri_osc_p[11] ));
 sg13g2_dfrbp_1 _7174_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net49),
    .D(_0221_),
    .Q_N(_3481_),
    .Q(\vgademo.soundtrack.tri_osc_p[12] ));
 sg13g2_dfrbp_1 _7175_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net48),
    .D(net319),
    .Q_N(_3480_),
    .Q(\vgademo.soundtrack.tri_osc_p[13] ));
 sg13g2_dfrbp_1 _7176_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net47),
    .D(net370),
    .Q_N(_3479_),
    .Q(\vgademo.soundtrack.tri_osc_p[14] ));
 sg13g2_dfrbp_1 _7177_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net46),
    .D(net432),
    .Q_N(_3478_),
    .Q(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_dfrbp_1 _7178_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net45),
    .D(_0225_),
    .Q_N(_3477_),
    .Q(\vgademo.plane_dx_div.d[16] ));
 sg13g2_dfrbp_1 _7179_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net44),
    .D(_0226_),
    .Q_N(_0070_),
    .Q(\vgademo.plane_dx_div.d[17] ));
 sg13g2_dfrbp_1 _7180_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net43),
    .D(_0227_),
    .Q_N(_0073_),
    .Q(\vgademo.plane_dx_div.d[18] ));
 sg13g2_dfrbp_1 _7181_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net42),
    .D(_0228_),
    .Q_N(_0076_),
    .Q(\vgademo.plane_dx_div.d[19] ));
 sg13g2_dfrbp_1 _7182_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net41),
    .D(_0229_),
    .Q_N(_0079_),
    .Q(\vgademo.plane_dx_div.d[20] ));
 sg13g2_dfrbp_1 _7183_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net40),
    .D(_0230_),
    .Q_N(_0013_),
    .Q(\vgademo.plane_dx_div.d[21] ));
 sg13g2_dfrbp_1 _7184_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net39),
    .D(_0231_),
    .Q_N(_0014_),
    .Q(\vgademo.plane_dx_div.d[22] ));
 sg13g2_dfrbp_1 _7185_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net38),
    .D(_0232_),
    .Q_N(_0018_),
    .Q(\vgademo.plane_dx_div.d[23] ));
 sg13g2_dfrbp_1 _7186_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net80),
    .D(_0233_),
    .Q_N(_0021_),
    .Q(\vgademo.plane_dx_div.d[24] ));
 sg13g2_dfrbp_1 _7187_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net81),
    .D(_0012_),
    .Q_N(_3573_),
    .Q(\vgademo.vsync ));
 sg13g2_dfrbp_1 _7188_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net82),
    .D(_0011_),
    .Q_N(_3574_),
    .Q(hsync));
 sg13g2_dfrbp_1 _7189_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1069),
    .D(_0000_),
    .Q_N(_3575_),
    .Q(\vgademo.h_count[0] ));
 sg13g2_dfrbp_1 _7190_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1069),
    .D(_0002_),
    .Q_N(_3576_),
    .Q(\vgademo.h_count[1] ));
 sg13g2_dfrbp_1 _7191_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1073),
    .D(_0003_),
    .Q_N(_0033_),
    .Q(\vgademo.h_count[2] ));
 sg13g2_dfrbp_1 _7192_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1078),
    .D(_0004_),
    .Q_N(_0034_),
    .Q(\vgademo.h_count[3] ));
 sg13g2_dfrbp_1 _7193_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(_0005_),
    .Q_N(_0044_),
    .Q(\vgademo.h_count[4] ));
 sg13g2_dfrbp_1 _7194_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(net294),
    .Q_N(_0035_),
    .Q(\vgademo.h_count[5] ));
 sg13g2_dfrbp_1 _7195_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1078),
    .D(net591),
    .Q_N(_0036_),
    .Q(\vgademo.h_count[6] ));
 sg13g2_dfrbp_1 _7196_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1078),
    .D(net557),
    .Q_N(_0037_),
    .Q(\vgademo.h_count[7] ));
 sg13g2_dfrbp_1 _7197_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(_0009_),
    .Q_N(_0038_),
    .Q(\vgademo.h_count[8] ));
 sg13g2_dfrbp_1 _7198_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(net257),
    .Q_N(_0039_),
    .Q(\vgademo.h_count[9] ));
 sg13g2_dfrbp_1 _7199_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1078),
    .D(_0001_),
    .Q_N(_0061_),
    .Q(\vgademo.h_count[10] ));
 sg13g2_dfrbp_1 _7200_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1078),
    .D(_0234_),
    .Q_N(_0064_),
    .Q(\vgademo.a_scrolly[3] ));
 sg13g2_dfrbp_1 _7201_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1078),
    .D(_0235_),
    .Q_N(_0069_),
    .Q(\vgademo.a_scrolly[4] ));
 sg13g2_dfrbp_1 _7202_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1078),
    .D(_0236_),
    .Q_N(_0056_),
    .Q(\vgademo.a_scrolly[5] ));
 sg13g2_dfrbp_1 _7203_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1076),
    .D(net596),
    .Q_N(_0075_),
    .Q(\vgademo.a_scrolly[6] ));
 sg13g2_dfrbp_1 _7204_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(net549),
    .Q_N(_0078_),
    .Q(\vgademo.a_scrolly[7] ));
 sg13g2_dfrbp_1 _7205_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(_0239_),
    .Q_N(_0080_),
    .Q(\vgademo.a_scrolly[8] ));
 sg13g2_dfrbp_1 _7206_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1077),
    .D(_0240_),
    .Q_N(_0065_),
    .Q(\vgademo.a_scrolly[9] ));
 sg13g2_dfrbp_1 _7207_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1077),
    .D(_0241_),
    .Q_N(_0016_),
    .Q(\vgademo.a_scrolly[10] ));
 sg13g2_dfrbp_1 _7208_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1077),
    .D(net528),
    .Q_N(_0020_),
    .Q(\vgademo.a_scrolly[11] ));
 sg13g2_dfrbp_1 _7209_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1076),
    .D(net519),
    .Q_N(_0067_),
    .Q(\vgademo.a_scrolly[12] ));
 sg13g2_dfrbp_1 _7210_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1077),
    .D(_0244_),
    .Q_N(_0066_),
    .Q(\vgademo.a_scrolly[13] ));
 sg13g2_dfrbp_1 _7211_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1079),
    .D(_0245_),
    .Q_N(_3476_),
    .Q(\vgademo.bayer_j[0] ));
 sg13g2_dfrbp_1 _7212_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net1092),
    .D(_0246_),
    .Q_N(_0072_),
    .Q(\vgademo.bayer_j[1] ));
 sg13g2_dfrbp_1 _7213_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1092),
    .D(net417),
    .Q_N(_0071_),
    .Q(\vgademo.v_count[2] ));
 sg13g2_dfrbp_1 _7214_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1092),
    .D(net461),
    .Q_N(_0074_),
    .Q(\vgademo.v_count[3] ));
 sg13g2_dfrbp_1 _7215_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1091),
    .D(_0249_),
    .Q_N(_0077_),
    .Q(\vgademo.v_count[4] ));
 sg13g2_dfrbp_1 _7216_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1091),
    .D(_0250_),
    .Q_N(_0063_),
    .Q(\vgademo.v_count[5] ));
 sg13g2_dfrbp_1 _7217_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1091),
    .D(net536),
    .Q_N(_0017_),
    .Q(\vgademo.v_count[6] ));
 sg13g2_dfrbp_1 _7218_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1091),
    .D(net498),
    .Q_N(_0015_),
    .Q(\vgademo.v_count[7] ));
 sg13g2_dfrbp_1 _7219_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1091),
    .D(net500),
    .Q_N(_0019_),
    .Q(\vgademo.v_count[8] ));
 sg13g2_dfrbp_1 _7220_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1091),
    .D(net391),
    .Q_N(_0022_),
    .Q(\vgademo.v_count[9] ));
 sg13g2_dfrbp_1 _7221_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net37),
    .D(_0255_),
    .Q_N(_3475_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7222_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net36),
    .D(_0256_),
    .Q_N(_3474_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7223_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1090),
    .D(net250),
    .Q_N(_3473_),
    .Q(\vgademo.a_cos[0] ));
 sg13g2_dfrbp_1 _7224_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1090),
    .D(net325),
    .Q_N(_3472_),
    .Q(\vgademo.a_cos[1] ));
 sg13g2_dfrbp_1 _7225_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1089),
    .D(_0259_),
    .Q_N(_3471_),
    .Q(\vgademo.a_cos[2] ));
 sg13g2_dfrbp_1 _7226_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1089),
    .D(_0260_),
    .Q_N(_3470_),
    .Q(\vgademo.a_cos[3] ));
 sg13g2_dfrbp_1 _7227_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1089),
    .D(_0261_),
    .Q_N(_3469_),
    .Q(\vgademo.a_cos[4] ));
 sg13g2_dfrbp_1 _7228_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1093),
    .D(_0262_),
    .Q_N(_3468_),
    .Q(\vgademo.a_cos[5] ));
 sg13g2_dfrbp_1 _7229_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1093),
    .D(net526),
    .Q_N(_3467_),
    .Q(\vgademo.a_cos[6] ));
 sg13g2_dfrbp_1 _7230_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1093),
    .D(_0264_),
    .Q_N(_3466_),
    .Q(\vgademo.a_cos[7] ));
 sg13g2_dfrbp_1 _7231_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1090),
    .D(_0265_),
    .Q_N(_3465_),
    .Q(\vgademo.a_cos[8] ));
 sg13g2_dfrbp_1 _7232_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1086),
    .D(_0266_),
    .Q_N(_3464_),
    .Q(\vgademo.a_cos[9] ));
 sg13g2_dfrbp_1 _7233_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1086),
    .D(_0267_),
    .Q_N(_3463_),
    .Q(\vgademo.a_cos[10] ));
 sg13g2_dfrbp_1 _7234_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1086),
    .D(_0268_),
    .Q_N(_3462_),
    .Q(\vgademo.a_cos[11] ));
 sg13g2_dfrbp_1 _7235_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1086),
    .D(_0269_),
    .Q_N(_3461_),
    .Q(\vgademo.a_cos[12] ));
 sg13g2_dfrbp_1 _7236_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1085),
    .D(_0270_),
    .Q_N(\vgademo.a_cos[13] ),
    .Q(_0110_));
 sg13g2_dfrbp_1 _7237_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1086),
    .D(_0271_),
    .Q_N(_3460_),
    .Q(\vgademo.a_cos[14] ));
 sg13g2_dfrbp_1 _7238_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1093),
    .D(_0272_),
    .Q_N(_3459_),
    .Q(\vgademo.a_sin[0] ));
 sg13g2_dfrbp_1 _7239_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1090),
    .D(_0273_),
    .Q_N(_3458_),
    .Q(\vgademo.a_sin[1] ));
 sg13g2_dfrbp_1 _7240_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1090),
    .D(_0274_),
    .Q_N(_3457_),
    .Q(\vgademo.a_sin[2] ));
 sg13g2_dfrbp_1 _7241_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1087),
    .D(_0275_),
    .Q_N(_3456_),
    .Q(\vgademo.a_sin[3] ));
 sg13g2_dfrbp_1 _7242_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1087),
    .D(_0276_),
    .Q_N(_3455_),
    .Q(\vgademo.a_sin[4] ));
 sg13g2_dfrbp_1 _7243_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1087),
    .D(_0277_),
    .Q_N(_3454_),
    .Q(\vgademo.a_sin[5] ));
 sg13g2_dfrbp_1 _7244_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1090),
    .D(_0278_),
    .Q_N(_3453_),
    .Q(\vgademo.a_sin[6] ));
 sg13g2_dfrbp_1 _7245_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1090),
    .D(_0279_),
    .Q_N(_3452_),
    .Q(\vgademo.a_sin[7] ));
 sg13g2_dfrbp_1 _7246_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1089),
    .D(net470),
    .Q_N(_3451_),
    .Q(\vgademo.a_sin[8] ));
 sg13g2_dfrbp_1 _7247_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1089),
    .D(_0281_),
    .Q_N(_3450_),
    .Q(\vgademo.a_sin[9] ));
 sg13g2_dfrbp_1 _7248_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1089),
    .D(_0282_),
    .Q_N(_3449_),
    .Q(\vgademo.a_sin[10] ));
 sg13g2_dfrbp_1 _7249_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1094),
    .D(_0283_),
    .Q_N(_3448_),
    .Q(\vgademo.a_sin[11] ));
 sg13g2_dfrbp_1 _7250_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1089),
    .D(_0284_),
    .Q_N(_3447_),
    .Q(\vgademo.a_sin[12] ));
 sg13g2_dfrbp_1 _7251_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1089),
    .D(_0285_),
    .Q_N(_3446_),
    .Q(\vgademo.a_sin[13] ));
 sg13g2_dfrbp_1 _7252_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1087),
    .D(_0286_),
    .Q_N(_3445_),
    .Q(\vgademo.a_sin[14] ));
 sg13g2_dfrbp_1 _7253_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net32),
    .D(_0287_),
    .Q_N(_3444_),
    .Q(\vgademo.scanline_audio_sample[0] ));
 sg13g2_dfrbp_1 _7254_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net30),
    .D(_0288_),
    .Q_N(_3443_),
    .Q(\vgademo.scanline_audio_sample[1] ));
 sg13g2_dfrbp_1 _7255_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net28),
    .D(_0289_),
    .Q_N(_3442_),
    .Q(\vgademo.scanline_audio_sample[2] ));
 sg13g2_dfrbp_1 _7256_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net26),
    .D(_0290_),
    .Q_N(_3441_),
    .Q(\vgademo.scanline_audio_sample[3] ));
 sg13g2_dfrbp_1 _7257_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net24),
    .D(_0291_),
    .Q_N(_3440_),
    .Q(\vgademo.scanline_audio_sample[4] ));
 sg13g2_dfrbp_1 _7258_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net22),
    .D(_0292_),
    .Q_N(_0043_),
    .Q(\vgademo.scanline_audio_sample[5] ));
 sg13g2_dfrbp_1 _7259_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net20),
    .D(_0293_),
    .Q_N(_3439_),
    .Q(\vgademo.scanline_audio_sample[6] ));
 sg13g2_dfrbp_1 _7260_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net18),
    .D(net309),
    .Q_N(_3438_),
    .Q(\vgademo.b_cos[0] ));
 sg13g2_dfrbp_1 _7261_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net16),
    .D(net344),
    .Q_N(_3437_),
    .Q(\vgademo.b_cos[1] ));
 sg13g2_dfrbp_1 _7262_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net163),
    .D(_0296_),
    .Q_N(_3436_),
    .Q(\vgademo.b_cos[2] ));
 sg13g2_dfrbp_1 _7263_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net161),
    .D(net386),
    .Q_N(_3435_),
    .Q(\vgademo.b_cos[3] ));
 sg13g2_dfrbp_1 _7264_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net159),
    .D(net408),
    .Q_N(_3434_),
    .Q(\vgademo.b_cos[4] ));
 sg13g2_dfrbp_1 _7265_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net157),
    .D(_0299_),
    .Q_N(_3433_),
    .Q(\vgademo.b_cos[5] ));
 sg13g2_dfrbp_1 _7266_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net156),
    .D(_0300_),
    .Q_N(_3432_),
    .Q(\vgademo.b_cos[6] ));
 sg13g2_dfrbp_1 _7267_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net155),
    .D(net489),
    .Q_N(_3431_),
    .Q(\vgademo.b_cos[7] ));
 sg13g2_dfrbp_1 _7268_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net154),
    .D(_0302_),
    .Q_N(_3430_),
    .Q(\vgademo.b_cos[8] ));
 sg13g2_dfrbp_1 _7269_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net153),
    .D(net516),
    .Q_N(_3429_),
    .Q(\vgademo.b_cos[9] ));
 sg13g2_dfrbp_1 _7270_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net152),
    .D(_0304_),
    .Q_N(_3428_),
    .Q(\vgademo.b_cos[10] ));
 sg13g2_dfrbp_1 _7271_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net151),
    .D(_0305_),
    .Q_N(_3427_),
    .Q(\vgademo.b_cos[11] ));
 sg13g2_dfrbp_1 _7272_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net150),
    .D(net341),
    .Q_N(_3426_),
    .Q(\vgademo.plane_dx_div.r[16] ));
 sg13g2_dfrbp_1 _7273_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net149),
    .D(_0307_),
    .Q_N(_3425_),
    .Q(\vgademo.plane_dx_div.r[17] ));
 sg13g2_dfrbp_1 _7274_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net148),
    .D(net359),
    .Q_N(_3424_),
    .Q(\vgademo.plane_dx_div.r[18] ));
 sg13g2_dfrbp_1 _7275_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net147),
    .D(_0309_),
    .Q_N(_3423_),
    .Q(\vgademo.plane_dx_div.r[19] ));
 sg13g2_dfrbp_1 _7276_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net146),
    .D(net279),
    .Q_N(_3422_),
    .Q(\vgademo.plane_dx_div.r[20] ));
 sg13g2_dfrbp_1 _7277_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net145),
    .D(_0311_),
    .Q_N(_3421_),
    .Q(\vgademo.plane_dx_div.r[21] ));
 sg13g2_dfrbp_1 _7278_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0312_),
    .Q_N(_3420_),
    .Q(\vgademo.plane_dx_div.r[22] ));
 sg13g2_dfrbp_1 _7279_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net143),
    .D(_0313_),
    .Q_N(_3419_),
    .Q(\vgademo.plane_dx_div.r[23] ));
 sg13g2_dfrbp_1 _7280_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net142),
    .D(_0314_),
    .Q_N(_3418_),
    .Q(\vgademo.plane_dx_div.r[24] ));
 sg13g2_dfrbp_1 _7281_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net141),
    .D(net346),
    .Q_N(\vgademo.plane_dx[0] ),
    .Q(\vgademo.plane_dx_div.r[25] ));
 sg13g2_dfrbp_1 _7282_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net139),
    .D(_0316_),
    .Q_N(_3417_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7283_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0317_),
    .Q_N(_3416_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7284_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net135),
    .D(net384),
    .Q_N(_3415_),
    .Q(\vgademo.b_sin[0] ));
 sg13g2_dfrbp_1 _7285_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net133),
    .D(net314),
    .Q_N(_3414_),
    .Q(\vgademo.b_sin[1] ));
 sg13g2_dfrbp_1 _7286_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net131),
    .D(net351),
    .Q_N(_3413_),
    .Q(\vgademo.b_sin[2] ));
 sg13g2_dfrbp_1 _7287_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net129),
    .D(net435),
    .Q_N(_3412_),
    .Q(\vgademo.b_sin[3] ));
 sg13g2_dfrbp_1 _7288_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net127),
    .D(net445),
    .Q_N(_3411_),
    .Q(\vgademo.b_sin[4] ));
 sg13g2_dfrbp_1 _7289_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net125),
    .D(net285),
    .Q_N(_3410_),
    .Q(\vgademo.b_sin[5] ));
 sg13g2_dfrbp_1 _7290_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net123),
    .D(_0324_),
    .Q_N(_3409_),
    .Q(\vgademo.b_sin[6] ));
 sg13g2_dfrbp_1 _7291_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net121),
    .D(net305),
    .Q_N(_3408_),
    .Q(\vgademo.b_sin[7] ));
 sg13g2_dfrbp_1 _7292_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net119),
    .D(_0326_),
    .Q_N(_3407_),
    .Q(\vgademo.b_sin[8] ));
 sg13g2_dfrbp_1 _7293_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net117),
    .D(_0327_),
    .Q_N(_3406_),
    .Q(\vgademo.b_sin[9] ));
 sg13g2_dfrbp_1 _7294_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net115),
    .D(_0328_),
    .Q_N(_3405_),
    .Q(\vgademo.b_sin[10] ));
 sg13g2_dfrbp_1 _7295_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net114),
    .D(net542),
    .Q_N(_3404_),
    .Q(\vgademo.b_sin[11] ));
 sg13g2_dfrbp_1 _7296_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net112),
    .D(net296),
    .Q_N(_3403_),
    .Q(\vgademo.plane_u[1] ));
 sg13g2_dfrbp_1 _7297_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net111),
    .D(_0331_),
    .Q_N(_3402_),
    .Q(\vgademo.plane_u[2] ));
 sg13g2_dfrbp_1 _7298_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net110),
    .D(_0332_),
    .Q_N(_3401_),
    .Q(\vgademo.plane_u[3] ));
 sg13g2_dfrbp_1 _7299_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net109),
    .D(_0333_),
    .Q_N(_3400_),
    .Q(\vgademo.plane_u[4] ));
 sg13g2_dfrbp_1 _7300_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net108),
    .D(_0334_),
    .Q_N(_3399_),
    .Q(\vgademo.plane_u[5] ));
 sg13g2_dfrbp_1 _7301_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net107),
    .D(_0335_),
    .Q_N(_3398_),
    .Q(\vgademo.plane_u[6] ));
 sg13g2_dfrbp_1 _7302_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net106),
    .D(_0336_),
    .Q_N(_3397_),
    .Q(\vgademo.plane_u[7] ));
 sg13g2_dfrbp_1 _7303_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net105),
    .D(_0337_),
    .Q_N(_3396_),
    .Q(\vgademo.plane_u[8] ));
 sg13g2_dfrbp_1 _7304_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net104),
    .D(_0338_),
    .Q_N(_3395_),
    .Q(\vgademo.plane_u[9] ));
 sg13g2_dfrbp_1 _7305_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net103),
    .D(_0339_),
    .Q_N(_3394_),
    .Q(\vgademo.plane_u[10] ));
 sg13g2_dfrbp_1 _7306_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net102),
    .D(net283),
    .Q_N(_0027_),
    .Q(\vgademo.plane_u[11] ));
 sg13g2_dfrbp_1 _7307_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net101),
    .D(net421),
    .Q_N(_0028_),
    .Q(\vgademo.plane_u[12] ));
 sg13g2_dfrbp_1 _7308_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net100),
    .D(_0342_),
    .Q_N(_0048_),
    .Q(\vgademo.plane_u[13] ));
 sg13g2_dfrbp_1 _7309_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net99),
    .D(_0343_),
    .Q_N(_0029_),
    .Q(\vgademo.plane_u[14] ));
 sg13g2_dfrbp_1 _7310_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net98),
    .D(_0344_),
    .Q_N(_0047_),
    .Q(\vgademo.plane_u[15] ));
 sg13g2_dfrbp_1 _7311_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net97),
    .D(_0345_),
    .Q_N(_0030_),
    .Q(\vgademo.plane_u[16] ));
 sg13g2_dfrbp_1 _7312_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net96),
    .D(net388),
    .Q_N(_0046_),
    .Q(\vgademo.plane_u[17] ));
 sg13g2_dfrbp_1 _7313_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net95),
    .D(_0347_),
    .Q_N(_0031_),
    .Q(\vgademo.plane_u[18] ));
 sg13g2_dfrbp_1 _7314_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net94),
    .D(net449),
    .Q_N(_0045_),
    .Q(\vgademo.plane_u[19] ));
 sg13g2_dfrbp_1 _7315_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net93),
    .D(_0349_),
    .Q_N(_0032_),
    .Q(\vgademo.plane_u[20] ));
 sg13g2_dfrbp_1 _7316_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net92),
    .D(net447),
    .Q_N(_3393_),
    .Q(\vgademo.plane_u[21] ));
 sg13g2_dfrbp_1 _7317_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net91),
    .D(_0351_),
    .Q_N(_3392_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _7318_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net90),
    .D(_0352_),
    .Q_N(_3391_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _7319_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net89),
    .D(net281),
    .Q_N(_3390_),
    .Q(\vgademo.plane_du[0] ));
 sg13g2_dfrbp_1 _7320_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net88),
    .D(net338),
    .Q_N(_3389_),
    .Q(\vgademo.plane_du[1] ));
 sg13g2_dfrbp_1 _7321_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net87),
    .D(net440),
    .Q_N(_3388_),
    .Q(\vgademo.plane_du[2] ));
 sg13g2_dfrbp_1 _7322_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net69),
    .D(net487),
    .Q_N(_0050_),
    .Q(\vgademo.plane_du[3] ));
 sg13g2_dfrbp_1 _7323_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net68),
    .D(net560),
    .Q_N(_0049_),
    .Q(\vgademo.plane_du[4] ));
 sg13g2_dfrbp_1 _7324_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net67),
    .D(_0358_),
    .Q_N(_0051_),
    .Q(\vgademo.plane_du[5] ));
 sg13g2_dfrbp_1 _7325_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net66),
    .D(_0359_),
    .Q_N(_0052_),
    .Q(\vgademo.plane_du[6] ));
 sg13g2_dfrbp_1 _7326_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net65),
    .D(_0360_),
    .Q_N(_0053_),
    .Q(\vgademo.plane_du[7] ));
 sg13g2_dfrbp_1 _7327_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net64),
    .D(_0361_),
    .Q_N(_0054_),
    .Q(\vgademo.plane_du[8] ));
 sg13g2_dfrbp_1 _7328_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net63),
    .D(_0362_),
    .Q_N(_3387_),
    .Q(\vgademo.plane_du[9] ));
 sg13g2_dfrbp_1 _7329_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net62),
    .D(net414),
    .Q_N(_3386_),
    .Q(\vgademo.plane_du[10] ));
 sg13g2_dfrbp_1 _7330_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net35),
    .D(net260),
    .Q_N(_3385_),
    .Q(\vgademo.plane_u[0] ));
 sg13g2_tiehi _7261__16 (.L_HI(net16));
 sg13g2_tiehi _7046__17 (.L_HI(net17));
 sg13g2_tiehi _7260__18 (.L_HI(net18));
 sg13g2_tiehi _7045__19 (.L_HI(net19));
 sg13g2_tiehi _7259__20 (.L_HI(net20));
 sg13g2_tiehi _7044__21 (.L_HI(net21));
 sg13g2_tiehi _7258__22 (.L_HI(net22));
 sg13g2_tiehi _7043__23 (.L_HI(net23));
 sg13g2_tiehi _7257__24 (.L_HI(net24));
 sg13g2_tiehi _7042__25 (.L_HI(net25));
 sg13g2_tiehi _7256__26 (.L_HI(net26));
 sg13g2_tiehi _7041__27 (.L_HI(net27));
 sg13g2_tiehi _7255__28 (.L_HI(net28));
 sg13g2_tiehi _7040__29 (.L_HI(net29));
 sg13g2_tiehi _7254__30 (.L_HI(net30));
 sg13g2_tiehi _7039__31 (.L_HI(net31));
 sg13g2_tiehi _7253__32 (.L_HI(net32));
 sg13g2_tiehi _7038__33 (.L_HI(net33));
 sg13g2_tiehi _7072__34 (.L_HI(net34));
 sg13g2_tiehi _7330__35 (.L_HI(net35));
 sg13g2_tiehi _7222__36 (.L_HI(net36));
 sg13g2_tiehi _7221__37 (.L_HI(net37));
 sg13g2_tiehi _7185__38 (.L_HI(net38));
 sg13g2_tiehi _7184__39 (.L_HI(net39));
 sg13g2_tiehi _7183__40 (.L_HI(net40));
 sg13g2_tiehi _7182__41 (.L_HI(net41));
 sg13g2_tiehi _7181__42 (.L_HI(net42));
 sg13g2_tiehi _7180__43 (.L_HI(net43));
 sg13g2_tiehi _7179__44 (.L_HI(net44));
 sg13g2_tiehi _7178__45 (.L_HI(net45));
 sg13g2_tiehi _7177__46 (.L_HI(net46));
 sg13g2_tiehi _7176__47 (.L_HI(net47));
 sg13g2_tiehi _7175__48 (.L_HI(net48));
 sg13g2_tiehi _7174__49 (.L_HI(net49));
 sg13g2_tiehi _7173__50 (.L_HI(net50));
 sg13g2_tiehi _7172__51 (.L_HI(net51));
 sg13g2_tiehi _7171__52 (.L_HI(net52));
 sg13g2_tiehi _7170__53 (.L_HI(net53));
 sg13g2_tiehi _7169__54 (.L_HI(net54));
 sg13g2_tiehi _7168__55 (.L_HI(net55));
 sg13g2_tiehi _7167__56 (.L_HI(net56));
 sg13g2_tiehi _7166__57 (.L_HI(net57));
 sg13g2_tiehi _7165__58 (.L_HI(net58));
 sg13g2_tiehi _7164__59 (.L_HI(net59));
 sg13g2_tiehi _7163__60 (.L_HI(net60));
 sg13g2_tiehi _7162__61 (.L_HI(net61));
 sg13g2_tiehi _7329__62 (.L_HI(net62));
 sg13g2_tiehi _7328__63 (.L_HI(net63));
 sg13g2_tiehi _7327__64 (.L_HI(net64));
 sg13g2_tiehi _7326__65 (.L_HI(net65));
 sg13g2_tiehi _7325__66 (.L_HI(net66));
 sg13g2_tiehi _7324__67 (.L_HI(net67));
 sg13g2_tiehi _7323__68 (.L_HI(net68));
 sg13g2_tiehi _7322__69 (.L_HI(net69));
 sg13g2_tiehi _7144__70 (.L_HI(net70));
 sg13g2_tiehi _7143__71 (.L_HI(net71));
 sg13g2_tiehi _7142__72 (.L_HI(net72));
 sg13g2_tiehi _7141__73 (.L_HI(net73));
 sg13g2_tiehi _7140__74 (.L_HI(net74));
 sg13g2_tiehi _7139__75 (.L_HI(net75));
 sg13g2_tiehi _7138__76 (.L_HI(net76));
 sg13g2_tiehi _7137__77 (.L_HI(net77));
 sg13g2_tiehi _7136__78 (.L_HI(net78));
 sg13g2_tiehi _7135__79 (.L_HI(net79));
 sg13g2_tiehi _7186__80 (.L_HI(net80));
 sg13g2_tiehi _7187__81 (.L_HI(net81));
 sg13g2_tiehi _7188__82 (.L_HI(net82));
 sg13g2_tiehi _7134__83 (.L_HI(net83));
 sg13g2_tiehi _7133__84 (.L_HI(net84));
 sg13g2_tiehi _7132__85 (.L_HI(net85));
 sg13g2_tiehi _7131__86 (.L_HI(net86));
 sg13g2_tiehi _7321__87 (.L_HI(net87));
 sg13g2_tiehi _7320__88 (.L_HI(net88));
 sg13g2_tiehi _7319__89 (.L_HI(net89));
 sg13g2_tiehi _7318__90 (.L_HI(net90));
 sg13g2_tiehi _7317__91 (.L_HI(net91));
 sg13g2_tiehi _7316__92 (.L_HI(net92));
 sg13g2_tiehi _7315__93 (.L_HI(net93));
 sg13g2_tiehi _7314__94 (.L_HI(net94));
 sg13g2_tiehi _7313__95 (.L_HI(net95));
 sg13g2_tiehi _7312__96 (.L_HI(net96));
 sg13g2_tiehi _7311__97 (.L_HI(net97));
 sg13g2_tiehi _7310__98 (.L_HI(net98));
 sg13g2_tiehi _7309__99 (.L_HI(net99));
 sg13g2_tiehi _7308__100 (.L_HI(net100));
 sg13g2_tiehi _7307__101 (.L_HI(net101));
 sg13g2_tiehi _7306__102 (.L_HI(net102));
 sg13g2_tiehi _7305__103 (.L_HI(net103));
 sg13g2_tiehi _7304__104 (.L_HI(net104));
 sg13g2_tiehi _7303__105 (.L_HI(net105));
 sg13g2_tiehi _7302__106 (.L_HI(net106));
 sg13g2_tiehi _7301__107 (.L_HI(net107));
 sg13g2_tiehi _7300__108 (.L_HI(net108));
 sg13g2_tiehi _7299__109 (.L_HI(net109));
 sg13g2_tiehi _7298__110 (.L_HI(net110));
 sg13g2_tiehi _7297__111 (.L_HI(net111));
 sg13g2_tiehi _7296__112 (.L_HI(net112));
 sg13g2_tiehi _7103__113 (.L_HI(net113));
 sg13g2_tiehi _7295__114 (.L_HI(net114));
 sg13g2_tiehi _7294__115 (.L_HI(net115));
 sg13g2_tiehi _7071__116 (.L_HI(net116));
 sg13g2_tiehi _7293__117 (.L_HI(net117));
 sg13g2_tiehi _7070__118 (.L_HI(net118));
 sg13g2_tiehi _7292__119 (.L_HI(net119));
 sg13g2_tiehi _7069__120 (.L_HI(net120));
 sg13g2_tiehi _7291__121 (.L_HI(net121));
 sg13g2_tiehi _7068__122 (.L_HI(net122));
 sg13g2_tiehi _7290__123 (.L_HI(net123));
 sg13g2_tiehi _7067__124 (.L_HI(net124));
 sg13g2_tiehi _7289__125 (.L_HI(net125));
 sg13g2_tiehi _7066__126 (.L_HI(net126));
 sg13g2_tiehi _7288__127 (.L_HI(net127));
 sg13g2_tiehi _7065__128 (.L_HI(net128));
 sg13g2_tiehi _7287__129 (.L_HI(net129));
 sg13g2_tiehi _7064__130 (.L_HI(net130));
 sg13g2_tiehi _7286__131 (.L_HI(net131));
 sg13g2_tiehi _7063__132 (.L_HI(net132));
 sg13g2_tiehi _7285__133 (.L_HI(net133));
 sg13g2_tiehi _7062__134 (.L_HI(net134));
 sg13g2_tiehi _7284__135 (.L_HI(net135));
 sg13g2_tiehi _7061__136 (.L_HI(net136));
 sg13g2_tiehi _7283__137 (.L_HI(net137));
 sg13g2_tiehi _7060__138 (.L_HI(net138));
 sg13g2_tiehi _7282__139 (.L_HI(net139));
 sg13g2_tiehi _7059__140 (.L_HI(net140));
 sg13g2_tiehi _7281__141 (.L_HI(net141));
 sg13g2_tiehi _7280__142 (.L_HI(net142));
 sg13g2_tiehi _7279__143 (.L_HI(net143));
 sg13g2_tiehi _7278__144 (.L_HI(net144));
 sg13g2_tiehi _7277__145 (.L_HI(net145));
 sg13g2_tiehi _7276__146 (.L_HI(net146));
 sg13g2_tiehi _7275__147 (.L_HI(net147));
 sg13g2_tiehi _7274__148 (.L_HI(net148));
 sg13g2_tiehi _7273__149 (.L_HI(net149));
 sg13g2_tiehi _7272__150 (.L_HI(net150));
 sg13g2_tiehi _7271__151 (.L_HI(net151));
 sg13g2_tiehi _7270__152 (.L_HI(net152));
 sg13g2_tiehi _7269__153 (.L_HI(net153));
 sg13g2_tiehi _7268__154 (.L_HI(net154));
 sg13g2_tiehi _7267__155 (.L_HI(net155));
 sg13g2_tiehi _7266__156 (.L_HI(net156));
 sg13g2_tiehi _7265__157 (.L_HI(net157));
 sg13g2_tiehi _7050__158 (.L_HI(net158));
 sg13g2_tiehi _7264__159 (.L_HI(net159));
 sg13g2_tiehi _7049__160 (.L_HI(net160));
 sg13g2_tiehi _7263__161 (.L_HI(net161));
 sg13g2_tiehi _7048__162 (.L_HI(net162));
 sg13g2_tiehi _7262__163 (.L_HI(net163));
 sg13g2_tiehi tt_um_a1k0n_demo_164 (.L_HI(net164));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_a1k0n_demo_2 (.L_LO(net2));
 sg13g2_tielo tt_um_a1k0n_demo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_a1k0n_demo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_a1k0n_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_a1k0n_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_a1k0n_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_a1k0n_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_a1k0n_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_a1k0n_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_a1k0n_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_a1k0n_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_a1k0n_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_a1k0n_demo_14 (.L_LO(net14));
 sg13g2_tiehi _7047__15 (.L_HI(net15));
 sg13g2_buf_2 _7495_ (.A(audio),
    .X(uio_out[7]));
 sg13g2_buf_2 _7496_ (.A(\vgademo.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _7497_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout826 (.A(_1717_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_1683_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(net829),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_1652_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(net832),
    .X(net830));
 sg13g2_buf_1 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_1651_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net834),
    .X(net833));
 sg13g2_buf_1 fanout834 (.A(net835),
    .X(net834));
 sg13g2_buf_1 fanout835 (.A(_1492_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_2458_),
    .X(net837));
 sg13g2_buf_4 fanout838 (.X(net838),
    .A(_2314_));
 sg13g2_buf_2 fanout839 (.A(_1430_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_1430_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net843),
    .X(net841));
 sg13g2_buf_1 fanout842 (.A(net843),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_1428_),
    .X(net843));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(_1772_));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(_1348_));
 sg13g2_buf_2 fanout846 (.A(_1347_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_0699_),
    .X(net847));
 sg13g2_buf_1 fanout848 (.A(_0699_),
    .X(net848));
 sg13g2_buf_4 fanout849 (.X(net849),
    .A(net850));
 sg13g2_buf_2 fanout850 (.A(_0630_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_0625_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_1716_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_1715_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(net856),
    .X(net855));
 sg13g2_buf_1 fanout856 (.A(net857),
    .X(net856));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(_1315_));
 sg13g2_buf_2 fanout858 (.A(net859),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_1314_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_1294_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_1293_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_0859_),
    .X(net864));
 sg13g2_buf_4 fanout865 (.X(net865),
    .A(_0828_));
 sg13g2_buf_2 fanout866 (.A(net867),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_0827_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_0827_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_0573_),
    .X(net870));
 sg13g2_buf_1 fanout871 (.A(_0573_),
    .X(net871));
 sg13g2_buf_4 fanout872 (.X(net872),
    .A(net873));
 sg13g2_buf_4 fanout873 (.X(net873),
    .A(_0572_));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net876),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_2701_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(net880),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(net880),
    .X(net879));
 sg13g2_buf_4 fanout880 (.X(net880),
    .A(_2701_));
 sg13g2_buf_4 fanout881 (.X(net881),
    .A(_1208_));
 sg13g2_buf_2 fanout882 (.A(net883),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_0592_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_0592_),
    .X(net884));
 sg13g2_buf_1 fanout885 (.A(_0592_),
    .X(net885));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(net887));
 sg13g2_buf_4 fanout887 (.X(net887),
    .A(_2393_));
 sg13g2_buf_2 fanout888 (.A(_1362_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_0709_),
    .X(net889));
 sg13g2_buf_1 fanout890 (.A(_0709_),
    .X(net890));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(net894));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(net893));
 sg13g2_buf_2 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_0580_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(net899),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net898),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(net898),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(_2387_));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(_0662_));
 sg13g2_buf_2 fanout901 (.A(_0662_),
    .X(net901));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(_0661_));
 sg13g2_buf_2 fanout903 (.A(_0661_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_0644_),
    .X(net904));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(net908));
 sg13g2_buf_2 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(net908));
 sg13g2_buf_2 fanout908 (.A(_0591_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(net912),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_4 fanout912 (.X(net912),
    .A(_0590_));
 sg13g2_buf_2 fanout913 (.A(net915),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(net915),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_0589_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(net918),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net918),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_0579_),
    .X(net918));
 sg13g2_buf_4 fanout919 (.X(net919),
    .A(_0578_));
 sg13g2_buf_2 fanout920 (.A(_0578_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(net922),
    .X(net921));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(net928));
 sg13g2_buf_1 fanout923 (.A(net928),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net928),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(net928),
    .X(net925));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(net927));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(net928));
 sg13g2_buf_2 fanout928 (.A(_0577_),
    .X(net928));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(net930));
 sg13g2_buf_2 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(_0576_));
 sg13g2_buf_2 fanout933 (.A(_1052_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_1052_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_0659_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_0659_),
    .X(net936));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_0658_));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(net939));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_3199_),
    .X(net940));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(_3198_));
 sg13g2_buf_2 fanout942 (.A(_2223_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_0702_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_0701_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_0628_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_3098_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_3098_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_3096_),
    .X(net948));
 sg13g2_buf_4 fanout949 (.X(net949),
    .A(_3090_));
 sg13g2_buf_4 fanout950 (.X(net950),
    .A(net579));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(net952));
 sg13g2_buf_2 fanout952 (.A(net541),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(net955),
    .X(net953));
 sg13g2_buf_1 fanout954 (.A(net955),
    .X(net954));
 sg13g2_buf_4 fanout955 (.X(net955),
    .A(\vgademo.plane_dx_div.r[25] ));
 sg13g2_buf_4 fanout956 (.X(net956),
    .A(\vgademo.b_cos[10] ));
 sg13g2_buf_4 fanout957 (.X(net957),
    .A(\vgademo.b_cos[9] ));
 sg13g2_buf_4 fanout958 (.X(net958),
    .A(net574));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(\vgademo.b_cos[6] ));
 sg13g2_buf_4 fanout960 (.X(net960),
    .A(net961));
 sg13g2_buf_2 fanout961 (.A(\vgademo.a_sin[14] ),
    .X(net961));
 sg13g2_buf_4 fanout962 (.X(net962),
    .A(\vgademo.v_count[9] ));
 sg13g2_buf_2 fanout963 (.A(\vgademo.v_count[7] ),
    .X(net963));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(\vgademo.v_count[6] ));
 sg13g2_buf_2 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(\vgademo.v_count[5] ),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(net562),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(\vgademo.v_count[2] ),
    .X(net968));
 sg13g2_buf_4 fanout969 (.X(net969),
    .A(net554));
 sg13g2_buf_2 fanout970 (.A(net971),
    .X(net970));
 sg13g2_buf_4 fanout971 (.X(net971),
    .A(\vgademo.a_scrolly[10] ));
 sg13g2_buf_2 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(net975),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(net975),
    .X(net974));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(\vgademo.a_scrolly[9] ));
 sg13g2_buf_4 fanout976 (.X(net976),
    .A(net978));
 sg13g2_buf_2 fanout977 (.A(net978),
    .X(net977));
 sg13g2_buf_4 fanout978 (.X(net978),
    .A(\vgademo.a_scrolly[8] ));
 sg13g2_buf_4 fanout979 (.X(net979),
    .A(net980));
 sg13g2_buf_4 fanout980 (.X(net980),
    .A(net548));
 sg13g2_buf_4 fanout981 (.X(net981),
    .A(net983));
 sg13g2_buf_2 fanout982 (.A(net983),
    .X(net982));
 sg13g2_buf_4 fanout983 (.X(net983),
    .A(\vgademo.a_scrolly[6] ));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(net987));
 sg13g2_buf_2 fanout985 (.A(net987),
    .X(net985));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(net987));
 sg13g2_buf_2 fanout987 (.A(net584),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_4 fanout989 (.X(net989),
    .A(net990));
 sg13g2_buf_2 fanout990 (.A(net576),
    .X(net990));
 sg13g2_buf_4 fanout991 (.X(net991),
    .A(\vgademo.a_scrolly[3] ));
 sg13g2_buf_2 fanout992 (.A(\vgademo.a_scrolly[3] ),
    .X(net992));
 sg13g2_buf_4 fanout993 (.X(net993),
    .A(net994));
 sg13g2_buf_2 fanout994 (.A(net552),
    .X(net994));
 sg13g2_buf_4 fanout995 (.X(net995),
    .A(net592));
 sg13g2_buf_2 fanout996 (.A(\vgademo.h_count[6] ),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(\vgademo.h_count[5] ),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(net593),
    .X(net998));
 sg13g2_buf_1 fanout999 (.A(\vgademo.h_count[4] ),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(\vgademo.h_count[3] ),
    .X(net1000));
 sg13g2_buf_1 fanout1001 (.A(\vgademo.h_count[3] ),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(\vgademo.h_count[2] ),
    .X(net1002));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(net1004));
 sg13g2_buf_4 fanout1004 (.X(net1004),
    .A(\vgademo.h_count[1] ));
 sg13g2_buf_2 fanout1005 (.A(\vgademo.h_count[0] ),
    .X(net1005));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_buf_2 fanout1008 (.A(\vgademo.soundtrack.pulse_vol[3] ),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(\vgademo.soundtrack.pulse_vol[3] ),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(\vgademo.soundtrack.pulse_vol[2] ),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(\vgademo.soundtrack.pulse_vol[1] ),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(\vgademo.soundtrack.pulse_vol[0] ),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(net1015),
    .X(net1014));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(\vgademo.audio_snare_frames[3] ));
 sg13g2_buf_2 fanout1016 (.A(net1018),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_buf_4 fanout1019 (.X(net1019),
    .A(\vgademo.audio_snare_frames[2] ));
 sg13g2_buf_2 fanout1020 (.A(net1021),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_1 fanout1022 (.A(net1023),
    .X(net1022));
 sg13g2_buf_1 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(\vgademo.audio_snare_frames[1] ),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(net1027),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(net1028),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(\vgademo.audio_snare_frames[0] ),
    .X(net1028));
 sg13g2_buf_4 fanout1029 (.X(net1029),
    .A(net545));
 sg13g2_buf_2 fanout1030 (.A(net413),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(net1032),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net573),
    .X(net1032));
 sg13g2_buf_4 fanout1033 (.X(net1033),
    .A(net355));
 sg13g2_buf_2 fanout1034 (.A(net581),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(\vgademo.plane_dx_div.q[6] ),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(\vgademo.plane_dx_div.q[5] ),
    .X(net1036));
 sg13g2_buf_4 fanout1037 (.X(net1037),
    .A(net315));
 sg13g2_buf_2 fanout1038 (.A(\vgademo.plane_dx_div.q[4] ),
    .X(net1038));
 sg13g2_buf_4 fanout1039 (.X(net1039),
    .A(net559));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(\vgademo.plane_dx[1] ));
 sg13g2_buf_4 fanout1041 (.X(net1041),
    .A(\vgademo.audio_songpos[7] ));
 sg13g2_buf_2 fanout1042 (.A(\vgademo.audio_songpos[6] ),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(net1046),
    .X(net1043));
 sg13g2_buf_1 fanout1044 (.A(net1046),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(net1046),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(\vgademo.audio_songpos[5] ),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(net1048),
    .X(net1047));
 sg13g2_buf_1 fanout1048 (.A(net1050),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(net1050),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(\vgademo.audio_songpos[4] ),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1054),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(net1054),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(\vgademo.audio_songpos[3] ),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(net1057),
    .X(net1055));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(net1057));
 sg13g2_buf_2 fanout1057 (.A(\vgademo.audio_songpos[2] ),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net1060),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(net1061),
    .X(net1059));
 sg13g2_buf_1 fanout1060 (.A(net1061),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(\vgademo.audio_songpos[1] ),
    .X(net1061));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(net1063));
 sg13g2_buf_2 fanout1063 (.A(\vgademo.audio_songpos[0] ),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(\vgademo.linelfsr[1] ),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(\vgademo.linelfsr[1] ),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(net1067),
    .X(net1066));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(\vgademo.linelfsr[0] ));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(net1071));
 sg13g2_buf_4 fanout1069 (.X(net1069),
    .A(net1071));
 sg13g2_buf_2 fanout1070 (.A(net1071),
    .X(net1070));
 sg13g2_buf_4 fanout1071 (.X(net1071),
    .A(net1095));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(net1075));
 sg13g2_buf_4 fanout1073 (.X(net1073),
    .A(net1075));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(net1075));
 sg13g2_buf_2 fanout1075 (.A(net1095),
    .X(net1075));
 sg13g2_buf_4 fanout1076 (.X(net1076),
    .A(net1079));
 sg13g2_buf_4 fanout1077 (.X(net1077),
    .A(net1079));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(net1079));
 sg13g2_buf_4 fanout1079 (.X(net1079),
    .A(net1095));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1081));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(net1088));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(net1084));
 sg13g2_buf_2 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(net1088));
 sg13g2_buf_4 fanout1085 (.X(net1085),
    .A(net1087));
 sg13g2_buf_2 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_4 fanout1087 (.X(net1087),
    .A(net1088));
 sg13g2_buf_2 fanout1088 (.A(net1094),
    .X(net1088));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(net1090));
 sg13g2_buf_4 fanout1090 (.X(net1090),
    .A(net1094));
 sg13g2_buf_4 fanout1091 (.X(net1091),
    .A(net1092));
 sg13g2_buf_4 fanout1092 (.X(net1092),
    .A(net1093));
 sg13g2_buf_2 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(rst_n),
    .X(net1095));
 sg13g2_tielo tt_um_a1k0n_demo_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_2_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_47_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_40_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_41_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_43_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_3_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_12_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_13_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_15_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_35_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_37_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_16_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_23_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_24_clk));
 sg13g2_inv_2 clkload33 (.A(clknet_leaf_30_clk));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_31_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vgademo.soundtrack.sample_div_[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold2 (.A(\vgademo.soundtrack.noise_lfsr[1] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0169_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold4 (.A(\vgademo.soundtrack.noise_lfsr[3] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0171_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold6 (.A(\vgademo.soundtrack.noise_lfsr[10] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0178_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0084_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0142_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold10 (.A(\vgademo.soundtrack.noise_lfsr[2] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0170_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold12 (.A(\vgademo.soundtrack.noise_lfsr[12] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0180_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0082_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0176_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold16 (.A(\vgademo.soundtrack.tick_div_[0] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0161_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0081_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0181_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0083_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0174_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0099_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0179_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0102_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0184_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0089_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0092_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0131_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0090_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0103_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0185_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0087_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0105_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold34 (.A(\vgademo.soundtrack.tick_div[6] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0796_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0167_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold37 (.A(\vgademo.linelfsr[0] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0593_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0086_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0125_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold41 (.A(\vgademo.soundtrack.sample_div[4] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold42 (.A(\vgademo.soundtrack.sample_div_[4] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold43 (.A(\vgademo.soundtrack.sample_div[8] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold44 (.A(\vgademo.soundtrack.sample_div_[8] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold45 (.A(\vgademo.plane_dx_div.q[3] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0666_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0109_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0208_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0104_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0186_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0110_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold52 (.A(\vgademo.soundtrack.tick_div[4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0165_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold54 (.A(\vgademo.soundtrack.noise_lfsr[13] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0182_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold56 (.A(\vgademo.soundtrack.sample_div[0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold57 (.A(\vgademo.soundtrack.sample_div_[1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0096_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0172_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold60 (.A(\vgademo.soundtrack.pulse_osc_p[10] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0198_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0106_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0107_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold64 (.A(\vgademo.soundtrack.sigma_delta_accum[0] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold65 (.A(\vgademo.soundtrack.noise_lfsr[4] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0173_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold67 (.A(\vgademo.soundtrack.tick_div[3] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0164_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold69 (.A(\vgademo.soundtrack.pulse_osc_p[9] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0941_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0197_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold72 (.A(\vgademo.soundtrack.tri_osc_p[0] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0209_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold74 (.A(\vgademo.soundtrack.sample_div[7] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold75 (.A(\vgademo.soundtrack.sample_div_[7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold76 (.A(\vgademo.soundtrack.tick_div[2] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0163_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0108_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold79 (.A(\vgademo.soundtrack.pulse_osc_p[13] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0201_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold81 (.A(\vgademo.soundtrack.sample_div[3] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold82 (.A(\vgademo.soundtrack.sample_div_[3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold83 (.A(\vgademo.soundtrack.noise_lfsr[7] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0175_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold85 (.A(\vgademo.a_cos[0] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0257_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold87 (.A(\vgademo.soundtrack.pulse_osc_p[8] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0196_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold89 (.A(\vgademo.a_sin[0] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold90 (.A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0192_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0039_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0010_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold94 (.A(\vgademo.plane_u[0] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold95 (.A(_3077_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0364_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold97 (.A(audio),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0160_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold99 (.A(\vgademo.soundtrack.tick_div[5] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0166_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold101 (.A(\vgademo.soundtrack.pulse_osc_p[1] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0189_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold103 (.A(\vgademo.soundtrack.pulse_osc_p[11] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold104 (.A(\vgademo.soundtrack.sample_div[9] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold105 (.A(\vgademo.soundtrack.sample_div[5] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold106 (.A(\vgademo.soundtrack.tick_div[7] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold107 (.A(\vgademo.soundtrack.pulse_osc_p[0] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold108 (.A(\vgademo.plane_u[4] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0091_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold110 (.A(\vgademo.plane_dx_div.r[24] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0085_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0124_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0088_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold114 (.A(\vgademo.plane_dx_div.r[20] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0310_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold116 (.A(\vgademo.plane_du[0] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0353_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold118 (.A(\vgademo.plane_u[11] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0340_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold120 (.A(\vgademo.b_sin[5] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0323_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold122 (.A(\vgademo.soundtrack.tri_osc_p[10] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0219_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold124 (.A(\vgademo.a_sin[2] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold125 (.A(\vgademo.plane_u[8] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold126 (.A(\vgademo.plane_u[5] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold127 (.A(\vgademo.soundtrack.noise_lfsr[0] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0183_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0035_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0006_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold131 (.A(\vgademo.plane_u[1] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0330_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold133 (.A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0193_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold135 (.A(\vgademo.a_sin[1] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold136 (.A(\vgademo.soundtrack.noise_lfsr[8] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0177_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold138 (.A(\vgademo.linelfsr[5] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0116_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold140 (.A(\vgademo.b_sin[7] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0325_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold142 (.A(\vgademo.a_cos[2] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold143 (.A(\vgademo.plane_dx_div.d[24] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold144 (.A(\vgademo.b_cos[0] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0294_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold146 (.A(\vgademo.linelfsr[11] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0121_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold148 (.A(\vgademo.a_sin[4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold149 (.A(_2636_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0319_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold151 (.A(\vgademo.plane_dx_div.q[4] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold152 (.A(\vgademo.soundtrack.sigma_delta_accum[2] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold153 (.A(\vgademo.soundtrack.sigma_delta_accum_[3] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold154 (.A(\vgademo.soundtrack.tri_osc_p[13] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0222_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold156 (.A(\vgademo.soundtrack.pulse_osc_p[7] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold157 (.A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold158 (.A(\vgademo.audio_beat_out[0] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0146_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold160 (.A(\vgademo.a_cos[1] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0258_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold162 (.A(\vgademo.linelfsr[3] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0113_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold164 (.A(\vgademo.soundtrack.pulse_osc_p[2] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0190_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold166 (.A(\vgademo.soundtrack.tri_osc_p[1] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0210_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold168 (.A(\vgademo.plane_dx_div.i[0] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0654_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0143_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold171 (.A(\vgademo.plane_u[20] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold172 (.A(\vgademo.plane_dx_div.r[23] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold173 (.A(\vgademo.plane_du[1] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0354_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold175 (.A(\vgademo.plane_dx_div.d[23] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold176 (.A(\vgademo.plane_dx_div.r[16] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0306_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold178 (.A(\vgademo.plane_dx_div.d[22] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold179 (.A(\vgademo.b_cos[1] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0295_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold181 (.A(\vgademo.plane_dx_div.r[25] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0315_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold183 (.A(\vgademo.plane_dx_div.d[20] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold184 (.A(\vgademo.linelfsr[4] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold185 (.A(\vgademo.a_sin[5] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold186 (.A(_2641_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0320_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold188 (.A(\vgademo.soundtrack.pulse_osc_p[6] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0062_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0149_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold191 (.A(\vgademo.plane_dx_div.q[7] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0671_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold193 (.A(\vgademo.plane_u[6] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold194 (.A(\vgademo.plane_dx_div.r[18] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0308_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold196 (.A(\vgademo.plane_dx_div.r[22] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold197 (.A(\vgademo.plane_dx_div.d[19] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold198 (.A(\vgademo.scanline_audio_sample[2] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold199 (.A(\vgademo.plane_dx_div.r[21] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold200 (.A(\vgademo.plane_dx_div.d[18] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold201 (.A(\vgademo.plane_dx_div.r[19] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0034_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold203 (.A(_3203_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold204 (.A(\vgademo.audio_kick_frames[1] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold205 (.A(\vgademo.soundtrack.tri_osc_p[14] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0223_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold207 (.A(\vgademo.audio_beat_out[1] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0147_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold209 (.A(\vgademo.linelfsr[12] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold210 (.A(\vgademo.linelfsr[6] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0117_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold212 (.A(\vgademo.plane_u[2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold213 (.A(\vgademo.plane_u[7] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold214 (.A(\vgademo.audio_kick_frames[2] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold215 (.A(\vgademo.scanline_audio_sample[1] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold216 (.A(\vgademo.soundtrack.tri_osc_p[4] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold217 (.A(\vgademo.plane_u[3] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold218 (.A(\vgademo.a_sin[3] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold219 (.A(_2632_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0318_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold221 (.A(\vgademo.b_cos[3] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0297_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold223 (.A(\vgademo.plane_u[17] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0346_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0022_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold226 (.A(_1265_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0254_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold228 (.A(\vgademo.plane_dx_div.q[5] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0041_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold230 (.A(_1025_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0218_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold232 (.A(\vgademo.scanline_audio_sample[0] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold233 (.A(\vgademo.soundtrack.tri_osc_p[11] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold234 (.A(\vgademo.soundtrack.sigma_delta_accum[1] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold235 (.A(\vgademo.plane_u[9] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold236 (.A(\vgademo.soundtrack.tri_osc_p[3] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0212_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold238 (.A(\vgademo.linelfsr[9] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0120_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold240 (.A(\vgademo.plane_u[10] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold241 (.A(\vgademo.plane_dx_div.d[17] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold242 (.A(\vgademo.plane_u[13] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold243 (.A(\vgademo.b_cos[4] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0298_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold245 (.A(\vgademo.plane_u[16] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold246 (.A(_2946_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold247 (.A(\vgademo.soundtrack.tri_osc_p[2] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0211_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold249 (.A(\vgademo.plane_dx_div.q[9] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0363_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold251 (.A(\vgademo.bayer_j[1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold252 (.A(_1245_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0247_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold254 (.A(\vgademo.plane_dx_div.i[3] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0676_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold256 (.A(\vgademo.plane_u[12] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0341_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold258 (.A(\vgademo.soundtrack.tri_osc_p[5] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0214_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold260 (.A(\vgademo.soundtrack.tri_osc_p[7] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold261 (.A(\vgademo.scanline_audio_sample[5] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold262 (.A(\vgademo.linelfsr[7] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0118_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold264 (.A(\vgademo.soundtrack.tri_osc_p[6] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold265 (.A(\vgademo.b_cos[2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold266 (.A(_2405_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold267 (.A(\vgademo.soundtrack.tri_osc_p[12] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0224_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold269 (.A(\vgademo.a_sin[6] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold270 (.A(_2648_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0321_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold272 (.A(\vgademo.a_cos[3] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold273 (.A(\vgademo.a_cos[5] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold274 (.A(_2266_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold275 (.A(\vgademo.plane_du[2] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0355_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold277 (.A(\vgademo.a_scrolly[13] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold278 (.A(\vgademo.soundtrack.tri_osc_p[8] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold279 (.A(\vgademo.b_sin[4] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold280 (.A(_2653_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0322_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold282 (.A(\vgademo.plane_u[21] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0350_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold284 (.A(\vgademo.plane_u[19] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0348_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold286 (.A(\vgademo.b_cos[5] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold287 (.A(\vgademo.plane_dx_div.i[2] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0675_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0016_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold290 (.A(_1229_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold291 (.A(\vgademo.b_sin[6] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold292 (.A(_2667_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold293 (.A(\vgademo.plane_du[8] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold294 (.A(\vgademo.plane_u[14] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold295 (.A(\vgademo.a_cos[14] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold296 (.A(\vgademo.v_count[3] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0248_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold298 (.A(\vgademo.b_sin[10] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold299 (.A(_2693_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold300 (.A(\vgademo.plane_dx_div.d[21] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold301 (.A(\vgademo.plane_dx_div.d[16] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold302 (.A(\vgademo.soundtrack.sample_div[6] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold303 (.A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold304 (.A(\vgademo.scanline_audio_sample[6] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold305 (.A(\vgademo.a_sin[8] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0280_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold307 (.A(\vgademo.soundtrack.sample_div[2] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0565_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold309 (.A(\vgademo.soundtrack.sample_div_[2] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold310 (.A(\vgademo.b_sin[8] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold311 (.A(_2682_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0065_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0033_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold314 (.A(_3201_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold315 (.A(\vgademo.b_cos[11] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold316 (.A(\vgademo.soundtrack.tri_osc_i[2] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold317 (.A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold318 (.A(\vgademo.soundtrack.tick_div[1] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0795_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0162_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold321 (.A(\vgademo.scanline_audio_sample[4] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold322 (.A(\vgademo.plane_du[3] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0356_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold324 (.A(\vgademo.a_cos[10] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0301_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold326 (.A(\vgademo.audio_beat_out[4] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0689_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0150_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold329 (.A(\vgademo.linelfsr[8] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0063_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold331 (.A(_1253_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0015_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold333 (.A(_1259_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0252_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold335 (.A(\vgademo.v_count[8] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0253_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold337 (.A(\vgademo.a_sin[9] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold338 (.A(\vgademo.soundtrack.sigma_delta_accum[7] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold339 (.A(\vgademo.soundtrack.sigma_delta_accum_[7] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold340 (.A(\vgademo.plane_u[18] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold341 (.A(\vgademo.a_cos[4] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold342 (.A(\vgademo.linelfsr[2] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0112_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold344 (.A(\vgademo.plane_dx_div.r[17] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold345 (.A(\vgademo.a_sin[7] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold346 (.A(\vgademo.plane_dx[2] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0664_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold348 (.A(\vgademo.soundtrack.sigma_delta_accum[13] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold349 (.A(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold350 (.A(\vgademo.soundtrack.sigma_delta_accum[8] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold351 (.A(\vgademo.a_cos[12] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0303_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0067_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold354 (.A(_1235_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0243_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold356 (.A(\vgademo.soundtrack.sigma_delta_accum[9] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold357 (.A(\vgademo.a_sin[10] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold358 (.A(\vgademo.soundtrack.sigma_delta_accum[12] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold359 (.A(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold360 (.A(\vgademo.soundtrack.tri_osc_i[4] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold361 (.A(\vgademo.a_cos[6] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0263_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold363 (.A(\vgademo.a_scrolly[11] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0242_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold365 (.A(\vgademo.soundtrack.sigma_delta_accum[11] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold366 (.A(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold367 (.A(\vgademo.a_sin[11] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold368 (.A(\vgademo.a_cos[11] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold369 (.A(\vgademo.soundtrack.sigma_delta_accum[10] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0017_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold371 (.A(_1257_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0251_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold373 (.A(\vgademo.b_sin[9] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold374 (.A(_2688_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold375 (.A(\vgademo.bayer_j[1] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold376 (.A(\vgademo.plane_u[15] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold377 (.A(\vgademo.b_sin[11] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0329_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold379 (.A(\vgademo.soundtrack.pulse_osc_p[12] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold380 (.A(\vgademo.a_sin[12] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold381 (.A(\vgademo.audio_beat_out[2] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold382 (.A(\vgademo.soundtrack.sigma_delta_accum[6] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold383 (.A(\vgademo.soundtrack.sigma_delta_accum_[6] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold384 (.A(\vgademo.a_scrolly[7] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0238_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold386 (.A(\vgademo.soundtrack.sigma_delta_accum[4] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold387 (.A(\vgademo.soundtrack.sigma_delta_accum_[4] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold388 (.A(\vgademo.a_scrolly[3] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold389 (.A(\vgademo.plane_dx[3] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold390 (.A(\vgademo.bayer_j[0] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0037_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold392 (.A(_3212_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0008_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold394 (.A(\vgademo.soundtrack.tri_osc_i[3] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0024_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0357_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold397 (.A(\vgademo.a_sin[13] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold398 (.A(\vgademo.v_count[4] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0077_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold400 (.A(\vgademo.plane_dx[0] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0132_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold402 (.A(\vgademo.soundtrack.sigma_delta_accum[5] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold403 (.A(\vgademo.a_cos[7] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold404 (.A(\vgademo.a_cos[9] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold405 (.A(_2427_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold406 (.A(\vgademo.a_cos[8] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold407 (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold408 (.A(\vgademo.soundtrack.sigma_delta_accum[14] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold409 (.A(\vgademo.plane_dx_div.q[8] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold410 (.A(\vgademo.b_cos[8] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold411 (.A(\vgademo.scanline_audio_sample[3] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold412 (.A(\vgademo.a_scrolly[4] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0038_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold414 (.A(\vgademo.plane_du[5] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold415 (.A(\vgademo.plane_du[9] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold416 (.A(\vgademo.a_cos[13] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold417 (.A(\vgademo.plane_dx_div.q[6] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold418 (.A(\vgademo.soundtrack.sigma_delta_accum[15] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold419 (.A(\vgademo.audio_kick_frames[0] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold420 (.A(\vgademo.a_scrolly[5] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0080_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold422 (.A(_1223_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold423 (.A(\vgademo.soundtrack.tri_osc_i[8] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold424 (.A(\vgademo.plane_du[7] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0036_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold426 (.A(_3209_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0007_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0061_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold429 (.A(\vgademo.h_count[4] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold430 (.A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0075_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0237_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold433 (.A(\vgademo.plane_du[6] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold434 (.A(\vgademo.soundtrack.tri_osc_i[6] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold435 (.A(\vgademo.soundtrack.tick_div[7] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold436 (.A(\vgademo.a_sin[1] ),
    .X(net600));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_4 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_264 ();
 sg13g2_decap_8 FILLER_13_271 ();
 sg13g2_decap_8 FILLER_13_278 ();
 sg13g2_decap_8 FILLER_13_285 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_decap_8 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_8 FILLER_13_404 ();
 sg13g2_decap_8 FILLER_13_411 ();
 sg13g2_decap_8 FILLER_13_418 ();
 sg13g2_decap_8 FILLER_13_425 ();
 sg13g2_decap_8 FILLER_13_432 ();
 sg13g2_decap_8 FILLER_13_439 ();
 sg13g2_decap_8 FILLER_13_446 ();
 sg13g2_decap_8 FILLER_13_453 ();
 sg13g2_decap_8 FILLER_13_460 ();
 sg13g2_decap_8 FILLER_13_467 ();
 sg13g2_decap_8 FILLER_13_474 ();
 sg13g2_decap_8 FILLER_13_481 ();
 sg13g2_decap_8 FILLER_13_488 ();
 sg13g2_decap_8 FILLER_13_495 ();
 sg13g2_decap_8 FILLER_13_502 ();
 sg13g2_decap_8 FILLER_13_509 ();
 sg13g2_decap_8 FILLER_13_516 ();
 sg13g2_decap_8 FILLER_13_523 ();
 sg13g2_decap_8 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_537 ();
 sg13g2_decap_8 FILLER_13_544 ();
 sg13g2_decap_8 FILLER_13_551 ();
 sg13g2_decap_8 FILLER_13_558 ();
 sg13g2_decap_8 FILLER_13_565 ();
 sg13g2_decap_8 FILLER_13_572 ();
 sg13g2_decap_8 FILLER_13_579 ();
 sg13g2_decap_8 FILLER_13_586 ();
 sg13g2_decap_8 FILLER_13_593 ();
 sg13g2_decap_8 FILLER_13_600 ();
 sg13g2_decap_8 FILLER_13_607 ();
 sg13g2_decap_8 FILLER_13_614 ();
 sg13g2_decap_8 FILLER_13_621 ();
 sg13g2_decap_8 FILLER_13_628 ();
 sg13g2_decap_8 FILLER_13_635 ();
 sg13g2_decap_8 FILLER_13_642 ();
 sg13g2_decap_8 FILLER_13_649 ();
 sg13g2_decap_8 FILLER_13_656 ();
 sg13g2_decap_8 FILLER_13_663 ();
 sg13g2_decap_8 FILLER_13_670 ();
 sg13g2_decap_8 FILLER_13_677 ();
 sg13g2_decap_8 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_691 ();
 sg13g2_decap_8 FILLER_13_698 ();
 sg13g2_decap_8 FILLER_13_705 ();
 sg13g2_decap_8 FILLER_13_712 ();
 sg13g2_decap_8 FILLER_13_719 ();
 sg13g2_decap_8 FILLER_13_726 ();
 sg13g2_decap_8 FILLER_13_733 ();
 sg13g2_decap_8 FILLER_13_740 ();
 sg13g2_decap_8 FILLER_13_747 ();
 sg13g2_decap_8 FILLER_13_754 ();
 sg13g2_decap_8 FILLER_13_761 ();
 sg13g2_decap_8 FILLER_13_768 ();
 sg13g2_decap_8 FILLER_13_775 ();
 sg13g2_decap_8 FILLER_13_782 ();
 sg13g2_decap_8 FILLER_13_789 ();
 sg13g2_decap_8 FILLER_13_796 ();
 sg13g2_decap_8 FILLER_13_803 ();
 sg13g2_decap_8 FILLER_13_810 ();
 sg13g2_decap_8 FILLER_13_817 ();
 sg13g2_decap_8 FILLER_13_824 ();
 sg13g2_decap_8 FILLER_13_831 ();
 sg13g2_decap_8 FILLER_13_838 ();
 sg13g2_decap_8 FILLER_13_845 ();
 sg13g2_decap_8 FILLER_13_852 ();
 sg13g2_fill_2 FILLER_13_859 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_fill_2 FILLER_14_70 ();
 sg13g2_fill_1 FILLER_14_72 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_4 FILLER_14_210 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_223 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_260 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_4 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_decap_4 FILLER_14_307 ();
 sg13g2_fill_2 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_92 ();
 sg13g2_decap_4 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_117 ();
 sg13g2_decap_8 FILLER_15_124 ();
 sg13g2_decap_8 FILLER_15_131 ();
 sg13g2_decap_8 FILLER_15_138 ();
 sg13g2_decap_8 FILLER_15_145 ();
 sg13g2_decap_8 FILLER_15_152 ();
 sg13g2_fill_2 FILLER_15_159 ();
 sg13g2_fill_2 FILLER_15_191 ();
 sg13g2_fill_1 FILLER_15_193 ();
 sg13g2_decap_4 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_fill_2 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_348 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_fill_2 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_fill_2 FILLER_15_383 ();
 sg13g2_fill_1 FILLER_15_385 ();
 sg13g2_decap_4 FILLER_15_399 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_15_414 ();
 sg13g2_fill_1 FILLER_15_421 ();
 sg13g2_decap_8 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_15_433 ();
 sg13g2_decap_8 FILLER_15_440 ();
 sg13g2_decap_8 FILLER_15_447 ();
 sg13g2_decap_8 FILLER_15_454 ();
 sg13g2_decap_8 FILLER_15_461 ();
 sg13g2_decap_8 FILLER_15_468 ();
 sg13g2_decap_8 FILLER_15_475 ();
 sg13g2_decap_8 FILLER_15_482 ();
 sg13g2_decap_8 FILLER_15_489 ();
 sg13g2_decap_8 FILLER_15_496 ();
 sg13g2_decap_8 FILLER_15_503 ();
 sg13g2_decap_8 FILLER_15_510 ();
 sg13g2_decap_8 FILLER_15_517 ();
 sg13g2_decap_8 FILLER_15_524 ();
 sg13g2_decap_8 FILLER_15_531 ();
 sg13g2_decap_8 FILLER_15_538 ();
 sg13g2_decap_8 FILLER_15_545 ();
 sg13g2_decap_8 FILLER_15_552 ();
 sg13g2_decap_8 FILLER_15_559 ();
 sg13g2_decap_8 FILLER_15_566 ();
 sg13g2_decap_8 FILLER_15_573 ();
 sg13g2_decap_8 FILLER_15_580 ();
 sg13g2_decap_8 FILLER_15_587 ();
 sg13g2_decap_8 FILLER_15_594 ();
 sg13g2_decap_8 FILLER_15_601 ();
 sg13g2_decap_8 FILLER_15_608 ();
 sg13g2_decap_8 FILLER_15_615 ();
 sg13g2_decap_8 FILLER_15_622 ();
 sg13g2_decap_8 FILLER_15_629 ();
 sg13g2_decap_8 FILLER_15_636 ();
 sg13g2_decap_8 FILLER_15_643 ();
 sg13g2_decap_8 FILLER_15_650 ();
 sg13g2_decap_8 FILLER_15_657 ();
 sg13g2_decap_8 FILLER_15_664 ();
 sg13g2_decap_8 FILLER_15_671 ();
 sg13g2_decap_8 FILLER_15_678 ();
 sg13g2_decap_8 FILLER_15_685 ();
 sg13g2_decap_8 FILLER_15_692 ();
 sg13g2_decap_8 FILLER_15_699 ();
 sg13g2_decap_8 FILLER_15_706 ();
 sg13g2_decap_8 FILLER_15_713 ();
 sg13g2_decap_8 FILLER_15_720 ();
 sg13g2_decap_8 FILLER_15_727 ();
 sg13g2_decap_8 FILLER_15_734 ();
 sg13g2_decap_8 FILLER_15_741 ();
 sg13g2_decap_8 FILLER_15_748 ();
 sg13g2_decap_8 FILLER_15_755 ();
 sg13g2_decap_8 FILLER_15_762 ();
 sg13g2_decap_8 FILLER_15_769 ();
 sg13g2_decap_8 FILLER_15_776 ();
 sg13g2_decap_8 FILLER_15_783 ();
 sg13g2_decap_8 FILLER_15_790 ();
 sg13g2_decap_8 FILLER_15_797 ();
 sg13g2_decap_8 FILLER_15_804 ();
 sg13g2_decap_8 FILLER_15_811 ();
 sg13g2_decap_8 FILLER_15_818 ();
 sg13g2_decap_8 FILLER_15_825 ();
 sg13g2_decap_8 FILLER_15_832 ();
 sg13g2_decap_8 FILLER_15_839 ();
 sg13g2_decap_8 FILLER_15_846 ();
 sg13g2_decap_8 FILLER_15_853 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_47 ();
 sg13g2_fill_2 FILLER_16_83 ();
 sg13g2_fill_2 FILLER_16_99 ();
 sg13g2_decap_4 FILLER_16_135 ();
 sg13g2_fill_2 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_193 ();
 sg13g2_fill_2 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_227 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_250 ();
 sg13g2_fill_1 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_257 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_293 ();
 sg13g2_fill_2 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_fill_1 FILLER_16_316 ();
 sg13g2_fill_1 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_370 ();
 sg13g2_decap_4 FILLER_16_375 ();
 sg13g2_fill_2 FILLER_16_405 ();
 sg13g2_fill_1 FILLER_16_407 ();
 sg13g2_fill_2 FILLER_16_438 ();
 sg13g2_fill_1 FILLER_16_445 ();
 sg13g2_fill_1 FILLER_16_458 ();
 sg13g2_decap_8 FILLER_16_472 ();
 sg13g2_decap_8 FILLER_16_479 ();
 sg13g2_decap_8 FILLER_16_486 ();
 sg13g2_decap_8 FILLER_16_493 ();
 sg13g2_fill_1 FILLER_16_500 ();
 sg13g2_decap_8 FILLER_16_521 ();
 sg13g2_decap_8 FILLER_16_528 ();
 sg13g2_decap_8 FILLER_16_535 ();
 sg13g2_decap_8 FILLER_16_542 ();
 sg13g2_decap_8 FILLER_16_549 ();
 sg13g2_decap_8 FILLER_16_556 ();
 sg13g2_decap_8 FILLER_16_563 ();
 sg13g2_decap_8 FILLER_16_570 ();
 sg13g2_decap_8 FILLER_16_577 ();
 sg13g2_decap_8 FILLER_16_584 ();
 sg13g2_decap_8 FILLER_16_591 ();
 sg13g2_decap_8 FILLER_16_598 ();
 sg13g2_decap_8 FILLER_16_605 ();
 sg13g2_decap_8 FILLER_16_612 ();
 sg13g2_decap_8 FILLER_16_619 ();
 sg13g2_decap_8 FILLER_16_626 ();
 sg13g2_decap_8 FILLER_16_633 ();
 sg13g2_decap_8 FILLER_16_640 ();
 sg13g2_decap_8 FILLER_16_647 ();
 sg13g2_decap_8 FILLER_16_654 ();
 sg13g2_decap_8 FILLER_16_661 ();
 sg13g2_decap_8 FILLER_16_668 ();
 sg13g2_decap_8 FILLER_16_675 ();
 sg13g2_decap_8 FILLER_16_682 ();
 sg13g2_decap_8 FILLER_16_689 ();
 sg13g2_decap_8 FILLER_16_696 ();
 sg13g2_decap_8 FILLER_16_703 ();
 sg13g2_decap_8 FILLER_16_710 ();
 sg13g2_decap_8 FILLER_16_717 ();
 sg13g2_decap_8 FILLER_16_724 ();
 sg13g2_decap_8 FILLER_16_731 ();
 sg13g2_decap_8 FILLER_16_738 ();
 sg13g2_decap_8 FILLER_16_745 ();
 sg13g2_decap_8 FILLER_16_752 ();
 sg13g2_decap_8 FILLER_16_759 ();
 sg13g2_decap_8 FILLER_16_766 ();
 sg13g2_decap_8 FILLER_16_773 ();
 sg13g2_decap_8 FILLER_16_780 ();
 sg13g2_decap_8 FILLER_16_787 ();
 sg13g2_decap_8 FILLER_16_794 ();
 sg13g2_decap_8 FILLER_16_801 ();
 sg13g2_decap_8 FILLER_16_808 ();
 sg13g2_decap_8 FILLER_16_815 ();
 sg13g2_decap_8 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_16_829 ();
 sg13g2_decap_8 FILLER_16_836 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_850 ();
 sg13g2_decap_4 FILLER_16_857 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_4 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_32 ();
 sg13g2_decap_8 FILLER_17_110 ();
 sg13g2_fill_2 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_decap_4 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_128 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_146 ();
 sg13g2_decap_4 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_fill_2 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_286 ();
 sg13g2_fill_2 FILLER_17_383 ();
 sg13g2_fill_2 FILLER_17_432 ();
 sg13g2_fill_1 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_478 ();
 sg13g2_decap_8 FILLER_17_485 ();
 sg13g2_fill_2 FILLER_17_492 ();
 sg13g2_fill_2 FILLER_17_499 ();
 sg13g2_fill_1 FILLER_17_522 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_18 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_fill_1 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_74 ();
 sg13g2_fill_1 FILLER_18_76 ();
 sg13g2_fill_2 FILLER_18_82 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_131 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_fill_2 FILLER_18_207 ();
 sg13g2_fill_1 FILLER_18_209 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_330 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_376 ();
 sg13g2_fill_2 FILLER_18_412 ();
 sg13g2_fill_1 FILLER_18_466 ();
 sg13g2_fill_1 FILLER_18_510 ();
 sg13g2_decap_8 FILLER_18_542 ();
 sg13g2_decap_8 FILLER_18_549 ();
 sg13g2_decap_8 FILLER_18_556 ();
 sg13g2_decap_8 FILLER_18_563 ();
 sg13g2_decap_8 FILLER_18_570 ();
 sg13g2_decap_8 FILLER_18_577 ();
 sg13g2_decap_8 FILLER_18_584 ();
 sg13g2_decap_8 FILLER_18_591 ();
 sg13g2_decap_8 FILLER_18_598 ();
 sg13g2_decap_8 FILLER_18_605 ();
 sg13g2_decap_8 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_633 ();
 sg13g2_decap_8 FILLER_18_640 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_decap_8 FILLER_18_654 ();
 sg13g2_decap_8 FILLER_18_661 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_decap_8 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_696 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_decap_8 FILLER_18_710 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_decap_8 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_decap_8 FILLER_18_738 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_780 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_decap_8 FILLER_18_850 ();
 sg13g2_decap_4 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_58 ();
 sg13g2_fill_1 FILLER_19_60 ();
 sg13g2_decap_4 FILLER_19_82 ();
 sg13g2_fill_2 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_fill_2 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_117 ();
 sg13g2_decap_4 FILLER_19_178 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_decap_4 FILLER_19_193 ();
 sg13g2_fill_1 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_decap_4 FILLER_19_227 ();
 sg13g2_fill_1 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_237 ();
 sg13g2_fill_1 FILLER_19_239 ();
 sg13g2_decap_4 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_264 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_fill_2 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_fill_1 FILLER_19_397 ();
 sg13g2_fill_2 FILLER_19_412 ();
 sg13g2_fill_2 FILLER_19_527 ();
 sg13g2_decap_8 FILLER_19_545 ();
 sg13g2_decap_8 FILLER_19_552 ();
 sg13g2_decap_8 FILLER_19_559 ();
 sg13g2_decap_8 FILLER_19_566 ();
 sg13g2_decap_8 FILLER_19_573 ();
 sg13g2_decap_8 FILLER_19_580 ();
 sg13g2_decap_8 FILLER_19_587 ();
 sg13g2_decap_8 FILLER_19_594 ();
 sg13g2_decap_8 FILLER_19_601 ();
 sg13g2_decap_8 FILLER_19_608 ();
 sg13g2_decap_8 FILLER_19_615 ();
 sg13g2_decap_8 FILLER_19_622 ();
 sg13g2_decap_8 FILLER_19_629 ();
 sg13g2_decap_8 FILLER_19_636 ();
 sg13g2_decap_8 FILLER_19_643 ();
 sg13g2_decap_8 FILLER_19_650 ();
 sg13g2_decap_8 FILLER_19_657 ();
 sg13g2_decap_8 FILLER_19_664 ();
 sg13g2_decap_8 FILLER_19_671 ();
 sg13g2_decap_8 FILLER_19_678 ();
 sg13g2_decap_8 FILLER_19_685 ();
 sg13g2_decap_8 FILLER_19_692 ();
 sg13g2_decap_8 FILLER_19_699 ();
 sg13g2_decap_8 FILLER_19_706 ();
 sg13g2_decap_8 FILLER_19_713 ();
 sg13g2_decap_8 FILLER_19_720 ();
 sg13g2_decap_8 FILLER_19_727 ();
 sg13g2_decap_8 FILLER_19_734 ();
 sg13g2_decap_8 FILLER_19_741 ();
 sg13g2_decap_8 FILLER_19_748 ();
 sg13g2_decap_8 FILLER_19_755 ();
 sg13g2_decap_8 FILLER_19_762 ();
 sg13g2_decap_8 FILLER_19_769 ();
 sg13g2_decap_8 FILLER_19_776 ();
 sg13g2_decap_8 FILLER_19_783 ();
 sg13g2_decap_8 FILLER_19_790 ();
 sg13g2_decap_8 FILLER_19_797 ();
 sg13g2_decap_8 FILLER_19_804 ();
 sg13g2_decap_8 FILLER_19_811 ();
 sg13g2_decap_8 FILLER_19_818 ();
 sg13g2_decap_8 FILLER_19_825 ();
 sg13g2_decap_8 FILLER_19_832 ();
 sg13g2_decap_8 FILLER_19_839 ();
 sg13g2_decap_8 FILLER_19_846 ();
 sg13g2_decap_8 FILLER_19_853 ();
 sg13g2_fill_2 FILLER_19_860 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_18 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_fill_1 FILLER_20_56 ();
 sg13g2_fill_1 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_106 ();
 sg13g2_decap_8 FILLER_20_113 ();
 sg13g2_decap_8 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_decap_4 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_decap_4 FILLER_20_223 ();
 sg13g2_fill_2 FILLER_20_227 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_fill_1 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_357 ();
 sg13g2_decap_4 FILLER_20_373 ();
 sg13g2_decap_4 FILLER_20_467 ();
 sg13g2_fill_2 FILLER_20_471 ();
 sg13g2_fill_1 FILLER_20_483 ();
 sg13g2_fill_1 FILLER_20_515 ();
 sg13g2_decap_8 FILLER_20_542 ();
 sg13g2_decap_8 FILLER_20_549 ();
 sg13g2_decap_8 FILLER_20_556 ();
 sg13g2_decap_8 FILLER_20_563 ();
 sg13g2_decap_8 FILLER_20_570 ();
 sg13g2_decap_8 FILLER_20_577 ();
 sg13g2_decap_8 FILLER_20_584 ();
 sg13g2_decap_8 FILLER_20_591 ();
 sg13g2_decap_8 FILLER_20_598 ();
 sg13g2_decap_8 FILLER_20_605 ();
 sg13g2_decap_8 FILLER_20_612 ();
 sg13g2_decap_8 FILLER_20_619 ();
 sg13g2_decap_8 FILLER_20_626 ();
 sg13g2_decap_8 FILLER_20_633 ();
 sg13g2_decap_8 FILLER_20_640 ();
 sg13g2_decap_8 FILLER_20_647 ();
 sg13g2_decap_8 FILLER_20_654 ();
 sg13g2_decap_8 FILLER_20_661 ();
 sg13g2_decap_8 FILLER_20_668 ();
 sg13g2_decap_8 FILLER_20_675 ();
 sg13g2_decap_8 FILLER_20_682 ();
 sg13g2_decap_8 FILLER_20_689 ();
 sg13g2_decap_8 FILLER_20_696 ();
 sg13g2_decap_8 FILLER_20_703 ();
 sg13g2_decap_8 FILLER_20_710 ();
 sg13g2_decap_8 FILLER_20_717 ();
 sg13g2_decap_8 FILLER_20_724 ();
 sg13g2_decap_8 FILLER_20_731 ();
 sg13g2_decap_8 FILLER_20_738 ();
 sg13g2_decap_8 FILLER_20_745 ();
 sg13g2_decap_8 FILLER_20_752 ();
 sg13g2_decap_8 FILLER_20_759 ();
 sg13g2_decap_8 FILLER_20_766 ();
 sg13g2_decap_8 FILLER_20_773 ();
 sg13g2_decap_8 FILLER_20_780 ();
 sg13g2_decap_8 FILLER_20_787 ();
 sg13g2_decap_8 FILLER_20_794 ();
 sg13g2_decap_8 FILLER_20_801 ();
 sg13g2_decap_8 FILLER_20_808 ();
 sg13g2_decap_8 FILLER_20_815 ();
 sg13g2_decap_8 FILLER_20_822 ();
 sg13g2_decap_8 FILLER_20_829 ();
 sg13g2_decap_8 FILLER_20_836 ();
 sg13g2_decap_8 FILLER_20_843 ();
 sg13g2_decap_8 FILLER_20_850 ();
 sg13g2_decap_4 FILLER_20_857 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_75 ();
 sg13g2_decap_8 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_decap_8 FILLER_21_155 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_181 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_4 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_246 ();
 sg13g2_fill_1 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_334 ();
 sg13g2_decap_4 FILLER_21_347 ();
 sg13g2_fill_1 FILLER_21_351 ();
 sg13g2_fill_1 FILLER_21_395 ();
 sg13g2_fill_1 FILLER_21_405 ();
 sg13g2_fill_2 FILLER_21_411 ();
 sg13g2_fill_1 FILLER_21_413 ();
 sg13g2_decap_4 FILLER_21_433 ();
 sg13g2_fill_2 FILLER_21_437 ();
 sg13g2_fill_2 FILLER_21_502 ();
 sg13g2_fill_1 FILLER_21_504 ();
 sg13g2_fill_1 FILLER_21_519 ();
 sg13g2_fill_1 FILLER_21_529 ();
 sg13g2_decap_8 FILLER_21_544 ();
 sg13g2_decap_8 FILLER_21_551 ();
 sg13g2_decap_8 FILLER_21_558 ();
 sg13g2_decap_8 FILLER_21_565 ();
 sg13g2_decap_8 FILLER_21_572 ();
 sg13g2_decap_8 FILLER_21_579 ();
 sg13g2_decap_8 FILLER_21_586 ();
 sg13g2_decap_8 FILLER_21_593 ();
 sg13g2_decap_8 FILLER_21_600 ();
 sg13g2_decap_8 FILLER_21_607 ();
 sg13g2_decap_8 FILLER_21_614 ();
 sg13g2_decap_8 FILLER_21_621 ();
 sg13g2_decap_8 FILLER_21_628 ();
 sg13g2_decap_8 FILLER_21_635 ();
 sg13g2_decap_8 FILLER_21_642 ();
 sg13g2_decap_8 FILLER_21_649 ();
 sg13g2_decap_8 FILLER_21_656 ();
 sg13g2_decap_8 FILLER_21_663 ();
 sg13g2_decap_8 FILLER_21_670 ();
 sg13g2_decap_8 FILLER_21_677 ();
 sg13g2_decap_8 FILLER_21_684 ();
 sg13g2_decap_8 FILLER_21_691 ();
 sg13g2_decap_8 FILLER_21_698 ();
 sg13g2_decap_8 FILLER_21_705 ();
 sg13g2_decap_8 FILLER_21_712 ();
 sg13g2_decap_8 FILLER_21_719 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_733 ();
 sg13g2_decap_8 FILLER_21_740 ();
 sg13g2_decap_8 FILLER_21_747 ();
 sg13g2_decap_8 FILLER_21_754 ();
 sg13g2_decap_8 FILLER_21_761 ();
 sg13g2_decap_8 FILLER_21_768 ();
 sg13g2_decap_8 FILLER_21_775 ();
 sg13g2_decap_8 FILLER_21_782 ();
 sg13g2_decap_8 FILLER_21_789 ();
 sg13g2_decap_8 FILLER_21_796 ();
 sg13g2_decap_8 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_810 ();
 sg13g2_decap_8 FILLER_21_817 ();
 sg13g2_decap_8 FILLER_21_824 ();
 sg13g2_decap_8 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_838 ();
 sg13g2_decap_8 FILLER_21_845 ();
 sg13g2_decap_8 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_859 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_16 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_4 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_185 ();
 sg13g2_fill_2 FILLER_22_192 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_decap_4 FILLER_22_208 ();
 sg13g2_fill_2 FILLER_22_212 ();
 sg13g2_decap_4 FILLER_22_227 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_fill_1 FILLER_22_317 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_decap_4 FILLER_22_364 ();
 sg13g2_fill_1 FILLER_22_373 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_fill_1 FILLER_22_394 ();
 sg13g2_decap_4 FILLER_22_415 ();
 sg13g2_decap_4 FILLER_22_473 ();
 sg13g2_fill_2 FILLER_22_477 ();
 sg13g2_decap_8 FILLER_22_545 ();
 sg13g2_decap_8 FILLER_22_552 ();
 sg13g2_decap_8 FILLER_22_559 ();
 sg13g2_decap_8 FILLER_22_566 ();
 sg13g2_decap_8 FILLER_22_573 ();
 sg13g2_decap_8 FILLER_22_580 ();
 sg13g2_decap_8 FILLER_22_587 ();
 sg13g2_decap_8 FILLER_22_594 ();
 sg13g2_decap_8 FILLER_22_601 ();
 sg13g2_decap_8 FILLER_22_608 ();
 sg13g2_decap_8 FILLER_22_615 ();
 sg13g2_decap_8 FILLER_22_622 ();
 sg13g2_decap_8 FILLER_22_629 ();
 sg13g2_decap_8 FILLER_22_636 ();
 sg13g2_decap_8 FILLER_22_643 ();
 sg13g2_decap_8 FILLER_22_650 ();
 sg13g2_decap_8 FILLER_22_657 ();
 sg13g2_decap_8 FILLER_22_664 ();
 sg13g2_decap_8 FILLER_22_671 ();
 sg13g2_decap_8 FILLER_22_678 ();
 sg13g2_decap_8 FILLER_22_685 ();
 sg13g2_decap_8 FILLER_22_692 ();
 sg13g2_decap_8 FILLER_22_699 ();
 sg13g2_decap_8 FILLER_22_706 ();
 sg13g2_decap_8 FILLER_22_713 ();
 sg13g2_decap_8 FILLER_22_720 ();
 sg13g2_decap_8 FILLER_22_727 ();
 sg13g2_decap_8 FILLER_22_734 ();
 sg13g2_decap_8 FILLER_22_741 ();
 sg13g2_decap_8 FILLER_22_748 ();
 sg13g2_decap_8 FILLER_22_755 ();
 sg13g2_decap_8 FILLER_22_762 ();
 sg13g2_decap_8 FILLER_22_769 ();
 sg13g2_decap_8 FILLER_22_776 ();
 sg13g2_decap_8 FILLER_22_783 ();
 sg13g2_decap_8 FILLER_22_790 ();
 sg13g2_decap_8 FILLER_22_797 ();
 sg13g2_decap_8 FILLER_22_804 ();
 sg13g2_decap_8 FILLER_22_811 ();
 sg13g2_decap_8 FILLER_22_818 ();
 sg13g2_decap_8 FILLER_22_825 ();
 sg13g2_decap_8 FILLER_22_832 ();
 sg13g2_decap_8 FILLER_22_839 ();
 sg13g2_decap_8 FILLER_22_846 ();
 sg13g2_decap_8 FILLER_22_853 ();
 sg13g2_fill_2 FILLER_22_860 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_23 ();
 sg13g2_fill_2 FILLER_23_37 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_fill_2 FILLER_23_64 ();
 sg13g2_fill_1 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_100 ();
 sg13g2_fill_1 FILLER_23_124 ();
 sg13g2_decap_4 FILLER_23_146 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_4 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_fill_2 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_342 ();
 sg13g2_fill_2 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_423 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_decap_4 FILLER_23_465 ();
 sg13g2_fill_2 FILLER_23_520 ();
 sg13g2_decap_8 FILLER_23_555 ();
 sg13g2_decap_8 FILLER_23_562 ();
 sg13g2_decap_8 FILLER_23_569 ();
 sg13g2_decap_8 FILLER_23_576 ();
 sg13g2_decap_8 FILLER_23_583 ();
 sg13g2_decap_8 FILLER_23_590 ();
 sg13g2_decap_8 FILLER_23_597 ();
 sg13g2_decap_8 FILLER_23_604 ();
 sg13g2_decap_8 FILLER_23_611 ();
 sg13g2_decap_8 FILLER_23_618 ();
 sg13g2_decap_8 FILLER_23_625 ();
 sg13g2_decap_8 FILLER_23_632 ();
 sg13g2_decap_8 FILLER_23_639 ();
 sg13g2_decap_8 FILLER_23_646 ();
 sg13g2_decap_8 FILLER_23_653 ();
 sg13g2_decap_8 FILLER_23_660 ();
 sg13g2_decap_8 FILLER_23_667 ();
 sg13g2_decap_8 FILLER_23_674 ();
 sg13g2_decap_8 FILLER_23_681 ();
 sg13g2_decap_8 FILLER_23_688 ();
 sg13g2_decap_8 FILLER_23_695 ();
 sg13g2_decap_8 FILLER_23_702 ();
 sg13g2_decap_8 FILLER_23_709 ();
 sg13g2_decap_8 FILLER_23_716 ();
 sg13g2_decap_8 FILLER_23_723 ();
 sg13g2_decap_8 FILLER_23_730 ();
 sg13g2_decap_8 FILLER_23_737 ();
 sg13g2_decap_8 FILLER_23_744 ();
 sg13g2_decap_8 FILLER_23_751 ();
 sg13g2_decap_8 FILLER_23_758 ();
 sg13g2_decap_8 FILLER_23_765 ();
 sg13g2_decap_8 FILLER_23_772 ();
 sg13g2_decap_8 FILLER_23_779 ();
 sg13g2_decap_8 FILLER_23_786 ();
 sg13g2_decap_8 FILLER_23_793 ();
 sg13g2_decap_8 FILLER_23_800 ();
 sg13g2_decap_8 FILLER_23_807 ();
 sg13g2_decap_8 FILLER_23_814 ();
 sg13g2_decap_8 FILLER_23_821 ();
 sg13g2_decap_8 FILLER_23_828 ();
 sg13g2_decap_8 FILLER_23_835 ();
 sg13g2_decap_8 FILLER_23_842 ();
 sg13g2_decap_8 FILLER_23_849 ();
 sg13g2_decap_4 FILLER_23_856 ();
 sg13g2_fill_2 FILLER_23_860 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_fill_1 FILLER_24_43 ();
 sg13g2_fill_2 FILLER_24_61 ();
 sg13g2_fill_1 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_144 ();
 sg13g2_decap_4 FILLER_24_171 ();
 sg13g2_fill_2 FILLER_24_175 ();
 sg13g2_decap_4 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_decap_4 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_decap_4 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_decap_4 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_331 ();
 sg13g2_decap_4 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_4 FILLER_24_395 ();
 sg13g2_fill_1 FILLER_24_482 ();
 sg13g2_fill_1 FILLER_24_509 ();
 sg13g2_fill_1 FILLER_24_519 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_11 ();
 sg13g2_fill_2 FILLER_25_45 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_decap_4 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_159 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_decap_4 FILLER_25_179 ();
 sg13g2_fill_2 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_decap_4 FILLER_25_234 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_decap_4 FILLER_25_369 ();
 sg13g2_decap_4 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_25_385 ();
 sg13g2_decap_4 FILLER_25_413 ();
 sg13g2_fill_1 FILLER_25_417 ();
 sg13g2_fill_1 FILLER_25_458 ();
 sg13g2_fill_2 FILLER_25_513 ();
 sg13g2_decap_8 FILLER_25_542 ();
 sg13g2_decap_8 FILLER_25_549 ();
 sg13g2_decap_8 FILLER_25_556 ();
 sg13g2_decap_8 FILLER_25_563 ();
 sg13g2_decap_8 FILLER_25_570 ();
 sg13g2_decap_8 FILLER_25_577 ();
 sg13g2_decap_8 FILLER_25_584 ();
 sg13g2_decap_8 FILLER_25_591 ();
 sg13g2_decap_8 FILLER_25_598 ();
 sg13g2_decap_8 FILLER_25_605 ();
 sg13g2_decap_8 FILLER_25_612 ();
 sg13g2_decap_8 FILLER_25_619 ();
 sg13g2_decap_8 FILLER_25_626 ();
 sg13g2_decap_8 FILLER_25_633 ();
 sg13g2_decap_8 FILLER_25_640 ();
 sg13g2_decap_8 FILLER_25_647 ();
 sg13g2_decap_8 FILLER_25_654 ();
 sg13g2_decap_8 FILLER_25_661 ();
 sg13g2_decap_8 FILLER_25_668 ();
 sg13g2_decap_8 FILLER_25_675 ();
 sg13g2_decap_8 FILLER_25_682 ();
 sg13g2_decap_8 FILLER_25_689 ();
 sg13g2_decap_8 FILLER_25_696 ();
 sg13g2_decap_8 FILLER_25_703 ();
 sg13g2_decap_8 FILLER_25_710 ();
 sg13g2_decap_8 FILLER_25_717 ();
 sg13g2_decap_8 FILLER_25_724 ();
 sg13g2_decap_8 FILLER_25_731 ();
 sg13g2_decap_8 FILLER_25_738 ();
 sg13g2_decap_8 FILLER_25_745 ();
 sg13g2_decap_8 FILLER_25_752 ();
 sg13g2_decap_8 FILLER_25_759 ();
 sg13g2_decap_8 FILLER_25_766 ();
 sg13g2_decap_8 FILLER_25_773 ();
 sg13g2_decap_8 FILLER_25_780 ();
 sg13g2_decap_8 FILLER_25_787 ();
 sg13g2_decap_8 FILLER_25_794 ();
 sg13g2_decap_8 FILLER_25_801 ();
 sg13g2_decap_8 FILLER_25_808 ();
 sg13g2_decap_8 FILLER_25_815 ();
 sg13g2_decap_8 FILLER_25_822 ();
 sg13g2_decap_8 FILLER_25_829 ();
 sg13g2_decap_8 FILLER_25_836 ();
 sg13g2_decap_8 FILLER_25_843 ();
 sg13g2_decap_8 FILLER_25_850 ();
 sg13g2_decap_4 FILLER_25_857 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_fill_2 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_decap_4 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_decap_4 FILLER_26_262 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_decap_4 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_decap_4 FILLER_26_428 ();
 sg13g2_fill_1 FILLER_26_432 ();
 sg13g2_fill_1 FILLER_26_452 ();
 sg13g2_fill_2 FILLER_26_479 ();
 sg13g2_fill_1 FILLER_26_481 ();
 sg13g2_fill_2 FILLER_26_519 ();
 sg13g2_decap_8 FILLER_26_530 ();
 sg13g2_decap_8 FILLER_26_537 ();
 sg13g2_decap_8 FILLER_26_544 ();
 sg13g2_decap_8 FILLER_26_551 ();
 sg13g2_decap_8 FILLER_26_558 ();
 sg13g2_decap_8 FILLER_26_565 ();
 sg13g2_decap_8 FILLER_26_572 ();
 sg13g2_decap_8 FILLER_26_579 ();
 sg13g2_decap_8 FILLER_26_586 ();
 sg13g2_decap_8 FILLER_26_593 ();
 sg13g2_decap_8 FILLER_26_600 ();
 sg13g2_decap_8 FILLER_26_607 ();
 sg13g2_decap_8 FILLER_26_614 ();
 sg13g2_decap_8 FILLER_26_621 ();
 sg13g2_decap_8 FILLER_26_628 ();
 sg13g2_decap_8 FILLER_26_635 ();
 sg13g2_decap_8 FILLER_26_642 ();
 sg13g2_decap_8 FILLER_26_649 ();
 sg13g2_decap_8 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_decap_8 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_698 ();
 sg13g2_decap_8 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_712 ();
 sg13g2_decap_8 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_747 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_fill_2 FILLER_26_859 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_110 ();
 sg13g2_decap_8 FILLER_27_117 ();
 sg13g2_decap_8 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_decap_4 FILLER_27_162 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_decap_4 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_fill_2 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_decap_4 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_320 ();
 sg13g2_decap_8 FILLER_27_327 ();
 sg13g2_fill_2 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_4 FILLER_27_414 ();
 sg13g2_fill_2 FILLER_27_418 ();
 sg13g2_fill_1 FILLER_27_462 ();
 sg13g2_fill_1 FILLER_27_477 ();
 sg13g2_fill_1 FILLER_27_495 ();
 sg13g2_fill_1 FILLER_27_513 ();
 sg13g2_decap_8 FILLER_27_524 ();
 sg13g2_decap_8 FILLER_27_531 ();
 sg13g2_decap_8 FILLER_27_538 ();
 sg13g2_decap_8 FILLER_27_545 ();
 sg13g2_decap_8 FILLER_27_552 ();
 sg13g2_decap_8 FILLER_27_559 ();
 sg13g2_decap_8 FILLER_27_566 ();
 sg13g2_decap_8 FILLER_27_573 ();
 sg13g2_decap_8 FILLER_27_580 ();
 sg13g2_decap_8 FILLER_27_587 ();
 sg13g2_decap_8 FILLER_27_594 ();
 sg13g2_decap_8 FILLER_27_601 ();
 sg13g2_decap_8 FILLER_27_608 ();
 sg13g2_decap_8 FILLER_27_615 ();
 sg13g2_decap_8 FILLER_27_622 ();
 sg13g2_decap_8 FILLER_27_629 ();
 sg13g2_decap_8 FILLER_27_636 ();
 sg13g2_decap_8 FILLER_27_643 ();
 sg13g2_decap_8 FILLER_27_650 ();
 sg13g2_decap_8 FILLER_27_657 ();
 sg13g2_decap_8 FILLER_27_664 ();
 sg13g2_decap_8 FILLER_27_671 ();
 sg13g2_decap_8 FILLER_27_678 ();
 sg13g2_decap_8 FILLER_27_685 ();
 sg13g2_decap_8 FILLER_27_692 ();
 sg13g2_decap_8 FILLER_27_699 ();
 sg13g2_decap_8 FILLER_27_706 ();
 sg13g2_decap_8 FILLER_27_713 ();
 sg13g2_decap_8 FILLER_27_720 ();
 sg13g2_decap_8 FILLER_27_727 ();
 sg13g2_decap_8 FILLER_27_734 ();
 sg13g2_decap_8 FILLER_27_741 ();
 sg13g2_decap_8 FILLER_27_748 ();
 sg13g2_decap_8 FILLER_27_755 ();
 sg13g2_decap_8 FILLER_27_762 ();
 sg13g2_decap_8 FILLER_27_769 ();
 sg13g2_decap_8 FILLER_27_776 ();
 sg13g2_decap_8 FILLER_27_783 ();
 sg13g2_decap_8 FILLER_27_790 ();
 sg13g2_decap_8 FILLER_27_797 ();
 sg13g2_decap_8 FILLER_27_804 ();
 sg13g2_decap_8 FILLER_27_811 ();
 sg13g2_decap_8 FILLER_27_818 ();
 sg13g2_decap_8 FILLER_27_825 ();
 sg13g2_decap_8 FILLER_27_832 ();
 sg13g2_decap_8 FILLER_27_839 ();
 sg13g2_decap_8 FILLER_27_846 ();
 sg13g2_decap_8 FILLER_27_853 ();
 sg13g2_fill_2 FILLER_27_860 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_11 ();
 sg13g2_fill_1 FILLER_28_34 ();
 sg13g2_fill_1 FILLER_28_92 ();
 sg13g2_fill_2 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_182 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_4 FILLER_28_321 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_348 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_decap_4 FILLER_28_411 ();
 sg13g2_decap_4 FILLER_28_424 ();
 sg13g2_fill_1 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_28_510 ();
 sg13g2_decap_8 FILLER_28_517 ();
 sg13g2_decap_8 FILLER_28_524 ();
 sg13g2_decap_8 FILLER_28_531 ();
 sg13g2_decap_8 FILLER_28_538 ();
 sg13g2_decap_8 FILLER_28_545 ();
 sg13g2_decap_8 FILLER_28_552 ();
 sg13g2_decap_8 FILLER_28_559 ();
 sg13g2_decap_8 FILLER_28_566 ();
 sg13g2_decap_8 FILLER_28_573 ();
 sg13g2_decap_8 FILLER_28_580 ();
 sg13g2_decap_8 FILLER_28_587 ();
 sg13g2_decap_8 FILLER_28_594 ();
 sg13g2_decap_8 FILLER_28_601 ();
 sg13g2_decap_8 FILLER_28_608 ();
 sg13g2_decap_8 FILLER_28_615 ();
 sg13g2_decap_8 FILLER_28_622 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_decap_8 FILLER_28_636 ();
 sg13g2_decap_8 FILLER_28_643 ();
 sg13g2_decap_8 FILLER_28_650 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_decap_8 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_671 ();
 sg13g2_decap_8 FILLER_28_678 ();
 sg13g2_decap_8 FILLER_28_685 ();
 sg13g2_decap_8 FILLER_28_692 ();
 sg13g2_decap_8 FILLER_28_699 ();
 sg13g2_decap_8 FILLER_28_706 ();
 sg13g2_decap_8 FILLER_28_713 ();
 sg13g2_decap_8 FILLER_28_720 ();
 sg13g2_decap_8 FILLER_28_727 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_decap_8 FILLER_28_741 ();
 sg13g2_decap_8 FILLER_28_748 ();
 sg13g2_decap_8 FILLER_28_755 ();
 sg13g2_decap_8 FILLER_28_762 ();
 sg13g2_decap_8 FILLER_28_769 ();
 sg13g2_decap_8 FILLER_28_776 ();
 sg13g2_decap_8 FILLER_28_783 ();
 sg13g2_decap_8 FILLER_28_790 ();
 sg13g2_decap_8 FILLER_28_797 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_8 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_818 ();
 sg13g2_decap_8 FILLER_28_825 ();
 sg13g2_decap_8 FILLER_28_832 ();
 sg13g2_decap_8 FILLER_28_839 ();
 sg13g2_decap_8 FILLER_28_846 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_134 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_decap_4 FILLER_29_212 ();
 sg13g2_fill_2 FILLER_29_221 ();
 sg13g2_decap_4 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_decap_4 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_4 FILLER_29_349 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_fill_1 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_415 ();
 sg13g2_fill_1 FILLER_29_433 ();
 sg13g2_decap_8 FILLER_29_443 ();
 sg13g2_decap_8 FILLER_29_450 ();
 sg13g2_decap_8 FILLER_29_457 ();
 sg13g2_decap_4 FILLER_29_464 ();
 sg13g2_fill_1 FILLER_29_484 ();
 sg13g2_decap_8 FILLER_29_494 ();
 sg13g2_decap_8 FILLER_29_501 ();
 sg13g2_decap_8 FILLER_29_508 ();
 sg13g2_decap_8 FILLER_29_515 ();
 sg13g2_decap_8 FILLER_29_522 ();
 sg13g2_decap_8 FILLER_29_529 ();
 sg13g2_decap_8 FILLER_29_536 ();
 sg13g2_decap_8 FILLER_29_543 ();
 sg13g2_decap_8 FILLER_29_550 ();
 sg13g2_decap_8 FILLER_29_557 ();
 sg13g2_decap_8 FILLER_29_564 ();
 sg13g2_decap_8 FILLER_29_571 ();
 sg13g2_decap_8 FILLER_29_578 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_decap_8 FILLER_29_592 ();
 sg13g2_decap_8 FILLER_29_599 ();
 sg13g2_decap_8 FILLER_29_606 ();
 sg13g2_decap_8 FILLER_29_613 ();
 sg13g2_decap_8 FILLER_29_620 ();
 sg13g2_decap_8 FILLER_29_627 ();
 sg13g2_decap_8 FILLER_29_634 ();
 sg13g2_decap_8 FILLER_29_641 ();
 sg13g2_decap_8 FILLER_29_648 ();
 sg13g2_decap_8 FILLER_29_655 ();
 sg13g2_decap_8 FILLER_29_662 ();
 sg13g2_decap_8 FILLER_29_669 ();
 sg13g2_decap_8 FILLER_29_676 ();
 sg13g2_decap_8 FILLER_29_683 ();
 sg13g2_decap_8 FILLER_29_690 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_decap_8 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_711 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_725 ();
 sg13g2_decap_8 FILLER_29_732 ();
 sg13g2_decap_8 FILLER_29_739 ();
 sg13g2_decap_8 FILLER_29_746 ();
 sg13g2_decap_8 FILLER_29_753 ();
 sg13g2_decap_8 FILLER_29_760 ();
 sg13g2_decap_8 FILLER_29_767 ();
 sg13g2_decap_8 FILLER_29_774 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_decap_8 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_802 ();
 sg13g2_decap_8 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_823 ();
 sg13g2_decap_8 FILLER_29_830 ();
 sg13g2_decap_8 FILLER_29_837 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_4 FILLER_29_858 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_33 ();
 sg13g2_fill_1 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_47 ();
 sg13g2_decap_8 FILLER_30_64 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_decap_4 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_decap_4 FILLER_30_113 ();
 sg13g2_fill_2 FILLER_30_117 ();
 sg13g2_decap_8 FILLER_30_148 ();
 sg13g2_decap_8 FILLER_30_155 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_171 ();
 sg13g2_decap_4 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_decap_4 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_233 ();
 sg13g2_decap_4 FILLER_30_240 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_fill_1 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_decap_4 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_fill_2 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_404 ();
 sg13g2_decap_4 FILLER_30_411 ();
 sg13g2_fill_2 FILLER_30_415 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_485 ();
 sg13g2_decap_8 FILLER_30_492 ();
 sg13g2_decap_8 FILLER_30_499 ();
 sg13g2_decap_8 FILLER_30_506 ();
 sg13g2_decap_8 FILLER_30_513 ();
 sg13g2_decap_8 FILLER_30_520 ();
 sg13g2_decap_8 FILLER_30_527 ();
 sg13g2_decap_8 FILLER_30_534 ();
 sg13g2_decap_8 FILLER_30_541 ();
 sg13g2_decap_8 FILLER_30_548 ();
 sg13g2_decap_8 FILLER_30_555 ();
 sg13g2_decap_8 FILLER_30_562 ();
 sg13g2_decap_8 FILLER_30_569 ();
 sg13g2_decap_8 FILLER_30_576 ();
 sg13g2_decap_8 FILLER_30_583 ();
 sg13g2_decap_8 FILLER_30_590 ();
 sg13g2_decap_8 FILLER_30_597 ();
 sg13g2_decap_8 FILLER_30_604 ();
 sg13g2_decap_8 FILLER_30_611 ();
 sg13g2_decap_8 FILLER_30_618 ();
 sg13g2_decap_8 FILLER_30_625 ();
 sg13g2_decap_8 FILLER_30_632 ();
 sg13g2_decap_8 FILLER_30_639 ();
 sg13g2_decap_8 FILLER_30_646 ();
 sg13g2_decap_8 FILLER_30_653 ();
 sg13g2_decap_8 FILLER_30_660 ();
 sg13g2_decap_8 FILLER_30_667 ();
 sg13g2_decap_8 FILLER_30_674 ();
 sg13g2_decap_8 FILLER_30_681 ();
 sg13g2_decap_8 FILLER_30_688 ();
 sg13g2_decap_8 FILLER_30_695 ();
 sg13g2_decap_8 FILLER_30_702 ();
 sg13g2_decap_8 FILLER_30_709 ();
 sg13g2_decap_8 FILLER_30_716 ();
 sg13g2_decap_8 FILLER_30_723 ();
 sg13g2_decap_8 FILLER_30_730 ();
 sg13g2_decap_8 FILLER_30_737 ();
 sg13g2_decap_8 FILLER_30_744 ();
 sg13g2_decap_8 FILLER_30_751 ();
 sg13g2_decap_8 FILLER_30_758 ();
 sg13g2_decap_8 FILLER_30_765 ();
 sg13g2_decap_8 FILLER_30_772 ();
 sg13g2_decap_8 FILLER_30_779 ();
 sg13g2_decap_8 FILLER_30_786 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_4 FILLER_30_856 ();
 sg13g2_fill_2 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_95 ();
 sg13g2_fill_2 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_139 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_fill_2 FILLER_31_269 ();
 sg13g2_decap_4 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_fill_1 FILLER_31_299 ();
 sg13g2_fill_2 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_fill_1 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_fill_1 FILLER_31_418 ();
 sg13g2_fill_2 FILLER_31_446 ();
 sg13g2_decap_8 FILLER_31_453 ();
 sg13g2_fill_2 FILLER_31_460 ();
 sg13g2_fill_2 FILLER_31_471 ();
 sg13g2_fill_1 FILLER_31_473 ();
 sg13g2_fill_2 FILLER_31_482 ();
 sg13g2_fill_1 FILLER_31_484 ();
 sg13g2_decap_8 FILLER_31_493 ();
 sg13g2_decap_8 FILLER_31_500 ();
 sg13g2_decap_8 FILLER_31_507 ();
 sg13g2_decap_8 FILLER_31_514 ();
 sg13g2_decap_8 FILLER_31_521 ();
 sg13g2_decap_8 FILLER_31_528 ();
 sg13g2_decap_8 FILLER_31_535 ();
 sg13g2_decap_8 FILLER_31_542 ();
 sg13g2_decap_8 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_556 ();
 sg13g2_decap_8 FILLER_31_563 ();
 sg13g2_decap_8 FILLER_31_570 ();
 sg13g2_decap_8 FILLER_31_577 ();
 sg13g2_decap_8 FILLER_31_584 ();
 sg13g2_fill_2 FILLER_31_591 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_43 ();
 sg13g2_fill_2 FILLER_32_54 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_74 ();
 sg13g2_fill_2 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_decap_4 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_197 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_264 ();
 sg13g2_fill_2 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_decap_4 FILLER_32_295 ();
 sg13g2_fill_2 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_311 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_decap_4 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_380 ();
 sg13g2_fill_1 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_406 ();
 sg13g2_fill_2 FILLER_32_410 ();
 sg13g2_fill_2 FILLER_32_438 ();
 sg13g2_fill_2 FILLER_32_474 ();
 sg13g2_fill_1 FILLER_32_476 ();
 sg13g2_fill_2 FILLER_32_495 ();
 sg13g2_fill_1 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_507 ();
 sg13g2_decap_8 FILLER_32_514 ();
 sg13g2_decap_8 FILLER_32_521 ();
 sg13g2_decap_8 FILLER_32_528 ();
 sg13g2_decap_4 FILLER_32_535 ();
 sg13g2_fill_1 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_556 ();
 sg13g2_decap_8 FILLER_32_563 ();
 sg13g2_decap_4 FILLER_32_570 ();
 sg13g2_fill_1 FILLER_32_574 ();
 sg13g2_decap_8 FILLER_32_610 ();
 sg13g2_decap_8 FILLER_32_617 ();
 sg13g2_decap_8 FILLER_32_624 ();
 sg13g2_decap_8 FILLER_32_631 ();
 sg13g2_decap_8 FILLER_32_638 ();
 sg13g2_decap_8 FILLER_32_645 ();
 sg13g2_decap_8 FILLER_32_652 ();
 sg13g2_decap_8 FILLER_32_659 ();
 sg13g2_decap_8 FILLER_32_666 ();
 sg13g2_decap_8 FILLER_32_673 ();
 sg13g2_decap_8 FILLER_32_680 ();
 sg13g2_decap_8 FILLER_32_687 ();
 sg13g2_decap_8 FILLER_32_694 ();
 sg13g2_decap_8 FILLER_32_701 ();
 sg13g2_decap_8 FILLER_32_708 ();
 sg13g2_decap_8 FILLER_32_715 ();
 sg13g2_decap_8 FILLER_32_722 ();
 sg13g2_decap_8 FILLER_32_729 ();
 sg13g2_decap_8 FILLER_32_736 ();
 sg13g2_decap_8 FILLER_32_743 ();
 sg13g2_decap_8 FILLER_32_750 ();
 sg13g2_decap_8 FILLER_32_757 ();
 sg13g2_decap_8 FILLER_32_764 ();
 sg13g2_decap_8 FILLER_32_771 ();
 sg13g2_decap_8 FILLER_32_778 ();
 sg13g2_decap_8 FILLER_32_785 ();
 sg13g2_decap_8 FILLER_32_792 ();
 sg13g2_decap_8 FILLER_32_799 ();
 sg13g2_decap_8 FILLER_32_806 ();
 sg13g2_decap_8 FILLER_32_813 ();
 sg13g2_decap_8 FILLER_32_820 ();
 sg13g2_decap_8 FILLER_32_827 ();
 sg13g2_decap_8 FILLER_32_834 ();
 sg13g2_decap_8 FILLER_32_841 ();
 sg13g2_decap_8 FILLER_32_848 ();
 sg13g2_decap_8 FILLER_32_855 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_53 ();
 sg13g2_decap_4 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_90 ();
 sg13g2_decap_4 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_99 ();
 sg13g2_decap_4 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_170 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_fill_1 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_decap_4 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_284 ();
 sg13g2_fill_1 FILLER_33_286 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_decap_8 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_364 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_fill_1 FILLER_33_442 ();
 sg13g2_fill_2 FILLER_33_456 ();
 sg13g2_fill_1 FILLER_33_458 ();
 sg13g2_fill_2 FILLER_33_480 ();
 sg13g2_fill_2 FILLER_33_508 ();
 sg13g2_fill_1 FILLER_33_510 ();
 sg13g2_fill_2 FILLER_33_541 ();
 sg13g2_fill_2 FILLER_33_569 ();
 sg13g2_fill_1 FILLER_33_571 ();
 sg13g2_fill_1 FILLER_33_575 ();
 sg13g2_decap_4 FILLER_33_597 ();
 sg13g2_decap_8 FILLER_33_610 ();
 sg13g2_fill_1 FILLER_33_617 ();
 sg13g2_decap_8 FILLER_33_627 ();
 sg13g2_decap_8 FILLER_33_634 ();
 sg13g2_decap_8 FILLER_33_641 ();
 sg13g2_decap_8 FILLER_33_648 ();
 sg13g2_decap_8 FILLER_33_655 ();
 sg13g2_decap_8 FILLER_33_662 ();
 sg13g2_decap_8 FILLER_33_669 ();
 sg13g2_decap_8 FILLER_33_676 ();
 sg13g2_decap_8 FILLER_33_683 ();
 sg13g2_decap_8 FILLER_33_690 ();
 sg13g2_decap_8 FILLER_33_697 ();
 sg13g2_decap_8 FILLER_33_704 ();
 sg13g2_decap_8 FILLER_33_711 ();
 sg13g2_decap_8 FILLER_33_718 ();
 sg13g2_decap_8 FILLER_33_725 ();
 sg13g2_decap_8 FILLER_33_732 ();
 sg13g2_decap_8 FILLER_33_739 ();
 sg13g2_decap_8 FILLER_33_746 ();
 sg13g2_decap_8 FILLER_33_753 ();
 sg13g2_decap_8 FILLER_33_760 ();
 sg13g2_decap_8 FILLER_33_767 ();
 sg13g2_decap_8 FILLER_33_774 ();
 sg13g2_decap_8 FILLER_33_781 ();
 sg13g2_decap_8 FILLER_33_788 ();
 sg13g2_decap_8 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_decap_8 FILLER_33_809 ();
 sg13g2_decap_8 FILLER_33_816 ();
 sg13g2_decap_8 FILLER_33_823 ();
 sg13g2_decap_8 FILLER_33_830 ();
 sg13g2_decap_8 FILLER_33_837 ();
 sg13g2_decap_8 FILLER_33_844 ();
 sg13g2_decap_8 FILLER_33_851 ();
 sg13g2_decap_4 FILLER_33_858 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_4 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_decap_8 FILLER_34_139 ();
 sg13g2_fill_2 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_decap_4 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_168 ();
 sg13g2_fill_2 FILLER_34_183 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_fill_2 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_decap_8 FILLER_34_247 ();
 sg13g2_decap_4 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_fill_2 FILLER_34_331 ();
 sg13g2_fill_2 FILLER_34_362 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_decap_4 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_4 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_441 ();
 sg13g2_fill_1 FILLER_34_443 ();
 sg13g2_fill_2 FILLER_34_505 ();
 sg13g2_fill_1 FILLER_34_507 ();
 sg13g2_fill_1 FILLER_34_544 ();
 sg13g2_decap_4 FILLER_34_554 ();
 sg13g2_fill_2 FILLER_34_558 ();
 sg13g2_fill_2 FILLER_34_573 ();
 sg13g2_fill_2 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_628 ();
 sg13g2_decap_8 FILLER_34_635 ();
 sg13g2_decap_8 FILLER_34_642 ();
 sg13g2_decap_8 FILLER_34_649 ();
 sg13g2_decap_8 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_663 ();
 sg13g2_decap_8 FILLER_34_670 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_691 ();
 sg13g2_decap_8 FILLER_34_698 ();
 sg13g2_decap_8 FILLER_34_705 ();
 sg13g2_decap_8 FILLER_34_712 ();
 sg13g2_decap_8 FILLER_34_719 ();
 sg13g2_decap_8 FILLER_34_726 ();
 sg13g2_decap_8 FILLER_34_733 ();
 sg13g2_decap_8 FILLER_34_740 ();
 sg13g2_decap_8 FILLER_34_747 ();
 sg13g2_decap_8 FILLER_34_754 ();
 sg13g2_decap_8 FILLER_34_761 ();
 sg13g2_decap_8 FILLER_34_768 ();
 sg13g2_decap_8 FILLER_34_775 ();
 sg13g2_decap_8 FILLER_34_782 ();
 sg13g2_decap_8 FILLER_34_789 ();
 sg13g2_decap_8 FILLER_34_796 ();
 sg13g2_decap_8 FILLER_34_803 ();
 sg13g2_decap_8 FILLER_34_810 ();
 sg13g2_decap_8 FILLER_34_817 ();
 sg13g2_decap_8 FILLER_34_824 ();
 sg13g2_decap_8 FILLER_34_831 ();
 sg13g2_decap_8 FILLER_34_838 ();
 sg13g2_decap_8 FILLER_34_845 ();
 sg13g2_decap_8 FILLER_34_852 ();
 sg13g2_fill_2 FILLER_34_859 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_186 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_decap_4 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_304 ();
 sg13g2_decap_8 FILLER_35_324 ();
 sg13g2_decap_4 FILLER_35_331 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_439 ();
 sg13g2_decap_8 FILLER_35_467 ();
 sg13g2_fill_1 FILLER_35_474 ();
 sg13g2_fill_2 FILLER_35_511 ();
 sg13g2_fill_1 FILLER_35_513 ();
 sg13g2_fill_1 FILLER_35_528 ();
 sg13g2_fill_2 FILLER_35_542 ();
 sg13g2_fill_2 FILLER_35_560 ();
 sg13g2_fill_1 FILLER_35_562 ();
 sg13g2_fill_2 FILLER_35_568 ();
 sg13g2_fill_1 FILLER_35_599 ();
 sg13g2_fill_2 FILLER_35_605 ();
 sg13g2_fill_1 FILLER_35_607 ();
 sg13g2_decap_8 FILLER_35_634 ();
 sg13g2_decap_8 FILLER_35_641 ();
 sg13g2_decap_8 FILLER_35_648 ();
 sg13g2_decap_8 FILLER_35_655 ();
 sg13g2_decap_8 FILLER_35_662 ();
 sg13g2_decap_8 FILLER_35_669 ();
 sg13g2_decap_8 FILLER_35_676 ();
 sg13g2_decap_8 FILLER_35_683 ();
 sg13g2_decap_8 FILLER_35_690 ();
 sg13g2_decap_8 FILLER_35_697 ();
 sg13g2_decap_8 FILLER_35_704 ();
 sg13g2_decap_8 FILLER_35_711 ();
 sg13g2_decap_8 FILLER_35_718 ();
 sg13g2_decap_8 FILLER_35_725 ();
 sg13g2_decap_8 FILLER_35_732 ();
 sg13g2_decap_8 FILLER_35_739 ();
 sg13g2_decap_8 FILLER_35_746 ();
 sg13g2_decap_8 FILLER_35_753 ();
 sg13g2_decap_8 FILLER_35_760 ();
 sg13g2_decap_8 FILLER_35_767 ();
 sg13g2_decap_8 FILLER_35_774 ();
 sg13g2_decap_8 FILLER_35_781 ();
 sg13g2_decap_8 FILLER_35_788 ();
 sg13g2_decap_8 FILLER_35_795 ();
 sg13g2_decap_8 FILLER_35_802 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_decap_8 FILLER_35_823 ();
 sg13g2_decap_8 FILLER_35_830 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_decap_8 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_decap_4 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_130 ();
 sg13g2_fill_2 FILLER_36_134 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_155 ();
 sg13g2_decap_4 FILLER_36_170 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_decap_4 FILLER_36_211 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_decap_4 FILLER_36_243 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_decap_8 FILLER_36_284 ();
 sg13g2_decap_4 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_decap_4 FILLER_36_301 ();
 sg13g2_decap_4 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_fill_2 FILLER_36_349 ();
 sg13g2_decap_4 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_fill_2 FILLER_36_408 ();
 sg13g2_fill_2 FILLER_36_430 ();
 sg13g2_decap_8 FILLER_36_445 ();
 sg13g2_decap_8 FILLER_36_452 ();
 sg13g2_fill_2 FILLER_36_459 ();
 sg13g2_fill_2 FILLER_36_466 ();
 sg13g2_fill_1 FILLER_36_468 ();
 sg13g2_fill_2 FILLER_36_531 ();
 sg13g2_fill_1 FILLER_36_547 ();
 sg13g2_decap_4 FILLER_36_552 ();
 sg13g2_fill_2 FILLER_36_556 ();
 sg13g2_decap_8 FILLER_36_562 ();
 sg13g2_fill_1 FILLER_36_595 ();
 sg13g2_decap_8 FILLER_36_621 ();
 sg13g2_decap_8 FILLER_36_628 ();
 sg13g2_decap_8 FILLER_36_635 ();
 sg13g2_decap_8 FILLER_36_642 ();
 sg13g2_decap_8 FILLER_36_649 ();
 sg13g2_decap_8 FILLER_36_656 ();
 sg13g2_decap_8 FILLER_36_663 ();
 sg13g2_decap_8 FILLER_36_670 ();
 sg13g2_decap_8 FILLER_36_677 ();
 sg13g2_decap_8 FILLER_36_684 ();
 sg13g2_decap_8 FILLER_36_691 ();
 sg13g2_decap_8 FILLER_36_698 ();
 sg13g2_decap_8 FILLER_36_705 ();
 sg13g2_decap_8 FILLER_36_712 ();
 sg13g2_decap_8 FILLER_36_719 ();
 sg13g2_decap_8 FILLER_36_726 ();
 sg13g2_decap_8 FILLER_36_733 ();
 sg13g2_decap_8 FILLER_36_740 ();
 sg13g2_decap_8 FILLER_36_747 ();
 sg13g2_decap_8 FILLER_36_754 ();
 sg13g2_decap_8 FILLER_36_761 ();
 sg13g2_decap_8 FILLER_36_768 ();
 sg13g2_decap_8 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_782 ();
 sg13g2_decap_8 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_fill_2 FILLER_37_77 ();
 sg13g2_fill_1 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_111 ();
 sg13g2_decap_4 FILLER_37_155 ();
 sg13g2_fill_1 FILLER_37_159 ();
 sg13g2_fill_1 FILLER_37_170 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_fill_1 FILLER_37_211 ();
 sg13g2_decap_4 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_256 ();
 sg13g2_decap_4 FILLER_37_265 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_328 ();
 sg13g2_fill_2 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_346 ();
 sg13g2_fill_2 FILLER_37_379 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_fill_1 FILLER_37_417 ();
 sg13g2_fill_2 FILLER_37_434 ();
 sg13g2_fill_2 FILLER_37_470 ();
 sg13g2_fill_1 FILLER_37_477 ();
 sg13g2_decap_8 FILLER_37_491 ();
 sg13g2_decap_4 FILLER_37_498 ();
 sg13g2_fill_1 FILLER_37_528 ();
 sg13g2_fill_2 FILLER_37_565 ();
 sg13g2_decap_8 FILLER_37_586 ();
 sg13g2_decap_4 FILLER_37_593 ();
 sg13g2_fill_1 FILLER_37_597 ();
 sg13g2_decap_8 FILLER_37_647 ();
 sg13g2_decap_8 FILLER_37_654 ();
 sg13g2_decap_8 FILLER_37_661 ();
 sg13g2_decap_8 FILLER_37_668 ();
 sg13g2_decap_8 FILLER_37_675 ();
 sg13g2_decap_8 FILLER_37_682 ();
 sg13g2_decap_8 FILLER_37_689 ();
 sg13g2_decap_8 FILLER_37_696 ();
 sg13g2_decap_8 FILLER_37_703 ();
 sg13g2_decap_8 FILLER_37_710 ();
 sg13g2_decap_8 FILLER_37_717 ();
 sg13g2_decap_8 FILLER_37_724 ();
 sg13g2_decap_8 FILLER_37_731 ();
 sg13g2_decap_8 FILLER_37_738 ();
 sg13g2_decap_8 FILLER_37_745 ();
 sg13g2_decap_8 FILLER_37_752 ();
 sg13g2_decap_8 FILLER_37_759 ();
 sg13g2_decap_8 FILLER_37_766 ();
 sg13g2_decap_8 FILLER_37_773 ();
 sg13g2_decap_8 FILLER_37_780 ();
 sg13g2_decap_8 FILLER_37_787 ();
 sg13g2_decap_8 FILLER_37_794 ();
 sg13g2_decap_8 FILLER_37_801 ();
 sg13g2_decap_8 FILLER_37_808 ();
 sg13g2_decap_8 FILLER_37_815 ();
 sg13g2_decap_8 FILLER_37_822 ();
 sg13g2_decap_8 FILLER_37_829 ();
 sg13g2_decap_8 FILLER_37_836 ();
 sg13g2_decap_8 FILLER_37_843 ();
 sg13g2_decap_8 FILLER_37_850 ();
 sg13g2_decap_4 FILLER_37_857 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_77 ();
 sg13g2_fill_1 FILLER_38_79 ();
 sg13g2_decap_4 FILLER_38_114 ();
 sg13g2_fill_1 FILLER_38_118 ();
 sg13g2_decap_4 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_decap_4 FILLER_38_187 ();
 sg13g2_decap_4 FILLER_38_205 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_fill_2 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_341 ();
 sg13g2_fill_2 FILLER_38_347 ();
 sg13g2_fill_1 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_fill_2 FILLER_38_413 ();
 sg13g2_decap_4 FILLER_38_439 ();
 sg13g2_fill_1 FILLER_38_443 ();
 sg13g2_decap_8 FILLER_38_452 ();
 sg13g2_decap_8 FILLER_38_459 ();
 sg13g2_fill_2 FILLER_38_466 ();
 sg13g2_decap_4 FILLER_38_488 ();
 sg13g2_fill_2 FILLER_38_492 ();
 sg13g2_decap_8 FILLER_38_499 ();
 sg13g2_fill_1 FILLER_38_506 ();
 sg13g2_fill_1 FILLER_38_531 ();
 sg13g2_fill_2 FILLER_38_536 ();
 sg13g2_fill_1 FILLER_38_563 ();
 sg13g2_fill_2 FILLER_38_602 ();
 sg13g2_decap_8 FILLER_38_666 ();
 sg13g2_decap_8 FILLER_38_673 ();
 sg13g2_decap_8 FILLER_38_680 ();
 sg13g2_decap_8 FILLER_38_687 ();
 sg13g2_decap_8 FILLER_38_694 ();
 sg13g2_decap_8 FILLER_38_701 ();
 sg13g2_decap_8 FILLER_38_708 ();
 sg13g2_decap_8 FILLER_38_715 ();
 sg13g2_decap_8 FILLER_38_722 ();
 sg13g2_decap_8 FILLER_38_729 ();
 sg13g2_decap_8 FILLER_38_736 ();
 sg13g2_decap_8 FILLER_38_743 ();
 sg13g2_decap_8 FILLER_38_750 ();
 sg13g2_decap_8 FILLER_38_757 ();
 sg13g2_decap_8 FILLER_38_764 ();
 sg13g2_decap_8 FILLER_38_771 ();
 sg13g2_decap_8 FILLER_38_778 ();
 sg13g2_decap_8 FILLER_38_785 ();
 sg13g2_decap_8 FILLER_38_792 ();
 sg13g2_decap_8 FILLER_38_799 ();
 sg13g2_decap_8 FILLER_38_806 ();
 sg13g2_decap_8 FILLER_38_813 ();
 sg13g2_decap_8 FILLER_38_820 ();
 sg13g2_decap_8 FILLER_38_827 ();
 sg13g2_decap_8 FILLER_38_834 ();
 sg13g2_decap_8 FILLER_38_841 ();
 sg13g2_decap_8 FILLER_38_848 ();
 sg13g2_decap_8 FILLER_38_855 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_fill_2 FILLER_39_86 ();
 sg13g2_fill_1 FILLER_39_88 ();
 sg13g2_decap_4 FILLER_39_97 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_decap_4 FILLER_39_120 ();
 sg13g2_fill_1 FILLER_39_124 ();
 sg13g2_fill_2 FILLER_39_135 ();
 sg13g2_fill_1 FILLER_39_137 ();
 sg13g2_fill_2 FILLER_39_151 ();
 sg13g2_fill_1 FILLER_39_183 ();
 sg13g2_fill_1 FILLER_39_211 ();
 sg13g2_fill_2 FILLER_39_229 ();
 sg13g2_fill_1 FILLER_39_231 ();
 sg13g2_decap_4 FILLER_39_242 ();
 sg13g2_fill_2 FILLER_39_246 ();
 sg13g2_fill_2 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_277 ();
 sg13g2_fill_2 FILLER_39_287 ();
 sg13g2_fill_1 FILLER_39_294 ();
 sg13g2_decap_4 FILLER_39_300 ();
 sg13g2_fill_2 FILLER_39_347 ();
 sg13g2_fill_1 FILLER_39_349 ();
 sg13g2_fill_2 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_fill_1 FILLER_39_392 ();
 sg13g2_fill_2 FILLER_39_464 ();
 sg13g2_fill_1 FILLER_39_466 ();
 sg13g2_decap_8 FILLER_39_481 ();
 sg13g2_fill_2 FILLER_39_488 ();
 sg13g2_decap_4 FILLER_39_495 ();
 sg13g2_fill_2 FILLER_39_542 ();
 sg13g2_fill_2 FILLER_39_576 ();
 sg13g2_fill_1 FILLER_39_597 ();
 sg13g2_fill_2 FILLER_39_622 ();
 sg13g2_fill_2 FILLER_39_662 ();
 sg13g2_fill_2 FILLER_39_675 ();
 sg13g2_fill_1 FILLER_39_677 ();
 sg13g2_decap_8 FILLER_39_682 ();
 sg13g2_decap_8 FILLER_39_689 ();
 sg13g2_decap_8 FILLER_39_696 ();
 sg13g2_decap_8 FILLER_39_703 ();
 sg13g2_decap_8 FILLER_39_710 ();
 sg13g2_decap_8 FILLER_39_717 ();
 sg13g2_decap_8 FILLER_39_724 ();
 sg13g2_decap_8 FILLER_39_731 ();
 sg13g2_decap_8 FILLER_39_738 ();
 sg13g2_decap_8 FILLER_39_745 ();
 sg13g2_decap_8 FILLER_39_752 ();
 sg13g2_decap_8 FILLER_39_759 ();
 sg13g2_decap_8 FILLER_39_766 ();
 sg13g2_decap_8 FILLER_39_773 ();
 sg13g2_decap_8 FILLER_39_780 ();
 sg13g2_decap_8 FILLER_39_787 ();
 sg13g2_decap_8 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_801 ();
 sg13g2_decap_8 FILLER_39_808 ();
 sg13g2_decap_8 FILLER_39_815 ();
 sg13g2_decap_8 FILLER_39_822 ();
 sg13g2_decap_8 FILLER_39_829 ();
 sg13g2_decap_8 FILLER_39_836 ();
 sg13g2_decap_8 FILLER_39_843 ();
 sg13g2_decap_8 FILLER_39_850 ();
 sg13g2_decap_4 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_decap_8 FILLER_40_156 ();
 sg13g2_decap_4 FILLER_40_163 ();
 sg13g2_fill_1 FILLER_40_167 ();
 sg13g2_fill_2 FILLER_40_203 ();
 sg13g2_fill_1 FILLER_40_205 ();
 sg13g2_fill_2 FILLER_40_222 ();
 sg13g2_fill_1 FILLER_40_229 ();
 sg13g2_fill_2 FILLER_40_236 ();
 sg13g2_fill_1 FILLER_40_259 ();
 sg13g2_fill_2 FILLER_40_274 ();
 sg13g2_fill_1 FILLER_40_276 ();
 sg13g2_decap_8 FILLER_40_290 ();
 sg13g2_fill_1 FILLER_40_297 ();
 sg13g2_decap_8 FILLER_40_314 ();
 sg13g2_fill_2 FILLER_40_321 ();
 sg13g2_fill_1 FILLER_40_333 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_fill_2 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_406 ();
 sg13g2_decap_4 FILLER_40_412 ();
 sg13g2_fill_1 FILLER_40_416 ();
 sg13g2_decap_8 FILLER_40_438 ();
 sg13g2_decap_4 FILLER_40_445 ();
 sg13g2_decap_8 FILLER_40_454 ();
 sg13g2_decap_4 FILLER_40_461 ();
 sg13g2_fill_2 FILLER_40_487 ();
 sg13g2_fill_1 FILLER_40_489 ();
 sg13g2_decap_4 FILLER_40_521 ();
 sg13g2_fill_2 FILLER_40_551 ();
 sg13g2_fill_1 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_697 ();
 sg13g2_decap_8 FILLER_40_704 ();
 sg13g2_decap_8 FILLER_40_711 ();
 sg13g2_decap_8 FILLER_40_718 ();
 sg13g2_decap_8 FILLER_40_725 ();
 sg13g2_decap_8 FILLER_40_732 ();
 sg13g2_decap_8 FILLER_40_739 ();
 sg13g2_decap_8 FILLER_40_746 ();
 sg13g2_decap_8 FILLER_40_753 ();
 sg13g2_decap_8 FILLER_40_760 ();
 sg13g2_decap_8 FILLER_40_767 ();
 sg13g2_decap_8 FILLER_40_774 ();
 sg13g2_decap_8 FILLER_40_781 ();
 sg13g2_decap_8 FILLER_40_788 ();
 sg13g2_decap_8 FILLER_40_795 ();
 sg13g2_decap_8 FILLER_40_802 ();
 sg13g2_decap_8 FILLER_40_809 ();
 sg13g2_decap_8 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_40_823 ();
 sg13g2_decap_8 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_837 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_4 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_4 FILLER_41_70 ();
 sg13g2_decap_4 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_102 ();
 sg13g2_fill_2 FILLER_41_108 ();
 sg13g2_fill_1 FILLER_41_110 ();
 sg13g2_fill_2 FILLER_41_128 ();
 sg13g2_fill_1 FILLER_41_144 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_fill_1 FILLER_41_177 ();
 sg13g2_fill_2 FILLER_41_199 ();
 sg13g2_fill_1 FILLER_41_201 ();
 sg13g2_fill_2 FILLER_41_228 ();
 sg13g2_fill_2 FILLER_41_257 ();
 sg13g2_fill_1 FILLER_41_259 ();
 sg13g2_fill_2 FILLER_41_265 ();
 sg13g2_fill_1 FILLER_41_267 ();
 sg13g2_fill_2 FILLER_41_289 ();
 sg13g2_fill_1 FILLER_41_291 ();
 sg13g2_fill_2 FILLER_41_297 ();
 sg13g2_fill_1 FILLER_41_299 ();
 sg13g2_fill_2 FILLER_41_313 ();
 sg13g2_fill_1 FILLER_41_315 ();
 sg13g2_fill_2 FILLER_41_342 ();
 sg13g2_fill_1 FILLER_41_344 ();
 sg13g2_fill_2 FILLER_41_362 ();
 sg13g2_decap_8 FILLER_41_394 ();
 sg13g2_fill_2 FILLER_41_401 ();
 sg13g2_fill_2 FILLER_41_419 ();
 sg13g2_fill_1 FILLER_41_421 ();
 sg13g2_fill_2 FILLER_41_438 ();
 sg13g2_fill_2 FILLER_41_445 ();
 sg13g2_fill_2 FILLER_41_495 ();
 sg13g2_fill_2 FILLER_41_533 ();
 sg13g2_fill_1 FILLER_41_535 ();
 sg13g2_fill_2 FILLER_41_549 ();
 sg13g2_fill_2 FILLER_41_575 ();
 sg13g2_fill_2 FILLER_41_592 ();
 sg13g2_fill_2 FILLER_41_609 ();
 sg13g2_fill_1 FILLER_41_627 ();
 sg13g2_fill_2 FILLER_41_637 ();
 sg13g2_fill_1 FILLER_41_648 ();
 sg13g2_fill_2 FILLER_41_677 ();
 sg13g2_decap_8 FILLER_41_713 ();
 sg13g2_decap_8 FILLER_41_720 ();
 sg13g2_decap_8 FILLER_41_727 ();
 sg13g2_decap_8 FILLER_41_734 ();
 sg13g2_decap_8 FILLER_41_741 ();
 sg13g2_decap_8 FILLER_41_748 ();
 sg13g2_decap_8 FILLER_41_755 ();
 sg13g2_decap_8 FILLER_41_762 ();
 sg13g2_decap_8 FILLER_41_769 ();
 sg13g2_decap_8 FILLER_41_776 ();
 sg13g2_decap_8 FILLER_41_783 ();
 sg13g2_decap_8 FILLER_41_790 ();
 sg13g2_decap_8 FILLER_41_797 ();
 sg13g2_decap_8 FILLER_41_804 ();
 sg13g2_decap_8 FILLER_41_811 ();
 sg13g2_decap_8 FILLER_41_818 ();
 sg13g2_decap_8 FILLER_41_825 ();
 sg13g2_decap_8 FILLER_41_832 ();
 sg13g2_decap_8 FILLER_41_839 ();
 sg13g2_decap_8 FILLER_41_846 ();
 sg13g2_decap_8 FILLER_41_853 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_133 ();
 sg13g2_fill_1 FILLER_42_135 ();
 sg13g2_fill_2 FILLER_42_172 ();
 sg13g2_fill_1 FILLER_42_183 ();
 sg13g2_decap_4 FILLER_42_207 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_fill_2 FILLER_42_269 ();
 sg13g2_fill_1 FILLER_42_271 ();
 sg13g2_fill_1 FILLER_42_298 ();
 sg13g2_decap_8 FILLER_42_305 ();
 sg13g2_decap_4 FILLER_42_312 ();
 sg13g2_fill_2 FILLER_42_344 ();
 sg13g2_fill_2 FILLER_42_371 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_fill_1 FILLER_42_410 ();
 sg13g2_fill_2 FILLER_42_450 ();
 sg13g2_fill_1 FILLER_42_452 ();
 sg13g2_decap_4 FILLER_42_458 ();
 sg13g2_fill_1 FILLER_42_462 ();
 sg13g2_fill_2 FILLER_42_479 ();
 sg13g2_fill_1 FILLER_42_481 ();
 sg13g2_decap_4 FILLER_42_512 ();
 sg13g2_fill_1 FILLER_42_527 ();
 sg13g2_fill_2 FILLER_42_537 ();
 sg13g2_fill_1 FILLER_42_539 ();
 sg13g2_decap_4 FILLER_42_545 ();
 sg13g2_fill_2 FILLER_42_588 ();
 sg13g2_fill_2 FILLER_42_615 ();
 sg13g2_fill_1 FILLER_42_617 ();
 sg13g2_fill_1 FILLER_42_649 ();
 sg13g2_fill_2 FILLER_42_665 ();
 sg13g2_fill_1 FILLER_42_667 ();
 sg13g2_decap_8 FILLER_42_721 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_826 ();
 sg13g2_decap_8 FILLER_42_833 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_fill_2 FILLER_43_42 ();
 sg13g2_fill_2 FILLER_43_51 ();
 sg13g2_fill_2 FILLER_43_58 ();
 sg13g2_fill_1 FILLER_43_60 ();
 sg13g2_decap_4 FILLER_43_65 ();
 sg13g2_decap_8 FILLER_43_72 ();
 sg13g2_decap_8 FILLER_43_79 ();
 sg13g2_decap_4 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_116 ();
 sg13g2_fill_2 FILLER_43_122 ();
 sg13g2_fill_1 FILLER_43_124 ();
 sg13g2_fill_1 FILLER_43_131 ();
 sg13g2_decap_4 FILLER_43_144 ();
 sg13g2_fill_2 FILLER_43_148 ();
 sg13g2_fill_2 FILLER_43_155 ();
 sg13g2_decap_4 FILLER_43_161 ();
 sg13g2_decap_4 FILLER_43_210 ();
 sg13g2_fill_2 FILLER_43_240 ();
 sg13g2_fill_1 FILLER_43_248 ();
 sg13g2_fill_2 FILLER_43_263 ();
 sg13g2_fill_2 FILLER_43_302 ();
 sg13g2_fill_2 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_368 ();
 sg13g2_decap_4 FILLER_43_450 ();
 sg13g2_fill_2 FILLER_43_480 ();
 sg13g2_fill_1 FILLER_43_482 ();
 sg13g2_fill_2 FILLER_43_515 ();
 sg13g2_fill_1 FILLER_43_517 ();
 sg13g2_fill_1 FILLER_43_580 ();
 sg13g2_fill_2 FILLER_43_616 ();
 sg13g2_fill_1 FILLER_43_618 ();
 sg13g2_fill_2 FILLER_43_646 ();
 sg13g2_fill_2 FILLER_43_656 ();
 sg13g2_fill_1 FILLER_43_684 ();
 sg13g2_decap_8 FILLER_43_722 ();
 sg13g2_decap_8 FILLER_43_729 ();
 sg13g2_decap_8 FILLER_43_736 ();
 sg13g2_decap_8 FILLER_43_743 ();
 sg13g2_decap_8 FILLER_43_750 ();
 sg13g2_decap_8 FILLER_43_757 ();
 sg13g2_decap_8 FILLER_43_764 ();
 sg13g2_decap_8 FILLER_43_771 ();
 sg13g2_decap_8 FILLER_43_778 ();
 sg13g2_decap_8 FILLER_43_785 ();
 sg13g2_decap_8 FILLER_43_792 ();
 sg13g2_decap_8 FILLER_43_799 ();
 sg13g2_decap_8 FILLER_43_806 ();
 sg13g2_decap_8 FILLER_43_813 ();
 sg13g2_decap_8 FILLER_43_820 ();
 sg13g2_decap_8 FILLER_43_827 ();
 sg13g2_decap_8 FILLER_43_834 ();
 sg13g2_decap_8 FILLER_43_841 ();
 sg13g2_decap_8 FILLER_43_848 ();
 sg13g2_decap_8 FILLER_43_855 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_14 ();
 sg13g2_fill_1 FILLER_44_16 ();
 sg13g2_fill_2 FILLER_44_43 ();
 sg13g2_fill_1 FILLER_44_85 ();
 sg13g2_decap_4 FILLER_44_109 ();
 sg13g2_fill_2 FILLER_44_116 ();
 sg13g2_decap_8 FILLER_44_129 ();
 sg13g2_fill_2 FILLER_44_136 ();
 sg13g2_fill_1 FILLER_44_138 ();
 sg13g2_fill_2 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_4 FILLER_44_168 ();
 sg13g2_fill_2 FILLER_44_172 ();
 sg13g2_decap_4 FILLER_44_183 ();
 sg13g2_fill_2 FILLER_44_187 ();
 sg13g2_fill_1 FILLER_44_249 ();
 sg13g2_fill_1 FILLER_44_282 ();
 sg13g2_decap_4 FILLER_44_288 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_decap_8 FILLER_44_310 ();
 sg13g2_fill_1 FILLER_44_317 ();
 sg13g2_fill_1 FILLER_44_353 ();
 sg13g2_fill_1 FILLER_44_380 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_4 FILLER_44_392 ();
 sg13g2_fill_2 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_417 ();
 sg13g2_fill_2 FILLER_44_424 ();
 sg13g2_fill_1 FILLER_44_426 ();
 sg13g2_fill_2 FILLER_44_468 ();
 sg13g2_fill_1 FILLER_44_470 ();
 sg13g2_fill_2 FILLER_44_536 ();
 sg13g2_fill_1 FILLER_44_555 ();
 sg13g2_fill_1 FILLER_44_560 ();
 sg13g2_decap_4 FILLER_44_609 ();
 sg13g2_decap_4 FILLER_44_618 ();
 sg13g2_fill_1 FILLER_44_635 ();
 sg13g2_fill_2 FILLER_44_655 ();
 sg13g2_fill_1 FILLER_44_657 ();
 sg13g2_fill_2 FILLER_44_675 ();
 sg13g2_fill_1 FILLER_44_677 ();
 sg13g2_fill_1 FILLER_44_696 ();
 sg13g2_decap_8 FILLER_44_723 ();
 sg13g2_decap_8 FILLER_44_730 ();
 sg13g2_decap_8 FILLER_44_737 ();
 sg13g2_decap_8 FILLER_44_744 ();
 sg13g2_decap_8 FILLER_44_751 ();
 sg13g2_decap_8 FILLER_44_758 ();
 sg13g2_decap_8 FILLER_44_765 ();
 sg13g2_decap_8 FILLER_44_772 ();
 sg13g2_decap_8 FILLER_44_779 ();
 sg13g2_decap_8 FILLER_44_786 ();
 sg13g2_decap_8 FILLER_44_793 ();
 sg13g2_decap_8 FILLER_44_800 ();
 sg13g2_decap_8 FILLER_44_807 ();
 sg13g2_decap_8 FILLER_44_814 ();
 sg13g2_decap_8 FILLER_44_821 ();
 sg13g2_decap_8 FILLER_44_828 ();
 sg13g2_decap_8 FILLER_44_835 ();
 sg13g2_decap_8 FILLER_44_842 ();
 sg13g2_decap_8 FILLER_44_849 ();
 sg13g2_decap_4 FILLER_44_856 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_11 ();
 sg13g2_fill_2 FILLER_45_48 ();
 sg13g2_fill_2 FILLER_45_59 ();
 sg13g2_fill_1 FILLER_45_61 ();
 sg13g2_fill_2 FILLER_45_88 ();
 sg13g2_fill_1 FILLER_45_90 ();
 sg13g2_fill_2 FILLER_45_117 ();
 sg13g2_fill_1 FILLER_45_136 ();
 sg13g2_fill_1 FILLER_45_166 ();
 sg13g2_decap_8 FILLER_45_190 ();
 sg13g2_fill_1 FILLER_45_197 ();
 sg13g2_decap_8 FILLER_45_202 ();
 sg13g2_decap_8 FILLER_45_209 ();
 sg13g2_fill_2 FILLER_45_216 ();
 sg13g2_fill_1 FILLER_45_218 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_fill_2 FILLER_45_231 ();
 sg13g2_fill_1 FILLER_45_247 ();
 sg13g2_fill_2 FILLER_45_273 ();
 sg13g2_decap_4 FILLER_45_292 ();
 sg13g2_decap_4 FILLER_45_304 ();
 sg13g2_fill_1 FILLER_45_369 ();
 sg13g2_fill_2 FILLER_45_379 ();
 sg13g2_fill_1 FILLER_45_385 ();
 sg13g2_fill_2 FILLER_45_390 ();
 sg13g2_fill_1 FILLER_45_436 ();
 sg13g2_fill_1 FILLER_45_441 ();
 sg13g2_fill_1 FILLER_45_471 ();
 sg13g2_fill_2 FILLER_45_495 ();
 sg13g2_fill_1 FILLER_45_497 ();
 sg13g2_fill_2 FILLER_45_533 ();
 sg13g2_fill_2 FILLER_45_544 ();
 sg13g2_fill_1 FILLER_45_551 ();
 sg13g2_fill_1 FILLER_45_562 ();
 sg13g2_fill_2 FILLER_45_575 ();
 sg13g2_decap_8 FILLER_45_611 ();
 sg13g2_fill_2 FILLER_45_677 ();
 sg13g2_fill_2 FILLER_45_695 ();
 sg13g2_fill_1 FILLER_45_706 ();
 sg13g2_decap_8 FILLER_45_716 ();
 sg13g2_decap_8 FILLER_45_723 ();
 sg13g2_decap_8 FILLER_45_730 ();
 sg13g2_decap_8 FILLER_45_737 ();
 sg13g2_decap_8 FILLER_45_744 ();
 sg13g2_decap_8 FILLER_45_751 ();
 sg13g2_decap_8 FILLER_45_758 ();
 sg13g2_decap_8 FILLER_45_765 ();
 sg13g2_decap_8 FILLER_45_772 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_8 FILLER_45_786 ();
 sg13g2_decap_8 FILLER_45_793 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_decap_8 FILLER_45_807 ();
 sg13g2_decap_8 FILLER_45_814 ();
 sg13g2_decap_8 FILLER_45_821 ();
 sg13g2_decap_8 FILLER_45_828 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_4 FILLER_45_856 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_41 ();
 sg13g2_fill_1 FILLER_46_43 ();
 sg13g2_fill_1 FILLER_46_64 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_fill_2 FILLER_46_109 ();
 sg13g2_fill_1 FILLER_46_111 ();
 sg13g2_decap_4 FILLER_46_117 ();
 sg13g2_fill_1 FILLER_46_121 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_4 FILLER_46_133 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_4 FILLER_46_182 ();
 sg13g2_fill_1 FILLER_46_186 ();
 sg13g2_decap_8 FILLER_46_205 ();
 sg13g2_decap_8 FILLER_46_212 ();
 sg13g2_fill_2 FILLER_46_219 ();
 sg13g2_fill_1 FILLER_46_226 ();
 sg13g2_fill_1 FILLER_46_233 ();
 sg13g2_decap_8 FILLER_46_265 ();
 sg13g2_decap_4 FILLER_46_296 ();
 sg13g2_fill_2 FILLER_46_321 ();
 sg13g2_fill_1 FILLER_46_346 ();
 sg13g2_decap_4 FILLER_46_361 ();
 sg13g2_fill_1 FILLER_46_365 ();
 sg13g2_fill_2 FILLER_46_373 ();
 sg13g2_fill_1 FILLER_46_375 ();
 sg13g2_fill_1 FILLER_46_416 ();
 sg13g2_fill_1 FILLER_46_463 ();
 sg13g2_fill_2 FILLER_46_469 ();
 sg13g2_fill_2 FILLER_46_481 ();
 sg13g2_fill_2 FILLER_46_506 ();
 sg13g2_fill_2 FILLER_46_544 ();
 sg13g2_fill_1 FILLER_46_551 ();
 sg13g2_fill_2 FILLER_46_577 ();
 sg13g2_fill_2 FILLER_46_611 ();
 sg13g2_fill_1 FILLER_46_613 ();
 sg13g2_fill_2 FILLER_46_647 ();
 sg13g2_fill_2 FILLER_46_671 ();
 sg13g2_fill_1 FILLER_46_673 ();
 sg13g2_fill_2 FILLER_46_682 ();
 sg13g2_fill_1 FILLER_46_684 ();
 sg13g2_fill_1 FILLER_46_694 ();
 sg13g2_decap_8 FILLER_46_708 ();
 sg13g2_decap_8 FILLER_46_715 ();
 sg13g2_decap_8 FILLER_46_722 ();
 sg13g2_decap_8 FILLER_46_729 ();
 sg13g2_decap_8 FILLER_46_736 ();
 sg13g2_decap_8 FILLER_46_743 ();
 sg13g2_decap_8 FILLER_46_750 ();
 sg13g2_decap_8 FILLER_46_757 ();
 sg13g2_decap_8 FILLER_46_764 ();
 sg13g2_decap_8 FILLER_46_771 ();
 sg13g2_decap_8 FILLER_46_778 ();
 sg13g2_decap_8 FILLER_46_785 ();
 sg13g2_decap_8 FILLER_46_792 ();
 sg13g2_decap_8 FILLER_46_799 ();
 sg13g2_decap_8 FILLER_46_806 ();
 sg13g2_decap_8 FILLER_46_813 ();
 sg13g2_decap_8 FILLER_46_820 ();
 sg13g2_decap_8 FILLER_46_827 ();
 sg13g2_decap_8 FILLER_46_834 ();
 sg13g2_decap_8 FILLER_46_841 ();
 sg13g2_decap_8 FILLER_46_848 ();
 sg13g2_decap_8 FILLER_46_855 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_38 ();
 sg13g2_fill_2 FILLER_47_74 ();
 sg13g2_fill_2 FILLER_47_89 ();
 sg13g2_fill_1 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_113 ();
 sg13g2_fill_2 FILLER_47_132 ();
 sg13g2_fill_1 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_147 ();
 sg13g2_decap_4 FILLER_47_161 ();
 sg13g2_fill_2 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_214 ();
 sg13g2_decap_4 FILLER_47_240 ();
 sg13g2_fill_2 FILLER_47_244 ();
 sg13g2_decap_8 FILLER_47_250 ();
 sg13g2_decap_8 FILLER_47_267 ();
 sg13g2_fill_1 FILLER_47_274 ();
 sg13g2_decap_8 FILLER_47_295 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_decap_8 FILLER_47_316 ();
 sg13g2_fill_2 FILLER_47_347 ();
 sg13g2_fill_1 FILLER_47_365 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_fill_2 FILLER_47_392 ();
 sg13g2_fill_2 FILLER_47_403 ();
 sg13g2_fill_1 FILLER_47_422 ();
 sg13g2_fill_2 FILLER_47_434 ();
 sg13g2_fill_2 FILLER_47_444 ();
 sg13g2_fill_1 FILLER_47_477 ();
 sg13g2_fill_2 FILLER_47_494 ();
 sg13g2_fill_1 FILLER_47_506 ();
 sg13g2_fill_2 FILLER_47_521 ();
 sg13g2_fill_1 FILLER_47_523 ();
 sg13g2_fill_1 FILLER_47_532 ();
 sg13g2_fill_2 FILLER_47_542 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_decap_4 FILLER_47_579 ();
 sg13g2_fill_1 FILLER_47_609 ();
 sg13g2_fill_2 FILLER_47_613 ();
 sg13g2_fill_1 FILLER_47_615 ();
 sg13g2_decap_4 FILLER_47_659 ();
 sg13g2_fill_1 FILLER_47_663 ();
 sg13g2_fill_2 FILLER_47_683 ();
 sg13g2_decap_8 FILLER_47_711 ();
 sg13g2_decap_8 FILLER_47_718 ();
 sg13g2_decap_8 FILLER_47_725 ();
 sg13g2_decap_8 FILLER_47_732 ();
 sg13g2_decap_8 FILLER_47_739 ();
 sg13g2_decap_8 FILLER_47_746 ();
 sg13g2_decap_8 FILLER_47_753 ();
 sg13g2_decap_8 FILLER_47_760 ();
 sg13g2_decap_8 FILLER_47_767 ();
 sg13g2_decap_8 FILLER_47_774 ();
 sg13g2_decap_8 FILLER_47_781 ();
 sg13g2_decap_8 FILLER_47_788 ();
 sg13g2_decap_8 FILLER_47_795 ();
 sg13g2_decap_8 FILLER_47_802 ();
 sg13g2_decap_8 FILLER_47_809 ();
 sg13g2_decap_8 FILLER_47_816 ();
 sg13g2_decap_8 FILLER_47_823 ();
 sg13g2_decap_8 FILLER_47_830 ();
 sg13g2_decap_8 FILLER_47_837 ();
 sg13g2_decap_8 FILLER_47_844 ();
 sg13g2_decap_8 FILLER_47_851 ();
 sg13g2_decap_4 FILLER_47_858 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_27 ();
 sg13g2_fill_1 FILLER_48_29 ();
 sg13g2_decap_4 FILLER_48_56 ();
 sg13g2_fill_1 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_76 ();
 sg13g2_decap_4 FILLER_48_83 ();
 sg13g2_decap_8 FILLER_48_94 ();
 sg13g2_decap_8 FILLER_48_101 ();
 sg13g2_decap_4 FILLER_48_108 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_decap_4 FILLER_48_117 ();
 sg13g2_decap_4 FILLER_48_129 ();
 sg13g2_fill_1 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_fill_2 FILLER_48_161 ();
 sg13g2_decap_4 FILLER_48_183 ();
 sg13g2_decap_4 FILLER_48_214 ();
 sg13g2_fill_2 FILLER_48_218 ();
 sg13g2_fill_1 FILLER_48_223 ();
 sg13g2_decap_8 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_fill_2 FILLER_48_293 ();
 sg13g2_fill_1 FILLER_48_295 ();
 sg13g2_decap_4 FILLER_48_326 ();
 sg13g2_fill_1 FILLER_48_338 ();
 sg13g2_fill_2 FILLER_48_347 ();
 sg13g2_decap_8 FILLER_48_354 ();
 sg13g2_decap_4 FILLER_48_361 ();
 sg13g2_fill_2 FILLER_48_365 ();
 sg13g2_fill_1 FILLER_48_372 ();
 sg13g2_fill_2 FILLER_48_386 ();
 sg13g2_fill_1 FILLER_48_419 ();
 sg13g2_fill_1 FILLER_48_432 ();
 sg13g2_fill_2 FILLER_48_437 ();
 sg13g2_fill_1 FILLER_48_439 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_4 FILLER_48_483 ();
 sg13g2_fill_1 FILLER_48_508 ();
 sg13g2_decap_4 FILLER_48_585 ();
 sg13g2_fill_2 FILLER_48_589 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_fill_2 FILLER_48_602 ();
 sg13g2_fill_1 FILLER_48_624 ();
 sg13g2_fill_2 FILLER_48_650 ();
 sg13g2_decap_4 FILLER_48_668 ();
 sg13g2_fill_2 FILLER_48_677 ();
 sg13g2_fill_2 FILLER_48_687 ();
 sg13g2_fill_1 FILLER_48_689 ();
 sg13g2_fill_2 FILLER_48_694 ();
 sg13g2_decap_8 FILLER_48_705 ();
 sg13g2_decap_8 FILLER_48_712 ();
 sg13g2_decap_8 FILLER_48_719 ();
 sg13g2_decap_8 FILLER_48_726 ();
 sg13g2_decap_8 FILLER_48_733 ();
 sg13g2_decap_8 FILLER_48_740 ();
 sg13g2_decap_8 FILLER_48_747 ();
 sg13g2_decap_8 FILLER_48_754 ();
 sg13g2_decap_8 FILLER_48_761 ();
 sg13g2_decap_8 FILLER_48_768 ();
 sg13g2_decap_8 FILLER_48_775 ();
 sg13g2_decap_8 FILLER_48_782 ();
 sg13g2_decap_8 FILLER_48_789 ();
 sg13g2_decap_8 FILLER_48_796 ();
 sg13g2_decap_8 FILLER_48_803 ();
 sg13g2_decap_8 FILLER_48_810 ();
 sg13g2_decap_8 FILLER_48_817 ();
 sg13g2_decap_8 FILLER_48_824 ();
 sg13g2_decap_8 FILLER_48_831 ();
 sg13g2_decap_8 FILLER_48_838 ();
 sg13g2_decap_8 FILLER_48_845 ();
 sg13g2_decap_8 FILLER_48_852 ();
 sg13g2_fill_2 FILLER_48_859 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_4 ();
 sg13g2_fill_1 FILLER_49_53 ();
 sg13g2_fill_1 FILLER_49_87 ();
 sg13g2_fill_2 FILLER_49_117 ();
 sg13g2_decap_4 FILLER_49_124 ();
 sg13g2_fill_1 FILLER_49_128 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_decap_8 FILLER_49_156 ();
 sg13g2_fill_2 FILLER_49_163 ();
 sg13g2_fill_1 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_180 ();
 sg13g2_fill_2 FILLER_49_187 ();
 sg13g2_fill_2 FILLER_49_195 ();
 sg13g2_decap_8 FILLER_49_216 ();
 sg13g2_decap_4 FILLER_49_223 ();
 sg13g2_fill_2 FILLER_49_233 ();
 sg13g2_fill_1 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_262 ();
 sg13g2_decap_4 FILLER_49_269 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_300 ();
 sg13g2_decap_8 FILLER_49_307 ();
 sg13g2_fill_2 FILLER_49_319 ();
 sg13g2_fill_1 FILLER_49_345 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_2 FILLER_49_429 ();
 sg13g2_decap_8 FILLER_49_457 ();
 sg13g2_fill_1 FILLER_49_472 ();
 sg13g2_decap_4 FILLER_49_479 ();
 sg13g2_fill_1 FILLER_49_483 ();
 sg13g2_decap_4 FILLER_49_534 ();
 sg13g2_fill_1 FILLER_49_538 ();
 sg13g2_fill_1 FILLER_49_549 ();
 sg13g2_fill_2 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_587 ();
 sg13g2_decap_4 FILLER_49_594 ();
 sg13g2_fill_2 FILLER_49_598 ();
 sg13g2_fill_1 FILLER_49_626 ();
 sg13g2_fill_1 FILLER_49_649 ();
 sg13g2_decap_8 FILLER_49_731 ();
 sg13g2_decap_8 FILLER_49_738 ();
 sg13g2_decap_8 FILLER_49_745 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_decap_8 FILLER_49_759 ();
 sg13g2_decap_8 FILLER_49_766 ();
 sg13g2_decap_8 FILLER_49_773 ();
 sg13g2_decap_8 FILLER_49_780 ();
 sg13g2_decap_8 FILLER_49_787 ();
 sg13g2_decap_8 FILLER_49_794 ();
 sg13g2_decap_8 FILLER_49_801 ();
 sg13g2_decap_8 FILLER_49_808 ();
 sg13g2_decap_8 FILLER_49_815 ();
 sg13g2_decap_8 FILLER_49_822 ();
 sg13g2_decap_8 FILLER_49_829 ();
 sg13g2_decap_8 FILLER_49_836 ();
 sg13g2_decap_8 FILLER_49_843 ();
 sg13g2_decap_8 FILLER_49_850 ();
 sg13g2_decap_4 FILLER_49_857 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_58 ();
 sg13g2_fill_1 FILLER_50_63 ();
 sg13g2_fill_1 FILLER_50_81 ();
 sg13g2_fill_1 FILLER_50_105 ();
 sg13g2_decap_4 FILLER_50_127 ();
 sg13g2_fill_2 FILLER_50_131 ();
 sg13g2_fill_2 FILLER_50_163 ();
 sg13g2_fill_2 FILLER_50_189 ();
 sg13g2_fill_1 FILLER_50_191 ();
 sg13g2_decap_8 FILLER_50_263 ();
 sg13g2_fill_1 FILLER_50_270 ();
 sg13g2_fill_2 FILLER_50_296 ();
 sg13g2_fill_2 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_325 ();
 sg13g2_decap_8 FILLER_50_332 ();
 sg13g2_fill_2 FILLER_50_339 ();
 sg13g2_fill_2 FILLER_50_382 ();
 sg13g2_fill_1 FILLER_50_384 ();
 sg13g2_fill_2 FILLER_50_410 ();
 sg13g2_fill_1 FILLER_50_416 ();
 sg13g2_fill_2 FILLER_50_426 ();
 sg13g2_decap_4 FILLER_50_432 ();
 sg13g2_fill_2 FILLER_50_443 ();
 sg13g2_decap_4 FILLER_50_449 ();
 sg13g2_decap_4 FILLER_50_477 ();
 sg13g2_fill_1 FILLER_50_490 ();
 sg13g2_decap_8 FILLER_50_500 ();
 sg13g2_decap_4 FILLER_50_507 ();
 sg13g2_decap_4 FILLER_50_525 ();
 sg13g2_decap_4 FILLER_50_533 ();
 sg13g2_fill_2 FILLER_50_537 ();
 sg13g2_decap_8 FILLER_50_568 ();
 sg13g2_decap_4 FILLER_50_575 ();
 sg13g2_fill_2 FILLER_50_614 ();
 sg13g2_fill_1 FILLER_50_616 ();
 sg13g2_decap_4 FILLER_50_634 ();
 sg13g2_fill_2 FILLER_50_661 ();
 sg13g2_decap_8 FILLER_50_692 ();
 sg13g2_decap_4 FILLER_50_699 ();
 sg13g2_fill_1 FILLER_50_708 ();
 sg13g2_fill_1 FILLER_50_712 ();
 sg13g2_decap_4 FILLER_50_717 ();
 sg13g2_decap_8 FILLER_50_730 ();
 sg13g2_decap_8 FILLER_50_737 ();
 sg13g2_decap_8 FILLER_50_744 ();
 sg13g2_decap_8 FILLER_50_751 ();
 sg13g2_decap_8 FILLER_50_758 ();
 sg13g2_decap_8 FILLER_50_765 ();
 sg13g2_decap_8 FILLER_50_772 ();
 sg13g2_decap_8 FILLER_50_779 ();
 sg13g2_decap_8 FILLER_50_786 ();
 sg13g2_decap_8 FILLER_50_793 ();
 sg13g2_decap_8 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_807 ();
 sg13g2_decap_8 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_821 ();
 sg13g2_decap_8 FILLER_50_828 ();
 sg13g2_decap_8 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_842 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_fill_2 FILLER_51_34 ();
 sg13g2_fill_1 FILLER_51_36 ();
 sg13g2_fill_2 FILLER_51_72 ();
 sg13g2_decap_8 FILLER_51_95 ();
 sg13g2_decap_8 FILLER_51_115 ();
 sg13g2_decap_8 FILLER_51_122 ();
 sg13g2_decap_8 FILLER_51_129 ();
 sg13g2_fill_1 FILLER_51_136 ();
 sg13g2_decap_8 FILLER_51_158 ();
 sg13g2_decap_4 FILLER_51_165 ();
 sg13g2_fill_2 FILLER_51_169 ();
 sg13g2_fill_1 FILLER_51_176 ();
 sg13g2_fill_1 FILLER_51_253 ();
 sg13g2_fill_2 FILLER_51_267 ();
 sg13g2_decap_8 FILLER_51_273 ();
 sg13g2_fill_2 FILLER_51_280 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_fill_2 FILLER_51_287 ();
 sg13g2_fill_2 FILLER_51_301 ();
 sg13g2_fill_1 FILLER_51_303 ();
 sg13g2_fill_2 FILLER_51_309 ();
 sg13g2_fill_1 FILLER_51_311 ();
 sg13g2_decap_4 FILLER_51_317 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_decap_8 FILLER_51_376 ();
 sg13g2_decap_4 FILLER_51_383 ();
 sg13g2_fill_1 FILLER_51_394 ();
 sg13g2_fill_1 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_414 ();
 sg13g2_fill_1 FILLER_51_416 ();
 sg13g2_fill_2 FILLER_51_443 ();
 sg13g2_decap_8 FILLER_51_448 ();
 sg13g2_decap_4 FILLER_51_484 ();
 sg13g2_fill_1 FILLER_51_518 ();
 sg13g2_fill_2 FILLER_51_603 ();
 sg13g2_fill_2 FILLER_51_617 ();
 sg13g2_fill_2 FILLER_51_645 ();
 sg13g2_fill_1 FILLER_51_655 ();
 sg13g2_fill_2 FILLER_51_675 ();
 sg13g2_fill_2 FILLER_51_693 ();
 sg13g2_fill_1 FILLER_51_700 ();
 sg13g2_fill_2 FILLER_51_729 ();
 sg13g2_fill_1 FILLER_51_731 ();
 sg13g2_decap_8 FILLER_51_740 ();
 sg13g2_decap_8 FILLER_51_747 ();
 sg13g2_decap_8 FILLER_51_754 ();
 sg13g2_decap_8 FILLER_51_761 ();
 sg13g2_decap_8 FILLER_51_768 ();
 sg13g2_decap_8 FILLER_51_775 ();
 sg13g2_decap_8 FILLER_51_782 ();
 sg13g2_decap_8 FILLER_51_789 ();
 sg13g2_decap_8 FILLER_51_796 ();
 sg13g2_decap_8 FILLER_51_803 ();
 sg13g2_decap_8 FILLER_51_810 ();
 sg13g2_decap_8 FILLER_51_817 ();
 sg13g2_decap_8 FILLER_51_824 ();
 sg13g2_decap_8 FILLER_51_831 ();
 sg13g2_decap_8 FILLER_51_838 ();
 sg13g2_decap_8 FILLER_51_845 ();
 sg13g2_decap_8 FILLER_51_852 ();
 sg13g2_fill_2 FILLER_51_859 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_24 ();
 sg13g2_fill_2 FILLER_52_53 ();
 sg13g2_fill_1 FILLER_52_55 ();
 sg13g2_decap_4 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_decap_4 FILLER_52_100 ();
 sg13g2_decap_4 FILLER_52_136 ();
 sg13g2_fill_2 FILLER_52_153 ();
 sg13g2_fill_1 FILLER_52_155 ();
 sg13g2_fill_2 FILLER_52_244 ();
 sg13g2_fill_1 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_251 ();
 sg13g2_decap_4 FILLER_52_258 ();
 sg13g2_fill_1 FILLER_52_262 ();
 sg13g2_decap_4 FILLER_52_283 ();
 sg13g2_fill_1 FILLER_52_287 ();
 sg13g2_decap_4 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_315 ();
 sg13g2_fill_2 FILLER_52_358 ();
 sg13g2_fill_1 FILLER_52_370 ();
 sg13g2_fill_2 FILLER_52_400 ();
 sg13g2_fill_1 FILLER_52_421 ();
 sg13g2_decap_8 FILLER_52_426 ();
 sg13g2_decap_4 FILLER_52_433 ();
 sg13g2_fill_1 FILLER_52_437 ();
 sg13g2_fill_2 FILLER_52_446 ();
 sg13g2_decap_8 FILLER_52_462 ();
 sg13g2_decap_8 FILLER_52_474 ();
 sg13g2_decap_4 FILLER_52_481 ();
 sg13g2_fill_2 FILLER_52_485 ();
 sg13g2_decap_8 FILLER_52_492 ();
 sg13g2_decap_8 FILLER_52_503 ();
 sg13g2_fill_2 FILLER_52_510 ();
 sg13g2_fill_1 FILLER_52_553 ();
 sg13g2_fill_1 FILLER_52_559 ();
 sg13g2_fill_2 FILLER_52_575 ();
 sg13g2_fill_1 FILLER_52_577 ();
 sg13g2_fill_2 FILLER_52_586 ();
 sg13g2_fill_1 FILLER_52_588 ();
 sg13g2_fill_1 FILLER_52_630 ();
 sg13g2_fill_2 FILLER_52_645 ();
 sg13g2_fill_2 FILLER_52_664 ();
 sg13g2_fill_1 FILLER_52_666 ();
 sg13g2_fill_2 FILLER_52_688 ();
 sg13g2_decap_4 FILLER_52_695 ();
 sg13g2_fill_1 FILLER_52_699 ();
 sg13g2_decap_4 FILLER_52_712 ();
 sg13g2_fill_2 FILLER_52_716 ();
 sg13g2_fill_2 FILLER_52_732 ();
 sg13g2_fill_1 FILLER_52_734 ();
 sg13g2_decap_8 FILLER_52_768 ();
 sg13g2_decap_8 FILLER_52_775 ();
 sg13g2_decap_8 FILLER_52_782 ();
 sg13g2_decap_8 FILLER_52_789 ();
 sg13g2_decap_8 FILLER_52_796 ();
 sg13g2_decap_8 FILLER_52_803 ();
 sg13g2_decap_8 FILLER_52_810 ();
 sg13g2_decap_8 FILLER_52_817 ();
 sg13g2_decap_8 FILLER_52_824 ();
 sg13g2_decap_8 FILLER_52_831 ();
 sg13g2_decap_8 FILLER_52_838 ();
 sg13g2_decap_8 FILLER_52_845 ();
 sg13g2_decap_8 FILLER_52_852 ();
 sg13g2_fill_2 FILLER_52_859 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_fill_2 FILLER_53_31 ();
 sg13g2_fill_1 FILLER_53_33 ();
 sg13g2_fill_2 FILLER_53_53 ();
 sg13g2_fill_1 FILLER_53_55 ();
 sg13g2_fill_2 FILLER_53_64 ();
 sg13g2_fill_1 FILLER_53_66 ();
 sg13g2_fill_2 FILLER_53_80 ();
 sg13g2_fill_1 FILLER_53_82 ();
 sg13g2_decap_4 FILLER_53_101 ();
 sg13g2_fill_2 FILLER_53_105 ();
 sg13g2_fill_1 FILLER_53_115 ();
 sg13g2_fill_1 FILLER_53_129 ();
 sg13g2_fill_2 FILLER_53_138 ();
 sg13g2_fill_1 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_156 ();
 sg13g2_fill_2 FILLER_53_172 ();
 sg13g2_fill_1 FILLER_53_193 ();
 sg13g2_fill_2 FILLER_53_256 ();
 sg13g2_fill_1 FILLER_53_258 ();
 sg13g2_fill_2 FILLER_53_264 ();
 sg13g2_decap_8 FILLER_53_284 ();
 sg13g2_fill_2 FILLER_53_291 ();
 sg13g2_fill_1 FILLER_53_293 ();
 sg13g2_decap_8 FILLER_53_299 ();
 sg13g2_decap_8 FILLER_53_306 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_fill_2 FILLER_53_337 ();
 sg13g2_fill_1 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_353 ();
 sg13g2_fill_1 FILLER_53_360 ();
 sg13g2_fill_2 FILLER_53_396 ();
 sg13g2_fill_1 FILLER_53_437 ();
 sg13g2_fill_2 FILLER_53_473 ();
 sg13g2_fill_1 FILLER_53_475 ();
 sg13g2_fill_2 FILLER_53_488 ();
 sg13g2_fill_2 FILLER_53_507 ();
 sg13g2_fill_1 FILLER_53_509 ();
 sg13g2_fill_2 FILLER_53_541 ();
 sg13g2_fill_2 FILLER_53_552 ();
 sg13g2_fill_2 FILLER_53_567 ();
 sg13g2_fill_1 FILLER_53_569 ();
 sg13g2_fill_1 FILLER_53_588 ();
 sg13g2_fill_2 FILLER_53_598 ();
 sg13g2_fill_1 FILLER_53_604 ();
 sg13g2_fill_2 FILLER_53_610 ();
 sg13g2_fill_2 FILLER_53_620 ();
 sg13g2_decap_8 FILLER_53_635 ();
 sg13g2_fill_1 FILLER_53_642 ();
 sg13g2_fill_2 FILLER_53_647 ();
 sg13g2_fill_1 FILLER_53_649 ();
 sg13g2_fill_2 FILLER_53_668 ();
 sg13g2_fill_1 FILLER_53_683 ();
 sg13g2_fill_2 FILLER_53_688 ();
 sg13g2_decap_8 FILLER_53_702 ();
 sg13g2_fill_1 FILLER_53_709 ();
 sg13g2_fill_2 FILLER_53_713 ();
 sg13g2_fill_1 FILLER_53_715 ();
 sg13g2_fill_2 FILLER_53_721 ();
 sg13g2_decap_8 FILLER_53_759 ();
 sg13g2_decap_8 FILLER_53_766 ();
 sg13g2_decap_8 FILLER_53_773 ();
 sg13g2_decap_8 FILLER_53_780 ();
 sg13g2_decap_8 FILLER_53_787 ();
 sg13g2_decap_8 FILLER_53_794 ();
 sg13g2_decap_8 FILLER_53_801 ();
 sg13g2_decap_8 FILLER_53_808 ();
 sg13g2_decap_8 FILLER_53_815 ();
 sg13g2_decap_8 FILLER_53_822 ();
 sg13g2_decap_8 FILLER_53_829 ();
 sg13g2_decap_8 FILLER_53_836 ();
 sg13g2_decap_8 FILLER_53_843 ();
 sg13g2_decap_8 FILLER_53_850 ();
 sg13g2_decap_4 FILLER_53_857 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_19 ();
 sg13g2_fill_1 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_77 ();
 sg13g2_fill_1 FILLER_54_79 ();
 sg13g2_decap_8 FILLER_54_85 ();
 sg13g2_decap_8 FILLER_54_110 ();
 sg13g2_fill_2 FILLER_54_117 ();
 sg13g2_fill_1 FILLER_54_119 ();
 sg13g2_decap_4 FILLER_54_133 ();
 sg13g2_fill_2 FILLER_54_173 ();
 sg13g2_fill_2 FILLER_54_189 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_1 FILLER_54_246 ();
 sg13g2_fill_2 FILLER_54_285 ();
 sg13g2_fill_1 FILLER_54_333 ();
 sg13g2_fill_1 FILLER_54_367 ();
 sg13g2_fill_2 FILLER_54_374 ();
 sg13g2_fill_2 FILLER_54_398 ();
 sg13g2_fill_2 FILLER_54_406 ();
 sg13g2_fill_2 FILLER_54_421 ();
 sg13g2_fill_1 FILLER_54_431 ();
 sg13g2_fill_2 FILLER_54_442 ();
 sg13g2_decap_8 FILLER_54_461 ();
 sg13g2_fill_2 FILLER_54_468 ();
 sg13g2_fill_1 FILLER_54_470 ();
 sg13g2_fill_2 FILLER_54_484 ();
 sg13g2_fill_1 FILLER_54_486 ();
 sg13g2_fill_2 FILLER_54_499 ();
 sg13g2_fill_2 FILLER_54_518 ();
 sg13g2_fill_1 FILLER_54_520 ();
 sg13g2_decap_4 FILLER_54_534 ();
 sg13g2_fill_2 FILLER_54_538 ();
 sg13g2_decap_8 FILLER_54_560 ();
 sg13g2_decap_8 FILLER_54_567 ();
 sg13g2_fill_2 FILLER_54_574 ();
 sg13g2_fill_1 FILLER_54_576 ();
 sg13g2_fill_1 FILLER_54_587 ();
 sg13g2_decap_4 FILLER_54_592 ();
 sg13g2_fill_1 FILLER_54_596 ();
 sg13g2_fill_2 FILLER_54_620 ();
 sg13g2_fill_1 FILLER_54_622 ();
 sg13g2_fill_1 FILLER_54_631 ();
 sg13g2_decap_8 FILLER_54_670 ();
 sg13g2_decap_8 FILLER_54_677 ();
 sg13g2_decap_4 FILLER_54_697 ();
 sg13g2_fill_2 FILLER_54_701 ();
 sg13g2_decap_4 FILLER_54_726 ();
 sg13g2_fill_1 FILLER_54_730 ();
 sg13g2_fill_2 FILLER_54_748 ();
 sg13g2_fill_1 FILLER_54_759 ();
 sg13g2_decap_8 FILLER_54_767 ();
 sg13g2_decap_8 FILLER_54_774 ();
 sg13g2_decap_8 FILLER_54_781 ();
 sg13g2_decap_8 FILLER_54_788 ();
 sg13g2_decap_8 FILLER_54_795 ();
 sg13g2_decap_8 FILLER_54_802 ();
 sg13g2_decap_8 FILLER_54_809 ();
 sg13g2_decap_8 FILLER_54_816 ();
 sg13g2_decap_8 FILLER_54_823 ();
 sg13g2_decap_8 FILLER_54_830 ();
 sg13g2_decap_8 FILLER_54_837 ();
 sg13g2_decap_8 FILLER_54_844 ();
 sg13g2_decap_8 FILLER_54_851 ();
 sg13g2_decap_4 FILLER_54_858 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_43 ();
 sg13g2_fill_2 FILLER_55_57 ();
 sg13g2_decap_4 FILLER_55_92 ();
 sg13g2_fill_2 FILLER_55_96 ();
 sg13g2_decap_8 FILLER_55_111 ();
 sg13g2_fill_2 FILLER_55_118 ();
 sg13g2_fill_1 FILLER_55_120 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_fill_2 FILLER_55_154 ();
 sg13g2_fill_2 FILLER_55_255 ();
 sg13g2_fill_2 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_268 ();
 sg13g2_fill_1 FILLER_55_270 ();
 sg13g2_fill_2 FILLER_55_284 ();
 sg13g2_fill_1 FILLER_55_286 ();
 sg13g2_decap_4 FILLER_55_300 ();
 sg13g2_fill_2 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_328 ();
 sg13g2_fill_1 FILLER_55_342 ();
 sg13g2_fill_1 FILLER_55_351 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_fill_2 FILLER_55_426 ();
 sg13g2_fill_1 FILLER_55_428 ();
 sg13g2_fill_2 FILLER_55_448 ();
 sg13g2_fill_1 FILLER_55_463 ();
 sg13g2_fill_1 FILLER_55_498 ();
 sg13g2_decap_8 FILLER_55_507 ();
 sg13g2_decap_4 FILLER_55_538 ();
 sg13g2_fill_2 FILLER_55_571 ();
 sg13g2_decap_4 FILLER_55_589 ();
 sg13g2_decap_4 FILLER_55_613 ();
 sg13g2_fill_2 FILLER_55_617 ();
 sg13g2_fill_2 FILLER_55_641 ();
 sg13g2_decap_8 FILLER_55_647 ();
 sg13g2_fill_2 FILLER_55_654 ();
 sg13g2_fill_1 FILLER_55_656 ();
 sg13g2_decap_4 FILLER_55_665 ();
 sg13g2_fill_2 FILLER_55_669 ();
 sg13g2_decap_4 FILLER_55_683 ();
 sg13g2_fill_1 FILLER_55_692 ();
 sg13g2_decap_8 FILLER_55_698 ();
 sg13g2_fill_2 FILLER_55_705 ();
 sg13g2_fill_2 FILLER_55_712 ();
 sg13g2_fill_1 FILLER_55_714 ();
 sg13g2_fill_2 FILLER_55_728 ();
 sg13g2_fill_1 FILLER_55_730 ();
 sg13g2_decap_8 FILLER_55_775 ();
 sg13g2_decap_8 FILLER_55_782 ();
 sg13g2_decap_8 FILLER_55_789 ();
 sg13g2_decap_8 FILLER_55_796 ();
 sg13g2_decap_8 FILLER_55_803 ();
 sg13g2_decap_8 FILLER_55_810 ();
 sg13g2_decap_8 FILLER_55_817 ();
 sg13g2_decap_8 FILLER_55_824 ();
 sg13g2_decap_8 FILLER_55_831 ();
 sg13g2_decap_8 FILLER_55_838 ();
 sg13g2_decap_8 FILLER_55_845 ();
 sg13g2_decap_8 FILLER_55_852 ();
 sg13g2_fill_2 FILLER_55_859 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_decap_8 FILLER_56_72 ();
 sg13g2_fill_2 FILLER_56_79 ();
 sg13g2_fill_1 FILLER_56_81 ();
 sg13g2_fill_2 FILLER_56_87 ();
 sg13g2_fill_1 FILLER_56_89 ();
 sg13g2_decap_4 FILLER_56_107 ();
 sg13g2_fill_1 FILLER_56_111 ();
 sg13g2_fill_2 FILLER_56_118 ();
 sg13g2_fill_1 FILLER_56_120 ();
 sg13g2_fill_2 FILLER_56_147 ();
 sg13g2_fill_1 FILLER_56_159 ();
 sg13g2_decap_4 FILLER_56_204 ();
 sg13g2_decap_4 FILLER_56_212 ();
 sg13g2_fill_1 FILLER_56_232 ();
 sg13g2_decap_8 FILLER_56_251 ();
 sg13g2_fill_2 FILLER_56_282 ();
 sg13g2_fill_2 FILLER_56_289 ();
 sg13g2_fill_1 FILLER_56_296 ();
 sg13g2_fill_2 FILLER_56_307 ();
 sg13g2_fill_2 FILLER_56_374 ();
 sg13g2_fill_2 FILLER_56_381 ();
 sg13g2_decap_4 FILLER_56_416 ();
 sg13g2_decap_8 FILLER_56_424 ();
 sg13g2_decap_4 FILLER_56_431 ();
 sg13g2_fill_2 FILLER_56_440 ();
 sg13g2_decap_8 FILLER_56_446 ();
 sg13g2_decap_8 FILLER_56_453 ();
 sg13g2_decap_8 FILLER_56_460 ();
 sg13g2_fill_1 FILLER_56_467 ();
 sg13g2_decap_8 FILLER_56_472 ();
 sg13g2_decap_4 FILLER_56_479 ();
 sg13g2_fill_1 FILLER_56_483 ();
 sg13g2_decap_8 FILLER_56_510 ();
 sg13g2_decap_4 FILLER_56_517 ();
 sg13g2_fill_1 FILLER_56_521 ();
 sg13g2_decap_8 FILLER_56_543 ();
 sg13g2_fill_1 FILLER_56_550 ();
 sg13g2_fill_2 FILLER_56_564 ();
 sg13g2_decap_8 FILLER_56_613 ();
 sg13g2_fill_2 FILLER_56_620 ();
 sg13g2_fill_2 FILLER_56_630 ();
 sg13g2_fill_1 FILLER_56_646 ();
 sg13g2_fill_1 FILLER_56_663 ();
 sg13g2_decap_8 FILLER_56_720 ();
 sg13g2_decap_8 FILLER_56_727 ();
 sg13g2_fill_2 FILLER_56_734 ();
 sg13g2_fill_1 FILLER_56_748 ();
 sg13g2_decap_8 FILLER_56_757 ();
 sg13g2_decap_8 FILLER_56_768 ();
 sg13g2_decap_8 FILLER_56_775 ();
 sg13g2_decap_8 FILLER_56_782 ();
 sg13g2_decap_8 FILLER_56_789 ();
 sg13g2_decap_8 FILLER_56_796 ();
 sg13g2_decap_8 FILLER_56_803 ();
 sg13g2_decap_8 FILLER_56_810 ();
 sg13g2_decap_8 FILLER_56_817 ();
 sg13g2_decap_8 FILLER_56_824 ();
 sg13g2_decap_8 FILLER_56_831 ();
 sg13g2_decap_8 FILLER_56_838 ();
 sg13g2_decap_8 FILLER_56_845 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_4 ();
 sg13g2_fill_2 FILLER_57_49 ();
 sg13g2_fill_1 FILLER_57_51 ();
 sg13g2_fill_1 FILLER_57_64 ();
 sg13g2_fill_2 FILLER_57_78 ();
 sg13g2_fill_1 FILLER_57_80 ();
 sg13g2_fill_2 FILLER_57_94 ();
 sg13g2_fill_1 FILLER_57_96 ();
 sg13g2_fill_2 FILLER_57_114 ();
 sg13g2_fill_1 FILLER_57_124 ();
 sg13g2_decap_4 FILLER_57_148 ();
 sg13g2_fill_1 FILLER_57_152 ();
 sg13g2_decap_8 FILLER_57_177 ();
 sg13g2_decap_4 FILLER_57_184 ();
 sg13g2_decap_4 FILLER_57_192 ();
 sg13g2_fill_2 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_206 ();
 sg13g2_decap_8 FILLER_57_213 ();
 sg13g2_fill_1 FILLER_57_256 ();
 sg13g2_fill_1 FILLER_57_284 ();
 sg13g2_decap_8 FILLER_57_290 ();
 sg13g2_decap_8 FILLER_57_297 ();
 sg13g2_fill_2 FILLER_57_321 ();
 sg13g2_fill_1 FILLER_57_331 ();
 sg13g2_fill_1 FILLER_57_358 ();
 sg13g2_decap_4 FILLER_57_372 ();
 sg13g2_fill_1 FILLER_57_376 ();
 sg13g2_fill_2 FILLER_57_424 ();
 sg13g2_fill_2 FILLER_57_447 ();
 sg13g2_fill_1 FILLER_57_449 ();
 sg13g2_decap_8 FILLER_57_481 ();
 sg13g2_decap_4 FILLER_57_488 ();
 sg13g2_fill_1 FILLER_57_492 ();
 sg13g2_decap_8 FILLER_57_502 ();
 sg13g2_decap_4 FILLER_57_531 ();
 sg13g2_fill_1 FILLER_57_541 ();
 sg13g2_decap_4 FILLER_57_547 ();
 sg13g2_fill_1 FILLER_57_551 ();
 sg13g2_decap_4 FILLER_57_556 ();
 sg13g2_fill_2 FILLER_57_565 ();
 sg13g2_decap_4 FILLER_57_578 ();
 sg13g2_fill_2 FILLER_57_582 ();
 sg13g2_decap_8 FILLER_57_589 ();
 sg13g2_fill_2 FILLER_57_606 ();
 sg13g2_fill_2 FILLER_57_616 ();
 sg13g2_fill_2 FILLER_57_626 ();
 sg13g2_fill_1 FILLER_57_642 ();
 sg13g2_fill_1 FILLER_57_672 ();
 sg13g2_fill_2 FILLER_57_686 ();
 sg13g2_decap_8 FILLER_57_692 ();
 sg13g2_fill_1 FILLER_57_699 ();
 sg13g2_decap_4 FILLER_57_720 ();
 sg13g2_fill_1 FILLER_57_724 ();
 sg13g2_fill_1 FILLER_57_730 ();
 sg13g2_fill_1 FILLER_57_744 ();
 sg13g2_decap_8 FILLER_57_780 ();
 sg13g2_decap_8 FILLER_57_787 ();
 sg13g2_decap_8 FILLER_57_794 ();
 sg13g2_decap_8 FILLER_57_801 ();
 sg13g2_decap_8 FILLER_57_808 ();
 sg13g2_decap_8 FILLER_57_815 ();
 sg13g2_decap_8 FILLER_57_822 ();
 sg13g2_decap_8 FILLER_57_829 ();
 sg13g2_decap_8 FILLER_57_836 ();
 sg13g2_decap_8 FILLER_57_843 ();
 sg13g2_decap_8 FILLER_57_850 ();
 sg13g2_decap_4 FILLER_57_857 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_fill_1 FILLER_58_65 ();
 sg13g2_decap_8 FILLER_58_71 ();
 sg13g2_decap_8 FILLER_58_78 ();
 sg13g2_fill_1 FILLER_58_85 ();
 sg13g2_fill_2 FILLER_58_99 ();
 sg13g2_fill_1 FILLER_58_101 ();
 sg13g2_decap_8 FILLER_58_114 ();
 sg13g2_decap_8 FILLER_58_121 ();
 sg13g2_fill_2 FILLER_58_128 ();
 sg13g2_fill_2 FILLER_58_154 ();
 sg13g2_fill_1 FILLER_58_156 ();
 sg13g2_fill_2 FILLER_58_161 ();
 sg13g2_fill_2 FILLER_58_246 ();
 sg13g2_fill_1 FILLER_58_281 ();
 sg13g2_fill_2 FILLER_58_291 ();
 sg13g2_fill_1 FILLER_58_293 ();
 sg13g2_fill_2 FILLER_58_315 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_fill_2 FILLER_58_332 ();
 sg13g2_fill_2 FILLER_58_339 ();
 sg13g2_fill_2 FILLER_58_346 ();
 sg13g2_fill_1 FILLER_58_348 ();
 sg13g2_fill_2 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_374 ();
 sg13g2_fill_1 FILLER_58_380 ();
 sg13g2_decap_8 FILLER_58_386 ();
 sg13g2_fill_1 FILLER_58_393 ();
 sg13g2_decap_4 FILLER_58_402 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_decap_4 FILLER_58_418 ();
 sg13g2_fill_2 FILLER_58_422 ();
 sg13g2_decap_4 FILLER_58_453 ();
 sg13g2_fill_2 FILLER_58_457 ();
 sg13g2_fill_2 FILLER_58_505 ();
 sg13g2_fill_1 FILLER_58_507 ();
 sg13g2_fill_1 FILLER_58_534 ();
 sg13g2_fill_1 FILLER_58_602 ();
 sg13g2_fill_1 FILLER_58_608 ();
 sg13g2_fill_2 FILLER_58_617 ();
 sg13g2_fill_1 FILLER_58_685 ();
 sg13g2_fill_1 FILLER_58_694 ();
 sg13g2_decap_4 FILLER_58_705 ();
 sg13g2_fill_2 FILLER_58_714 ();
 sg13g2_fill_1 FILLER_58_716 ();
 sg13g2_decap_8 FILLER_58_721 ();
 sg13g2_decap_4 FILLER_58_728 ();
 sg13g2_fill_2 FILLER_58_754 ();
 sg13g2_fill_2 FILLER_58_769 ();
 sg13g2_fill_1 FILLER_58_771 ();
 sg13g2_decap_8 FILLER_58_781 ();
 sg13g2_decap_8 FILLER_58_788 ();
 sg13g2_decap_8 FILLER_58_795 ();
 sg13g2_decap_8 FILLER_58_802 ();
 sg13g2_decap_8 FILLER_58_809 ();
 sg13g2_decap_8 FILLER_58_816 ();
 sg13g2_decap_8 FILLER_58_823 ();
 sg13g2_decap_8 FILLER_58_830 ();
 sg13g2_decap_8 FILLER_58_837 ();
 sg13g2_decap_8 FILLER_58_844 ();
 sg13g2_decap_8 FILLER_58_851 ();
 sg13g2_decap_4 FILLER_58_858 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_4 ();
 sg13g2_fill_1 FILLER_59_46 ();
 sg13g2_fill_2 FILLER_59_51 ();
 sg13g2_fill_2 FILLER_59_74 ();
 sg13g2_decap_4 FILLER_59_89 ();
 sg13g2_fill_2 FILLER_59_93 ();
 sg13g2_fill_1 FILLER_59_108 ();
 sg13g2_fill_2 FILLER_59_173 ();
 sg13g2_decap_4 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_215 ();
 sg13g2_decap_4 FILLER_59_222 ();
 sg13g2_decap_4 FILLER_59_243 ();
 sg13g2_fill_1 FILLER_59_247 ();
 sg13g2_decap_8 FILLER_59_256 ();
 sg13g2_decap_8 FILLER_59_263 ();
 sg13g2_decap_4 FILLER_59_270 ();
 sg13g2_fill_2 FILLER_59_282 ();
 sg13g2_fill_1 FILLER_59_284 ();
 sg13g2_fill_2 FILLER_59_301 ();
 sg13g2_fill_2 FILLER_59_307 ();
 sg13g2_fill_1 FILLER_59_367 ();
 sg13g2_decap_8 FILLER_59_390 ();
 sg13g2_decap_4 FILLER_59_397 ();
 sg13g2_fill_1 FILLER_59_401 ();
 sg13g2_decap_4 FILLER_59_416 ();
 sg13g2_fill_2 FILLER_59_430 ();
 sg13g2_decap_4 FILLER_59_461 ();
 sg13g2_fill_1 FILLER_59_465 ();
 sg13g2_decap_8 FILLER_59_470 ();
 sg13g2_fill_2 FILLER_59_477 ();
 sg13g2_decap_8 FILLER_59_531 ();
 sg13g2_fill_1 FILLER_59_538 ();
 sg13g2_decap_4 FILLER_59_545 ();
 sg13g2_decap_8 FILLER_59_553 ();
 sg13g2_fill_2 FILLER_59_560 ();
 sg13g2_decap_8 FILLER_59_579 ();
 sg13g2_fill_1 FILLER_59_586 ();
 sg13g2_decap_4 FILLER_59_590 ();
 sg13g2_fill_2 FILLER_59_607 ();
 sg13g2_fill_1 FILLER_59_617 ();
 sg13g2_fill_2 FILLER_59_694 ();
 sg13g2_fill_1 FILLER_59_705 ();
 sg13g2_fill_2 FILLER_59_749 ();
 sg13g2_fill_1 FILLER_59_751 ();
 sg13g2_decap_8 FILLER_59_778 ();
 sg13g2_decap_8 FILLER_59_785 ();
 sg13g2_decap_8 FILLER_59_792 ();
 sg13g2_decap_8 FILLER_59_799 ();
 sg13g2_decap_8 FILLER_59_806 ();
 sg13g2_decap_8 FILLER_59_813 ();
 sg13g2_decap_8 FILLER_59_820 ();
 sg13g2_decap_8 FILLER_59_827 ();
 sg13g2_decap_8 FILLER_59_834 ();
 sg13g2_decap_8 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_855 ();
 sg13g2_fill_2 FILLER_60_48 ();
 sg13g2_fill_1 FILLER_60_50 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_fill_2 FILLER_60_63 ();
 sg13g2_fill_1 FILLER_60_65 ();
 sg13g2_decap_4 FILLER_60_71 ();
 sg13g2_fill_2 FILLER_60_102 ();
 sg13g2_fill_1 FILLER_60_104 ();
 sg13g2_decap_4 FILLER_60_128 ();
 sg13g2_fill_1 FILLER_60_132 ();
 sg13g2_fill_2 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_145 ();
 sg13g2_decap_4 FILLER_60_160 ();
 sg13g2_fill_1 FILLER_60_173 ();
 sg13g2_fill_2 FILLER_60_203 ();
 sg13g2_fill_1 FILLER_60_205 ();
 sg13g2_fill_2 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_234 ();
 sg13g2_fill_2 FILLER_60_269 ();
 sg13g2_fill_1 FILLER_60_271 ();
 sg13g2_fill_2 FILLER_60_302 ();
 sg13g2_fill_2 FILLER_60_339 ();
 sg13g2_fill_1 FILLER_60_341 ();
 sg13g2_fill_1 FILLER_60_365 ();
 sg13g2_decap_4 FILLER_60_381 ();
 sg13g2_fill_2 FILLER_60_393 ();
 sg13g2_fill_1 FILLER_60_395 ();
 sg13g2_fill_2 FILLER_60_399 ();
 sg13g2_decap_4 FILLER_60_420 ();
 sg13g2_fill_1 FILLER_60_424 ();
 sg13g2_fill_1 FILLER_60_449 ();
 sg13g2_fill_2 FILLER_60_473 ();
 sg13g2_fill_2 FILLER_60_500 ();
 sg13g2_fill_1 FILLER_60_502 ();
 sg13g2_decap_4 FILLER_60_512 ();
 sg13g2_fill_2 FILLER_60_516 ();
 sg13g2_decap_4 FILLER_60_528 ();
 sg13g2_fill_2 FILLER_60_532 ();
 sg13g2_fill_1 FILLER_60_564 ();
 sg13g2_fill_2 FILLER_60_626 ();
 sg13g2_fill_2 FILLER_60_654 ();
 sg13g2_fill_2 FILLER_60_670 ();
 sg13g2_fill_1 FILLER_60_680 ();
 sg13g2_fill_2 FILLER_60_689 ();
 sg13g2_fill_1 FILLER_60_691 ();
 sg13g2_fill_1 FILLER_60_710 ();
 sg13g2_fill_1 FILLER_60_724 ();
 sg13g2_fill_1 FILLER_60_733 ();
 sg13g2_fill_1 FILLER_60_742 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_decap_8 FILLER_60_801 ();
 sg13g2_decap_8 FILLER_60_808 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_822 ();
 sg13g2_decap_8 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_836 ();
 sg13g2_decap_8 FILLER_60_843 ();
 sg13g2_decap_8 FILLER_60_850 ();
 sg13g2_decap_4 FILLER_60_857 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_15 ();
 sg13g2_decap_8 FILLER_61_22 ();
 sg13g2_fill_2 FILLER_61_29 ();
 sg13g2_fill_1 FILLER_61_31 ();
 sg13g2_fill_1 FILLER_61_45 ();
 sg13g2_decap_4 FILLER_61_79 ();
 sg13g2_fill_1 FILLER_61_83 ();
 sg13g2_decap_4 FILLER_61_101 ();
 sg13g2_fill_1 FILLER_61_105 ();
 sg13g2_fill_1 FILLER_61_132 ();
 sg13g2_fill_2 FILLER_61_143 ();
 sg13g2_fill_1 FILLER_61_145 ();
 sg13g2_fill_1 FILLER_61_151 ();
 sg13g2_fill_2 FILLER_61_160 ();
 sg13g2_fill_1 FILLER_61_162 ();
 sg13g2_decap_4 FILLER_61_176 ();
 sg13g2_fill_2 FILLER_61_190 ();
 sg13g2_fill_1 FILLER_61_200 ();
 sg13g2_fill_2 FILLER_61_206 ();
 sg13g2_fill_1 FILLER_61_208 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_fill_2 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_226 ();
 sg13g2_decap_4 FILLER_61_247 ();
 sg13g2_fill_1 FILLER_61_251 ();
 sg13g2_decap_4 FILLER_61_274 ();
 sg13g2_fill_2 FILLER_61_278 ();
 sg13g2_fill_2 FILLER_61_366 ();
 sg13g2_fill_2 FILLER_61_390 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_decap_8 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_61_435 ();
 sg13g2_decap_4 FILLER_61_442 ();
 sg13g2_fill_2 FILLER_61_458 ();
 sg13g2_fill_1 FILLER_61_460 ();
 sg13g2_decap_4 FILLER_61_473 ();
 sg13g2_fill_1 FILLER_61_495 ();
 sg13g2_fill_2 FILLER_61_521 ();
 sg13g2_decap_4 FILLER_61_549 ();
 sg13g2_fill_2 FILLER_61_553 ();
 sg13g2_fill_2 FILLER_61_564 ();
 sg13g2_fill_1 FILLER_61_566 ();
 sg13g2_fill_1 FILLER_61_700 ();
 sg13g2_fill_2 FILLER_61_708 ();
 sg13g2_fill_2 FILLER_61_722 ();
 sg13g2_fill_1 FILLER_61_724 ();
 sg13g2_decap_8 FILLER_61_788 ();
 sg13g2_decap_8 FILLER_61_795 ();
 sg13g2_decap_8 FILLER_61_802 ();
 sg13g2_decap_8 FILLER_61_809 ();
 sg13g2_decap_8 FILLER_61_816 ();
 sg13g2_decap_8 FILLER_61_823 ();
 sg13g2_decap_8 FILLER_61_830 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_8 FILLER_61_851 ();
 sg13g2_decap_4 FILLER_61_858 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_fill_2 FILLER_62_21 ();
 sg13g2_fill_1 FILLER_62_36 ();
 sg13g2_fill_2 FILLER_62_50 ();
 sg13g2_fill_1 FILLER_62_52 ();
 sg13g2_fill_1 FILLER_62_68 ();
 sg13g2_decap_4 FILLER_62_78 ();
 sg13g2_decap_4 FILLER_62_93 ();
 sg13g2_fill_2 FILLER_62_123 ();
 sg13g2_fill_2 FILLER_62_140 ();
 sg13g2_fill_2 FILLER_62_158 ();
 sg13g2_fill_1 FILLER_62_160 ();
 sg13g2_fill_2 FILLER_62_170 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_decap_4 FILLER_62_181 ();
 sg13g2_fill_2 FILLER_62_195 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_decap_4 FILLER_62_214 ();
 sg13g2_decap_8 FILLER_62_232 ();
 sg13g2_decap_4 FILLER_62_239 ();
 sg13g2_fill_2 FILLER_62_243 ();
 sg13g2_decap_4 FILLER_62_253 ();
 sg13g2_fill_2 FILLER_62_257 ();
 sg13g2_fill_2 FILLER_62_264 ();
 sg13g2_fill_1 FILLER_62_266 ();
 sg13g2_fill_2 FILLER_62_284 ();
 sg13g2_fill_1 FILLER_62_286 ();
 sg13g2_fill_1 FILLER_62_299 ();
 sg13g2_fill_2 FILLER_62_335 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_fill_1 FILLER_62_361 ();
 sg13g2_decap_8 FILLER_62_383 ();
 sg13g2_decap_8 FILLER_62_439 ();
 sg13g2_decap_4 FILLER_62_446 ();
 sg13g2_fill_2 FILLER_62_503 ();
 sg13g2_decap_4 FILLER_62_517 ();
 sg13g2_fill_2 FILLER_62_521 ();
 sg13g2_fill_1 FILLER_62_536 ();
 sg13g2_decap_8 FILLER_62_541 ();
 sg13g2_fill_2 FILLER_62_548 ();
 sg13g2_fill_1 FILLER_62_581 ();
 sg13g2_fill_1 FILLER_62_617 ();
 sg13g2_decap_4 FILLER_62_643 ();
 sg13g2_fill_1 FILLER_62_647 ();
 sg13g2_fill_1 FILLER_62_673 ();
 sg13g2_fill_1 FILLER_62_688 ();
 sg13g2_fill_2 FILLER_62_740 ();
 sg13g2_fill_1 FILLER_62_742 ();
 sg13g2_decap_8 FILLER_62_782 ();
 sg13g2_decap_8 FILLER_62_789 ();
 sg13g2_decap_8 FILLER_62_796 ();
 sg13g2_decap_8 FILLER_62_803 ();
 sg13g2_decap_8 FILLER_62_810 ();
 sg13g2_decap_8 FILLER_62_817 ();
 sg13g2_decap_8 FILLER_62_824 ();
 sg13g2_decap_8 FILLER_62_831 ();
 sg13g2_decap_8 FILLER_62_838 ();
 sg13g2_decap_8 FILLER_62_845 ();
 sg13g2_decap_8 FILLER_62_852 ();
 sg13g2_fill_2 FILLER_62_859 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_71 ();
 sg13g2_fill_2 FILLER_63_75 ();
 sg13g2_fill_1 FILLER_63_77 ();
 sg13g2_fill_2 FILLER_63_94 ();
 sg13g2_fill_2 FILLER_63_100 ();
 sg13g2_fill_1 FILLER_63_102 ();
 sg13g2_fill_2 FILLER_63_111 ();
 sg13g2_fill_1 FILLER_63_148 ();
 sg13g2_decap_4 FILLER_63_172 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_fill_1 FILLER_63_187 ();
 sg13g2_fill_2 FILLER_63_193 ();
 sg13g2_fill_1 FILLER_63_195 ();
 sg13g2_decap_4 FILLER_63_228 ();
 sg13g2_fill_1 FILLER_63_232 ();
 sg13g2_fill_2 FILLER_63_258 ();
 sg13g2_fill_1 FILLER_63_260 ();
 sg13g2_fill_2 FILLER_63_274 ();
 sg13g2_fill_1 FILLER_63_276 ();
 sg13g2_fill_2 FILLER_63_292 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_decap_4 FILLER_63_314 ();
 sg13g2_fill_2 FILLER_63_363 ();
 sg13g2_decap_8 FILLER_63_435 ();
 sg13g2_fill_2 FILLER_63_488 ();
 sg13g2_decap_4 FILLER_63_513 ();
 sg13g2_fill_1 FILLER_63_525 ();
 sg13g2_fill_1 FILLER_63_552 ();
 sg13g2_fill_2 FILLER_63_558 ();
 sg13g2_fill_2 FILLER_63_573 ();
 sg13g2_fill_1 FILLER_63_575 ();
 sg13g2_fill_2 FILLER_63_586 ();
 sg13g2_fill_1 FILLER_63_588 ();
 sg13g2_fill_1 FILLER_63_602 ();
 sg13g2_fill_1 FILLER_63_663 ();
 sg13g2_decap_8 FILLER_63_690 ();
 sg13g2_fill_1 FILLER_63_697 ();
 sg13g2_fill_2 FILLER_63_702 ();
 sg13g2_fill_1 FILLER_63_704 ();
 sg13g2_fill_2 FILLER_63_724 ();
 sg13g2_fill_1 FILLER_63_726 ();
 sg13g2_fill_2 FILLER_63_761 ();
 sg13g2_fill_1 FILLER_63_763 ();
 sg13g2_decap_8 FILLER_63_773 ();
 sg13g2_decap_8 FILLER_63_780 ();
 sg13g2_decap_8 FILLER_63_787 ();
 sg13g2_decap_8 FILLER_63_794 ();
 sg13g2_decap_8 FILLER_63_801 ();
 sg13g2_decap_8 FILLER_63_808 ();
 sg13g2_decap_8 FILLER_63_815 ();
 sg13g2_decap_8 FILLER_63_822 ();
 sg13g2_decap_8 FILLER_63_829 ();
 sg13g2_decap_8 FILLER_63_836 ();
 sg13g2_decap_8 FILLER_63_843 ();
 sg13g2_decap_8 FILLER_63_850 ();
 sg13g2_decap_4 FILLER_63_857 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_18 ();
 sg13g2_fill_2 FILLER_64_44 ();
 sg13g2_fill_1 FILLER_64_46 ();
 sg13g2_fill_1 FILLER_64_57 ();
 sg13g2_fill_2 FILLER_64_89 ();
 sg13g2_fill_1 FILLER_64_100 ();
 sg13g2_fill_1 FILLER_64_113 ();
 sg13g2_decap_8 FILLER_64_118 ();
 sg13g2_fill_2 FILLER_64_131 ();
 sg13g2_decap_4 FILLER_64_141 ();
 sg13g2_fill_2 FILLER_64_145 ();
 sg13g2_fill_1 FILLER_64_156 ();
 sg13g2_fill_1 FILLER_64_165 ();
 sg13g2_decap_4 FILLER_64_205 ();
 sg13g2_fill_1 FILLER_64_209 ();
 sg13g2_fill_2 FILLER_64_234 ();
 sg13g2_decap_4 FILLER_64_252 ();
 sg13g2_fill_1 FILLER_64_256 ();
 sg13g2_fill_2 FILLER_64_269 ();
 sg13g2_decap_4 FILLER_64_285 ();
 sg13g2_decap_4 FILLER_64_297 ();
 sg13g2_fill_2 FILLER_64_306 ();
 sg13g2_fill_1 FILLER_64_308 ();
 sg13g2_decap_4 FILLER_64_317 ();
 sg13g2_fill_2 FILLER_64_321 ();
 sg13g2_fill_2 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_371 ();
 sg13g2_fill_1 FILLER_64_378 ();
 sg13g2_fill_2 FILLER_64_383 ();
 sg13g2_fill_2 FILLER_64_430 ();
 sg13g2_fill_1 FILLER_64_432 ();
 sg13g2_fill_2 FILLER_64_444 ();
 sg13g2_fill_2 FILLER_64_477 ();
 sg13g2_fill_2 FILLER_64_496 ();
 sg13g2_decap_8 FILLER_64_502 ();
 sg13g2_decap_4 FILLER_64_509 ();
 sg13g2_fill_1 FILLER_64_539 ();
 sg13g2_fill_2 FILLER_64_543 ();
 sg13g2_fill_1 FILLER_64_545 ();
 sg13g2_fill_1 FILLER_64_655 ();
 sg13g2_decap_4 FILLER_64_691 ();
 sg13g2_decap_8 FILLER_64_721 ();
 sg13g2_decap_8 FILLER_64_728 ();
 sg13g2_fill_2 FILLER_64_735 ();
 sg13g2_decap_8 FILLER_64_754 ();
 sg13g2_decap_8 FILLER_64_761 ();
 sg13g2_decap_8 FILLER_64_768 ();
 sg13g2_decap_8 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_782 ();
 sg13g2_decap_8 FILLER_64_789 ();
 sg13g2_decap_8 FILLER_64_796 ();
 sg13g2_decap_8 FILLER_64_803 ();
 sg13g2_decap_8 FILLER_64_810 ();
 sg13g2_decap_8 FILLER_64_817 ();
 sg13g2_decap_8 FILLER_64_824 ();
 sg13g2_decap_8 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_fill_1 FILLER_65_26 ();
 sg13g2_fill_1 FILLER_65_57 ();
 sg13g2_decap_8 FILLER_65_74 ();
 sg13g2_fill_2 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_83 ();
 sg13g2_decap_8 FILLER_65_94 ();
 sg13g2_fill_2 FILLER_65_101 ();
 sg13g2_decap_8 FILLER_65_121 ();
 sg13g2_decap_8 FILLER_65_128 ();
 sg13g2_decap_8 FILLER_65_148 ();
 sg13g2_decap_4 FILLER_65_155 ();
 sg13g2_decap_8 FILLER_65_167 ();
 sg13g2_decap_4 FILLER_65_179 ();
 sg13g2_fill_2 FILLER_65_183 ();
 sg13g2_fill_1 FILLER_65_218 ();
 sg13g2_fill_2 FILLER_65_228 ();
 sg13g2_fill_1 FILLER_65_230 ();
 sg13g2_fill_2 FILLER_65_257 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_fill_1 FILLER_65_285 ();
 sg13g2_decap_8 FILLER_65_291 ();
 sg13g2_fill_1 FILLER_65_304 ();
 sg13g2_fill_1 FILLER_65_320 ();
 sg13g2_fill_1 FILLER_65_330 ();
 sg13g2_fill_1 FILLER_65_343 ();
 sg13g2_fill_1 FILLER_65_353 ();
 sg13g2_decap_4 FILLER_65_388 ();
 sg13g2_fill_2 FILLER_65_451 ();
 sg13g2_fill_2 FILLER_65_490 ();
 sg13g2_fill_1 FILLER_65_492 ();
 sg13g2_fill_2 FILLER_65_510 ();
 sg13g2_fill_2 FILLER_65_579 ();
 sg13g2_decap_4 FILLER_65_586 ();
 sg13g2_fill_1 FILLER_65_590 ();
 sg13g2_fill_1 FILLER_65_605 ();
 sg13g2_fill_1 FILLER_65_622 ();
 sg13g2_fill_1 FILLER_65_651 ();
 sg13g2_fill_1 FILLER_65_660 ();
 sg13g2_decap_4 FILLER_65_701 ();
 sg13g2_fill_1 FILLER_65_705 ();
 sg13g2_decap_8 FILLER_65_710 ();
 sg13g2_decap_8 FILLER_65_717 ();
 sg13g2_decap_8 FILLER_65_724 ();
 sg13g2_decap_8 FILLER_65_731 ();
 sg13g2_decap_8 FILLER_65_738 ();
 sg13g2_decap_8 FILLER_65_745 ();
 sg13g2_decap_8 FILLER_65_752 ();
 sg13g2_decap_8 FILLER_65_759 ();
 sg13g2_decap_8 FILLER_65_766 ();
 sg13g2_decap_8 FILLER_65_773 ();
 sg13g2_decap_8 FILLER_65_780 ();
 sg13g2_decap_8 FILLER_65_787 ();
 sg13g2_decap_8 FILLER_65_794 ();
 sg13g2_decap_8 FILLER_65_801 ();
 sg13g2_decap_8 FILLER_65_808 ();
 sg13g2_decap_8 FILLER_65_815 ();
 sg13g2_decap_8 FILLER_65_822 ();
 sg13g2_decap_8 FILLER_65_829 ();
 sg13g2_decap_8 FILLER_65_836 ();
 sg13g2_decap_8 FILLER_65_843 ();
 sg13g2_decap_8 FILLER_65_850 ();
 sg13g2_decap_4 FILLER_65_857 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_4 ();
 sg13g2_decap_8 FILLER_66_24 ();
 sg13g2_fill_2 FILLER_66_31 ();
 sg13g2_fill_2 FILLER_66_74 ();
 sg13g2_fill_1 FILLER_66_103 ();
 sg13g2_fill_1 FILLER_66_109 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_fill_2 FILLER_66_126 ();
 sg13g2_fill_1 FILLER_66_157 ();
 sg13g2_fill_2 FILLER_66_166 ();
 sg13g2_decap_4 FILLER_66_194 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_decap_8 FILLER_66_204 ();
 sg13g2_decap_4 FILLER_66_211 ();
 sg13g2_decap_8 FILLER_66_228 ();
 sg13g2_decap_8 FILLER_66_235 ();
 sg13g2_decap_4 FILLER_66_242 ();
 sg13g2_fill_2 FILLER_66_246 ();
 sg13g2_decap_8 FILLER_66_251 ();
 sg13g2_decap_8 FILLER_66_258 ();
 sg13g2_fill_2 FILLER_66_265 ();
 sg13g2_decap_8 FILLER_66_276 ();
 sg13g2_decap_4 FILLER_66_283 ();
 sg13g2_decap_8 FILLER_66_296 ();
 sg13g2_decap_4 FILLER_66_303 ();
 sg13g2_fill_1 FILLER_66_307 ();
 sg13g2_decap_8 FILLER_66_317 ();
 sg13g2_fill_1 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_333 ();
 sg13g2_fill_2 FILLER_66_347 ();
 sg13g2_fill_1 FILLER_66_365 ();
 sg13g2_fill_1 FILLER_66_371 ();
 sg13g2_decap_4 FILLER_66_415 ();
 sg13g2_fill_2 FILLER_66_419 ();
 sg13g2_fill_1 FILLER_66_437 ();
 sg13g2_fill_2 FILLER_66_469 ();
 sg13g2_decap_4 FILLER_66_489 ();
 sg13g2_fill_1 FILLER_66_493 ();
 sg13g2_fill_1 FILLER_66_517 ();
 sg13g2_decap_8 FILLER_66_523 ();
 sg13g2_decap_8 FILLER_66_530 ();
 sg13g2_fill_2 FILLER_66_537 ();
 sg13g2_decap_4 FILLER_66_569 ();
 sg13g2_decap_8 FILLER_66_588 ();
 sg13g2_decap_8 FILLER_66_595 ();
 sg13g2_decap_8 FILLER_66_621 ();
 sg13g2_decap_8 FILLER_66_628 ();
 sg13g2_decap_4 FILLER_66_635 ();
 sg13g2_fill_1 FILLER_66_639 ();
 sg13g2_decap_8 FILLER_66_702 ();
 sg13g2_decap_8 FILLER_66_709 ();
 sg13g2_decap_8 FILLER_66_716 ();
 sg13g2_decap_8 FILLER_66_723 ();
 sg13g2_decap_8 FILLER_66_730 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_744 ();
 sg13g2_decap_8 FILLER_66_751 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_67_31 ();
 sg13g2_decap_4 FILLER_67_52 ();
 sg13g2_fill_1 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_81 ();
 sg13g2_fill_2 FILLER_67_101 ();
 sg13g2_fill_1 FILLER_67_134 ();
 sg13g2_decap_4 FILLER_67_154 ();
 sg13g2_fill_1 FILLER_67_158 ();
 sg13g2_decap_8 FILLER_67_163 ();
 sg13g2_fill_1 FILLER_67_170 ();
 sg13g2_fill_2 FILLER_67_191 ();
 sg13g2_fill_1 FILLER_67_209 ();
 sg13g2_fill_1 FILLER_67_213 ();
 sg13g2_decap_8 FILLER_67_223 ();
 sg13g2_fill_1 FILLER_67_230 ();
 sg13g2_decap_8 FILLER_67_250 ();
 sg13g2_fill_2 FILLER_67_265 ();
 sg13g2_fill_1 FILLER_67_267 ();
 sg13g2_fill_1 FILLER_67_303 ();
 sg13g2_decap_8 FILLER_67_309 ();
 sg13g2_fill_2 FILLER_67_316 ();
 sg13g2_fill_1 FILLER_67_318 ();
 sg13g2_fill_2 FILLER_67_323 ();
 sg13g2_fill_1 FILLER_67_325 ();
 sg13g2_fill_1 FILLER_67_338 ();
 sg13g2_fill_2 FILLER_67_344 ();
 sg13g2_fill_2 FILLER_67_355 ();
 sg13g2_fill_1 FILLER_67_357 ();
 sg13g2_decap_8 FILLER_67_363 ();
 sg13g2_decap_4 FILLER_67_370 ();
 sg13g2_fill_1 FILLER_67_374 ();
 sg13g2_fill_1 FILLER_67_379 ();
 sg13g2_decap_4 FILLER_67_391 ();
 sg13g2_fill_1 FILLER_67_395 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_67_406 ();
 sg13g2_decap_4 FILLER_67_413 ();
 sg13g2_fill_1 FILLER_67_417 ();
 sg13g2_decap_8 FILLER_67_433 ();
 sg13g2_fill_2 FILLER_67_440 ();
 sg13g2_decap_4 FILLER_67_476 ();
 sg13g2_decap_8 FILLER_67_506 ();
 sg13g2_decap_4 FILLER_67_513 ();
 sg13g2_decap_4 FILLER_67_532 ();
 sg13g2_fill_2 FILLER_67_567 ();
 sg13g2_fill_1 FILLER_67_621 ();
 sg13g2_decap_8 FILLER_67_686 ();
 sg13g2_decap_8 FILLER_67_693 ();
 sg13g2_decap_8 FILLER_67_700 ();
 sg13g2_decap_8 FILLER_67_707 ();
 sg13g2_decap_8 FILLER_67_714 ();
 sg13g2_decap_8 FILLER_67_721 ();
 sg13g2_decap_8 FILLER_67_728 ();
 sg13g2_decap_8 FILLER_67_735 ();
 sg13g2_decap_8 FILLER_67_742 ();
 sg13g2_decap_8 FILLER_67_749 ();
 sg13g2_decap_8 FILLER_67_756 ();
 sg13g2_decap_8 FILLER_67_763 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_decap_8 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_784 ();
 sg13g2_decap_8 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_798 ();
 sg13g2_decap_8 FILLER_67_805 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_854 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_16 ();
 sg13g2_fill_1 FILLER_68_21 ();
 sg13g2_fill_1 FILLER_68_31 ();
 sg13g2_decap_4 FILLER_68_55 ();
 sg13g2_fill_1 FILLER_68_59 ();
 sg13g2_fill_2 FILLER_68_82 ();
 sg13g2_fill_1 FILLER_68_84 ();
 sg13g2_decap_4 FILLER_68_107 ();
 sg13g2_fill_2 FILLER_68_111 ();
 sg13g2_fill_2 FILLER_68_118 ();
 sg13g2_fill_1 FILLER_68_120 ();
 sg13g2_fill_2 FILLER_68_126 ();
 sg13g2_fill_1 FILLER_68_128 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_4 FILLER_68_140 ();
 sg13g2_fill_1 FILLER_68_144 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_4 FILLER_68_168 ();
 sg13g2_fill_2 FILLER_68_172 ();
 sg13g2_fill_1 FILLER_68_184 ();
 sg13g2_decap_8 FILLER_68_190 ();
 sg13g2_fill_2 FILLER_68_197 ();
 sg13g2_fill_1 FILLER_68_199 ();
 sg13g2_fill_1 FILLER_68_205 ();
 sg13g2_fill_2 FILLER_68_226 ();
 sg13g2_fill_1 FILLER_68_228 ();
 sg13g2_fill_1 FILLER_68_258 ();
 sg13g2_decap_4 FILLER_68_269 ();
 sg13g2_fill_2 FILLER_68_293 ();
 sg13g2_decap_8 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_332 ();
 sg13g2_fill_2 FILLER_68_340 ();
 sg13g2_fill_1 FILLER_68_356 ();
 sg13g2_decap_4 FILLER_68_392 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_fill_1 FILLER_68_439 ();
 sg13g2_decap_8 FILLER_68_461 ();
 sg13g2_fill_2 FILLER_68_468 ();
 sg13g2_decap_8 FILLER_68_487 ();
 sg13g2_decap_8 FILLER_68_502 ();
 sg13g2_decap_4 FILLER_68_509 ();
 sg13g2_fill_2 FILLER_68_513 ();
 sg13g2_fill_2 FILLER_68_541 ();
 sg13g2_fill_1 FILLER_68_543 ();
 sg13g2_fill_2 FILLER_68_596 ();
 sg13g2_decap_8 FILLER_68_623 ();
 sg13g2_fill_1 FILLER_68_643 ();
 sg13g2_decap_4 FILLER_68_657 ();
 sg13g2_fill_1 FILLER_68_661 ();
 sg13g2_fill_1 FILLER_68_676 ();
 sg13g2_decap_8 FILLER_68_693 ();
 sg13g2_decap_8 FILLER_68_700 ();
 sg13g2_decap_8 FILLER_68_707 ();
 sg13g2_decap_8 FILLER_68_714 ();
 sg13g2_decap_8 FILLER_68_721 ();
 sg13g2_decap_8 FILLER_68_728 ();
 sg13g2_decap_8 FILLER_68_735 ();
 sg13g2_decap_8 FILLER_68_742 ();
 sg13g2_decap_8 FILLER_68_749 ();
 sg13g2_decap_8 FILLER_68_756 ();
 sg13g2_decap_8 FILLER_68_763 ();
 sg13g2_decap_8 FILLER_68_770 ();
 sg13g2_decap_8 FILLER_68_777 ();
 sg13g2_decap_8 FILLER_68_784 ();
 sg13g2_decap_8 FILLER_68_791 ();
 sg13g2_decap_8 FILLER_68_798 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_decap_8 FILLER_68_812 ();
 sg13g2_decap_8 FILLER_68_819 ();
 sg13g2_decap_8 FILLER_68_826 ();
 sg13g2_decap_8 FILLER_68_833 ();
 sg13g2_decap_8 FILLER_68_840 ();
 sg13g2_decap_8 FILLER_68_847 ();
 sg13g2_decap_8 FILLER_68_854 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_97 ();
 sg13g2_decap_4 FILLER_69_104 ();
 sg13g2_fill_2 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_125 ();
 sg13g2_fill_2 FILLER_69_134 ();
 sg13g2_fill_1 FILLER_69_136 ();
 sg13g2_fill_2 FILLER_69_142 ();
 sg13g2_decap_4 FILLER_69_159 ();
 sg13g2_decap_8 FILLER_69_169 ();
 sg13g2_fill_2 FILLER_69_176 ();
 sg13g2_fill_2 FILLER_69_211 ();
 sg13g2_decap_4 FILLER_69_228 ();
 sg13g2_fill_1 FILLER_69_232 ();
 sg13g2_fill_1 FILLER_69_243 ();
 sg13g2_fill_2 FILLER_69_254 ();
 sg13g2_fill_1 FILLER_69_256 ();
 sg13g2_decap_4 FILLER_69_289 ();
 sg13g2_fill_1 FILLER_69_293 ();
 sg13g2_decap_8 FILLER_69_313 ();
 sg13g2_decap_8 FILLER_69_320 ();
 sg13g2_fill_2 FILLER_69_327 ();
 sg13g2_fill_1 FILLER_69_329 ();
 sg13g2_decap_4 FILLER_69_355 ();
 sg13g2_fill_2 FILLER_69_359 ();
 sg13g2_decap_4 FILLER_69_374 ();
 sg13g2_fill_1 FILLER_69_378 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_fill_2 FILLER_69_422 ();
 sg13g2_fill_2 FILLER_69_429 ();
 sg13g2_fill_1 FILLER_69_443 ();
 sg13g2_fill_2 FILLER_69_459 ();
 sg13g2_decap_4 FILLER_69_474 ();
 sg13g2_fill_1 FILLER_69_478 ();
 sg13g2_decap_4 FILLER_69_487 ();
 sg13g2_fill_1 FILLER_69_491 ();
 sg13g2_fill_2 FILLER_69_553 ();
 sg13g2_fill_1 FILLER_69_568 ();
 sg13g2_fill_2 FILLER_69_598 ();
 sg13g2_fill_1 FILLER_69_600 ();
 sg13g2_fill_1 FILLER_69_640 ();
 sg13g2_fill_2 FILLER_69_654 ();
 sg13g2_fill_1 FILLER_69_656 ();
 sg13g2_decap_8 FILLER_69_709 ();
 sg13g2_decap_8 FILLER_69_716 ();
 sg13g2_decap_8 FILLER_69_723 ();
 sg13g2_decap_8 FILLER_69_730 ();
 sg13g2_decap_8 FILLER_69_737 ();
 sg13g2_decap_8 FILLER_69_744 ();
 sg13g2_decap_8 FILLER_69_751 ();
 sg13g2_decap_8 FILLER_69_758 ();
 sg13g2_decap_8 FILLER_69_765 ();
 sg13g2_decap_8 FILLER_69_772 ();
 sg13g2_decap_8 FILLER_69_779 ();
 sg13g2_decap_8 FILLER_69_786 ();
 sg13g2_decap_8 FILLER_69_793 ();
 sg13g2_decap_8 FILLER_69_800 ();
 sg13g2_decap_8 FILLER_69_807 ();
 sg13g2_decap_8 FILLER_69_814 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_decap_8 FILLER_69_835 ();
 sg13g2_decap_8 FILLER_69_842 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_4 FILLER_69_856 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_32 ();
 sg13g2_fill_2 FILLER_70_45 ();
 sg13g2_decap_4 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_137 ();
 sg13g2_decap_4 FILLER_70_148 ();
 sg13g2_fill_1 FILLER_70_174 ();
 sg13g2_fill_2 FILLER_70_197 ();
 sg13g2_fill_1 FILLER_70_212 ();
 sg13g2_decap_4 FILLER_70_223 ();
 sg13g2_fill_1 FILLER_70_227 ();
 sg13g2_decap_4 FILLER_70_236 ();
 sg13g2_decap_8 FILLER_70_257 ();
 sg13g2_decap_4 FILLER_70_264 ();
 sg13g2_fill_1 FILLER_70_268 ();
 sg13g2_fill_1 FILLER_70_281 ();
 sg13g2_fill_1 FILLER_70_286 ();
 sg13g2_decap_8 FILLER_70_291 ();
 sg13g2_decap_4 FILLER_70_298 ();
 sg13g2_fill_1 FILLER_70_302 ();
 sg13g2_fill_1 FILLER_70_311 ();
 sg13g2_decap_8 FILLER_70_320 ();
 sg13g2_fill_2 FILLER_70_327 ();
 sg13g2_decap_8 FILLER_70_365 ();
 sg13g2_decap_4 FILLER_70_372 ();
 sg13g2_fill_1 FILLER_70_391 ();
 sg13g2_fill_2 FILLER_70_395 ();
 sg13g2_decap_8 FILLER_70_424 ();
 sg13g2_decap_8 FILLER_70_431 ();
 sg13g2_decap_8 FILLER_70_438 ();
 sg13g2_fill_1 FILLER_70_445 ();
 sg13g2_decap_8 FILLER_70_450 ();
 sg13g2_fill_2 FILLER_70_457 ();
 sg13g2_decap_8 FILLER_70_480 ();
 sg13g2_decap_8 FILLER_70_487 ();
 sg13g2_decap_8 FILLER_70_494 ();
 sg13g2_fill_2 FILLER_70_501 ();
 sg13g2_fill_2 FILLER_70_507 ();
 sg13g2_decap_8 FILLER_70_542 ();
 sg13g2_decap_8 FILLER_70_585 ();
 sg13g2_decap_4 FILLER_70_592 ();
 sg13g2_fill_2 FILLER_70_596 ();
 sg13g2_decap_8 FILLER_70_630 ();
 sg13g2_decap_8 FILLER_70_637 ();
 sg13g2_fill_2 FILLER_70_644 ();
 sg13g2_fill_1 FILLER_70_656 ();
 sg13g2_decap_8 FILLER_70_708 ();
 sg13g2_decap_8 FILLER_70_715 ();
 sg13g2_decap_8 FILLER_70_722 ();
 sg13g2_decap_8 FILLER_70_729 ();
 sg13g2_decap_8 FILLER_70_736 ();
 sg13g2_decap_8 FILLER_70_743 ();
 sg13g2_decap_8 FILLER_70_750 ();
 sg13g2_decap_8 FILLER_70_757 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_decap_8 FILLER_70_771 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_decap_8 FILLER_70_785 ();
 sg13g2_decap_8 FILLER_70_792 ();
 sg13g2_decap_8 FILLER_70_799 ();
 sg13g2_decap_8 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_813 ();
 sg13g2_decap_8 FILLER_70_820 ();
 sg13g2_decap_8 FILLER_70_827 ();
 sg13g2_decap_8 FILLER_70_834 ();
 sg13g2_decap_8 FILLER_70_841 ();
 sg13g2_decap_8 FILLER_70_848 ();
 sg13g2_decap_8 FILLER_70_855 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_fill_1 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_34 ();
 sg13g2_decap_8 FILLER_71_41 ();
 sg13g2_decap_8 FILLER_71_48 ();
 sg13g2_decap_8 FILLER_71_55 ();
 sg13g2_decap_8 FILLER_71_62 ();
 sg13g2_decap_8 FILLER_71_69 ();
 sg13g2_fill_2 FILLER_71_76 ();
 sg13g2_decap_8 FILLER_71_81 ();
 sg13g2_decap_4 FILLER_71_88 ();
 sg13g2_decap_8 FILLER_71_101 ();
 sg13g2_fill_2 FILLER_71_108 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_4 FILLER_71_137 ();
 sg13g2_fill_2 FILLER_71_146 ();
 sg13g2_fill_2 FILLER_71_152 ();
 sg13g2_decap_8 FILLER_71_159 ();
 sg13g2_decap_8 FILLER_71_166 ();
 sg13g2_fill_1 FILLER_71_173 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_4 FILLER_71_211 ();
 sg13g2_fill_2 FILLER_71_231 ();
 sg13g2_fill_1 FILLER_71_233 ();
 sg13g2_fill_2 FILLER_71_252 ();
 sg13g2_fill_1 FILLER_71_254 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_fill_2 FILLER_71_266 ();
 sg13g2_fill_1 FILLER_71_280 ();
 sg13g2_decap_4 FILLER_71_296 ();
 sg13g2_decap_4 FILLER_71_313 ();
 sg13g2_fill_1 FILLER_71_317 ();
 sg13g2_fill_1 FILLER_71_324 ();
 sg13g2_fill_2 FILLER_71_339 ();
 sg13g2_fill_1 FILLER_71_350 ();
 sg13g2_decap_4 FILLER_71_355 ();
 sg13g2_fill_1 FILLER_71_372 ();
 sg13g2_fill_2 FILLER_71_391 ();
 sg13g2_fill_1 FILLER_71_393 ();
 sg13g2_decap_4 FILLER_71_400 ();
 sg13g2_fill_1 FILLER_71_404 ();
 sg13g2_fill_1 FILLER_71_420 ();
 sg13g2_fill_2 FILLER_71_430 ();
 sg13g2_fill_1 FILLER_71_432 ();
 sg13g2_fill_2 FILLER_71_460 ();
 sg13g2_fill_1 FILLER_71_462 ();
 sg13g2_decap_8 FILLER_71_467 ();
 sg13g2_fill_1 FILLER_71_539 ();
 sg13g2_fill_1 FILLER_71_568 ();
 sg13g2_fill_2 FILLER_71_640 ();
 sg13g2_fill_2 FILLER_71_668 ();
 sg13g2_fill_2 FILLER_71_684 ();
 sg13g2_decap_8 FILLER_71_709 ();
 sg13g2_decap_8 FILLER_71_716 ();
 sg13g2_decap_8 FILLER_71_723 ();
 sg13g2_decap_8 FILLER_71_730 ();
 sg13g2_decap_8 FILLER_71_737 ();
 sg13g2_decap_8 FILLER_71_744 ();
 sg13g2_decap_8 FILLER_71_751 ();
 sg13g2_decap_8 FILLER_71_758 ();
 sg13g2_decap_8 FILLER_71_765 ();
 sg13g2_decap_8 FILLER_71_772 ();
 sg13g2_decap_8 FILLER_71_779 ();
 sg13g2_decap_8 FILLER_71_786 ();
 sg13g2_decap_8 FILLER_71_793 ();
 sg13g2_decap_8 FILLER_71_800 ();
 sg13g2_decap_8 FILLER_71_807 ();
 sg13g2_decap_8 FILLER_71_814 ();
 sg13g2_decap_8 FILLER_71_821 ();
 sg13g2_decap_8 FILLER_71_828 ();
 sg13g2_decap_8 FILLER_71_835 ();
 sg13g2_decap_8 FILLER_71_842 ();
 sg13g2_decap_8 FILLER_71_849 ();
 sg13g2_decap_4 FILLER_71_856 ();
 sg13g2_fill_2 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_4 FILLER_72_105 ();
 sg13g2_fill_2 FILLER_72_109 ();
 sg13g2_fill_2 FILLER_72_137 ();
 sg13g2_fill_2 FILLER_72_155 ();
 sg13g2_fill_1 FILLER_72_157 ();
 sg13g2_decap_4 FILLER_72_169 ();
 sg13g2_fill_2 FILLER_72_173 ();
 sg13g2_decap_8 FILLER_72_180 ();
 sg13g2_decap_4 FILLER_72_187 ();
 sg13g2_fill_2 FILLER_72_191 ();
 sg13g2_decap_4 FILLER_72_205 ();
 sg13g2_fill_1 FILLER_72_209 ();
 sg13g2_decap_8 FILLER_72_222 ();
 sg13g2_decap_8 FILLER_72_229 ();
 sg13g2_fill_2 FILLER_72_268 ();
 sg13g2_fill_1 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_289 ();
 sg13g2_fill_2 FILLER_72_296 ();
 sg13g2_decap_4 FILLER_72_310 ();
 sg13g2_fill_2 FILLER_72_318 ();
 sg13g2_decap_4 FILLER_72_328 ();
 sg13g2_decap_4 FILLER_72_337 ();
 sg13g2_decap_8 FILLER_72_351 ();
 sg13g2_fill_1 FILLER_72_358 ();
 sg13g2_decap_4 FILLER_72_363 ();
 sg13g2_decap_8 FILLER_72_372 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_fill_1 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_415 ();
 sg13g2_decap_4 FILLER_72_442 ();
 sg13g2_fill_2 FILLER_72_446 ();
 sg13g2_fill_1 FILLER_72_468 ();
 sg13g2_decap_8 FILLER_72_485 ();
 sg13g2_fill_1 FILLER_72_492 ();
 sg13g2_fill_1 FILLER_72_497 ();
 sg13g2_fill_2 FILLER_72_511 ();
 sg13g2_fill_1 FILLER_72_550 ();
 sg13g2_fill_1 FILLER_72_564 ();
 sg13g2_fill_2 FILLER_72_581 ();
 sg13g2_fill_1 FILLER_72_583 ();
 sg13g2_decap_8 FILLER_72_589 ();
 sg13g2_fill_1 FILLER_72_608 ();
 sg13g2_fill_2 FILLER_72_622 ();
 sg13g2_fill_2 FILLER_72_641 ();
 sg13g2_fill_1 FILLER_72_643 ();
 sg13g2_decap_4 FILLER_72_654 ();
 sg13g2_fill_2 FILLER_72_671 ();
 sg13g2_fill_1 FILLER_72_673 ();
 sg13g2_decap_8 FILLER_72_700 ();
 sg13g2_decap_8 FILLER_72_707 ();
 sg13g2_decap_8 FILLER_72_714 ();
 sg13g2_decap_8 FILLER_72_721 ();
 sg13g2_decap_8 FILLER_72_728 ();
 sg13g2_decap_8 FILLER_72_735 ();
 sg13g2_decap_8 FILLER_72_742 ();
 sg13g2_decap_8 FILLER_72_749 ();
 sg13g2_decap_8 FILLER_72_756 ();
 sg13g2_decap_8 FILLER_72_763 ();
 sg13g2_decap_8 FILLER_72_770 ();
 sg13g2_decap_8 FILLER_72_777 ();
 sg13g2_decap_8 FILLER_72_784 ();
 sg13g2_decap_8 FILLER_72_791 ();
 sg13g2_decap_8 FILLER_72_798 ();
 sg13g2_decap_8 FILLER_72_805 ();
 sg13g2_decap_8 FILLER_72_812 ();
 sg13g2_decap_8 FILLER_72_819 ();
 sg13g2_decap_8 FILLER_72_826 ();
 sg13g2_decap_8 FILLER_72_833 ();
 sg13g2_decap_8 FILLER_72_840 ();
 sg13g2_decap_8 FILLER_72_847 ();
 sg13g2_decap_8 FILLER_72_854 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_fill_1 FILLER_73_140 ();
 sg13g2_fill_1 FILLER_73_146 ();
 sg13g2_decap_4 FILLER_73_152 ();
 sg13g2_fill_1 FILLER_73_156 ();
 sg13g2_decap_4 FILLER_73_165 ();
 sg13g2_decap_4 FILLER_73_178 ();
 sg13g2_fill_2 FILLER_73_182 ();
 sg13g2_fill_2 FILLER_73_202 ();
 sg13g2_decap_4 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_233 ();
 sg13g2_decap_4 FILLER_73_271 ();
 sg13g2_fill_2 FILLER_73_275 ();
 sg13g2_decap_4 FILLER_73_304 ();
 sg13g2_fill_2 FILLER_73_335 ();
 sg13g2_fill_1 FILLER_73_361 ();
 sg13g2_fill_2 FILLER_73_376 ();
 sg13g2_fill_1 FILLER_73_378 ();
 sg13g2_fill_1 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_4 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_410 ();
 sg13g2_decap_8 FILLER_73_431 ();
 sg13g2_fill_1 FILLER_73_438 ();
 sg13g2_fill_1 FILLER_73_465 ();
 sg13g2_decap_8 FILLER_73_478 ();
 sg13g2_fill_2 FILLER_73_485 ();
 sg13g2_fill_1 FILLER_73_487 ();
 sg13g2_fill_2 FILLER_73_523 ();
 sg13g2_fill_2 FILLER_73_606 ();
 sg13g2_decap_8 FILLER_73_634 ();
 sg13g2_decap_8 FILLER_73_641 ();
 sg13g2_decap_4 FILLER_73_648 ();
 sg13g2_fill_2 FILLER_73_652 ();
 sg13g2_decap_8 FILLER_73_659 ();
 sg13g2_decap_4 FILLER_73_666 ();
 sg13g2_fill_1 FILLER_73_670 ();
 sg13g2_decap_4 FILLER_73_680 ();
 sg13g2_fill_1 FILLER_73_684 ();
 sg13g2_fill_1 FILLER_73_689 ();
 sg13g2_decap_8 FILLER_73_699 ();
 sg13g2_decap_8 FILLER_73_706 ();
 sg13g2_decap_8 FILLER_73_713 ();
 sg13g2_decap_8 FILLER_73_720 ();
 sg13g2_decap_8 FILLER_73_727 ();
 sg13g2_decap_8 FILLER_73_734 ();
 sg13g2_decap_8 FILLER_73_741 ();
 sg13g2_decap_8 FILLER_73_748 ();
 sg13g2_decap_8 FILLER_73_755 ();
 sg13g2_decap_8 FILLER_73_762 ();
 sg13g2_decap_8 FILLER_73_769 ();
 sg13g2_decap_8 FILLER_73_776 ();
 sg13g2_decap_8 FILLER_73_783 ();
 sg13g2_decap_8 FILLER_73_790 ();
 sg13g2_decap_8 FILLER_73_797 ();
 sg13g2_decap_8 FILLER_73_804 ();
 sg13g2_decap_8 FILLER_73_811 ();
 sg13g2_decap_8 FILLER_73_818 ();
 sg13g2_decap_8 FILLER_73_825 ();
 sg13g2_decap_8 FILLER_73_832 ();
 sg13g2_decap_8 FILLER_73_839 ();
 sg13g2_decap_8 FILLER_73_846 ();
 sg13g2_decap_8 FILLER_73_853 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_fill_2 FILLER_74_133 ();
 sg13g2_fill_2 FILLER_74_159 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_2 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_fill_2 FILLER_74_222 ();
 sg13g2_fill_2 FILLER_74_256 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_decap_4 FILLER_74_264 ();
 sg13g2_fill_1 FILLER_74_268 ();
 sg13g2_decap_8 FILLER_74_278 ();
 sg13g2_fill_1 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_312 ();
 sg13g2_decap_4 FILLER_74_319 ();
 sg13g2_fill_1 FILLER_74_323 ();
 sg13g2_decap_4 FILLER_74_328 ();
 sg13g2_fill_1 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_349 ();
 sg13g2_decap_4 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_365 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_fill_1 FILLER_74_385 ();
 sg13g2_fill_2 FILLER_74_392 ();
 sg13g2_fill_1 FILLER_74_402 ();
 sg13g2_fill_1 FILLER_74_413 ();
 sg13g2_fill_1 FILLER_74_437 ();
 sg13g2_decap_4 FILLER_74_443 ();
 sg13g2_fill_2 FILLER_74_447 ();
 sg13g2_fill_2 FILLER_74_466 ();
 sg13g2_fill_1 FILLER_74_468 ();
 sg13g2_decap_8 FILLER_74_486 ();
 sg13g2_decap_8 FILLER_74_493 ();
 sg13g2_decap_4 FILLER_74_500 ();
 sg13g2_fill_2 FILLER_74_504 ();
 sg13g2_fill_1 FILLER_74_546 ();
 sg13g2_fill_1 FILLER_74_560 ();
 sg13g2_fill_2 FILLER_74_582 ();
 sg13g2_fill_1 FILLER_74_584 ();
 sg13g2_fill_1 FILLER_74_598 ();
 sg13g2_decap_8 FILLER_74_607 ();
 sg13g2_decap_8 FILLER_74_614 ();
 sg13g2_decap_8 FILLER_74_621 ();
 sg13g2_decap_8 FILLER_74_628 ();
 sg13g2_decap_8 FILLER_74_635 ();
 sg13g2_decap_8 FILLER_74_642 ();
 sg13g2_decap_8 FILLER_74_649 ();
 sg13g2_decap_8 FILLER_74_656 ();
 sg13g2_decap_8 FILLER_74_663 ();
 sg13g2_decap_8 FILLER_74_670 ();
 sg13g2_decap_8 FILLER_74_677 ();
 sg13g2_decap_8 FILLER_74_684 ();
 sg13g2_decap_8 FILLER_74_691 ();
 sg13g2_decap_8 FILLER_74_698 ();
 sg13g2_decap_8 FILLER_74_705 ();
 sg13g2_decap_8 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_719 ();
 sg13g2_decap_8 FILLER_74_726 ();
 sg13g2_decap_8 FILLER_74_733 ();
 sg13g2_decap_8 FILLER_74_740 ();
 sg13g2_decap_8 FILLER_74_747 ();
 sg13g2_decap_8 FILLER_74_754 ();
 sg13g2_decap_8 FILLER_74_761 ();
 sg13g2_decap_8 FILLER_74_768 ();
 sg13g2_decap_8 FILLER_74_775 ();
 sg13g2_decap_8 FILLER_74_782 ();
 sg13g2_decap_8 FILLER_74_789 ();
 sg13g2_decap_8 FILLER_74_796 ();
 sg13g2_decap_8 FILLER_74_803 ();
 sg13g2_decap_8 FILLER_74_810 ();
 sg13g2_decap_8 FILLER_74_817 ();
 sg13g2_decap_8 FILLER_74_824 ();
 sg13g2_decap_8 FILLER_74_831 ();
 sg13g2_decap_8 FILLER_74_838 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_8 FILLER_74_852 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_4 FILLER_75_126 ();
 sg13g2_fill_2 FILLER_75_130 ();
 sg13g2_fill_2 FILLER_75_150 ();
 sg13g2_fill_2 FILLER_75_174 ();
 sg13g2_fill_2 FILLER_75_186 ();
 sg13g2_fill_1 FILLER_75_188 ();
 sg13g2_fill_1 FILLER_75_204 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_fill_2 FILLER_75_259 ();
 sg13g2_fill_1 FILLER_75_266 ();
 sg13g2_fill_2 FILLER_75_273 ();
 sg13g2_fill_2 FILLER_75_311 ();
 sg13g2_fill_2 FILLER_75_329 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_decap_4 FILLER_75_361 ();
 sg13g2_fill_1 FILLER_75_383 ();
 sg13g2_fill_1 FILLER_75_388 ();
 sg13g2_decap_4 FILLER_75_394 ();
 sg13g2_fill_1 FILLER_75_398 ();
 sg13g2_fill_2 FILLER_75_409 ();
 sg13g2_decap_4 FILLER_75_433 ();
 sg13g2_fill_2 FILLER_75_437 ();
 sg13g2_fill_2 FILLER_75_481 ();
 sg13g2_fill_2 FILLER_75_514 ();
 sg13g2_fill_1 FILLER_75_516 ();
 sg13g2_decap_8 FILLER_75_526 ();
 sg13g2_decap_8 FILLER_75_533 ();
 sg13g2_decap_4 FILLER_75_540 ();
 sg13g2_fill_2 FILLER_75_544 ();
 sg13g2_decap_8 FILLER_75_572 ();
 sg13g2_decap_8 FILLER_75_579 ();
 sg13g2_decap_8 FILLER_75_586 ();
 sg13g2_decap_8 FILLER_75_593 ();
 sg13g2_decap_8 FILLER_75_600 ();
 sg13g2_decap_8 FILLER_75_607 ();
 sg13g2_decap_8 FILLER_75_614 ();
 sg13g2_decap_8 FILLER_75_621 ();
 sg13g2_decap_8 FILLER_75_628 ();
 sg13g2_decap_8 FILLER_75_635 ();
 sg13g2_decap_8 FILLER_75_642 ();
 sg13g2_decap_8 FILLER_75_649 ();
 sg13g2_decap_8 FILLER_75_656 ();
 sg13g2_decap_8 FILLER_75_663 ();
 sg13g2_decap_8 FILLER_75_670 ();
 sg13g2_decap_8 FILLER_75_677 ();
 sg13g2_decap_8 FILLER_75_684 ();
 sg13g2_decap_8 FILLER_75_691 ();
 sg13g2_decap_8 FILLER_75_698 ();
 sg13g2_decap_8 FILLER_75_705 ();
 sg13g2_decap_8 FILLER_75_712 ();
 sg13g2_decap_8 FILLER_75_719 ();
 sg13g2_decap_8 FILLER_75_726 ();
 sg13g2_decap_8 FILLER_75_733 ();
 sg13g2_decap_8 FILLER_75_740 ();
 sg13g2_decap_8 FILLER_75_747 ();
 sg13g2_decap_8 FILLER_75_754 ();
 sg13g2_decap_8 FILLER_75_761 ();
 sg13g2_decap_8 FILLER_75_768 ();
 sg13g2_decap_8 FILLER_75_775 ();
 sg13g2_decap_8 FILLER_75_782 ();
 sg13g2_decap_8 FILLER_75_789 ();
 sg13g2_decap_8 FILLER_75_796 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_4 FILLER_76_133 ();
 sg13g2_fill_1 FILLER_76_137 ();
 sg13g2_fill_2 FILLER_76_157 ();
 sg13g2_decap_8 FILLER_76_174 ();
 sg13g2_decap_8 FILLER_76_181 ();
 sg13g2_decap_4 FILLER_76_188 ();
 sg13g2_fill_1 FILLER_76_198 ();
 sg13g2_decap_8 FILLER_76_204 ();
 sg13g2_decap_4 FILLER_76_228 ();
 sg13g2_decap_4 FILLER_76_238 ();
 sg13g2_decap_4 FILLER_76_259 ();
 sg13g2_fill_2 FILLER_76_275 ();
 sg13g2_fill_1 FILLER_76_277 ();
 sg13g2_decap_8 FILLER_76_310 ();
 sg13g2_decap_4 FILLER_76_317 ();
 sg13g2_decap_4 FILLER_76_328 ();
 sg13g2_fill_1 FILLER_76_332 ();
 sg13g2_fill_2 FILLER_76_388 ();
 sg13g2_fill_2 FILLER_76_396 ();
 sg13g2_fill_1 FILLER_76_398 ();
 sg13g2_fill_2 FILLER_76_415 ();
 sg13g2_fill_1 FILLER_76_417 ();
 sg13g2_decap_8 FILLER_76_430 ();
 sg13g2_fill_2 FILLER_76_437 ();
 sg13g2_decap_8 FILLER_76_457 ();
 sg13g2_fill_2 FILLER_76_464 ();
 sg13g2_fill_1 FILLER_76_466 ();
 sg13g2_decap_8 FILLER_76_473 ();
 sg13g2_decap_8 FILLER_76_480 ();
 sg13g2_decap_8 FILLER_76_487 ();
 sg13g2_decap_8 FILLER_76_498 ();
 sg13g2_decap_8 FILLER_76_505 ();
 sg13g2_decap_8 FILLER_76_512 ();
 sg13g2_decap_8 FILLER_76_519 ();
 sg13g2_decap_8 FILLER_76_526 ();
 sg13g2_decap_8 FILLER_76_533 ();
 sg13g2_decap_8 FILLER_76_540 ();
 sg13g2_decap_8 FILLER_76_547 ();
 sg13g2_decap_8 FILLER_76_554 ();
 sg13g2_decap_8 FILLER_76_561 ();
 sg13g2_decap_8 FILLER_76_568 ();
 sg13g2_decap_8 FILLER_76_575 ();
 sg13g2_decap_8 FILLER_76_582 ();
 sg13g2_decap_8 FILLER_76_589 ();
 sg13g2_decap_8 FILLER_76_596 ();
 sg13g2_decap_8 FILLER_76_603 ();
 sg13g2_decap_8 FILLER_76_610 ();
 sg13g2_decap_8 FILLER_76_617 ();
 sg13g2_decap_8 FILLER_76_624 ();
 sg13g2_decap_8 FILLER_76_631 ();
 sg13g2_decap_8 FILLER_76_638 ();
 sg13g2_decap_8 FILLER_76_645 ();
 sg13g2_decap_8 FILLER_76_652 ();
 sg13g2_decap_8 FILLER_76_659 ();
 sg13g2_decap_8 FILLER_76_666 ();
 sg13g2_decap_8 FILLER_76_673 ();
 sg13g2_decap_8 FILLER_76_680 ();
 sg13g2_decap_8 FILLER_76_687 ();
 sg13g2_decap_8 FILLER_76_694 ();
 sg13g2_decap_8 FILLER_76_701 ();
 sg13g2_decap_8 FILLER_76_708 ();
 sg13g2_decap_8 FILLER_76_715 ();
 sg13g2_decap_8 FILLER_76_722 ();
 sg13g2_decap_8 FILLER_76_729 ();
 sg13g2_decap_8 FILLER_76_736 ();
 sg13g2_decap_8 FILLER_76_743 ();
 sg13g2_decap_8 FILLER_76_750 ();
 sg13g2_decap_8 FILLER_76_757 ();
 sg13g2_decap_8 FILLER_76_764 ();
 sg13g2_decap_8 FILLER_76_771 ();
 sg13g2_decap_8 FILLER_76_778 ();
 sg13g2_decap_8 FILLER_76_785 ();
 sg13g2_decap_8 FILLER_76_792 ();
 sg13g2_decap_8 FILLER_76_799 ();
 sg13g2_decap_8 FILLER_76_806 ();
 sg13g2_decap_8 FILLER_76_813 ();
 sg13g2_decap_8 FILLER_76_820 ();
 sg13g2_decap_8 FILLER_76_827 ();
 sg13g2_decap_8 FILLER_76_834 ();
 sg13g2_decap_8 FILLER_76_841 ();
 sg13g2_decap_8 FILLER_76_848 ();
 sg13g2_decap_8 FILLER_76_855 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_fill_1 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_181 ();
 sg13g2_decap_8 FILLER_77_188 ();
 sg13g2_decap_4 FILLER_77_195 ();
 sg13g2_fill_1 FILLER_77_199 ();
 sg13g2_fill_2 FILLER_77_205 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_4 FILLER_77_266 ();
 sg13g2_fill_1 FILLER_77_270 ();
 sg13g2_fill_2 FILLER_77_278 ();
 sg13g2_fill_1 FILLER_77_280 ();
 sg13g2_fill_2 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_4 FILLER_77_308 ();
 sg13g2_fill_2 FILLER_77_312 ();
 sg13g2_fill_2 FILLER_77_330 ();
 sg13g2_fill_2 FILLER_77_340 ();
 sg13g2_fill_2 FILLER_77_352 ();
 sg13g2_fill_1 FILLER_77_354 ();
 sg13g2_fill_1 FILLER_77_367 ();
 sg13g2_decap_4 FILLER_77_376 ();
 sg13g2_decap_4 FILLER_77_391 ();
 sg13g2_decap_4 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_77_417 ();
 sg13g2_fill_2 FILLER_77_429 ();
 sg13g2_fill_1 FILLER_77_431 ();
 sg13g2_decap_8 FILLER_77_477 ();
 sg13g2_decap_8 FILLER_77_484 ();
 sg13g2_decap_8 FILLER_77_491 ();
 sg13g2_decap_8 FILLER_77_498 ();
 sg13g2_decap_8 FILLER_77_505 ();
 sg13g2_decap_8 FILLER_77_512 ();
 sg13g2_decap_8 FILLER_77_519 ();
 sg13g2_decap_8 FILLER_77_526 ();
 sg13g2_decap_8 FILLER_77_533 ();
 sg13g2_decap_8 FILLER_77_540 ();
 sg13g2_decap_8 FILLER_77_547 ();
 sg13g2_decap_8 FILLER_77_554 ();
 sg13g2_decap_8 FILLER_77_561 ();
 sg13g2_decap_8 FILLER_77_568 ();
 sg13g2_decap_8 FILLER_77_575 ();
 sg13g2_decap_8 FILLER_77_582 ();
 sg13g2_decap_8 FILLER_77_589 ();
 sg13g2_decap_8 FILLER_77_596 ();
 sg13g2_decap_8 FILLER_77_603 ();
 sg13g2_decap_8 FILLER_77_610 ();
 sg13g2_decap_8 FILLER_77_617 ();
 sg13g2_decap_8 FILLER_77_624 ();
 sg13g2_decap_8 FILLER_77_631 ();
 sg13g2_decap_8 FILLER_77_638 ();
 sg13g2_decap_8 FILLER_77_645 ();
 sg13g2_decap_8 FILLER_77_652 ();
 sg13g2_decap_8 FILLER_77_659 ();
 sg13g2_decap_8 FILLER_77_666 ();
 sg13g2_decap_8 FILLER_77_673 ();
 sg13g2_decap_8 FILLER_77_680 ();
 sg13g2_decap_8 FILLER_77_687 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_decap_8 FILLER_77_701 ();
 sg13g2_decap_8 FILLER_77_708 ();
 sg13g2_decap_8 FILLER_77_715 ();
 sg13g2_decap_8 FILLER_77_722 ();
 sg13g2_decap_8 FILLER_77_729 ();
 sg13g2_decap_8 FILLER_77_736 ();
 sg13g2_decap_8 FILLER_77_743 ();
 sg13g2_decap_8 FILLER_77_750 ();
 sg13g2_decap_8 FILLER_77_757 ();
 sg13g2_decap_8 FILLER_77_764 ();
 sg13g2_decap_8 FILLER_77_771 ();
 sg13g2_decap_8 FILLER_77_778 ();
 sg13g2_decap_8 FILLER_77_785 ();
 sg13g2_decap_8 FILLER_77_792 ();
 sg13g2_decap_8 FILLER_77_799 ();
 sg13g2_decap_8 FILLER_77_806 ();
 sg13g2_decap_8 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_820 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_decap_8 FILLER_77_834 ();
 sg13g2_decap_8 FILLER_77_841 ();
 sg13g2_decap_8 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_855 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_fill_1 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_164 ();
 sg13g2_fill_2 FILLER_78_183 ();
 sg13g2_fill_1 FILLER_78_185 ();
 sg13g2_decap_8 FILLER_78_190 ();
 sg13g2_decap_4 FILLER_78_197 ();
 sg13g2_fill_2 FILLER_78_201 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_4 FILLER_78_245 ();
 sg13g2_fill_2 FILLER_78_254 ();
 sg13g2_decap_4 FILLER_78_269 ();
 sg13g2_fill_1 FILLER_78_283 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_fill_1 FILLER_78_322 ();
 sg13g2_decap_4 FILLER_78_328 ();
 sg13g2_fill_1 FILLER_78_332 ();
 sg13g2_fill_2 FILLER_78_338 ();
 sg13g2_fill_2 FILLER_78_351 ();
 sg13g2_fill_2 FILLER_78_364 ();
 sg13g2_fill_2 FILLER_78_387 ();
 sg13g2_fill_1 FILLER_78_398 ();
 sg13g2_fill_2 FILLER_78_412 ();
 sg13g2_fill_2 FILLER_78_419 ();
 sg13g2_fill_1 FILLER_78_431 ();
 sg13g2_decap_4 FILLER_78_437 ();
 sg13g2_decap_8 FILLER_78_454 ();
 sg13g2_decap_8 FILLER_78_461 ();
 sg13g2_decap_8 FILLER_78_468 ();
 sg13g2_decap_8 FILLER_78_475 ();
 sg13g2_decap_8 FILLER_78_482 ();
 sg13g2_decap_8 FILLER_78_489 ();
 sg13g2_decap_8 FILLER_78_496 ();
 sg13g2_decap_8 FILLER_78_503 ();
 sg13g2_decap_8 FILLER_78_510 ();
 sg13g2_decap_8 FILLER_78_517 ();
 sg13g2_decap_8 FILLER_78_524 ();
 sg13g2_decap_8 FILLER_78_531 ();
 sg13g2_decap_8 FILLER_78_538 ();
 sg13g2_decap_8 FILLER_78_545 ();
 sg13g2_decap_8 FILLER_78_552 ();
 sg13g2_decap_8 FILLER_78_559 ();
 sg13g2_decap_8 FILLER_78_566 ();
 sg13g2_decap_8 FILLER_78_573 ();
 sg13g2_decap_8 FILLER_78_580 ();
 sg13g2_decap_8 FILLER_78_587 ();
 sg13g2_decap_8 FILLER_78_594 ();
 sg13g2_decap_8 FILLER_78_601 ();
 sg13g2_decap_8 FILLER_78_608 ();
 sg13g2_decap_8 FILLER_78_615 ();
 sg13g2_decap_8 FILLER_78_622 ();
 sg13g2_decap_8 FILLER_78_629 ();
 sg13g2_decap_8 FILLER_78_636 ();
 sg13g2_decap_8 FILLER_78_643 ();
 sg13g2_decap_8 FILLER_78_650 ();
 sg13g2_decap_8 FILLER_78_657 ();
 sg13g2_decap_8 FILLER_78_664 ();
 sg13g2_decap_8 FILLER_78_671 ();
 sg13g2_decap_8 FILLER_78_678 ();
 sg13g2_decap_8 FILLER_78_685 ();
 sg13g2_decap_8 FILLER_78_692 ();
 sg13g2_decap_8 FILLER_78_699 ();
 sg13g2_decap_8 FILLER_78_706 ();
 sg13g2_decap_8 FILLER_78_713 ();
 sg13g2_decap_8 FILLER_78_720 ();
 sg13g2_decap_8 FILLER_78_727 ();
 sg13g2_decap_8 FILLER_78_734 ();
 sg13g2_decap_8 FILLER_78_741 ();
 sg13g2_decap_8 FILLER_78_748 ();
 sg13g2_decap_8 FILLER_78_755 ();
 sg13g2_decap_8 FILLER_78_762 ();
 sg13g2_decap_8 FILLER_78_769 ();
 sg13g2_decap_8 FILLER_78_776 ();
 sg13g2_decap_8 FILLER_78_783 ();
 sg13g2_decap_8 FILLER_78_790 ();
 sg13g2_decap_8 FILLER_78_797 ();
 sg13g2_decap_8 FILLER_78_804 ();
 sg13g2_decap_8 FILLER_78_811 ();
 sg13g2_decap_8 FILLER_78_818 ();
 sg13g2_decap_8 FILLER_78_825 ();
 sg13g2_decap_8 FILLER_78_832 ();
 sg13g2_decap_8 FILLER_78_839 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_853 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_4 FILLER_79_161 ();
 sg13g2_fill_1 FILLER_79_165 ();
 sg13g2_decap_4 FILLER_79_201 ();
 sg13g2_fill_1 FILLER_79_205 ();
 sg13g2_fill_1 FILLER_79_219 ();
 sg13g2_decap_8 FILLER_79_256 ();
 sg13g2_fill_2 FILLER_79_263 ();
 sg13g2_fill_1 FILLER_79_265 ();
 sg13g2_fill_1 FILLER_79_281 ();
 sg13g2_fill_2 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_307 ();
 sg13g2_decap_8 FILLER_79_314 ();
 sg13g2_fill_2 FILLER_79_321 ();
 sg13g2_fill_1 FILLER_79_323 ();
 sg13g2_fill_2 FILLER_79_338 ();
 sg13g2_fill_1 FILLER_79_340 ();
 sg13g2_decap_4 FILLER_79_350 ();
 sg13g2_fill_2 FILLER_79_390 ();
 sg13g2_fill_1 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_412 ();
 sg13g2_fill_2 FILLER_79_419 ();
 sg13g2_decap_8 FILLER_79_442 ();
 sg13g2_decap_8 FILLER_79_449 ();
 sg13g2_decap_8 FILLER_79_456 ();
 sg13g2_decap_8 FILLER_79_463 ();
 sg13g2_decap_8 FILLER_79_470 ();
 sg13g2_decap_8 FILLER_79_477 ();
 sg13g2_decap_8 FILLER_79_484 ();
 sg13g2_decap_8 FILLER_79_491 ();
 sg13g2_decap_8 FILLER_79_498 ();
 sg13g2_decap_8 FILLER_79_505 ();
 sg13g2_decap_8 FILLER_79_512 ();
 sg13g2_decap_8 FILLER_79_519 ();
 sg13g2_decap_8 FILLER_79_526 ();
 sg13g2_decap_8 FILLER_79_533 ();
 sg13g2_decap_8 FILLER_79_540 ();
 sg13g2_decap_8 FILLER_79_547 ();
 sg13g2_decap_8 FILLER_79_554 ();
 sg13g2_decap_8 FILLER_79_561 ();
 sg13g2_decap_8 FILLER_79_568 ();
 sg13g2_decap_8 FILLER_79_575 ();
 sg13g2_decap_8 FILLER_79_582 ();
 sg13g2_decap_8 FILLER_79_589 ();
 sg13g2_decap_8 FILLER_79_596 ();
 sg13g2_decap_8 FILLER_79_603 ();
 sg13g2_decap_8 FILLER_79_610 ();
 sg13g2_decap_8 FILLER_79_617 ();
 sg13g2_decap_8 FILLER_79_624 ();
 sg13g2_decap_8 FILLER_79_631 ();
 sg13g2_decap_8 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_645 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_8 FILLER_79_659 ();
 sg13g2_decap_8 FILLER_79_666 ();
 sg13g2_decap_8 FILLER_79_673 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_687 ();
 sg13g2_decap_8 FILLER_79_694 ();
 sg13g2_decap_8 FILLER_79_701 ();
 sg13g2_decap_8 FILLER_79_708 ();
 sg13g2_decap_8 FILLER_79_715 ();
 sg13g2_decap_8 FILLER_79_722 ();
 sg13g2_decap_8 FILLER_79_729 ();
 sg13g2_decap_8 FILLER_79_736 ();
 sg13g2_decap_8 FILLER_79_743 ();
 sg13g2_decap_8 FILLER_79_750 ();
 sg13g2_decap_8 FILLER_79_757 ();
 sg13g2_decap_8 FILLER_79_764 ();
 sg13g2_decap_8 FILLER_79_771 ();
 sg13g2_decap_8 FILLER_79_778 ();
 sg13g2_decap_8 FILLER_79_785 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_827 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_fill_1 FILLER_80_156 ();
 sg13g2_decap_8 FILLER_80_195 ();
 sg13g2_decap_8 FILLER_80_202 ();
 sg13g2_fill_2 FILLER_80_209 ();
 sg13g2_decap_8 FILLER_80_245 ();
 sg13g2_decap_4 FILLER_80_252 ();
 sg13g2_fill_1 FILLER_80_256 ();
 sg13g2_decap_4 FILLER_80_288 ();
 sg13g2_decap_8 FILLER_80_318 ();
 sg13g2_decap_8 FILLER_80_325 ();
 sg13g2_fill_1 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_338 ();
 sg13g2_fill_1 FILLER_80_342 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_fill_1 FILLER_80_355 ();
 sg13g2_fill_2 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_4 FILLER_80_397 ();
 sg13g2_fill_2 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_413 ();
 sg13g2_decap_8 FILLER_80_420 ();
 sg13g2_decap_8 FILLER_80_427 ();
 sg13g2_decap_8 FILLER_80_434 ();
 sg13g2_decap_8 FILLER_80_441 ();
 sg13g2_decap_8 FILLER_80_448 ();
 sg13g2_decap_8 FILLER_80_455 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_decap_8 FILLER_80_469 ();
 sg13g2_decap_8 FILLER_80_476 ();
 sg13g2_decap_8 FILLER_80_483 ();
 sg13g2_decap_8 FILLER_80_490 ();
 sg13g2_decap_8 FILLER_80_497 ();
 sg13g2_decap_8 FILLER_80_504 ();
 sg13g2_decap_8 FILLER_80_511 ();
 sg13g2_decap_8 FILLER_80_518 ();
 sg13g2_decap_8 FILLER_80_525 ();
 sg13g2_decap_8 FILLER_80_532 ();
 sg13g2_decap_8 FILLER_80_539 ();
 sg13g2_decap_8 FILLER_80_546 ();
 sg13g2_decap_8 FILLER_80_553 ();
 sg13g2_decap_8 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_567 ();
 sg13g2_decap_8 FILLER_80_574 ();
 sg13g2_decap_8 FILLER_80_581 ();
 sg13g2_decap_8 FILLER_80_588 ();
 sg13g2_decap_8 FILLER_80_595 ();
 sg13g2_decap_8 FILLER_80_602 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_decap_8 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_623 ();
 sg13g2_decap_8 FILLER_80_630 ();
 sg13g2_decap_8 FILLER_80_637 ();
 sg13g2_decap_8 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_651 ();
 sg13g2_decap_8 FILLER_80_658 ();
 sg13g2_decap_8 FILLER_80_665 ();
 sg13g2_decap_8 FILLER_80_672 ();
 sg13g2_decap_8 FILLER_80_679 ();
 sg13g2_decap_8 FILLER_80_686 ();
 sg13g2_decap_8 FILLER_80_693 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_8 FILLER_80_707 ();
 sg13g2_decap_8 FILLER_80_714 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net164;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule

module tt_um_multiplier_tt10 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire \mul_uut.C1.fa_1.sum ;
 wire \mul_uut.C1.fa_5.sum ;
 wire \mul_uut.C1.fa_6.sum ;
 wire \mul_uut.C1.ha_5.sum ;
 wire \mul_uut.C2.fa_4.sum ;
 wire \mul_uut.C2.fa_5.sum ;
 wire \mul_uut.C2.fa_6.sum ;
 wire \mul_uut.C2.fa_7.sum ;
 wire \mul_uut.C2.ha_1.sum ;
 wire \mul_uut.C2.ha_6.sum ;
 wire \mul_uut.C2.ha_8.sum ;
 wire \mul_uut.N1.C1.fa_1.sum ;
 wire \mul_uut.N1.C1.ha_3.sum ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;

 sg13g2_a22oi_1 _295_ (.Y(_227_),
    .B1(net71),
    .B2(net62),
    .A2(net72),
    .A1(net61));
 sg13g2_nand2_2 _296_ (.Y(_229_),
    .A(net62),
    .B(net72));
 sg13g2_nand2_1 _297_ (.Y(_230_),
    .A(net61),
    .B(net71));
 sg13g2_nor2_1 _298_ (.A(_229_),
    .B(_230_),
    .Y(_231_));
 sg13g2_nor2_1 _299_ (.A(_227_),
    .B(_231_),
    .Y(_232_));
 sg13g2_nand2_1 _300_ (.Y(_233_),
    .A(net75),
    .B(net62));
 sg13g2_nand4_1 _301_ (.B(net75),
    .C(net73),
    .A(net61),
    .Y(_234_),
    .D(net62));
 sg13g2_inv_1 _302_ (.Y(_235_),
    .A(_234_));
 sg13g2_nand2_1 _303_ (.Y(_236_),
    .A(net65),
    .B(net72));
 sg13g2_nand4_1 _304_ (.B(net63),
    .C(net72),
    .A(net65),
    .Y(_237_),
    .D(net71));
 sg13g2_inv_1 _305_ (.Y(_238_),
    .A(_237_));
 sg13g2_nand2_1 _306_ (.Y(_239_),
    .A(_235_),
    .B(_238_));
 sg13g2_nand2_1 _307_ (.Y(_240_),
    .A(_234_),
    .B(_237_));
 sg13g2_nand3_1 _308_ (.B(net73),
    .C(_233_),
    .A(net61),
    .Y(_241_));
 sg13g2_nand3_1 _309_ (.B(net71),
    .C(_236_),
    .A(net63),
    .Y(_242_));
 sg13g2_nor2_1 _310_ (.A(_241_),
    .B(_242_),
    .Y(_243_));
 sg13g2_a21oi_1 _311_ (.A1(_239_),
    .A2(_240_),
    .Y(_244_),
    .B1(_243_));
 sg13g2_a22oi_1 _312_ (.Y(_245_),
    .B1(net73),
    .B2(net62),
    .A2(net75),
    .A1(net61));
 sg13g2_nor2_1 _313_ (.A(_235_),
    .B(_245_),
    .Y(_246_));
 sg13g2_a22oi_1 _314_ (.Y(_247_),
    .B1(net71),
    .B2(net65),
    .A2(net72),
    .A1(net63));
 sg13g2_nor2_1 _315_ (.A(_238_),
    .B(_247_),
    .Y(_248_));
 sg13g2_nand2_1 _316_ (.Y(_249_),
    .A(net65),
    .B(net73));
 sg13g2_nand2_1 _317_ (.Y(_250_),
    .A(net75),
    .B(net63));
 sg13g2_nand2_2 _318_ (.Y(_251_),
    .A(net75),
    .B(net65));
 sg13g2_or2_1 _319_ (.X(_252_),
    .B(_250_),
    .A(_249_));
 sg13g2_xnor2_1 _320_ (.Y(_253_),
    .A(_246_),
    .B(_248_));
 sg13g2_nor2_1 _321_ (.A(_252_),
    .B(_253_),
    .Y(_254_));
 sg13g2_a21oi_1 _322_ (.A1(_246_),
    .A2(_248_),
    .Y(_255_),
    .B1(_254_));
 sg13g2_xnor2_1 _323_ (.Y(_256_),
    .A(_241_),
    .B(_242_));
 sg13g2_nor2_1 _324_ (.A(_255_),
    .B(_256_),
    .Y(_257_));
 sg13g2_xor2_1 _325_ (.B(_236_),
    .A(_233_),
    .X(_258_));
 sg13g2_nand3_1 _326_ (.B(net73),
    .C(_251_),
    .A(net63),
    .Y(_259_));
 sg13g2_nand4_1 _327_ (.B(net73),
    .C(_251_),
    .A(net63),
    .Y(_260_),
    .D(_258_));
 sg13g2_o21ai_1 _328_ (.B1(_260_),
    .Y(_261_),
    .A1(_229_),
    .A2(_251_));
 sg13g2_xor2_1 _329_ (.B(_253_),
    .A(_252_),
    .X(_262_));
 sg13g2_nand2_1 _330_ (.Y(_263_),
    .A(_261_),
    .B(_262_));
 sg13g2_xnor2_1 _331_ (.Y(_264_),
    .A(_255_),
    .B(_256_));
 sg13g2_nor2_1 _332_ (.A(_263_),
    .B(_264_),
    .Y(_265_));
 sg13g2_nor2_1 _333_ (.A(_257_),
    .B(_265_),
    .Y(_266_));
 sg13g2_xnor2_1 _334_ (.Y(_267_),
    .A(_244_),
    .B(_266_));
 sg13g2_or3_1 _335_ (.A(_227_),
    .B(_231_),
    .C(_267_),
    .X(_268_));
 sg13g2_xor2_1 _336_ (.B(_264_),
    .A(_263_),
    .X(_269_));
 sg13g2_nand2b_1 _337_ (.Y(_270_),
    .B(_269_),
    .A_N(_229_));
 sg13g2_xor2_1 _338_ (.B(_267_),
    .A(_232_),
    .X(_271_));
 sg13g2_o21ai_1 _339_ (.B1(_268_),
    .Y(_272_),
    .A1(_270_),
    .A2(_271_));
 sg13g2_nand2b_1 _340_ (.Y(_273_),
    .B(_229_),
    .A_N(_230_));
 sg13g2_o21ai_1 _341_ (.B1(_239_),
    .Y(_274_),
    .A1(_244_),
    .A2(_266_));
 sg13g2_nand2b_1 _342_ (.Y(_275_),
    .B(_274_),
    .A_N(_273_));
 sg13g2_xnor2_1 _343_ (.Y(_276_),
    .A(_273_),
    .B(_274_));
 sg13g2_xor2_1 _344_ (.B(_276_),
    .A(_272_),
    .X(_277_));
 sg13g2_xnor2_1 _345_ (.Y(_278_),
    .A(_229_),
    .B(_269_));
 sg13g2_nand2_2 _346_ (.Y(_279_),
    .A(net77),
    .B(net11));
 sg13g2_nand2_1 _347_ (.Y(_280_),
    .A(net12),
    .B(net76));
 sg13g2_nor2_1 _348_ (.A(_279_),
    .B(_280_),
    .Y(_281_));
 sg13g2_a22oi_1 _349_ (.Y(_282_),
    .B1(net11),
    .B2(net76),
    .A2(net77),
    .A1(net12));
 sg13g2_nor2_1 _350_ (.A(_281_),
    .B(_282_),
    .Y(_283_));
 sg13g2_inv_1 _351_ (.Y(_284_),
    .A(_283_));
 sg13g2_nand2_1 _352_ (.Y(_285_),
    .A(net80),
    .B(net62));
 sg13g2_nand4_1 _353_ (.B(net78),
    .C(net80),
    .A(net61),
    .Y(_286_),
    .D(net62));
 sg13g2_inv_1 _354_ (.Y(_287_),
    .A(_286_));
 sg13g2_nand2_1 _355_ (.Y(_288_),
    .A(net10),
    .B(net77));
 sg13g2_nand4_1 _356_ (.B(net76),
    .C(net77),
    .A(net10),
    .Y(_289_),
    .D(net64));
 sg13g2_inv_1 _357_ (.Y(_290_),
    .A(_289_));
 sg13g2_xor2_1 _358_ (.B(_289_),
    .A(_286_),
    .X(_291_));
 sg13g2_nand3_1 _359_ (.B(net78),
    .C(_285_),
    .A(net61),
    .Y(_292_));
 sg13g2_nand3_1 _360_ (.B(net64),
    .C(_288_),
    .A(net76),
    .Y(_293_));
 sg13g2_nor2_1 _361_ (.A(_292_),
    .B(_293_),
    .Y(_294_));
 sg13g2_nor2_1 _362_ (.A(_291_),
    .B(_294_),
    .Y(_000_));
 sg13g2_a22oi_1 _363_ (.Y(_001_),
    .B1(net62),
    .B2(net78),
    .A2(net80),
    .A1(net61));
 sg13g2_nor2_1 _364_ (.A(_287_),
    .B(_001_),
    .Y(_002_));
 sg13g2_a22oi_1 _365_ (.Y(_003_),
    .B1(net77),
    .B2(net64),
    .A2(net76),
    .A1(net65));
 sg13g2_nor2_1 _366_ (.A(_290_),
    .B(_003_),
    .Y(_004_));
 sg13g2_nand2_1 _367_ (.Y(_005_),
    .A(net78),
    .B(net65));
 sg13g2_nand2_1 _368_ (.Y(_006_),
    .A(net80),
    .B(net64));
 sg13g2_nand2_2 _369_ (.Y(_007_),
    .A(net80),
    .B(net65));
 sg13g2_or2_1 _370_ (.X(_008_),
    .B(_006_),
    .A(_005_));
 sg13g2_xnor2_1 _371_ (.Y(_009_),
    .A(_002_),
    .B(_004_));
 sg13g2_nor2_1 _372_ (.A(_008_),
    .B(_009_),
    .Y(_010_));
 sg13g2_a21oi_1 _373_ (.A1(_002_),
    .A2(_004_),
    .Y(_011_),
    .B1(_010_));
 sg13g2_xnor2_1 _374_ (.Y(_012_),
    .A(_292_),
    .B(_293_));
 sg13g2_nor2_1 _375_ (.A(_011_),
    .B(_012_),
    .Y(_013_));
 sg13g2_xor2_1 _376_ (.B(_288_),
    .A(_285_),
    .X(_014_));
 sg13g2_nand3_1 _377_ (.B(net63),
    .C(_007_),
    .A(net78),
    .Y(_015_));
 sg13g2_nand4_1 _378_ (.B(net63),
    .C(_007_),
    .A(net78),
    .Y(_016_),
    .D(_014_));
 sg13g2_o21ai_1 _379_ (.B1(_016_),
    .Y(_017_),
    .A1(_279_),
    .A2(_007_));
 sg13g2_xor2_1 _380_ (.B(_009_),
    .A(_008_),
    .X(_018_));
 sg13g2_nand2_1 _381_ (.Y(_019_),
    .A(_017_),
    .B(_018_));
 sg13g2_xnor2_1 _382_ (.Y(_020_),
    .A(_011_),
    .B(_012_));
 sg13g2_nor2_1 _383_ (.A(_019_),
    .B(_020_),
    .Y(_021_));
 sg13g2_nor2_1 _384_ (.A(_013_),
    .B(_021_),
    .Y(_022_));
 sg13g2_nor2_1 _385_ (.A(_000_),
    .B(_022_),
    .Y(_023_));
 sg13g2_xnor2_1 _386_ (.Y(_024_),
    .A(_000_),
    .B(_022_));
 sg13g2_nor2_1 _387_ (.A(_284_),
    .B(_024_),
    .Y(_025_));
 sg13g2_xor2_1 _388_ (.B(_020_),
    .A(_019_),
    .X(_026_));
 sg13g2_nand2b_1 _389_ (.Y(_027_),
    .B(_026_),
    .A_N(_279_));
 sg13g2_xnor2_1 _390_ (.Y(_028_),
    .A(_284_),
    .B(_024_));
 sg13g2_nor2_1 _391_ (.A(_027_),
    .B(_028_),
    .Y(_029_));
 sg13g2_nor2b_1 _392_ (.A(_280_),
    .B_N(_279_),
    .Y(_030_));
 sg13g2_a21oi_1 _393_ (.A1(_287_),
    .A2(_290_),
    .Y(_031_),
    .B1(_023_));
 sg13g2_xnor2_1 _394_ (.Y(_032_),
    .A(_030_),
    .B(_031_));
 sg13g2_o21ai_1 _395_ (.B1(_032_),
    .Y(_033_),
    .A1(_025_),
    .A2(_029_));
 sg13g2_a21oi_1 _396_ (.A1(_279_),
    .A2(_031_),
    .Y(_034_),
    .B1(_280_));
 sg13g2_nand2b_1 _397_ (.Y(_035_),
    .B(_033_),
    .A_N(_034_));
 sg13g2_nand2_2 _398_ (.Y(_036_),
    .A(net67),
    .B(net5));
 sg13g2_and4_1 _399_ (.A(net67),
    .B(net66),
    .C(net5),
    .D(net6),
    .X(_037_));
 sg13g2_a22oi_1 _400_ (.Y(_038_),
    .B1(net6),
    .B2(net67),
    .A2(net5),
    .A1(net66));
 sg13g2_nor2_1 _401_ (.A(_037_),
    .B(_038_),
    .Y(_039_));
 sg13g2_nand2_1 _402_ (.Y(_040_),
    .A(net4),
    .B(net67));
 sg13g2_nand4_1 _403_ (.B(net8),
    .C(net9),
    .A(net4),
    .Y(_041_),
    .D(net74));
 sg13g2_inv_1 _404_ (.Y(_042_),
    .A(_041_));
 sg13g2_nand2_1 _405_ (.Y(_043_),
    .A(net70),
    .B(net72));
 sg13g2_nand4_1 _406_ (.B(net68),
    .C(net72),
    .A(net70),
    .Y(_044_),
    .D(net6));
 sg13g2_inv_1 _407_ (.Y(_045_),
    .A(_044_));
 sg13g2_nand2_1 _408_ (.Y(_046_),
    .A(_042_),
    .B(_045_));
 sg13g2_nand2_1 _409_ (.Y(_047_),
    .A(_041_),
    .B(_044_));
 sg13g2_nand3_1 _410_ (.B(net74),
    .C(_040_),
    .A(net66),
    .Y(_048_));
 sg13g2_nand3_1 _411_ (.B(net71),
    .C(_043_),
    .A(net68),
    .Y(_049_));
 sg13g2_nor2_1 _412_ (.A(_048_),
    .B(_049_),
    .Y(_050_));
 sg13g2_a21oi_1 _413_ (.A1(_046_),
    .A2(_047_),
    .Y(_051_),
    .B1(_050_));
 sg13g2_a22oi_1 _414_ (.Y(_052_),
    .B1(net74),
    .B2(net67),
    .A2(net9),
    .A1(net75));
 sg13g2_nor2_1 _415_ (.A(_042_),
    .B(_052_),
    .Y(_053_));
 sg13g2_a22oi_1 _416_ (.Y(_054_),
    .B1(net71),
    .B2(net70),
    .A2(net72),
    .A1(net68));
 sg13g2_nor2_1 _417_ (.A(_045_),
    .B(_054_),
    .Y(_055_));
 sg13g2_nand2_1 _418_ (.Y(_056_),
    .A(net70),
    .B(net74));
 sg13g2_nand2_1 _419_ (.Y(_057_),
    .A(net75),
    .B(net69));
 sg13g2_nand2_2 _420_ (.Y(_058_),
    .A(net70),
    .B(net75));
 sg13g2_or2_1 _421_ (.X(_059_),
    .B(_057_),
    .A(_056_));
 sg13g2_xnor2_1 _422_ (.Y(_060_),
    .A(_053_),
    .B(_055_));
 sg13g2_nor2_1 _423_ (.A(_059_),
    .B(_060_),
    .Y(_061_));
 sg13g2_a21oi_1 _424_ (.A1(_053_),
    .A2(_055_),
    .Y(_062_),
    .B1(_061_));
 sg13g2_xnor2_1 _425_ (.Y(_063_),
    .A(_048_),
    .B(_049_));
 sg13g2_nor2_1 _426_ (.A(_062_),
    .B(_063_),
    .Y(_064_));
 sg13g2_xor2_1 _427_ (.B(_043_),
    .A(_040_),
    .X(_065_));
 sg13g2_nand3_1 _428_ (.B(net73),
    .C(_058_),
    .A(net68),
    .Y(_066_));
 sg13g2_nand4_1 _429_ (.B(net73),
    .C(_058_),
    .A(net68),
    .Y(_067_),
    .D(_065_));
 sg13g2_o21ai_1 _430_ (.B1(_067_),
    .Y(_068_),
    .A1(_036_),
    .A2(_058_));
 sg13g2_xor2_1 _431_ (.B(_060_),
    .A(_059_),
    .X(_069_));
 sg13g2_nand2_1 _432_ (.Y(_070_),
    .A(_068_),
    .B(_069_));
 sg13g2_xnor2_1 _433_ (.Y(_071_),
    .A(_062_),
    .B(_063_));
 sg13g2_nor2_1 _434_ (.A(_070_),
    .B(_071_),
    .Y(_072_));
 sg13g2_nor2_1 _435_ (.A(_064_),
    .B(_072_),
    .Y(_073_));
 sg13g2_xnor2_1 _436_ (.Y(_074_),
    .A(_051_),
    .B(_073_));
 sg13g2_or3_1 _437_ (.A(_037_),
    .B(_038_),
    .C(_074_),
    .X(_075_));
 sg13g2_xor2_1 _438_ (.B(_071_),
    .A(_070_),
    .X(_076_));
 sg13g2_nand2b_1 _439_ (.Y(_077_),
    .B(_076_),
    .A_N(_036_));
 sg13g2_xor2_1 _440_ (.B(_074_),
    .A(_039_),
    .X(_078_));
 sg13g2_o21ai_1 _441_ (.B1(_075_),
    .Y(_079_),
    .A1(_077_),
    .A2(_078_));
 sg13g2_nand3_1 _442_ (.B(net71),
    .C(_036_),
    .A(net66),
    .Y(_080_));
 sg13g2_o21ai_1 _443_ (.B1(_046_),
    .Y(_081_),
    .A1(_051_),
    .A2(_073_));
 sg13g2_nand2b_1 _444_ (.Y(_082_),
    .B(_081_),
    .A_N(_080_));
 sg13g2_xnor2_1 _445_ (.Y(_083_),
    .A(_080_),
    .B(_081_));
 sg13g2_a21oi_1 _446_ (.A1(_079_),
    .A2(_083_),
    .Y(_084_),
    .B1(_037_));
 sg13g2_nand2_1 _447_ (.Y(_085_),
    .A(_082_),
    .B(_084_));
 sg13g2_xor2_1 _448_ (.B(_085_),
    .A(_035_),
    .X(_086_));
 sg13g2_inv_1 _449_ (.Y(_087_),
    .A(_086_));
 sg13g2_or3_1 _450_ (.A(_025_),
    .B(_029_),
    .C(_032_),
    .X(_088_));
 sg13g2_nand2_1 _451_ (.Y(_089_),
    .A(_033_),
    .B(_088_));
 sg13g2_xnor2_1 _452_ (.Y(_090_),
    .A(_079_),
    .B(_083_));
 sg13g2_nor2_1 _453_ (.A(_089_),
    .B(_090_),
    .Y(_091_));
 sg13g2_xor2_1 _454_ (.B(_078_),
    .A(_077_),
    .X(_092_));
 sg13g2_xor2_1 _455_ (.B(_028_),
    .A(_027_),
    .X(_093_));
 sg13g2_nand2_1 _456_ (.Y(_094_),
    .A(_092_),
    .B(_093_));
 sg13g2_xnor2_1 _457_ (.Y(_095_),
    .A(_036_),
    .B(_076_));
 sg13g2_xnor2_1 _458_ (.Y(_096_),
    .A(_279_),
    .B(_026_));
 sg13g2_and2_1 _459_ (.A(_095_),
    .B(_096_),
    .X(_097_));
 sg13g2_xor2_1 _460_ (.B(_006_),
    .A(_005_),
    .X(_098_));
 sg13g2_xor2_1 _461_ (.B(_057_),
    .A(_056_),
    .X(_099_));
 sg13g2_and2_1 _462_ (.A(_098_),
    .B(_099_),
    .X(_100_));
 sg13g2_or2_1 _463_ (.X(_101_),
    .B(_099_),
    .A(_098_));
 sg13g2_nand2b_1 _464_ (.Y(_102_),
    .B(_101_),
    .A_N(_100_));
 sg13g2_nand2_2 _465_ (.Y(_103_),
    .A(net8),
    .B(net2));
 sg13g2_nand2_1 _466_ (.Y(_104_),
    .A(net7),
    .B(net1));
 sg13g2_inv_1 _467_ (.Y(uo_out[0]),
    .A(_104_));
 sg13g2_nand2_1 _468_ (.Y(_105_),
    .A(net1),
    .B(net8));
 sg13g2_nand2_1 _469_ (.Y(_106_),
    .A(net70),
    .B(net2));
 sg13g2_xor2_1 _470_ (.B(_106_),
    .A(_105_),
    .X(_107_));
 sg13g2_nand3_1 _471_ (.B(net69),
    .C(_104_),
    .A(net79),
    .Y(_108_));
 sg13g2_nand4_1 _472_ (.B(net69),
    .C(_104_),
    .A(net79),
    .Y(_109_),
    .D(_107_));
 sg13g2_o21ai_1 _473_ (.B1(_109_),
    .Y(_110_),
    .A1(_103_),
    .A2(_104_));
 sg13g2_and3_1 _474_ (.X(_111_),
    .A(net79),
    .B(net69),
    .C(uo_out[0]));
 sg13g2_a22oi_1 _475_ (.Y(_112_),
    .B1(net68),
    .B2(net77),
    .A2(net3),
    .A1(net70));
 sg13g2_nand4_1 _476_ (.B(net3),
    .C(net68),
    .A(net7),
    .Y(_113_),
    .D(net77));
 sg13g2_nand2b_1 _477_ (.Y(_114_),
    .B(_113_),
    .A_N(_112_));
 sg13g2_a22oi_1 _478_ (.Y(_115_),
    .B1(net9),
    .B2(net80),
    .A2(net67),
    .A1(net78));
 sg13g2_nand4_1 _479_ (.B(net80),
    .C(net67),
    .A(net79),
    .Y(_116_),
    .D(net66));
 sg13g2_nand2b_1 _480_ (.Y(_117_),
    .B(_116_),
    .A_N(_115_));
 sg13g2_nor2_1 _481_ (.A(_114_),
    .B(_117_),
    .Y(_118_));
 sg13g2_nand2_1 _482_ (.Y(_119_),
    .A(_114_),
    .B(_117_));
 sg13g2_xnor2_1 _483_ (.Y(_120_),
    .A(_114_),
    .B(_117_));
 sg13g2_xnor2_1 _484_ (.Y(_121_),
    .A(_111_),
    .B(_120_));
 sg13g2_and2_1 _485_ (.A(_110_),
    .B(_121_),
    .X(_122_));
 sg13g2_a21oi_2 _486_ (.B1(_118_),
    .Y(_123_),
    .A2(_119_),
    .A1(_111_));
 sg13g2_nand3_1 _487_ (.B(net66),
    .C(_105_),
    .A(net79),
    .Y(_124_));
 sg13g2_nand3_1 _488_ (.B(net69),
    .C(_106_),
    .A(net76),
    .Y(_125_));
 sg13g2_nor2_1 _489_ (.A(_124_),
    .B(_125_),
    .Y(_126_));
 sg13g2_xnor2_1 _490_ (.Y(_127_),
    .A(_124_),
    .B(_125_));
 sg13g2_nor2_1 _491_ (.A(_123_),
    .B(_127_),
    .Y(_128_));
 sg13g2_nand2_1 _492_ (.Y(_129_),
    .A(_123_),
    .B(_127_));
 sg13g2_xnor2_1 _493_ (.Y(_130_),
    .A(_123_),
    .B(_127_));
 sg13g2_xnor2_1 _494_ (.Y(_131_),
    .A(_122_),
    .B(_130_));
 sg13g2_nand2b_1 _495_ (.Y(_132_),
    .B(_131_),
    .A_N(_103_));
 sg13g2_inv_1 _496_ (.Y(_133_),
    .A(_132_));
 sg13g2_nand2_1 _497_ (.Y(_134_),
    .A(net67),
    .B(net76));
 sg13g2_nand2_1 _498_ (.Y(_135_),
    .A(net66),
    .B(net77));
 sg13g2_or2_1 _499_ (.X(_136_),
    .B(_135_),
    .A(_134_));
 sg13g2_xor2_1 _500_ (.B(_135_),
    .A(_134_),
    .X(_137_));
 sg13g2_inv_1 _501_ (.Y(_138_),
    .A(_137_));
 sg13g2_a21oi_1 _502_ (.A1(_122_),
    .A2(_129_),
    .Y(_139_),
    .B1(_128_));
 sg13g2_nand2_1 _503_ (.Y(_140_),
    .A(_113_),
    .B(_116_));
 sg13g2_or2_1 _504_ (.X(_141_),
    .B(_116_),
    .A(_113_));
 sg13g2_a21oi_1 _505_ (.A1(_140_),
    .A2(_141_),
    .Y(_142_),
    .B1(_126_));
 sg13g2_xnor2_1 _506_ (.Y(_143_),
    .A(_139_),
    .B(_142_));
 sg13g2_nor2_1 _507_ (.A(_138_),
    .B(_143_),
    .Y(_144_));
 sg13g2_xnor2_1 _508_ (.Y(_145_),
    .A(_137_),
    .B(_143_));
 sg13g2_xnor2_1 _509_ (.Y(_146_),
    .A(_132_),
    .B(_145_));
 sg13g2_xnor2_1 _510_ (.Y(_147_),
    .A(_102_),
    .B(_146_));
 sg13g2_xnor2_1 _511_ (.Y(_148_),
    .A(_103_),
    .B(_131_));
 sg13g2_xor2_1 _512_ (.B(_058_),
    .A(_007_),
    .X(_149_));
 sg13g2_nand2_1 _513_ (.Y(_150_),
    .A(_148_),
    .B(_149_));
 sg13g2_o21ai_1 _514_ (.B1(_150_),
    .Y(_151_),
    .A1(_007_),
    .A2(_058_));
 sg13g2_a21o_1 _515_ (.A2(_146_),
    .A1(_101_),
    .B1(_100_),
    .X(_152_));
 sg13g2_and3_1 _516_ (.X(_153_),
    .A(_147_),
    .B(_151_),
    .C(_152_));
 sg13g2_nand3_1 _517_ (.B(_151_),
    .C(_152_),
    .A(_147_),
    .Y(_154_));
 sg13g2_a21oi_1 _518_ (.A1(_133_),
    .A2(_145_),
    .Y(_155_),
    .B1(_144_));
 sg13g2_nand3_1 _519_ (.B(net76),
    .C(_103_),
    .A(net66),
    .Y(_156_));
 sg13g2_o21ai_1 _520_ (.B1(_141_),
    .Y(_157_),
    .A1(_139_),
    .A2(_142_));
 sg13g2_nand2b_1 _521_ (.Y(_158_),
    .B(_157_),
    .A_N(_156_));
 sg13g2_xnor2_1 _522_ (.Y(_159_),
    .A(_156_),
    .B(_157_));
 sg13g2_nand2b_1 _523_ (.Y(_160_),
    .B(_159_),
    .A_N(_155_));
 sg13g2_xnor2_1 _524_ (.Y(_161_),
    .A(_155_),
    .B(_159_));
 sg13g2_xor2_1 _525_ (.B(_015_),
    .A(_014_),
    .X(_162_));
 sg13g2_xor2_1 _526_ (.B(_066_),
    .A(_065_),
    .X(_163_));
 sg13g2_xor2_1 _527_ (.B(_163_),
    .A(_162_),
    .X(_164_));
 sg13g2_nand2_1 _528_ (.Y(_165_),
    .A(_161_),
    .B(_164_));
 sg13g2_xnor2_1 _529_ (.Y(_166_),
    .A(_161_),
    .B(_164_));
 sg13g2_a21oi_1 _530_ (.A1(_147_),
    .A2(_151_),
    .Y(_167_),
    .B1(_152_));
 sg13g2_nor2_1 _531_ (.A(_153_),
    .B(_167_),
    .Y(_168_));
 sg13g2_o21ai_1 _532_ (.B1(_154_),
    .Y(_169_),
    .A1(_166_),
    .A2(_167_));
 sg13g2_o21ai_1 _533_ (.B1(_165_),
    .Y(_170_),
    .A1(_162_),
    .A2(_163_));
 sg13g2_nand2_1 _534_ (.Y(_171_),
    .A(_169_),
    .B(_170_));
 sg13g2_xnor2_1 _535_ (.Y(_172_),
    .A(_169_),
    .B(_170_));
 sg13g2_nand3_1 _536_ (.B(_158_),
    .C(_160_),
    .A(_136_),
    .Y(_173_));
 sg13g2_xor2_1 _537_ (.B(_018_),
    .A(_017_),
    .X(_174_));
 sg13g2_xor2_1 _538_ (.B(_069_),
    .A(_068_),
    .X(_175_));
 sg13g2_and2_1 _539_ (.A(_174_),
    .B(_175_),
    .X(_176_));
 sg13g2_xor2_1 _540_ (.B(_175_),
    .A(_174_),
    .X(_177_));
 sg13g2_xnor2_1 _541_ (.Y(_178_),
    .A(_173_),
    .B(_177_));
 sg13g2_o21ai_1 _542_ (.B1(_171_),
    .Y(_179_),
    .A1(_172_),
    .A2(_178_));
 sg13g2_a21o_1 _543_ (.A2(_177_),
    .A1(_173_),
    .B1(_176_),
    .X(_180_));
 sg13g2_nand3_1 _544_ (.B(_179_),
    .C(_180_),
    .A(_097_),
    .Y(_181_));
 sg13g2_nor2_1 _545_ (.A(_094_),
    .B(_181_),
    .Y(_182_));
 sg13g2_xnor2_1 _546_ (.Y(_183_),
    .A(_091_),
    .B(_182_));
 sg13g2_xnor2_1 _547_ (.Y(_184_),
    .A(_089_),
    .B(_090_));
 sg13g2_xnor2_1 _548_ (.Y(_185_),
    .A(_092_),
    .B(_093_));
 sg13g2_inv_1 _549_ (.Y(_186_),
    .A(_185_));
 sg13g2_xnor2_1 _550_ (.Y(_187_),
    .A(_095_),
    .B(_096_));
 sg13g2_xnor2_1 _551_ (.Y(_188_),
    .A(_179_),
    .B(_180_));
 sg13g2_a21oi_1 _552_ (.A1(_179_),
    .A2(_180_),
    .Y(_189_),
    .B1(_097_));
 sg13g2_o21ai_1 _553_ (.B1(_189_),
    .Y(_190_),
    .A1(_187_),
    .A2(_188_));
 sg13g2_and3_1 _554_ (.X(_191_),
    .A(_181_),
    .B(_186_),
    .C(_190_));
 sg13g2_nand3_1 _555_ (.B(_186_),
    .C(_190_),
    .A(_181_),
    .Y(_192_));
 sg13g2_xnor2_1 _556_ (.Y(_193_),
    .A(_094_),
    .B(_181_));
 sg13g2_a21o_1 _557_ (.A2(_193_),
    .A1(_192_),
    .B1(_184_),
    .X(_194_));
 sg13g2_a21oi_1 _558_ (.A1(_183_),
    .A2(_194_),
    .Y(_195_),
    .B1(_087_));
 sg13g2_a221oi_1 _559_ (.B2(_182_),
    .C1(_195_),
    .B1(_091_),
    .A1(_035_),
    .Y(_196_),
    .A2(_085_));
 sg13g2_nand2b_1 _560_ (.Y(_197_),
    .B(_278_),
    .A_N(_196_));
 sg13g2_xnor2_1 _561_ (.Y(_198_),
    .A(_261_),
    .B(_262_));
 sg13g2_and3_1 _562_ (.X(_199_),
    .A(_087_),
    .B(_183_),
    .C(_194_));
 sg13g2_nor3_1 _563_ (.A(_195_),
    .B(_198_),
    .C(_199_),
    .Y(_200_));
 sg13g2_xnor2_1 _564_ (.Y(_201_),
    .A(_258_),
    .B(_259_));
 sg13g2_nand3_1 _565_ (.B(_192_),
    .C(_193_),
    .A(_184_),
    .Y(_202_));
 sg13g2_and3_1 _566_ (.X(_203_),
    .A(_194_),
    .B(_201_),
    .C(_202_));
 sg13g2_nand3_1 _567_ (.B(_201_),
    .C(_202_),
    .A(_194_),
    .Y(_204_));
 sg13g2_xnor2_1 _568_ (.Y(_205_),
    .A(_249_),
    .B(_250_));
 sg13g2_a21oi_1 _569_ (.A1(_181_),
    .A2(_190_),
    .Y(_206_),
    .B1(_186_));
 sg13g2_nor3_1 _570_ (.A(_191_),
    .B(_205_),
    .C(_206_),
    .Y(_207_));
 sg13g2_xor2_1 _571_ (.B(_188_),
    .A(_187_),
    .X(_208_));
 sg13g2_nand2b_1 _572_ (.Y(_209_),
    .B(_208_),
    .A_N(_251_));
 sg13g2_inv_1 _573_ (.Y(_210_),
    .A(_209_));
 sg13g2_o21ai_1 _574_ (.B1(_205_),
    .Y(_211_),
    .A1(_191_),
    .A2(_206_));
 sg13g2_nand2b_1 _575_ (.Y(_212_),
    .B(_211_),
    .A_N(_207_));
 sg13g2_a21oi_1 _576_ (.A1(_210_),
    .A2(_211_),
    .Y(_213_),
    .B1(_207_));
 sg13g2_a21oi_1 _577_ (.A1(_194_),
    .A2(_202_),
    .Y(_214_),
    .B1(_201_));
 sg13g2_nor2_1 _578_ (.A(_203_),
    .B(_214_),
    .Y(_215_));
 sg13g2_o21ai_1 _579_ (.B1(_204_),
    .Y(_216_),
    .A1(_213_),
    .A2(_214_));
 sg13g2_o21ai_1 _580_ (.B1(_198_),
    .Y(_217_),
    .A1(_195_),
    .A2(_199_));
 sg13g2_nand2b_1 _581_ (.Y(_218_),
    .B(_217_),
    .A_N(_200_));
 sg13g2_a21oi_1 _582_ (.A1(_216_),
    .A2(_217_),
    .Y(_219_),
    .B1(_200_));
 sg13g2_nor2b_1 _583_ (.A(_278_),
    .B_N(_196_),
    .Y(_220_));
 sg13g2_xnor2_1 _584_ (.Y(_221_),
    .A(_278_),
    .B(_196_));
 sg13g2_o21ai_1 _585_ (.B1(_197_),
    .Y(_222_),
    .A1(_219_),
    .A2(_220_));
 sg13g2_xor2_1 _586_ (.B(_271_),
    .A(_270_),
    .X(_223_));
 sg13g2_nand3_1 _587_ (.B(_222_),
    .C(_223_),
    .A(_277_),
    .Y(_224_));
 sg13g2_a21o_1 _588_ (.A2(_223_),
    .A1(_222_),
    .B1(_277_),
    .X(_225_));
 sg13g2_and2_1 _589_ (.A(_224_),
    .B(_225_),
    .X(\mul_uut.C2.ha_8.sum ));
 sg13g2_a21oi_1 _590_ (.A1(_272_),
    .A2(_276_),
    .Y(_226_),
    .B1(_231_));
 sg13g2_nand3_1 _591_ (.B(_224_),
    .C(_226_),
    .A(_275_),
    .Y(uio_out[7]));
 sg13g2_xnor2_1 _592_ (.Y(\mul_uut.C2.fa_4.sum ),
    .A(_213_),
    .B(_215_));
 sg13g2_xnor2_1 _593_ (.Y(\mul_uut.C2.fa_5.sum ),
    .A(_216_),
    .B(_218_));
 sg13g2_xnor2_1 _594_ (.Y(\mul_uut.C2.fa_6.sum ),
    .A(_219_),
    .B(_221_));
 sg13g2_xor2_1 _595_ (.B(_223_),
    .A(_222_),
    .X(\mul_uut.C2.fa_7.sum ));
 sg13g2_xor2_1 _596_ (.B(_151_),
    .A(_147_),
    .X(\mul_uut.C1.ha_5.sum ));
 sg13g2_xor2_1 _597_ (.B(_149_),
    .A(_148_),
    .X(\mul_uut.C1.fa_1.sum ));
 sg13g2_xnor2_1 _598_ (.Y(\mul_uut.C1.fa_5.sum ),
    .A(_166_),
    .B(_168_));
 sg13g2_xor2_1 _599_ (.B(_178_),
    .A(_172_),
    .X(\mul_uut.C1.fa_6.sum ));
 sg13g2_a22oi_1 _600_ (.Y(_228_),
    .B1(net80),
    .B2(net68),
    .A2(net78),
    .A1(net70));
 sg13g2_nor2_1 _601_ (.A(_111_),
    .B(_228_),
    .Y(uo_out[1]));
 sg13g2_xnor2_1 _602_ (.Y(\mul_uut.N1.C1.fa_1.sum ),
    .A(_107_),
    .B(_108_));
 sg13g2_xor2_1 _603_ (.B(_121_),
    .A(_110_),
    .X(\mul_uut.N1.C1.ha_3.sum ));
 sg13g2_xnor2_1 _604_ (.Y(\mul_uut.C2.ha_1.sum ),
    .A(_251_),
    .B(_208_));
 sg13g2_xnor2_1 _605_ (.Y(\mul_uut.C2.ha_6.sum ),
    .A(_210_),
    .B(_212_));
 sg13g2_tielo tt_um_multiplier_tt10_14 (.L_LO(net14));
 sg13g2_tielo tt_um_multiplier_tt10_15 (.L_LO(net15));
 sg13g2_tielo tt_um_multiplier_tt10_16 (.L_LO(net16));
 sg13g2_tielo tt_um_multiplier_tt10_17 (.L_LO(net17));
 sg13g2_tielo tt_um_multiplier_tt10_18 (.L_LO(net18));
 sg13g2_tielo tt_um_multiplier_tt10_19 (.L_LO(net19));
 sg13g2_tielo tt_um_multiplier_tt10_20 (.L_LO(net20));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _614_ (.A(\mul_uut.C2.ha_1.sum ),
    .X(uio_out[0]));
 sg13g2_buf_1 _615_ (.A(\mul_uut.C2.ha_6.sum ),
    .X(uio_out[1]));
 sg13g2_buf_1 _616_ (.A(\mul_uut.C2.fa_4.sum ),
    .X(uio_out[2]));
 sg13g2_buf_1 _617_ (.A(\mul_uut.C2.fa_5.sum ),
    .X(uio_out[3]));
 sg13g2_buf_1 _618_ (.A(\mul_uut.C2.fa_6.sum ),
    .X(uio_out[4]));
 sg13g2_buf_1 _619_ (.A(\mul_uut.C2.fa_7.sum ),
    .X(uio_out[5]));
 sg13g2_buf_1 _620_ (.A(\mul_uut.C2.ha_8.sum ),
    .X(uio_out[6]));
 sg13g2_buf_1 _621_ (.A(\mul_uut.N1.C1.fa_1.sum ),
    .X(uo_out[2]));
 sg13g2_buf_1 _622_ (.A(\mul_uut.N1.C1.ha_3.sum ),
    .X(uo_out[3]));
 sg13g2_buf_1 _623_ (.A(\mul_uut.C1.fa_1.sum ),
    .X(uo_out[4]));
 sg13g2_buf_1 _624_ (.A(\mul_uut.C1.ha_5.sum ),
    .X(uo_out[5]));
 sg13g2_buf_1 _625_ (.A(\mul_uut.C1.fa_5.sum ),
    .X(uo_out[6]));
 sg13g2_buf_1 _626_ (.A(\mul_uut.C1.fa_6.sum ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout61 (.A(net12),
    .X(net61));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(net11));
 sg13g2_buf_2 fanout63 (.A(uio_in[5]),
    .X(net63));
 sg13g2_buf_1 fanout64 (.A(uio_in[5]),
    .X(net64));
 sg13g2_buf_4 fanout65 (.X(net65),
    .A(net10));
 sg13g2_buf_2 fanout66 (.A(net9),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(net8),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(uio_in[1]),
    .X(net68));
 sg13g2_buf_1 fanout69 (.A(uio_in[1]),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(net7),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(net6),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(net5),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(ui_in[5]),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(ui_in[5]),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(net4),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net3),
    .X(net76));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(net2));
 sg13g2_buf_2 fanout78 (.A(ui_in[1]),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(ui_in[1]),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(net1),
    .X(net80));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[6]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[7]),
    .X(net12));
 sg13g2_tielo tt_um_multiplier_tt10_13 (.L_LO(net13));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_decap_8 FILLER_25_176 ();
 sg13g2_decap_8 FILLER_25_183 ();
 sg13g2_decap_8 FILLER_25_190 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_decap_8 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_decap_8 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_decap_8 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_303 ();
 sg13g2_decap_8 FILLER_25_310 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_decap_4 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_241 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_fill_2 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_fill_1 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_4 FILLER_27_154 ();
 sg13g2_decap_4 FILLER_27_170 ();
 sg13g2_fill_2 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_decap_4 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_242 ();
 sg13g2_decap_4 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_decap_4 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_195 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_decap_4 FILLER_28_240 ();
 sg13g2_fill_1 FILLER_28_244 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_265 ();
 sg13g2_decap_8 FILLER_28_270 ();
 sg13g2_decap_4 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_8 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_153 ();
 sg13g2_decap_4 FILLER_29_172 ();
 sg13g2_decap_4 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_243 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_306 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_352 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_decap_8 FILLER_29_366 ();
 sg13g2_decap_8 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_decap_4 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_decap_4 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_253 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_decap_8 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_decap_8 FILLER_31_144 ();
 sg13g2_decap_8 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_fill_2 FILLER_31_175 ();
 sg13g2_decap_4 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_217 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_decap_4 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_340 ();
 sg13g2_decap_8 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_354 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_decap_8 FILLER_31_368 ();
 sg13g2_decap_8 FILLER_31_375 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_31_389 ();
 sg13g2_decap_8 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_145 ();
 sg13g2_decap_4 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_198 ();
 sg13g2_decap_4 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_decap_8 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_decap_4 FILLER_32_299 ();
 sg13g2_decap_4 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_121 ();
 sg13g2_decap_4 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_decap_8 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_decap_4 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_decap_4 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_4 FILLER_34_126 ();
 sg13g2_decap_4 FILLER_34_138 ();
 sg13g2_fill_2 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_fill_2 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_decap_4 FILLER_34_184 ();
 sg13g2_decap_8 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_228 ();
 sg13g2_decap_4 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_264 ();
 sg13g2_decap_4 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_decap_4 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_decap_4 FILLER_34_320 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_decap_4 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_decap_8 FILLER_34_352 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_4 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_decap_8 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_decap_4 FILLER_35_175 ();
 sg13g2_fill_2 FILLER_35_179 ();
 sg13g2_decap_8 FILLER_35_187 ();
 sg13g2_fill_1 FILLER_35_205 ();
 sg13g2_decap_8 FILLER_35_239 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_257 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_321 ();
 sg13g2_decap_4 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_decap_4 FILLER_36_153 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_decap_4 FILLER_36_190 ();
 sg13g2_fill_1 FILLER_36_194 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_fill_2 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_decap_4 FILLER_36_258 ();
 sg13g2_fill_2 FILLER_36_267 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_4 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_157 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_187 ();
 sg13g2_fill_1 FILLER_37_206 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_decap_4 FILLER_37_241 ();
 sg13g2_fill_1 FILLER_37_245 ();
 sg13g2_fill_1 FILLER_37_252 ();
 sg13g2_fill_2 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_decap_8 FILLER_38_130 ();
 sg13g2_decap_4 FILLER_38_137 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_161 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_231 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
endmodule

module tt_um_htfab_caterpillar (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire \btn.button_state[0] ;
 wire \btn.button_state[1] ;
 wire \btn.button_state[2] ;
 wire \btn.button_state[3] ;
 wire \btn.change_timer[0] ;
 wire \btn.change_timer[1] ;
 wire \btn.change_timer[2] ;
 wire \btn.change_timer[3] ;
 wire \btn.change_timer[4] ;
 wire \btn.change_timer[5] ;
 wire \btn.change_timer[6] ;
 wire \btn.current_event[0] ;
 wire \btn.current_event[1] ;
 wire \btn.current_event[2] ;
 wire \btn.current_event[3] ;
 wire \btn.gate_200hz ;
 wire \btn.input_event[0] ;
 wire \btn.input_event[1] ;
 wire \btn.input_event[2] ;
 wire \btn.input_event[3] ;
 wire \btn.input_event[4] ;
 wire \btn.long_press ;
 wire \btn.sample_10ms[0] ;
 wire \btn.sample_10ms[1] ;
 wire \btn.sample_10ms[2] ;
 wire \btn.sample_10ms[3] ;
 wire \btn.sample_15ms[0] ;
 wire \btn.sample_15ms[1] ;
 wire \btn.sample_15ms[2] ;
 wire \btn.sample_15ms[3] ;
 wire \btn.sample_5ms[0] ;
 wire \btn.sample_5ms[1] ;
 wire \btn.sample_5ms[2] ;
 wire \btn.sample_5ms[3] ;
 wire \clk_div_counter[0] ;
 wire \clk_div_counter[1] ;
 wire \clk_div_counter[2] ;
 wire \clk_div_counter[3] ;
 wire \clk_div_counter[4] ;
 wire \clk_div_counter[5] ;
 wire \clk_div_counter[6] ;
 wire \clk_div_counter[7] ;
 wire display_graphical;
 wire \display_value[0] ;
 wire \display_value[1] ;
 wire \display_value[2] ;
 wire \display_value[3] ;
 wire \display_value[4] ;
 wire \dsp.digit ;
 wire \dsp.digit_sel_raw[1] ;
 wire \dsp.segments_raw[0] ;
 wire \dsp.segments_raw[1] ;
 wire \dsp.segments_raw[2] ;
 wire \dsp.segments_raw[3] ;
 wire \dsp.segments_raw[4] ;
 wire \dsp.segments_raw[5] ;
 wire \dsp.segments_raw[6] ;
 wire \game.challenge_mode ;
 wire \game.challenge_num[0] ;
 wire \game.challenge_num[1] ;
 wire \game.challenge_num[2] ;
 wire \game.challenge_num[3] ;
 wire \game.counter[0] ;
 wire \game.counter[1] ;
 wire \game.counter[2] ;
 wire \game.counter[3] ;
 wire \game.counter[4] ;
 wire \game.counter[5] ;
 wire \game.counter[6] ;
 wire \game.counter[7] ;
 wire \game.current_level[0] ;
 wire \game.current_level[1] ;
 wire \game.current_level[2] ;
 wire \game.current_level[3] ;
 wire \game.current_level[4] ;
 wire \game.fsm.block_len[0][0] ;
 wire \game.fsm.block_len[0][1] ;
 wire \game.fsm.block_len[0][2] ;
 wire \game.fsm.block_len[1][0] ;
 wire \game.fsm.block_len[1][1] ;
 wire \game.fsm.block_len[1][2] ;
 wire \game.fsm.block_len[2][0] ;
 wire \game.fsm.block_len[2][1] ;
 wire \game.fsm.block_len[2][2] ;
 wire \game.fsm.block_len[3][0] ;
 wire \game.fsm.block_len[3][1] ;
 wire \game.fsm.block_len[3][2] ;
 wire \game.fsm.block_len[4][0] ;
 wire \game.fsm.block_len[4][1] ;
 wire \game.fsm.block_len[4][2] ;
 wire \game.fsm.block_len[5][0] ;
 wire \game.fsm.block_len[5][1] ;
 wire \game.fsm.block_len[5][2] ;
 wire \game.fsm.block_len[6][0] ;
 wire \game.fsm.block_len[6][1] ;
 wire \game.fsm.block_len[6][2] ;
 wire \game.fsm.block_len[7][0] ;
 wire \game.fsm.block_len[7][1] ;
 wire \game.fsm.block_len[7][2] ;
 wire \game.fsm.color_count[0][0] ;
 wire \game.fsm.color_count[0][1] ;
 wire \game.fsm.color_count[0][2] ;
 wire \game.fsm.color_count[1][0] ;
 wire \game.fsm.color_count[1][1] ;
 wire \game.fsm.color_count[1][2] ;
 wire \game.fsm.color_count[2][0] ;
 wire \game.fsm.color_count[2][1] ;
 wire \game.fsm.color_count[2][2] ;
 wire \game.fsm.color_count[3][0] ;
 wire \game.fsm.color_count[3][1] ;
 wire \game.fsm.color_count[3][2] ;
 wire \game.fsm.green_block_count[0] ;
 wire \game.fsm.green_block_count[1] ;
 wire \game.fsm.green_block_count[2] ;
 wire \game.fsm.len1_block_count[0] ;
 wire \game.fsm.len1_block_count[1] ;
 wire \game.fsm.len1_block_count[2] ;
 wire \game.fsm.len1_color_count[0][0] ;
 wire \game.fsm.len1_color_count[0][1] ;
 wire \game.fsm.len1_color_count[0][2] ;
 wire \game.fsm.len1_color_count[1][0] ;
 wire \game.fsm.len1_color_count[1][1] ;
 wire \game.fsm.len1_color_count[1][2] ;
 wire \game.fsm.len1_color_count[2][0] ;
 wire \game.fsm.len1_color_count[2][1] ;
 wire \game.fsm.len1_color_count[2][2] ;
 wire \game.fsm.len1_color_count[3][0] ;
 wire \game.fsm.len1_color_count[3][1] ;
 wire \game.fsm.len1_color_count[3][2] ;
 wire \game.fsm.len2_block_count[0] ;
 wire \game.fsm.len2_block_count[1] ;
 wire \game.fsm.len2_color_count[0][0] ;
 wire \game.fsm.len2_color_count[0][1] ;
 wire \game.fsm.len2_color_count[1][0] ;
 wire \game.fsm.len2_color_count[1][1] ;
 wire \game.fsm.len2_color_count[2][0] ;
 wire \game.fsm.len2_color_count[2][1] ;
 wire \game.fsm.len2_color_count[3][0] ;
 wire \game.fsm.len2_color_count[3][1] ;
 wire \game.fsm.len3_block_count[0] ;
 wire \game.fsm.len3_block_count[1] ;
 wire \game.fsm.len3_color_count[0][0] ;
 wire \game.fsm.len3_color_count[0][1] ;
 wire \game.fsm.len3_color_count[1][0] ;
 wire \game.fsm.len3_color_count[1][1] ;
 wire \game.fsm.len3_color_count[2][0] ;
 wire \game.fsm.len3_color_count[2][1] ;
 wire \game.fsm.len3_color_count[3][0] ;
 wire \game.fsm.len3_color_count[3][1] ;
 wire \game.fsm.length[0] ;
 wire \game.fsm.length[1] ;
 wire \game.fsm.length[2] ;
 wire \game.fsm.num_blocks[0] ;
 wire \game.fsm.num_blocks[1] ;
 wire \game.fsm.num_blocks[2] ;
 wire \game.fsm.read_pos[0] ;
 wire \game.fsm.read_pos[1] ;
 wire \game.fsm.read_pos[2] ;
 wire \game.fsm.seq[0][0] ;
 wire \game.fsm.seq[0][1] ;
 wire \game.fsm.seq[1][0] ;
 wire \game.fsm.seq[1][1] ;
 wire \game.fsm.seq[2][0] ;
 wire \game.fsm.seq[2][1] ;
 wire \game.fsm.seq[3][0] ;
 wire \game.fsm.seq[3][1] ;
 wire \game.fsm.seq[4][0] ;
 wire \game.fsm.seq[4][1] ;
 wire \game.fsm.seq[5][0] ;
 wire \game.fsm.seq[5][1] ;
 wire \game.fsm.seq[6][0] ;
 wire \game.fsm.seq[6][1] ;
 wire \game.fsm.seq[7][0] ;
 wire \game.fsm.seq[7][1] ;
 wire \game.input_color[0] ;
 wire \game.input_color[1] ;
 wire \game.input_erase ;
 wire \game.input_reset ;
 wire \game.input_update ;
 wire \game.next_state[0] ;
 wire \game.next_state[2] ;
 wire \game.slv.fsm_color[0] ;
 wire \game.slv.fsm_color[1] ;
 wire \game.slv.fsm_reset ;
 wire \game.slv.fsm_update ;
 wire \game.slv.length[0] ;
 wire \game.slv.length[1] ;
 wire \game.slv.length[2] ;
 wire \game.slv.lfsr[0] ;
 wire \game.slv.lfsr[10] ;
 wire \game.slv.lfsr[11] ;
 wire \game.slv.lfsr[12] ;
 wire \game.slv.lfsr[13] ;
 wire \game.slv.lfsr[14] ;
 wire \game.slv.lfsr[15] ;
 wire \game.slv.lfsr[16] ;
 wire \game.slv.lfsr[17] ;
 wire \game.slv.lfsr[18] ;
 wire \game.slv.lfsr[19] ;
 wire \game.slv.lfsr[1] ;
 wire \game.slv.lfsr[20] ;
 wire \game.slv.lfsr[2] ;
 wire \game.slv.lfsr[3] ;
 wire \game.slv.lfsr[4] ;
 wire \game.slv.lfsr[5] ;
 wire \game.slv.lfsr[6] ;
 wire \game.slv.lfsr[7] ;
 wire \game.slv.lfsr[8] ;
 wire \game.slv.lfsr[9] ;
 wire \game.slv.pos[0] ;
 wire \game.slv.pos[1] ;
 wire \game.slv.pos[2] ;
 wire \game.slv.ready ;
 wire \game.slv.retries[0] ;
 wire \game.slv.retries[1] ;
 wire \game.slv.retries[2] ;
 wire \game.slv.saved_target ;
 wire \game.slv.state[1] ;
 wire \game.slv.state[2] ;
 wire \game.slv.state[3] ;
 wire \game.slv.target[0] ;
 wire \game.slv.target[1] ;
 wire \game.slv.trigger ;
 wire \game.solver_active ;
 wire \game.solver_trigger_delayed ;
 wire \game.sound_mode[0] ;
 wire \game.sound_mode[1] ;
 wire \game.sound_mode[2] ;
 wire \game.sound_on ;
 wire \game.state[0] ;
 wire \game.state[1] ;
 wire \game.state[2] ;
 wire \game.state[3] ;
 wire \game.tune[0] ;
 wire \game.tune[1] ;
 wire \snd.active_tune[0] ;
 wire \snd.active_tune[1] ;
 wire \snd.chord[0][0] ;
 wire \snd.chord[0][1] ;
 wire \snd.chord[0][2] ;
 wire \snd.chord[0][3] ;
 wire \snd.chord[0][4] ;
 wire \snd.chord[0][5] ;
 wire \snd.chord[1][0] ;
 wire \snd.chord[1][5] ;
 wire \snd.chord[2][2] ;
 wire \snd.chord[3][0] ;
 wire \snd.counter[0] ;
 wire \snd.counter[1] ;
 wire \snd.counter[2] ;
 wire \snd.counter[3] ;
 wire \snd.counter[4] ;
 wire \snd.counter[5] ;
 wire \snd.counter[6] ;
 wire \snd.counter[7] ;
 wire \snd.counter[8] ;
 wire \snd.next_note_sel[0] ;
 wire \snd.next_note_sel[1] ;
 wire \snd.next_note_timing[0] ;
 wire \snd.next_note_timing[1] ;
 wire \snd.next_note_timing[2] ;
 wire \snd.next_note_timing[3] ;
 wire \snd.next_note_timing[4] ;
 wire \snd.next_note_timing[5] ;
 wire \snd.next_note_timing[6] ;
 wire \snd.next_note_timing[7] ;
 wire \snd.next_note_timing[8] ;
 wire \snd.note_sel[0] ;
 wire \snd.note_sel[1] ;
 wire \snd.note_timing[0] ;
 wire \snd.note_timing[1] ;
 wire \snd.note_timing[2] ;
 wire \snd.note_timing[3] ;
 wire \snd.note_timing[4] ;
 wire \snd.note_timing[5] ;
 wire \snd.note_timing[6] ;
 wire \snd.note_timing[7] ;
 wire \snd.note_timing[8] ;
 wire \snd.sequencer_state[0] ;
 wire \snd.sequencer_state[1] ;
 wire \snd.sound ;
 wire \snd.tune_counter[0] ;
 wire \snd.tune_counter[1] ;
 wire \snd.tune_counter[2] ;
 wire \snd.tune_counter[3] ;
 wire \snd.tune_counter[4] ;
 wire \snd.tune_counter[5] ;
 wire \snd.tune_counter[6] ;
 wire \snd.tune_pos[0] ;
 wire \snd.tune_pos[1] ;
 wire \snd.tune_pos[2] ;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire clknet_leaf_0_clk;
 wire net7;
 wire net8;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;

 sg13g2_inv_1 _2613_ (.Y(_1776_),
    .A(net701));
 sg13g2_inv_1 _2614_ (.Y(_1777_),
    .A(\snd.active_tune[1] ));
 sg13g2_inv_1 _2615_ (.Y(_1778_),
    .A(\snd.chord[0][5] ));
 sg13g2_inv_1 _2616_ (.Y(_1779_),
    .A(\snd.chord[1][5] ));
 sg13g2_inv_1 _2617_ (.Y(_1780_),
    .A(\snd.chord[2][2] ));
 sg13g2_inv_1 _2618_ (.Y(_1781_),
    .A(net408));
 sg13g2_inv_1 _2619_ (.Y(_1782_),
    .A(net476));
 sg13g2_inv_1 _2620_ (.Y(_1783_),
    .A(net712));
 sg13g2_inv_1 _2621_ (.Y(_1784_),
    .A(net557));
 sg13g2_inv_1 _2622_ (.Y(_1785_),
    .A(net497));
 sg13g2_inv_1 _2623_ (.Y(_1786_),
    .A(net473));
 sg13g2_inv_1 _2624_ (.Y(_1787_),
    .A(net500));
 sg13g2_inv_1 _2625_ (.Y(_1788_),
    .A(net520));
 sg13g2_inv_1 _2626_ (.Y(_1789_),
    .A(net542));
 sg13g2_inv_1 _2627_ (.Y(_1790_),
    .A(net490));
 sg13g2_inv_1 _2628_ (.Y(_1791_),
    .A(net638));
 sg13g2_inv_1 _2629_ (.Y(_1792_),
    .A(net441));
 sg13g2_inv_1 _2630_ (.Y(_1793_),
    .A(net332));
 sg13g2_inv_1 _2631_ (.Y(_1794_),
    .A(net457));
 sg13g2_inv_1 _2632_ (.Y(_1795_),
    .A(net454));
 sg13g2_inv_1 _2633_ (.Y(_1796_),
    .A(net452));
 sg13g2_inv_1 _2634_ (.Y(_1797_),
    .A(net665));
 sg13g2_inv_1 _2635_ (.Y(_1798_),
    .A(net469));
 sg13g2_inv_1 _2636_ (.Y(_1799_),
    .A(net479));
 sg13g2_inv_1 _2637_ (.Y(_1800_),
    .A(\game.counter[7] ));
 sg13g2_inv_1 _2638_ (.Y(_1801_),
    .A(\game.counter[4] ));
 sg13g2_inv_2 _2639_ (.Y(_1802_),
    .A(net782));
 sg13g2_inv_2 _2640_ (.Y(_1803_),
    .A(\game.state[2] ));
 sg13g2_inv_1 _2641_ (.Y(_1804_),
    .A(net381));
 sg13g2_inv_1 _2642_ (.Y(_1805_),
    .A(net710));
 sg13g2_inv_1 _2643_ (.Y(_1806_),
    .A(\display_value[2] ));
 sg13g2_inv_1 _2644_ (.Y(_1807_),
    .A(\game.sound_mode[2] ));
 sg13g2_inv_1 _2645_ (.Y(_1808_),
    .A(net678));
 sg13g2_inv_1 _2646_ (.Y(_1809_),
    .A(\game.current_level[4] ));
 sg13g2_inv_1 _2647_ (.Y(_1810_),
    .A(\game.current_level[3] ));
 sg13g2_inv_1 _2648_ (.Y(_1811_),
    .A(net463));
 sg13g2_inv_1 _2649_ (.Y(_1812_),
    .A(\game.challenge_num[3] ));
 sg13g2_inv_1 _2650_ (.Y(_1813_),
    .A(net496));
 sg13g2_inv_1 _2651_ (.Y(_1814_),
    .A(\game.fsm.green_block_count[1] ));
 sg13g2_inv_1 _2652_ (.Y(_1815_),
    .A(net442));
 sg13g2_inv_1 _2653_ (.Y(_1816_),
    .A(net328));
 sg13g2_inv_1 _2654_ (.Y(_1817_),
    .A(net326));
 sg13g2_inv_2 _2655_ (.Y(_1818_),
    .A(\game.fsm.num_blocks[2] ));
 sg13g2_inv_2 _2656_ (.Y(_1819_),
    .A(\game.fsm.num_blocks[1] ));
 sg13g2_inv_4 _2657_ (.A(\game.fsm.length[2] ),
    .Y(_1820_));
 sg13g2_inv_1 _2658_ (.Y(_1821_),
    .A(net397));
 sg13g2_inv_2 _2659_ (.Y(_1822_),
    .A(net401));
 sg13g2_inv_1 _2660_ (.Y(_1823_),
    .A(net743));
 sg13g2_inv_1 _2661_ (.Y(_1824_),
    .A(net661));
 sg13g2_inv_1 _2662_ (.Y(_1825_),
    .A(net735));
 sg13g2_inv_1 _2663_ (.Y(_1826_),
    .A(net656));
 sg13g2_inv_1 _2664_ (.Y(_1827_),
    .A(net662));
 sg13g2_inv_1 _2665_ (.Y(_1828_),
    .A(\snd.chord[3][0] ));
 sg13g2_inv_1 _2666_ (.Y(_1829_),
    .A(net624));
 sg13g2_inv_1 _2667_ (.Y(_1830_),
    .A(net585));
 sg13g2_inv_1 _2668_ (.Y(_1831_),
    .A(net583));
 sg13g2_inv_1 _2669_ (.Y(_1832_),
    .A(net575));
 sg13g2_inv_1 _2670_ (.Y(_1833_),
    .A(net609));
 sg13g2_inv_1 _2671_ (.Y(_1834_),
    .A(net580));
 sg13g2_inv_1 _2672_ (.Y(_1835_),
    .A(net650));
 sg13g2_inv_1 _2673_ (.Y(_1836_),
    .A(net551));
 sg13g2_inv_1 _2674_ (.Y(_1837_),
    .A(\snd.note_timing[2] ));
 sg13g2_inv_1 _2675_ (.Y(_1838_),
    .A(net532));
 sg13g2_inv_1 _2676_ (.Y(_1839_),
    .A(net470));
 sg13g2_inv_1 _2677_ (.Y(_1840_),
    .A(\snd.note_sel[1] ));
 sg13g2_inv_1 _2678_ (.Y(_1841_),
    .A(net510));
 sg13g2_inv_1 _2679_ (.Y(_1842_),
    .A(\game.fsm.seq[4][0] ));
 sg13g2_inv_1 _2680_ (.Y(_1843_),
    .A(\game.fsm.block_len[1][0] ));
 sg13g2_inv_1 _2681_ (.Y(_1844_),
    .A(\game.fsm.block_len[3][0] ));
 sg13g2_inv_1 _2682_ (.Y(_1845_),
    .A(_0069_));
 sg13g2_inv_1 _2683_ (.Y(_1846_),
    .A(\game.fsm.block_len[5][0] ));
 sg13g2_inv_1 _2684_ (.Y(_1847_),
    .A(\game.fsm.block_len[4][0] ));
 sg13g2_inv_1 _2685_ (.Y(_1848_),
    .A(net503));
 sg13g2_inv_1 _2686_ (.Y(_1849_),
    .A(\game.fsm.block_len[1][1] ));
 sg13g2_inv_1 _2687_ (.Y(_1850_),
    .A(\game.fsm.block_len[3][1] ));
 sg13g2_inv_1 _2688_ (.Y(_1851_),
    .A(\game.fsm.block_len[2][1] ));
 sg13g2_inv_1 _2689_ (.Y(_1852_),
    .A(\game.fsm.block_len[1][2] ));
 sg13g2_inv_1 _2690_ (.Y(_1853_),
    .A(\game.fsm.block_len[3][2] ));
 sg13g2_inv_1 _2691_ (.Y(_1854_),
    .A(\game.fsm.block_len[2][2] ));
 sg13g2_inv_1 _2692_ (.Y(_1855_),
    .A(\game.fsm.block_len[5][2] ));
 sg13g2_inv_1 _2693_ (.Y(_1856_),
    .A(_0076_));
 sg13g2_inv_1 _2694_ (.Y(_1857_),
    .A(_0077_));
 sg13g2_inv_1 _2695_ (.Y(_1858_),
    .A(\game.input_erase ));
 sg13g2_inv_1 _2696_ (.Y(_1859_),
    .A(_0078_));
 sg13g2_inv_1 _2697_ (.Y(_1860_),
    .A(_0080_));
 sg13g2_inv_1 _2698_ (.Y(_1861_),
    .A(net753));
 sg13g2_inv_1 _2699_ (.Y(_1862_),
    .A(\game.fsm.color_count[1][1] ));
 sg13g2_inv_1 _2700_ (.Y(_1863_),
    .A(\game.fsm.color_count[1][0] ));
 sg13g2_inv_1 _2701_ (.Y(_1864_),
    .A(net410));
 sg13g2_inv_1 _2702_ (.Y(_1865_),
    .A(net795));
 sg13g2_inv_1 _2703_ (.Y(_1866_),
    .A(net723));
 sg13g2_inv_1 _2704_ (.Y(_1867_),
    .A(net786));
 sg13g2_inv_1 _2705_ (.Y(_1868_),
    .A(_0024_));
 sg13g2_inv_1 _2706_ (.Y(_1869_),
    .A(net731));
 sg13g2_inv_1 _2707_ (.Y(_1870_),
    .A(\game.fsm.color_count[2][1] ));
 sg13g2_inv_1 _2708_ (.Y(_1871_),
    .A(\game.fsm.color_count[2][0] ));
 sg13g2_inv_1 _2709_ (.Y(_1872_),
    .A(_0025_));
 sg13g2_inv_1 _2710_ (.Y(_1873_),
    .A(_0034_));
 sg13g2_inv_1 _2711_ (.Y(_1874_),
    .A(_0035_));
 sg13g2_inv_1 _2712_ (.Y(_1875_),
    .A(_0036_));
 sg13g2_inv_1 _2713_ (.Y(_1876_),
    .A(net601));
 sg13g2_inv_1 _2714_ (.Y(_1877_),
    .A(_0038_));
 sg13g2_inv_1 _2715_ (.Y(_1878_),
    .A(_0083_));
 sg13g2_inv_1 _2716_ (.Y(_1879_),
    .A(net403));
 sg13g2_inv_2 _2717_ (.Y(_1880_),
    .A(net424));
 sg13g2_inv_2 _2718_ (.Y(_1881_),
    .A(\btn.input_event[0] ));
 sg13g2_inv_2 _2719_ (.Y(_1882_),
    .A(\btn.input_event[2] ));
 sg13g2_inv_1 _2720_ (.Y(_1883_),
    .A(\game.slv.ready ));
 sg13g2_inv_1 _2721_ (.Y(_1884_),
    .A(\snd.counter[7] ));
 sg13g2_inv_1 _2722_ (.Y(_1885_),
    .A(\snd.counter[6] ));
 sg13g2_inv_1 _2723_ (.Y(_1886_),
    .A(\snd.counter[5] ));
 sg13g2_inv_1 _2724_ (.Y(_1887_),
    .A(\snd.counter[4] ));
 sg13g2_inv_1 _2725_ (.Y(_1888_),
    .A(\snd.counter[2] ));
 sg13g2_inv_1 _2726_ (.Y(_1889_),
    .A(\snd.counter[1] ));
 sg13g2_inv_1 _2727_ (.Y(_1890_),
    .A(_0053_));
 sg13g2_inv_1 _2728_ (.Y(_1891_),
    .A(\dsp.digit ));
 sg13g2_inv_1 _2729_ (.Y(_1892_),
    .A(net768));
 sg13g2_inv_1 _2730_ (.Y(_1893_),
    .A(net323));
 sg13g2_nand2_1 _2731_ (.Y(_1894_),
    .A(\game.slv.lfsr[1] ),
    .B(\game.slv.lfsr[0] ));
 sg13g2_nor2_1 _2732_ (.A(\game.slv.lfsr[1] ),
    .B(\game.slv.lfsr[0] ),
    .Y(_1895_));
 sg13g2_nor2_1 _2733_ (.A(\game.slv.lfsr[2] ),
    .B(_1895_),
    .Y(_1896_));
 sg13g2_a21oi_1 _2734_ (.A1(\game.slv.lfsr[2] ),
    .A2(_1894_),
    .Y(_1897_),
    .B1(_1896_));
 sg13g2_a21oi_1 _2735_ (.A1(net402),
    .A2(_1897_),
    .Y(_1898_),
    .B1(net720));
 sg13g2_nor2_1 _2736_ (.A(net412),
    .B(_1898_),
    .Y(_0012_));
 sg13g2_nor2_2 _2737_ (.A(net720),
    .B(net412),
    .Y(_1899_));
 sg13g2_nor2_1 _2738_ (.A(\game.fsm.len2_color_count[0][1] ),
    .B(\game.fsm.len2_color_count[0][0] ),
    .Y(_1900_));
 sg13g2_or2_1 _2739_ (.X(_1901_),
    .B(\game.fsm.len3_color_count[3][0] ),
    .A(\game.fsm.len3_color_count[3][1] ));
 sg13g2_nor2_2 _2740_ (.A(\game.fsm.len2_color_count[2][1] ),
    .B(\game.fsm.len2_color_count[2][0] ),
    .Y(_1902_));
 sg13g2_nor2_1 _2741_ (.A(\game.fsm.len3_color_count[2][1] ),
    .B(\game.fsm.len3_color_count[2][0] ),
    .Y(_1903_));
 sg13g2_nor2_1 _2742_ (.A(\game.fsm.len3_color_count[0][1] ),
    .B(\game.fsm.len3_color_count[0][0] ),
    .Y(_1904_));
 sg13g2_nor2_1 _2743_ (.A(\game.fsm.len3_color_count[1][1] ),
    .B(\game.fsm.len3_color_count[1][0] ),
    .Y(_1905_));
 sg13g2_nor2_1 _2744_ (.A(\game.fsm.len2_color_count[1][1] ),
    .B(\game.fsm.len2_color_count[1][0] ),
    .Y(_1906_));
 sg13g2_nor2_1 _2745_ (.A(\game.fsm.len2_color_count[3][1] ),
    .B(\game.fsm.len2_color_count[3][0] ),
    .Y(_1907_));
 sg13g2_xor2_1 _2746_ (.B(_1907_),
    .A(_1906_),
    .X(_1908_));
 sg13g2_nand2b_1 _2747_ (.Y(_1909_),
    .B(_1908_),
    .A_N(_1905_));
 sg13g2_xnor2_1 _2748_ (.Y(_1910_),
    .A(_1905_),
    .B(_1908_));
 sg13g2_and2_1 _2749_ (.A(\game.fsm.num_blocks[1] ),
    .B(net394),
    .X(_1911_));
 sg13g2_nor2_2 _2750_ (.A(\game.fsm.num_blocks[2] ),
    .B(net373),
    .Y(_1912_));
 sg13g2_or2_1 _2751_ (.X(_1913_),
    .B(net373),
    .A(\game.fsm.num_blocks[2] ));
 sg13g2_a21o_1 _2752_ (.A2(net373),
    .A1(_0069_),
    .B1(_1818_),
    .X(_1914_));
 sg13g2_a22oi_1 _2753_ (.Y(_1915_),
    .B1(_1853_),
    .B2(\game.fsm.block_len[2][2] ),
    .A2(\game.fsm.block_len[2][1] ),
    .A1(_1850_));
 sg13g2_nand2b_1 _2754_ (.Y(_1916_),
    .B(\game.fsm.block_len[3][1] ),
    .A_N(\game.fsm.block_len[2][1] ));
 sg13g2_o21ai_1 _2755_ (.B1(_1916_),
    .Y(_1917_),
    .A1(_1844_),
    .A2(\game.fsm.block_len[2][0] ));
 sg13g2_a22oi_1 _2756_ (.Y(_1918_),
    .B1(_1915_),
    .B2(_1917_),
    .A2(_1854_),
    .A1(\game.fsm.block_len[3][2] ));
 sg13g2_or2_2 _2757_ (.X(_1919_),
    .B(_1918_),
    .A(_1914_));
 sg13g2_mux2_1 _2758_ (.A0(_0074_),
    .A1(_0075_),
    .S(_1919_),
    .X(_1920_));
 sg13g2_nor2_1 _2759_ (.A(_1912_),
    .B(_1920_),
    .Y(_1921_));
 sg13g2_or2_1 _2760_ (.X(_1922_),
    .B(\game.fsm.num_blocks[1] ),
    .A(\game.fsm.num_blocks[2] ));
 sg13g2_a21oi_2 _2761_ (.B1(\game.fsm.block_len[0][2] ),
    .Y(_1923_),
    .A2(_1922_),
    .A1(\game.fsm.block_len[1][2] ));
 sg13g2_nor2b_1 _2762_ (.A(_1921_),
    .B_N(_1923_),
    .Y(_1924_));
 sg13g2_o21ai_1 _2763_ (.B1(_1923_),
    .Y(_1925_),
    .A1(_1912_),
    .A2(_1920_));
 sg13g2_nor2_1 _2764_ (.A(_1818_),
    .B(_1819_),
    .Y(_1926_));
 sg13g2_nor2_1 _2765_ (.A(_1855_),
    .B(\game.fsm.block_len[4][2] ),
    .Y(_1927_));
 sg13g2_nor2b_1 _2766_ (.A(\game.fsm.block_len[5][1] ),
    .B_N(\game.fsm.block_len[4][1] ),
    .Y(_1928_));
 sg13g2_nand2b_1 _2767_ (.Y(_1929_),
    .B(\game.fsm.block_len[5][0] ),
    .A_N(\game.fsm.block_len[4][0] ));
 sg13g2_nand2b_1 _2768_ (.Y(_1930_),
    .B(\game.fsm.block_len[5][1] ),
    .A_N(\game.fsm.block_len[4][1] ));
 sg13g2_a221oi_1 _2769_ (.B2(_1930_),
    .C1(_1928_),
    .B1(_1929_),
    .A1(_1855_),
    .Y(_1931_),
    .A2(\game.fsm.block_len[4][2] ));
 sg13g2_o21ai_1 _2770_ (.B1(_1926_),
    .Y(_1932_),
    .A1(_1927_),
    .A2(_1931_));
 sg13g2_mux2_1 _2771_ (.A0(_1856_),
    .A1(_1857_),
    .S(_1932_),
    .X(_1933_));
 sg13g2_mux2_1 _2772_ (.A0(_0027_),
    .A1(_0028_),
    .S(_1932_),
    .X(_1934_));
 sg13g2_nor2_1 _2773_ (.A(\game.fsm.block_len[6][1] ),
    .B(_1934_),
    .Y(_1935_));
 sg13g2_mux2_1 _2774_ (.A0(_1846_),
    .A1(_1847_),
    .S(_1932_),
    .X(_1936_));
 sg13g2_nor2_1 _2775_ (.A(_1830_),
    .B(_0026_),
    .Y(_1937_));
 sg13g2_nand2b_1 _2776_ (.Y(_1938_),
    .B(\game.fsm.block_len[6][0] ),
    .A_N(_0026_));
 sg13g2_xnor2_1 _2777_ (.Y(_1939_),
    .A(\game.fsm.block_len[6][2] ),
    .B(_1933_));
 sg13g2_a22oi_1 _2778_ (.Y(_1940_),
    .B1(_1936_),
    .B2(_1937_),
    .A2(_1934_),
    .A1(\game.fsm.block_len[6][1] ));
 sg13g2_o21ai_1 _2779_ (.B1(_1939_),
    .Y(_1941_),
    .A1(_1935_),
    .A2(_1940_));
 sg13g2_o21ai_1 _2780_ (.B1(_1926_),
    .Y(_1942_),
    .A1(net394),
    .A2(_0069_));
 sg13g2_nor2_1 _2781_ (.A(_0029_),
    .B(_1942_),
    .Y(_1943_));
 sg13g2_a21oi_2 _2782_ (.B1(_1933_),
    .Y(_1944_),
    .A2(_1943_),
    .A1(_1941_));
 sg13g2_nor2_2 _2783_ (.A(\game.fsm.num_blocks[1] ),
    .B(net395),
    .Y(_1945_));
 sg13g2_o21ai_1 _2784_ (.B1(\game.fsm.num_blocks[2] ),
    .Y(_1946_),
    .A1(\game.fsm.num_blocks[1] ),
    .A2(net394));
 sg13g2_o21ai_1 _2785_ (.B1(_1924_),
    .Y(_1947_),
    .A1(_1944_),
    .A2(_1946_));
 sg13g2_nor2_1 _2786_ (.A(\game.fsm.len1_color_count[3][1] ),
    .B(\game.fsm.len1_color_count[3][0] ),
    .Y(_1948_));
 sg13g2_nand2_1 _2787_ (.Y(_1949_),
    .A(_0037_),
    .B(_1948_));
 sg13g2_nor3_2 _2788_ (.A(\game.fsm.len1_color_count[0][1] ),
    .B(\game.fsm.len1_color_count[0][0] ),
    .C(_1874_),
    .Y(_1950_));
 sg13g2_nor3_1 _2789_ (.A(\game.fsm.len1_color_count[1][1] ),
    .B(\game.fsm.len1_color_count[1][0] ),
    .C(_1875_),
    .Y(_1951_));
 sg13g2_xor2_1 _2790_ (.B(_1951_),
    .A(_1950_),
    .X(_1952_));
 sg13g2_nand2_1 _2791_ (.Y(_1953_),
    .A(_1949_),
    .B(_1952_));
 sg13g2_xor2_1 _2792_ (.B(_1952_),
    .A(_1949_),
    .X(_1954_));
 sg13g2_and2_1 _2793_ (.A(_1947_),
    .B(_1954_),
    .X(_1955_));
 sg13g2_xor2_1 _2794_ (.B(_1954_),
    .A(_1947_),
    .X(_1956_));
 sg13g2_xnor2_1 _2795_ (.Y(_1957_),
    .A(_1910_),
    .B(_1956_));
 sg13g2_xor2_1 _2796_ (.B(_1957_),
    .A(_1904_),
    .X(_1958_));
 sg13g2_nand2b_1 _2797_ (.Y(_1959_),
    .B(_1958_),
    .A_N(_1903_));
 sg13g2_xnor2_1 _2798_ (.Y(_1960_),
    .A(_1903_),
    .B(_1958_));
 sg13g2_nor2b_1 _2799_ (.A(_1902_),
    .B_N(_1960_),
    .Y(_1961_));
 sg13g2_xnor2_1 _2800_ (.Y(_1962_),
    .A(_1902_),
    .B(_1960_));
 sg13g2_xor2_1 _2801_ (.B(_1962_),
    .A(_1901_),
    .X(_1963_));
 sg13g2_nand2b_1 _2802_ (.Y(_1964_),
    .B(_1963_),
    .A_N(_1900_));
 sg13g2_a21oi_1 _2803_ (.A1(_1901_),
    .A2(_1962_),
    .Y(_1965_),
    .B1(_1961_));
 sg13g2_o21ai_1 _2804_ (.B1(_1959_),
    .Y(_1966_),
    .A1(_1904_),
    .A2(_1957_));
 sg13g2_a21oi_1 _2805_ (.A1(_1910_),
    .A2(_1956_),
    .Y(_1967_),
    .B1(_1955_));
 sg13g2_o21ai_1 _2806_ (.B1(_1953_),
    .Y(_1968_),
    .A1(_1950_),
    .A2(_1951_));
 sg13g2_o21ai_1 _2807_ (.B1(_1909_),
    .Y(_1969_),
    .A1(_1906_),
    .A2(_1907_));
 sg13g2_xnor2_1 _2808_ (.Y(_1970_),
    .A(_1968_),
    .B(_1969_));
 sg13g2_xnor2_1 _2809_ (.Y(_1971_),
    .A(_1967_),
    .B(_1970_));
 sg13g2_xnor2_1 _2810_ (.Y(_1972_),
    .A(_1966_),
    .B(_1971_));
 sg13g2_xnor2_1 _2811_ (.Y(_1973_),
    .A(_1965_),
    .B(_1972_));
 sg13g2_xnor2_1 _2812_ (.Y(_1974_),
    .A(_1964_),
    .B(_1973_));
 sg13g2_nor3_1 _2813_ (.A(\game.fsm.len1_color_count[2][1] ),
    .B(\game.fsm.len1_color_count[2][0] ),
    .C(_1877_),
    .Y(_1975_));
 sg13g2_xor2_1 _2814_ (.B(_1963_),
    .A(_1900_),
    .X(_1976_));
 sg13g2_nand2_1 _2815_ (.Y(_1977_),
    .A(_1975_),
    .B(_1976_));
 sg13g2_o21ai_1 _2816_ (.B1(\game.current_level[0] ),
    .Y(_1978_),
    .A1(_1975_),
    .A2(_1976_));
 sg13g2_nand3b_1 _2817_ (.B(_1977_),
    .C(_1974_),
    .Y(_1979_),
    .A_N(_1978_));
 sg13g2_nor2b_2 _2818_ (.A(net391),
    .B_N(net392),
    .Y(_1980_));
 sg13g2_nand2b_1 _2819_ (.Y(_1981_),
    .B(\game.fsm.block_len[1][2] ),
    .A_N(\game.fsm.block_len[0][2] ));
 sg13g2_a22oi_1 _2820_ (.Y(_1982_),
    .B1(_1852_),
    .B2(\game.fsm.block_len[0][2] ),
    .A2(\game.fsm.block_len[0][1] ),
    .A1(_1849_));
 sg13g2_nand2b_1 _2821_ (.Y(_1983_),
    .B(\game.fsm.block_len[1][1] ),
    .A_N(\game.fsm.block_len[0][1] ));
 sg13g2_o21ai_1 _2822_ (.B1(_1983_),
    .Y(_1984_),
    .A1(_1843_),
    .A2(\game.fsm.block_len[0][0] ));
 sg13g2_nand2_1 _2823_ (.Y(_1985_),
    .A(_1982_),
    .B(_1984_));
 sg13g2_a22oi_1 _2824_ (.Y(_1986_),
    .B1(_1981_),
    .B2(_1985_),
    .A2(_1819_),
    .A1(_1818_));
 sg13g2_mux2_1 _2825_ (.A0(_0031_),
    .A1(_0030_),
    .S(_1986_),
    .X(_1987_));
 sg13g2_inv_1 _2826_ (.Y(_1988_),
    .A(_1987_));
 sg13g2_nand2b_1 _2827_ (.Y(_1989_),
    .B(_1919_),
    .A_N(_0033_));
 sg13g2_o21ai_1 _2828_ (.B1(_1989_),
    .Y(_1990_),
    .A1(_0032_),
    .A2(_1919_));
 sg13g2_nand2b_1 _2829_ (.Y(_1991_),
    .B(_1919_),
    .A_N(_0068_));
 sg13g2_o21ai_1 _2830_ (.B1(_1991_),
    .Y(_1992_),
    .A1(_0067_),
    .A2(_1919_));
 sg13g2_mux2_1 _2831_ (.A0(_0066_),
    .A1(_0065_),
    .S(_1986_),
    .X(_1993_));
 sg13g2_inv_1 _2832_ (.Y(_1994_),
    .A(_1993_));
 sg13g2_a22oi_1 _2833_ (.Y(_1995_),
    .B1(_1992_),
    .B2(_1993_),
    .A2(_1990_),
    .A1(_1987_));
 sg13g2_nor2_1 _2834_ (.A(_1987_),
    .B(_1990_),
    .Y(_1996_));
 sg13g2_a21oi_1 _2835_ (.A1(_1913_),
    .A2(_1923_),
    .Y(_1997_),
    .B1(_1921_));
 sg13g2_nor3_1 _2836_ (.A(_1995_),
    .B(_1996_),
    .C(_1997_),
    .Y(_1998_));
 sg13g2_a21oi_1 _2837_ (.A1(_1921_),
    .A2(_1923_),
    .Y(_1999_),
    .B1(_1998_));
 sg13g2_mux2_1 _2838_ (.A0(_1990_),
    .A1(_1988_),
    .S(_1999_),
    .X(_2000_));
 sg13g2_a21oi_1 _2839_ (.A1(_0029_),
    .A2(_1933_),
    .Y(_2001_),
    .B1(_1942_));
 sg13g2_nand2_1 _2840_ (.Y(_2002_),
    .A(_1941_),
    .B(_2001_));
 sg13g2_nand2_1 _2841_ (.Y(_2003_),
    .A(_1934_),
    .B(_2002_));
 sg13g2_o21ai_1 _2842_ (.B1(_2003_),
    .Y(_2004_),
    .A1(_1873_),
    .A2(_2002_));
 sg13g2_nand2b_1 _2843_ (.Y(_2005_),
    .B(_2002_),
    .A_N(_1936_));
 sg13g2_or2_1 _2844_ (.X(_2006_),
    .B(_2002_),
    .A(_0026_));
 sg13g2_mux2_1 _2845_ (.A0(_1992_),
    .A1(_1994_),
    .S(_1999_),
    .X(_2007_));
 sg13g2_a221oi_1 _2846_ (.B2(_2006_),
    .C1(_2007_),
    .B1(_2005_),
    .A1(_2000_),
    .Y(_2008_),
    .A2(_2004_));
 sg13g2_nand2b_1 _2847_ (.Y(_2009_),
    .B(_1924_),
    .A_N(_1944_));
 sg13g2_o21ai_1 _2848_ (.B1(_2009_),
    .Y(_2010_),
    .A1(_2000_),
    .A2(_2004_));
 sg13g2_a21oi_1 _2849_ (.A1(_1925_),
    .A2(_1944_),
    .Y(_2011_),
    .B1(_1946_));
 sg13g2_o21ai_1 _2850_ (.B1(_2011_),
    .Y(_2012_),
    .A1(_2008_),
    .A2(_2010_));
 sg13g2_nand2_1 _2851_ (.Y(_2013_),
    .A(_2000_),
    .B(_2012_));
 sg13g2_o21ai_1 _2852_ (.B1(_2013_),
    .Y(_2014_),
    .A1(_2004_),
    .A2(_2012_));
 sg13g2_nor2_1 _2853_ (.A(\game.fsm.len1_block_count[2] ),
    .B(\game.fsm.len1_block_count[1] ),
    .Y(_2015_));
 sg13g2_nand2_2 _2854_ (.Y(_2016_),
    .A(\game.fsm.len1_block_count[0] ),
    .B(_2015_));
 sg13g2_nor2b_1 _2855_ (.A(_2014_),
    .B_N(_2016_),
    .Y(_2017_));
 sg13g2_nand2b_1 _2856_ (.Y(_2018_),
    .B(\game.fsm.len3_block_count[0] ),
    .A_N(\game.fsm.len3_block_count[1] ));
 sg13g2_a21oi_1 _2857_ (.A1(_2005_),
    .A2(_2006_),
    .Y(_2019_),
    .B1(_2012_));
 sg13g2_a21oi_2 _2858_ (.B1(_2019_),
    .Y(_2020_),
    .A2(_2012_),
    .A1(_2007_));
 sg13g2_a21oi_1 _2859_ (.A1(_2014_),
    .A2(_2018_),
    .Y(_2021_),
    .B1(_2020_));
 sg13g2_nor2b_1 _2860_ (.A(_2017_),
    .B_N(_2021_),
    .Y(_2022_));
 sg13g2_nor2b_1 _2861_ (.A(\game.fsm.len2_block_count[1] ),
    .B_N(\game.fsm.len2_block_count[0] ),
    .Y(_2023_));
 sg13g2_nand2_1 _2862_ (.Y(_2024_),
    .A(_2014_),
    .B(_2020_));
 sg13g2_and3_1 _2863_ (.X(_2025_),
    .A(_2014_),
    .B(_2020_),
    .C(_2023_));
 sg13g2_nor4_1 _2864_ (.A(net391),
    .B(_1947_),
    .C(_2022_),
    .D(_2025_),
    .Y(_2026_));
 sg13g2_o21ai_1 _2865_ (.B1(_1979_),
    .Y(_2027_),
    .A1(_1980_),
    .A2(_2026_));
 sg13g2_nor2b_1 _2866_ (.A(\game.fsm.block_len[5][0] ),
    .B_N(\game.fsm.block_len[4][0] ),
    .Y(_2028_));
 sg13g2_a221oi_1 _2867_ (.B2(_2028_),
    .C1(_1928_),
    .B1(_1930_),
    .A1(_1855_),
    .Y(_2029_),
    .A2(\game.fsm.block_len[4][2] ));
 sg13g2_nor4_2 _2868_ (.A(_1818_),
    .B(_1819_),
    .C(_1927_),
    .Y(_2030_),
    .D(_2029_));
 sg13g2_mux2_1 _2869_ (.A0(_0071_),
    .A1(_0070_),
    .S(_2030_),
    .X(_2031_));
 sg13g2_nand2_1 _2870_ (.Y(_2032_),
    .A(_0076_),
    .B(_2030_));
 sg13g2_o21ai_1 _2871_ (.B1(_2032_),
    .Y(_2033_),
    .A1(_1857_),
    .A2(_2030_));
 sg13g2_nor2_1 _2872_ (.A(\game.fsm.block_len[6][2] ),
    .B(_2033_),
    .Y(_2034_));
 sg13g2_mux2_2 _2873_ (.A0(_0028_),
    .A1(_0027_),
    .S(_2030_),
    .X(_2035_));
 sg13g2_nand2b_1 _2874_ (.Y(_2036_),
    .B(_0034_),
    .A_N(_2035_));
 sg13g2_xnor2_1 _2875_ (.Y(_2037_),
    .A(_0026_),
    .B(_2031_));
 sg13g2_or2_1 _2876_ (.X(_2038_),
    .B(_2035_),
    .A(\game.fsm.block_len[6][1] ));
 sg13g2_and2_1 _2877_ (.A(_1873_),
    .B(_2035_),
    .X(_2039_));
 sg13g2_o21ai_1 _2878_ (.B1(_1938_),
    .Y(_2040_),
    .A1(_1873_),
    .A2(_2035_));
 sg13g2_a221oi_1 _2879_ (.B2(_2040_),
    .C1(_2039_),
    .B1(_2038_),
    .A1(_2036_),
    .Y(_2041_),
    .A2(_2037_));
 sg13g2_a21oi_1 _2880_ (.A1(\game.fsm.block_len[6][2] ),
    .A2(_2033_),
    .Y(_2042_),
    .B1(_1942_));
 sg13g2_o21ai_1 _2881_ (.B1(_2042_),
    .Y(_2043_),
    .A1(_2034_),
    .A2(_2041_));
 sg13g2_mux2_1 _2882_ (.A0(_0026_),
    .A1(_2031_),
    .S(_2043_),
    .X(_2044_));
 sg13g2_nand2_1 _2883_ (.Y(_2045_),
    .A(_1922_),
    .B(_1981_));
 sg13g2_nand3_1 _2884_ (.B(\game.fsm.block_len[0][0] ),
    .C(_1983_),
    .A(_1843_),
    .Y(_2046_));
 sg13g2_a21oi_2 _2885_ (.B1(_2045_),
    .Y(_2047_),
    .A2(_2046_),
    .A1(_1982_));
 sg13g2_mux2_1 _2886_ (.A0(_0031_),
    .A1(_0030_),
    .S(_2047_),
    .X(_2048_));
 sg13g2_nand3_1 _2887_ (.B(\game.fsm.block_len[2][0] ),
    .C(_1916_),
    .A(_1844_),
    .Y(_2049_));
 sg13g2_a221oi_1 _2888_ (.B2(_2049_),
    .C1(_1914_),
    .B1(_1915_),
    .A1(\game.fsm.block_len[3][2] ),
    .Y(_2050_),
    .A2(_1854_));
 sg13g2_mux2_1 _2889_ (.A0(_0075_),
    .A1(_0074_),
    .S(_2050_),
    .X(_2051_));
 sg13g2_inv_1 _2890_ (.Y(_2052_),
    .A(_2051_));
 sg13g2_mux2_1 _2891_ (.A0(_0073_),
    .A1(_0072_),
    .S(_2047_),
    .X(_2053_));
 sg13g2_nor2_1 _2892_ (.A(_2052_),
    .B(_2053_),
    .Y(_2054_));
 sg13g2_mux2_1 _2893_ (.A0(_0033_),
    .A1(_0032_),
    .S(_2050_),
    .X(_2055_));
 sg13g2_nor2b_1 _2894_ (.A(_2055_),
    .B_N(_2048_),
    .Y(_2056_));
 sg13g2_nand2b_1 _2895_ (.Y(_2057_),
    .B(_2055_),
    .A_N(_2048_));
 sg13g2_mux2_1 _2896_ (.A0(_0066_),
    .A1(_0065_),
    .S(_2047_),
    .X(_2058_));
 sg13g2_mux2_1 _2897_ (.A0(_0068_),
    .A1(_0067_),
    .S(_2050_),
    .X(_2059_));
 sg13g2_nor2b_1 _2898_ (.A(_2059_),
    .B_N(_2058_),
    .Y(_2060_));
 sg13g2_o21ai_1 _2899_ (.B1(_2057_),
    .Y(_2061_),
    .A1(_2056_),
    .A2(_2060_));
 sg13g2_a21oi_1 _2900_ (.A1(_2052_),
    .A2(_2053_),
    .Y(_2062_),
    .B1(_1912_));
 sg13g2_o21ai_1 _2901_ (.B1(_2062_),
    .Y(_2063_),
    .A1(_2054_),
    .A2(_2061_));
 sg13g2_nand2b_1 _2902_ (.Y(_2064_),
    .B(_2063_),
    .A_N(_2048_));
 sg13g2_o21ai_1 _2903_ (.B1(_2064_),
    .Y(_2065_),
    .A1(_2055_),
    .A2(_2063_));
 sg13g2_nor2_1 _2904_ (.A(_1873_),
    .B(_2043_),
    .Y(_2066_));
 sg13g2_a21oi_2 _2905_ (.B1(_2066_),
    .Y(_2067_),
    .A2(_2043_),
    .A1(_2035_));
 sg13g2_inv_1 _2906_ (.Y(_2068_),
    .A(_2067_));
 sg13g2_nand2b_1 _2907_ (.Y(_2069_),
    .B(_2067_),
    .A_N(_2065_));
 sg13g2_mux2_1 _2908_ (.A0(_2059_),
    .A1(_2058_),
    .S(_2063_),
    .X(_2070_));
 sg13g2_inv_1 _2909_ (.Y(_2071_),
    .A(_2070_));
 sg13g2_nand3_1 _2910_ (.B(_2069_),
    .C(_2071_),
    .A(_2044_),
    .Y(_2072_));
 sg13g2_a21oi_1 _2911_ (.A1(_1913_),
    .A2(_2051_),
    .Y(_2073_),
    .B1(_2053_));
 sg13g2_mux2_1 _2912_ (.A0(_0029_),
    .A1(_2033_),
    .S(_2043_),
    .X(_2074_));
 sg13g2_a22oi_1 _2913_ (.Y(_2075_),
    .B1(_2073_),
    .B2(_2074_),
    .A2(_2068_),
    .A1(_2065_));
 sg13g2_nand2b_1 _2914_ (.Y(_0388_),
    .B(_2074_),
    .A_N(_1946_));
 sg13g2_nand2b_1 _2915_ (.Y(_0389_),
    .B(_2073_),
    .A_N(_1946_));
 sg13g2_a22oi_1 _2916_ (.Y(_0390_),
    .B1(_0388_),
    .B2(_0389_),
    .A2(_2075_),
    .A1(_2072_));
 sg13g2_nand2_1 _2917_ (.Y(_0391_),
    .A(_2044_),
    .B(_0390_));
 sg13g2_o21ai_1 _2918_ (.B1(_0391_),
    .Y(_0392_),
    .A1(_2071_),
    .A2(_0390_));
 sg13g2_nor2_1 _2919_ (.A(_2065_),
    .B(_0390_),
    .Y(_0393_));
 sg13g2_a21oi_1 _2920_ (.A1(_2068_),
    .A2(_0390_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_nand2b_1 _2921_ (.Y(_0395_),
    .B(_0394_),
    .A_N(_0392_));
 sg13g2_nand2_1 _2922_ (.Y(_0396_),
    .A(_2023_),
    .B(_0394_));
 sg13g2_o21ai_1 _2923_ (.B1(_0396_),
    .Y(_0397_),
    .A1(_2016_),
    .A2(_0392_));
 sg13g2_nor2b_1 _2924_ (.A(net392),
    .B_N(net391),
    .Y(_0398_));
 sg13g2_nand2b_1 _2925_ (.Y(_0399_),
    .B(net391),
    .A_N(net392));
 sg13g2_a21oi_1 _2926_ (.A1(_2073_),
    .A2(_0388_),
    .Y(_0400_),
    .B1(_0399_));
 sg13g2_o21ai_1 _2927_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_2018_),
    .A2(_0395_));
 sg13g2_a21o_1 _2928_ (.A2(_0397_),
    .A1(_0395_),
    .B1(_0401_),
    .X(_0402_));
 sg13g2_and2_2 _2929_ (.A(net391),
    .B(\game.current_level[0] ),
    .X(_0403_));
 sg13g2_nand2_2 _2930_ (.Y(_0404_),
    .A(\game.current_level[1] ),
    .B(net392));
 sg13g2_nor4_1 _2931_ (.A(\game.fsm.len1_color_count[3][2] ),
    .B(\game.fsm.len1_color_count[3][1] ),
    .C(\game.fsm.len2_color_count[1][1] ),
    .D(\game.fsm.len2_color_count[3][1] ),
    .Y(_0405_));
 sg13g2_nor4_1 _2932_ (.A(\game.fsm.len1_color_count[0][2] ),
    .B(\game.fsm.len1_color_count[0][1] ),
    .C(\game.fsm.len1_color_count[1][2] ),
    .D(\game.fsm.len1_color_count[1][1] ),
    .Y(_0406_));
 sg13g2_nor4_1 _2933_ (.A(\game.fsm.len3_color_count[3][1] ),
    .B(\game.fsm.len2_color_count[0][1] ),
    .C(\game.fsm.len1_color_count[2][2] ),
    .D(\game.fsm.len1_color_count[2][1] ),
    .Y(_0407_));
 sg13g2_nor2_1 _2934_ (.A(\game.fsm.len3_color_count[1][1] ),
    .B(\game.fsm.len2_color_count[2][1] ),
    .Y(_0408_));
 sg13g2_nand4_1 _2935_ (.B(_0406_),
    .C(_0407_),
    .A(_0405_),
    .Y(_0409_),
    .D(_0408_));
 sg13g2_nor3_1 _2936_ (.A(\game.fsm.len3_color_count[0][1] ),
    .B(\game.fsm.len3_color_count[2][1] ),
    .C(_0409_),
    .Y(_0410_));
 sg13g2_nor3_2 _2937_ (.A(_1809_),
    .B(\game.current_level[3] ),
    .C(\game.current_level[2] ),
    .Y(_0411_));
 sg13g2_o21ai_1 _2938_ (.B1(_0411_),
    .Y(_0412_),
    .A1(_0404_),
    .A2(_0410_));
 sg13g2_nor2b_1 _2939_ (.A(_0412_),
    .B_N(_0402_),
    .Y(_0413_));
 sg13g2_o21ai_1 _2940_ (.B1(_1980_),
    .Y(_0414_),
    .A1(_1947_),
    .A2(_2024_));
 sg13g2_a22oi_1 _2941_ (.Y(_0415_),
    .B1(\game.fsm.block_len[1][2] ),
    .B2(_1854_),
    .A2(_1851_),
    .A1(\game.fsm.block_len[1][1] ));
 sg13g2_nand2_1 _2942_ (.Y(_0416_),
    .A(_1843_),
    .B(\game.fsm.block_len[2][0] ));
 sg13g2_o21ai_1 _2943_ (.B1(_0416_),
    .Y(_0417_),
    .A1(\game.fsm.block_len[1][1] ),
    .A2(_1851_));
 sg13g2_a22oi_1 _2944_ (.Y(_0418_),
    .B1(_0415_),
    .B2(_0417_),
    .A2(\game.fsm.block_len[2][2] ),
    .A1(_1852_));
 sg13g2_nor2_1 _2945_ (.A(_1912_),
    .B(_0418_),
    .Y(_0419_));
 sg13g2_nand2_1 _2946_ (.Y(_0420_),
    .A(_1850_),
    .B(\game.fsm.block_len[4][1] ));
 sg13g2_o21ai_1 _2947_ (.B1(_0420_),
    .Y(_0421_),
    .A1(\game.fsm.block_len[3][0] ),
    .A2(_1847_));
 sg13g2_nand2b_1 _2948_ (.Y(_0422_),
    .B(\game.fsm.block_len[3][2] ),
    .A_N(\game.fsm.block_len[4][2] ));
 sg13g2_o21ai_1 _2949_ (.B1(_0422_),
    .Y(_0423_),
    .A1(_1850_),
    .A2(\game.fsm.block_len[4][1] ));
 sg13g2_nand2b_1 _2950_ (.Y(_0424_),
    .B(_0421_),
    .A_N(_0423_));
 sg13g2_nand2_1 _2951_ (.Y(_0425_),
    .A(_1853_),
    .B(\game.fsm.block_len[4][2] ));
 sg13g2_a21oi_1 _2952_ (.A1(_0424_),
    .A2(_0425_),
    .Y(_0426_),
    .B1(_1946_));
 sg13g2_nor3_1 _2953_ (.A(_1986_),
    .B(_0419_),
    .C(_0426_),
    .Y(_0427_));
 sg13g2_nand3_1 _2954_ (.B(_1932_),
    .C(_0427_),
    .A(_1919_),
    .Y(_0428_));
 sg13g2_o21ai_1 _2955_ (.B1(_0415_),
    .Y(_0429_),
    .A1(_1843_),
    .A2(\game.fsm.block_len[2][0] ));
 sg13g2_and2_1 _2956_ (.A(_1913_),
    .B(_0418_),
    .X(_0430_));
 sg13g2_o21ai_1 _2957_ (.B1(_0430_),
    .Y(_0431_),
    .A1(_0417_),
    .A2(_0429_));
 sg13g2_nor2_1 _2958_ (.A(_1844_),
    .B(\game.fsm.block_len[4][0] ),
    .Y(_0432_));
 sg13g2_nor3_1 _2959_ (.A(_0421_),
    .B(_0423_),
    .C(_0432_),
    .Y(_0433_));
 sg13g2_nor2_1 _2960_ (.A(_1946_),
    .B(_0433_),
    .Y(_0434_));
 sg13g2_nand3_1 _2961_ (.B(_0425_),
    .C(_0434_),
    .A(_0424_),
    .Y(_0435_));
 sg13g2_nor3_1 _2962_ (.A(_2030_),
    .B(_2047_),
    .C(_2050_),
    .Y(_0436_));
 sg13g2_and2_1 _2963_ (.A(_0435_),
    .B(_0436_),
    .X(_0437_));
 sg13g2_a21oi_1 _2964_ (.A1(_0431_),
    .A2(_0437_),
    .Y(_0438_),
    .B1(_0399_));
 sg13g2_nor3_1 _2965_ (.A(\game.fsm.color_count[2][1] ),
    .B(\game.fsm.color_count[2][0] ),
    .C(_1872_),
    .Y(_0439_));
 sg13g2_nor2_1 _2966_ (.A(\game.fsm.color_count[1][1] ),
    .B(\game.fsm.color_count[1][0] ),
    .Y(_0440_));
 sg13g2_and2_1 _2967_ (.A(_0023_),
    .B(_0440_),
    .X(_0441_));
 sg13g2_nand2_1 _2968_ (.Y(_0442_),
    .A(_0023_),
    .B(_0440_));
 sg13g2_xnor2_1 _2969_ (.Y(_0443_),
    .A(\game.fsm.color_count[1][2] ),
    .B(\game.fsm.color_count[2][2] ));
 sg13g2_a22oi_1 _2970_ (.Y(_0444_),
    .B1(_1871_),
    .B2(\game.fsm.color_count[1][0] ),
    .A2(_1870_),
    .A1(\game.fsm.color_count[1][1] ));
 sg13g2_a22oi_1 _2971_ (.Y(_0445_),
    .B1(\game.fsm.color_count[2][0] ),
    .B2(_1863_),
    .A2(\game.fsm.color_count[2][1] ),
    .A1(_1862_));
 sg13g2_nand3_1 _2972_ (.B(_0444_),
    .C(_0445_),
    .A(_0443_),
    .Y(_0446_));
 sg13g2_nor3_1 _2973_ (.A(\game.fsm.color_count[3][1] ),
    .B(\game.fsm.color_count[3][0] ),
    .C(_1868_),
    .Y(_0447_));
 sg13g2_nand3b_1 _2974_ (.B(_1867_),
    .C(_0024_),
    .Y(_0448_),
    .A_N(net404));
 sg13g2_a22oi_1 _2975_ (.Y(_0449_),
    .B1(_1870_),
    .B2(net404),
    .A2(_1869_),
    .A1(\game.fsm.color_count[3][2] ));
 sg13g2_nand2_1 _2976_ (.Y(_0450_),
    .A(\game.fsm.color_count[3][0] ),
    .B(_1871_));
 sg13g2_nor2_1 _2977_ (.A(net404),
    .B(_1870_),
    .Y(_0451_));
 sg13g2_nand2_1 _2978_ (.Y(_0452_),
    .A(_1866_),
    .B(\game.fsm.color_count[2][2] ));
 sg13g2_a21oi_1 _2979_ (.A1(_1867_),
    .A2(\game.fsm.color_count[2][0] ),
    .Y(_0453_),
    .B1(_0451_));
 sg13g2_nand4_1 _2980_ (.B(_0450_),
    .C(_0452_),
    .A(_0449_),
    .Y(_0454_),
    .D(_0453_));
 sg13g2_a22oi_1 _2981_ (.Y(_0455_),
    .B1(_0448_),
    .B2(_0454_),
    .A2(_0446_),
    .A1(_0442_));
 sg13g2_nor3_2 _2982_ (.A(\game.fsm.color_count[0][0] ),
    .B(\game.fsm.color_count[0][1] ),
    .C(\game.fsm.color_count[0][2] ),
    .Y(_0456_));
 sg13g2_xnor2_1 _2983_ (.Y(_0457_),
    .A(net410),
    .B(\game.fsm.color_count[3][0] ));
 sg13g2_nor2_1 _2984_ (.A(net409),
    .B(net404),
    .Y(_0458_));
 sg13g2_xnor2_1 _2985_ (.Y(_0459_),
    .A(net409),
    .B(net404));
 sg13g2_xnor2_1 _2986_ (.Y(_0460_),
    .A(\game.fsm.color_count[0][2] ),
    .B(\game.fsm.color_count[3][2] ));
 sg13g2_inv_1 _2987_ (.Y(_0461_),
    .A(_0460_));
 sg13g2_nand3_1 _2988_ (.B(_0459_),
    .C(_0460_),
    .A(_0457_),
    .Y(_0462_));
 sg13g2_xnor2_1 _2989_ (.Y(_0463_),
    .A(\game.fsm.color_count[1][2] ),
    .B(\game.fsm.color_count[0][2] ));
 sg13g2_xnor2_1 _2990_ (.Y(_0464_),
    .A(\game.fsm.color_count[1][1] ),
    .B(net409));
 sg13g2_xnor2_1 _2991_ (.Y(_0465_),
    .A(\game.fsm.color_count[1][0] ),
    .B(net410));
 sg13g2_nand3_1 _2992_ (.B(_0464_),
    .C(_0465_),
    .A(_0463_),
    .Y(_0466_));
 sg13g2_a22oi_1 _2993_ (.Y(_0467_),
    .B1(_0466_),
    .B2(_0442_),
    .A2(_0462_),
    .A1(_0448_));
 sg13g2_nor2_1 _2994_ (.A(_0456_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_nand2_1 _2995_ (.Y(_0469_),
    .A(_0442_),
    .B(_0448_));
 sg13g2_xor2_1 _2996_ (.B(net404),
    .A(\game.fsm.color_count[1][1] ),
    .X(_0470_));
 sg13g2_a22oi_1 _2997_ (.Y(_0471_),
    .B1(\game.fsm.color_count[3][0] ),
    .B2(_1863_),
    .A2(\game.fsm.color_count[3][2] ),
    .A1(_1861_));
 sg13g2_a221oi_1 _2998_ (.B2(\game.fsm.color_count[1][0] ),
    .C1(_0470_),
    .B1(_1867_),
    .A1(\game.fsm.color_count[1][2] ),
    .Y(_0472_),
    .A2(_1866_));
 sg13g2_a21oi_1 _2999_ (.A1(_0471_),
    .A2(_0472_),
    .Y(_0473_),
    .B1(_0469_));
 sg13g2_or2_1 _3000_ (.X(_0474_),
    .B(_0456_),
    .A(_0439_));
 sg13g2_a22oi_1 _3001_ (.Y(_0475_),
    .B1(\game.fsm.color_count[2][0] ),
    .B2(_1864_),
    .A2(\game.fsm.color_count[2][2] ),
    .A1(_1865_));
 sg13g2_xor2_1 _3002_ (.B(\game.fsm.color_count[2][1] ),
    .A(net409),
    .X(_0476_));
 sg13g2_a221oi_1 _3003_ (.B2(net410),
    .C1(_0476_),
    .B1(_1871_),
    .A1(\game.fsm.color_count[0][2] ),
    .Y(_0477_),
    .A2(_1869_));
 sg13g2_a21oi_1 _3004_ (.A1(_0475_),
    .A2(_0477_),
    .Y(_0478_),
    .B1(_0474_));
 sg13g2_nor3_1 _3005_ (.A(_0468_),
    .B(_0473_),
    .C(_0478_),
    .Y(_0479_));
 sg13g2_o21ai_1 _3006_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0439_),
    .A2(_0455_));
 sg13g2_or2_2 _3007_ (.X(_0481_),
    .B(net392),
    .A(net391));
 sg13g2_nor2b_1 _3008_ (.A(\game.fsm.len2_block_count[0] ),
    .B_N(\game.fsm.len2_block_count[1] ),
    .Y(_0482_));
 sg13g2_o21ai_1 _3009_ (.B1(net390),
    .Y(_0483_),
    .A1(_0481_),
    .A2(_0482_));
 sg13g2_a221oi_1 _3010_ (.B2(_0403_),
    .C1(_0483_),
    .B1(_0480_),
    .A1(_0428_),
    .Y(_0484_),
    .A2(_0438_));
 sg13g2_nand2_1 _3011_ (.Y(_0485_),
    .A(_0414_),
    .B(_0484_));
 sg13g2_a21oi_1 _3012_ (.A1(net409),
    .A2(net404),
    .Y(_0486_),
    .B1(_0461_));
 sg13g2_nor2_1 _3013_ (.A(_0458_),
    .B(_0460_),
    .Y(_0487_));
 sg13g2_nor4_1 _3014_ (.A(net392),
    .B(_0457_),
    .C(_0486_),
    .D(_0487_),
    .Y(_0488_));
 sg13g2_or2_1 _3015_ (.X(_0489_),
    .B(\game.fsm.len1_block_count[0] ),
    .A(\game.fsm.len1_block_count[1] ));
 sg13g2_o21ai_1 _3016_ (.B1(net392),
    .Y(_0490_),
    .A1(\game.fsm.len2_block_count[1] ),
    .A2(\game.fsm.len2_block_count[0] ));
 sg13g2_nor3_2 _3017_ (.A(\game.fsm.len1_block_count[2] ),
    .B(_0489_),
    .C(_0490_),
    .Y(_0491_));
 sg13g2_nor3_1 _3018_ (.A(net391),
    .B(_0488_),
    .C(_0491_),
    .Y(_0492_));
 sg13g2_nor3_1 _3019_ (.A(\game.fsm.green_block_count[2] ),
    .B(_1814_),
    .C(\game.fsm.green_block_count[0] ),
    .Y(_0493_));
 sg13g2_a21oi_1 _3020_ (.A1(\game.fsm.num_blocks[2] ),
    .A2(_1945_),
    .Y(_0494_),
    .B1(_0399_));
 sg13g2_nor3_1 _3021_ (.A(net390),
    .B(_0492_),
    .C(_0494_),
    .Y(_0495_));
 sg13g2_o21ai_1 _3022_ (.B1(_0495_),
    .Y(_0496_),
    .A1(_0404_),
    .A2(_0493_));
 sg13g2_nand3_1 _3023_ (.B(_0485_),
    .C(_0496_),
    .A(\game.current_level[3] ),
    .Y(_0497_));
 sg13g2_nor2_2 _3024_ (.A(net397),
    .B(net401),
    .Y(_0498_));
 sg13g2_nand2_2 _3025_ (.Y(_0499_),
    .A(\game.fsm.length[1] ),
    .B(net401));
 sg13g2_nor2b_2 _3026_ (.A(_0498_),
    .B_N(_0499_),
    .Y(_0500_));
 sg13g2_nand2b_2 _3027_ (.Y(_0501_),
    .B(_0499_),
    .A_N(_0498_));
 sg13g2_mux2_1 _3028_ (.A0(\game.fsm.seq[3][1] ),
    .A1(\game.fsm.seq[2][1] ),
    .S(net400),
    .X(_0502_));
 sg13g2_xnor2_1 _3029_ (.Y(_0503_),
    .A(_0064_),
    .B(_0498_));
 sg13g2_inv_1 _3030_ (.Y(_0504_),
    .A(_0503_));
 sg13g2_mux2_1 _3031_ (.A0(\game.fsm.seq[1][1] ),
    .A1(\game.fsm.seq[0][1] ),
    .S(net400),
    .X(_0505_));
 sg13g2_mux2_1 _3032_ (.A0(\game.fsm.seq[5][1] ),
    .A1(\game.fsm.seq[4][1] ),
    .S(net398),
    .X(_0506_));
 sg13g2_nor2_1 _3033_ (.A(net398),
    .B(\game.fsm.seq[7][1] ),
    .Y(_0507_));
 sg13g2_a21oi_2 _3034_ (.B1(_0507_),
    .Y(_0508_),
    .A2(_1823_),
    .A1(net398));
 sg13g2_mux4_1 _3035_ (.S0(_0500_),
    .A0(_0502_),
    .A1(_0505_),
    .A2(_0508_),
    .A3(_0506_),
    .S1(_0503_),
    .X(_0509_));
 sg13g2_inv_2 _3036_ (.Y(_0510_),
    .A(_0509_));
 sg13g2_xor2_1 _3037_ (.B(net354),
    .A(\game.fsm.seq[0][1] ),
    .X(_0511_));
 sg13g2_mux2_1 _3038_ (.A0(\game.fsm.seq[3][0] ),
    .A1(\game.fsm.seq[2][0] ),
    .S(net400),
    .X(_0512_));
 sg13g2_and2_1 _3039_ (.A(net400),
    .B(_0063_),
    .X(_0513_));
 sg13g2_a21oi_1 _3040_ (.A1(_1822_),
    .A2(_0062_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_nor2_1 _3041_ (.A(net399),
    .B(\game.fsm.seq[5][0] ),
    .Y(_0515_));
 sg13g2_a21oi_1 _3042_ (.A1(net399),
    .A2(_1842_),
    .Y(_0516_),
    .B1(_0515_));
 sg13g2_nor2_1 _3043_ (.A(net399),
    .B(\game.fsm.seq[7][0] ),
    .Y(_0517_));
 sg13g2_a21oi_1 _3044_ (.A1(net399),
    .A2(_1824_),
    .Y(_0518_),
    .B1(_0517_));
 sg13g2_mux4_1 _3045_ (.S0(_0500_),
    .A0(_0512_),
    .A1(_0514_),
    .A2(_0518_),
    .A3(_0516_),
    .S1(_0503_),
    .X(_0519_));
 sg13g2_inv_2 _3046_ (.Y(_0520_),
    .A(net353));
 sg13g2_xnor2_1 _3047_ (.Y(_0521_),
    .A(_0063_),
    .B(net353));
 sg13g2_nor2_1 _3048_ (.A(_0511_),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_nand2_1 _3049_ (.Y(_0523_),
    .A(net396),
    .B(net397));
 sg13g2_nor2_1 _3050_ (.A(net396),
    .B(net397),
    .Y(_0524_));
 sg13g2_xor2_1 _3051_ (.B(net397),
    .A(net396),
    .X(_0525_));
 sg13g2_mux2_1 _3052_ (.A0(\game.fsm.seq[2][1] ),
    .A1(\game.fsm.seq[3][1] ),
    .S(net398),
    .X(_0526_));
 sg13g2_mux2_1 _3053_ (.A0(\game.fsm.seq[0][1] ),
    .A1(\game.fsm.seq[1][1] ),
    .S(net398),
    .X(_0527_));
 sg13g2_mux2_1 _3054_ (.A0(\game.fsm.seq[4][1] ),
    .A1(\game.fsm.seq[5][1] ),
    .S(net398),
    .X(_0528_));
 sg13g2_mux2_1 _3055_ (.A0(\game.fsm.seq[6][1] ),
    .A1(\game.fsm.seq[7][1] ),
    .S(net398),
    .X(_0529_));
 sg13g2_mux4_1 _3056_ (.S0(net397),
    .A0(_0526_),
    .A1(_0528_),
    .A2(_0529_),
    .A3(_0527_),
    .S1(_1820_),
    .X(_0530_));
 sg13g2_xnor2_1 _3057_ (.Y(_0531_),
    .A(\game.fsm.seq[1][1] ),
    .B(_0530_));
 sg13g2_mux4_1 _3058_ (.S0(net396),
    .A0(\game.fsm.seq[0][0] ),
    .A1(\game.fsm.seq[2][0] ),
    .A2(\game.fsm.seq[1][0] ),
    .A3(\game.fsm.seq[3][0] ),
    .S1(net398),
    .X(_0532_));
 sg13g2_mux2_1 _3059_ (.A0(\game.fsm.seq[6][0] ),
    .A1(\game.fsm.seq[7][0] ),
    .S(net399),
    .X(_0533_));
 sg13g2_nor2_1 _3060_ (.A(net399),
    .B(\game.fsm.seq[4][0] ),
    .Y(_0534_));
 sg13g2_nor2_1 _3061_ (.A(_1822_),
    .B(\game.fsm.seq[5][0] ),
    .Y(_0535_));
 sg13g2_nor3_1 _3062_ (.A(_0523_),
    .B(_0534_),
    .C(_0535_),
    .Y(_0536_));
 sg13g2_a221oi_1 _3063_ (.B2(_0524_),
    .C1(_0536_),
    .B1(_0533_),
    .A1(_0525_),
    .Y(_0537_),
    .A2(_0532_));
 sg13g2_xnor2_1 _3064_ (.Y(_0538_),
    .A(_0062_),
    .B(_0537_));
 sg13g2_nand2_1 _3065_ (.Y(_0539_),
    .A(_0531_),
    .B(_0538_));
 sg13g2_xnor2_1 _3066_ (.Y(_0540_),
    .A(_1820_),
    .B(_0499_));
 sg13g2_mux4_1 _3067_ (.S0(_0501_),
    .A0(_0512_),
    .A1(_0514_),
    .A2(_0518_),
    .A3(_0516_),
    .S1(_0540_),
    .X(_0541_));
 sg13g2_xnor2_1 _3068_ (.Y(_0542_),
    .A(\game.fsm.seq[2][0] ),
    .B(_0541_));
 sg13g2_mux4_1 _3069_ (.S0(_0501_),
    .A0(_0502_),
    .A1(_0505_),
    .A2(_0508_),
    .A3(_0506_),
    .S1(_0540_),
    .X(_0543_));
 sg13g2_xnor2_1 _3070_ (.Y(_0544_),
    .A(\game.fsm.seq[2][1] ),
    .B(_0543_));
 sg13g2_a21oi_1 _3071_ (.A1(_0542_),
    .A2(_0544_),
    .Y(_0545_),
    .B1(_1821_));
 sg13g2_o21ai_1 _3072_ (.B1(net396),
    .Y(_0546_),
    .A1(_0539_),
    .A2(_0545_));
 sg13g2_a221oi_1 _3073_ (.B2(_0546_),
    .C1(_0481_),
    .B1(_0522_),
    .A1(_1820_),
    .Y(_0547_),
    .A2(_1821_));
 sg13g2_nor3_1 _3074_ (.A(_0404_),
    .B(_0447_),
    .C(_0456_),
    .Y(_0548_));
 sg13g2_a21oi_1 _3075_ (.A1(_0398_),
    .A2(_0441_),
    .Y(_0549_),
    .B1(_0548_));
 sg13g2_a21oi_1 _3076_ (.A1(_1980_),
    .A2(_0522_),
    .Y(_0550_),
    .B1(_0547_));
 sg13g2_a21o_1 _3077_ (.A2(_0550_),
    .A1(_0549_),
    .B1(net390),
    .X(_0551_));
 sg13g2_a21oi_1 _3078_ (.A1(_0439_),
    .A2(_0456_),
    .Y(_0552_),
    .B1(_0469_));
 sg13g2_nand2_1 _3079_ (.Y(_0553_),
    .A(_0441_),
    .B(_0447_));
 sg13g2_nor2b_1 _3080_ (.A(_0474_),
    .B_N(_0469_),
    .Y(_0554_));
 sg13g2_a22oi_1 _3081_ (.Y(_0555_),
    .B1(_0553_),
    .B2(_0554_),
    .A2(_0552_),
    .A1(_0474_));
 sg13g2_nor2_1 _3082_ (.A(_0481_),
    .B(_0555_),
    .Y(_0556_));
 sg13g2_o21ai_1 _3083_ (.B1(_0449_),
    .Y(_0557_),
    .A1(_0450_),
    .A2(_0451_));
 sg13g2_nand3_1 _3084_ (.B(_0452_),
    .C(_0557_),
    .A(_0398_),
    .Y(_0558_));
 sg13g2_nand4_1 _3085_ (.B(net409),
    .C(_1865_),
    .A(net410),
    .Y(_0559_),
    .D(_1980_));
 sg13g2_nor2_1 _3086_ (.A(\game.fsm.seq[1][1] ),
    .B(\game.fsm.seq[2][1] ),
    .Y(_0560_));
 sg13g2_nor2_1 _3087_ (.A(\game.fsm.seq[1][0] ),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_a22oi_1 _3088_ (.Y(_0562_),
    .B1(_0499_),
    .B2(_0064_),
    .A2(\game.fsm.seq[2][1] ),
    .A1(\game.fsm.seq[1][1] ));
 sg13g2_nor2_1 _3089_ (.A(_1820_),
    .B(\game.fsm.seq[3][0] ),
    .Y(_0563_));
 sg13g2_xor2_1 _3090_ (.B(\game.fsm.seq[2][1] ),
    .A(\game.fsm.seq[3][1] ),
    .X(_0564_));
 sg13g2_a22oi_1 _3091_ (.Y(_0565_),
    .B1(_0563_),
    .B2(_0564_),
    .A2(_0562_),
    .A1(_0561_));
 sg13g2_nor2_1 _3092_ (.A(_0092_),
    .B(\game.fsm.seq[6][0] ),
    .Y(_0566_));
 sg13g2_o21ai_1 _3093_ (.B1(\game.fsm.seq[5][1] ),
    .Y(_0567_),
    .A1(\game.fsm.seq[4][0] ),
    .A2(\game.fsm.seq[4][1] ));
 sg13g2_a21oi_1 _3094_ (.A1(_1823_),
    .A2(_0566_),
    .Y(_0568_),
    .B1(_0567_));
 sg13g2_a221oi_1 _3095_ (.B2(\game.fsm.seq[6][1] ),
    .C1(\game.fsm.seq[5][1] ),
    .B1(_0566_),
    .A1(_1842_),
    .Y(_0569_),
    .A2(\game.fsm.seq[4][1] ));
 sg13g2_nor4_1 _3096_ (.A(\game.fsm.seq[5][0] ),
    .B(_0523_),
    .C(_0568_),
    .D(_0569_),
    .Y(_0570_));
 sg13g2_or2_1 _3097_ (.X(_0571_),
    .B(\game.fsm.seq[4][0] ),
    .A(\game.fsm.seq[3][0] ));
 sg13g2_xnor2_1 _3098_ (.Y(_0572_),
    .A(\game.fsm.seq[3][1] ),
    .B(\game.fsm.seq[4][1] ));
 sg13g2_nor4_1 _3099_ (.A(_0064_),
    .B(_0498_),
    .C(_0571_),
    .D(_0572_),
    .Y(_0573_));
 sg13g2_xnor2_1 _3100_ (.Y(_0574_),
    .A(\game.fsm.seq[1][1] ),
    .B(\game.fsm.seq[0][1] ));
 sg13g2_nor4_1 _3101_ (.A(\game.fsm.seq[1][0] ),
    .B(\game.fsm.seq[0][0] ),
    .C(_0524_),
    .D(_0574_),
    .Y(_0575_));
 sg13g2_nor4_1 _3102_ (.A(_0404_),
    .B(_0570_),
    .C(_0573_),
    .D(_0575_),
    .Y(_0576_));
 sg13g2_o21ai_1 _3103_ (.B1(_0576_),
    .Y(_0577_),
    .A1(\game.fsm.seq[2][0] ),
    .A2(_0565_));
 sg13g2_nand4_1 _3104_ (.B(_0558_),
    .C(_0559_),
    .A(net390),
    .Y(_0578_),
    .D(_0577_));
 sg13g2_o21ai_1 _3105_ (.B1(_0551_),
    .Y(_0579_),
    .A1(_0556_),
    .A2(_0578_));
 sg13g2_a21oi_1 _3106_ (.A1(_1810_),
    .A2(_0579_),
    .Y(_0580_),
    .B1(\game.current_level[4] ));
 sg13g2_a22oi_1 _3107_ (.Y(_0581_),
    .B1(_0497_),
    .B2(_0580_),
    .A2(_0413_),
    .A1(_2027_));
 sg13g2_xor2_1 _3108_ (.B(_0581_),
    .A(\game.slv.saved_target ),
    .X(_0582_));
 sg13g2_nand2b_1 _3109_ (.Y(_0583_),
    .B(net481),
    .A_N(_0582_));
 sg13g2_nand2b_1 _3110_ (.Y(_0584_),
    .B(net402),
    .A_N(_1897_));
 sg13g2_nor3_1 _3111_ (.A(net680),
    .B(\game.slv.pos[1] ),
    .C(\game.slv.pos[0] ),
    .Y(_0585_));
 sg13g2_or3_1 _3112_ (.A(\game.slv.pos[2] ),
    .B(\game.slv.pos[1] ),
    .C(\game.slv.pos[0] ),
    .X(_0586_));
 sg13g2_nand2_1 _3113_ (.Y(_0587_),
    .A(net682),
    .B(_0586_));
 sg13g2_nand3_1 _3114_ (.B(_0584_),
    .C(_0587_),
    .A(_0583_),
    .Y(_0588_));
 sg13g2_and2_1 _3115_ (.A(_1899_),
    .B(_0588_),
    .X(_0011_));
 sg13g2_nor2_2 _3116_ (.A(\game.state[3] ),
    .B(\game.state[2] ),
    .Y(_0589_));
 sg13g2_nand2_2 _3117_ (.Y(_0590_),
    .A(_1802_),
    .B(_1803_));
 sg13g2_nor2_1 _3118_ (.A(net381),
    .B(net383),
    .Y(_0591_));
 sg13g2_nor2_1 _3119_ (.A(net381),
    .B(_0590_),
    .Y(_0592_));
 sg13g2_nand2_1 _3120_ (.Y(_0593_),
    .A(_1804_),
    .B(_0589_));
 sg13g2_nor2_1 _3121_ (.A(net383),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_nand2_2 _3122_ (.Y(_0595_),
    .A(_0589_),
    .B(_0591_));
 sg13g2_nor2b_2 _3123_ (.A(\btn.input_event[0] ),
    .B_N(\btn.input_event[1] ),
    .Y(_0596_));
 sg13g2_nor2_1 _3124_ (.A(\btn.input_event[3] ),
    .B(\btn.input_event[2] ),
    .Y(_0597_));
 sg13g2_nand2_1 _3125_ (.Y(_0598_),
    .A(\btn.input_event[4] ),
    .B(_0597_));
 sg13g2_nand3_1 _3126_ (.B(_0596_),
    .C(_0597_),
    .A(\btn.input_event[4] ),
    .Y(_0599_));
 sg13g2_and2_2 _3127_ (.A(net351),
    .B(_0599_),
    .X(_0600_));
 sg13g2_nand2_2 _3128_ (.Y(_0601_),
    .A(net351),
    .B(_0599_));
 sg13g2_nand3_1 _3129_ (.B(\game.current_level[2] ),
    .C(_0403_),
    .A(\game.current_level[3] ),
    .Y(_0602_));
 sg13g2_xor2_1 _3130_ (.B(_0602_),
    .A(_0084_),
    .X(_0603_));
 sg13g2_nand3_1 _3131_ (.B(\game.challenge_num[2] ),
    .C(\game.challenge_num[1] ),
    .A(\game.challenge_num[3] ),
    .Y(_0604_));
 sg13g2_nor2_2 _3132_ (.A(net393),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_nor2_2 _3133_ (.A(\game.state[3] ),
    .B(_1803_),
    .Y(_0606_));
 sg13g2_nand2_1 _3134_ (.Y(_0607_),
    .A(_1802_),
    .B(\game.state[2] ));
 sg13g2_nor3_1 _3135_ (.A(_1804_),
    .B(net384),
    .C(_0607_),
    .Y(_0608_));
 sg13g2_nand2_1 _3136_ (.Y(_0609_),
    .A(_0605_),
    .B(_0608_));
 sg13g2_nand2_2 _3137_ (.Y(_0610_),
    .A(net382),
    .B(net383));
 sg13g2_nand2_2 _3138_ (.Y(_0611_),
    .A(_0606_),
    .B(_0610_));
 sg13g2_nand2_1 _3139_ (.Y(_0612_),
    .A(_0590_),
    .B(_0611_));
 sg13g2_nand3_1 _3140_ (.B(net384),
    .C(_0606_),
    .A(_1804_),
    .Y(_0613_));
 sg13g2_nor2_1 _3141_ (.A(_0590_),
    .B(_0591_),
    .Y(_0614_));
 sg13g2_o21ai_1 _3142_ (.B1(_0613_),
    .Y(_0615_),
    .A1(_0590_),
    .A2(_0591_));
 sg13g2_nand2_1 _3143_ (.Y(_0616_),
    .A(net371),
    .B(_0611_));
 sg13g2_and3_2 _3144_ (.X(_0617_),
    .A(_0609_),
    .B(_0613_),
    .C(_0616_));
 sg13g2_nor3_2 _3145_ (.A(\game.state[3] ),
    .B(net381),
    .C(net384),
    .Y(_0618_));
 sg13g2_nand2_1 _3146_ (.Y(_0619_),
    .A(\game.challenge_num[1] ),
    .B(net393));
 sg13g2_nor3_1 _3147_ (.A(_1813_),
    .B(_0604_),
    .C(net372),
    .Y(_0620_));
 sg13g2_a21oi_1 _3148_ (.A1(_0600_),
    .A2(_0603_),
    .Y(_0621_),
    .B1(_0620_));
 sg13g2_o21ai_1 _3149_ (.B1(net430),
    .Y(_0622_),
    .A1(\display_value[4] ),
    .A2(net346));
 sg13g2_a21o_2 _3150_ (.A2(_0621_),
    .A1(_0617_),
    .B1(_0622_),
    .X(_0623_));
 sg13g2_inv_1 _3151_ (.Y(_0239_),
    .A(_0623_));
 sg13g2_and2_1 _3152_ (.A(\game.state[2] ),
    .B(net372),
    .X(_0624_));
 sg13g2_nand2_1 _3153_ (.Y(_0625_),
    .A(\game.state[2] ),
    .B(net372));
 sg13g2_nor2_1 _3154_ (.A(_0054_),
    .B(_0619_),
    .Y(_0626_));
 sg13g2_xor2_1 _3155_ (.B(_0619_),
    .A(_0054_),
    .X(_0627_));
 sg13g2_o21ai_1 _3156_ (.B1(net371),
    .Y(_0628_),
    .A1(net370),
    .A2(_0627_));
 sg13g2_a21oi_1 _3157_ (.A1(_0054_),
    .A2(net370),
    .Y(_0629_),
    .B1(_0628_));
 sg13g2_nor2_1 _3158_ (.A(_0086_),
    .B(_0404_),
    .Y(_0630_));
 sg13g2_xnor2_1 _3159_ (.Y(_0631_),
    .A(_0086_),
    .B(_0403_));
 sg13g2_a21oi_1 _3160_ (.A1(_0600_),
    .A2(_0631_),
    .Y(_0632_),
    .B1(_0629_));
 sg13g2_nand2b_1 _3161_ (.Y(_0633_),
    .B(_0617_),
    .A_N(_0632_));
 sg13g2_o21ai_1 _3162_ (.B1(_0633_),
    .Y(_0634_),
    .A1(_0057_),
    .A2(_0617_));
 sg13g2_nand2_1 _3163_ (.Y(_0635_),
    .A(net430),
    .B(_0634_));
 sg13g2_nand2_1 _3164_ (.Y(_0636_),
    .A(_0022_),
    .B(_0600_));
 sg13g2_nor2_1 _3165_ (.A(net393),
    .B(net372),
    .Y(_0637_));
 sg13g2_a21oi_1 _3166_ (.A1(net393),
    .A2(net370),
    .Y(_0638_),
    .B1(_0637_));
 sg13g2_nand3_1 _3167_ (.B(_0636_),
    .C(_0638_),
    .A(net346),
    .Y(_0639_));
 sg13g2_o21ai_1 _3168_ (.B1(_0639_),
    .Y(_0640_),
    .A1(\display_value[0] ),
    .A2(net346));
 sg13g2_inv_1 _3169_ (.Y(_0641_),
    .A(_0640_));
 sg13g2_nand2_1 _3170_ (.Y(_0235_),
    .A(net430),
    .B(_0640_));
 sg13g2_nand2_2 _3171_ (.Y(_0642_),
    .A(_0404_),
    .B(_0481_));
 sg13g2_nor2_1 _3172_ (.A(\game.challenge_num[1] ),
    .B(net393),
    .Y(_0643_));
 sg13g2_xnor2_1 _3173_ (.Y(_0644_),
    .A(\game.challenge_num[1] ),
    .B(net393));
 sg13g2_a21oi_1 _3174_ (.A1(_0625_),
    .A2(_0644_),
    .Y(_0645_),
    .B1(net351));
 sg13g2_o21ai_1 _3175_ (.B1(_0645_),
    .Y(_0646_),
    .A1(_1890_),
    .A2(net369));
 sg13g2_o21ai_1 _3176_ (.B1(_0646_),
    .Y(_0647_),
    .A1(_0601_),
    .A2(_0642_));
 sg13g2_mux2_1 _3177_ (.A0(\display_value[1] ),
    .A1(_0647_),
    .S(net346),
    .X(_0648_));
 sg13g2_or2_2 _3178_ (.X(_0649_),
    .B(_0648_),
    .A(_0235_));
 sg13g2_nand2b_2 _3179_ (.Y(_0650_),
    .B(_0649_),
    .A_N(_0635_));
 sg13g2_xor2_1 _3180_ (.B(_0626_),
    .A(_0055_),
    .X(_0651_));
 sg13g2_or2_1 _3181_ (.X(_0652_),
    .B(_0651_),
    .A(net372));
 sg13g2_xnor2_1 _3182_ (.Y(_0653_),
    .A(net773),
    .B(_0630_));
 sg13g2_nand2_1 _3183_ (.Y(_0654_),
    .A(_0600_),
    .B(_0653_));
 sg13g2_nand2b_1 _3184_ (.Y(_0655_),
    .B(net370),
    .A_N(_0055_));
 sg13g2_and3_1 _3185_ (.X(_0656_),
    .A(net346),
    .B(_0652_),
    .C(_0654_));
 sg13g2_nor2_1 _3186_ (.A(net386),
    .B(net346),
    .Y(_0657_));
 sg13g2_a21oi_2 _3187_ (.B1(_0657_),
    .Y(_0658_),
    .A2(_0656_),
    .A1(_0655_));
 sg13g2_nand2_1 _3188_ (.Y(_0659_),
    .A(net430),
    .B(_0658_));
 sg13g2_inv_1 _3189_ (.Y(_0238_),
    .A(_0659_));
 sg13g2_a21oi_1 _3190_ (.A1(_0650_),
    .A2(_0659_),
    .Y(_0660_),
    .B1(_0623_));
 sg13g2_nand2_1 _3191_ (.Y(_0661_),
    .A(net430),
    .B(_0648_));
 sg13g2_inv_1 _3192_ (.Y(_0236_),
    .A(_0661_));
 sg13g2_nor2_1 _3193_ (.A(_0641_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_and2_1 _3194_ (.A(_0235_),
    .B(_0648_),
    .X(_0663_));
 sg13g2_a22oi_1 _3195_ (.Y(_0664_),
    .B1(_0663_),
    .B2(_0635_),
    .A2(_0662_),
    .A1(_0634_));
 sg13g2_nand2_1 _3196_ (.Y(_0665_),
    .A(_0238_),
    .B(_0664_));
 sg13g2_nand2_1 _3197_ (.Y(_0666_),
    .A(_0623_),
    .B(_0238_));
 sg13g2_nor2_2 _3198_ (.A(_0634_),
    .B(_0661_),
    .Y(_0667_));
 sg13g2_inv_1 _3199_ (.Y(_0668_),
    .A(_0667_));
 sg13g2_nand3_1 _3200_ (.B(_0650_),
    .C(_0668_),
    .A(_0623_),
    .Y(_0669_));
 sg13g2_nand2_1 _3201_ (.Y(_0670_),
    .A(_0666_),
    .B(_0669_));
 sg13g2_a21oi_1 _3202_ (.A1(_0665_),
    .A2(_0670_),
    .Y(_0000_),
    .B1(_0660_));
 sg13g2_nor2_1 _3203_ (.A(_0650_),
    .B(_0663_),
    .Y(_0671_));
 sg13g2_inv_1 _3204_ (.Y(_0672_),
    .A(_0671_));
 sg13g2_o21ai_1 _3205_ (.B1(_0672_),
    .Y(_0673_),
    .A1(_0634_),
    .A2(_0649_));
 sg13g2_nor2b_1 _3206_ (.A(_0635_),
    .B_N(_0658_),
    .Y(_0674_));
 sg13g2_a221oi_1 _3207_ (.B2(_0663_),
    .C1(_0660_),
    .B1(_0674_),
    .A1(_0659_),
    .Y(_0001_),
    .A2(_0673_));
 sg13g2_nand2b_1 _3208_ (.Y(_0675_),
    .B(_0239_),
    .A_N(_0658_));
 sg13g2_nand2b_1 _3209_ (.Y(_0676_),
    .B(_0650_),
    .A_N(_0675_));
 sg13g2_or2_1 _3210_ (.X(_0677_),
    .B(_0235_),
    .A(_0634_));
 sg13g2_nand3b_1 _3211_ (.B(_0658_),
    .C(_0634_),
    .Y(_0678_),
    .A_N(_0649_));
 sg13g2_o21ai_1 _3212_ (.B1(_0678_),
    .Y(_0679_),
    .A1(_0658_),
    .A2(_0677_));
 sg13g2_o21ai_1 _3213_ (.B1(_0676_),
    .Y(_0002_),
    .A1(_0239_),
    .A2(_0679_));
 sg13g2_a21oi_1 _3214_ (.A1(_0649_),
    .A2(_0668_),
    .Y(_0680_),
    .B1(_0675_));
 sg13g2_o21ai_1 _3215_ (.B1(_0659_),
    .Y(_0681_),
    .A1(_0667_),
    .A2(_0671_));
 sg13g2_a21oi_1 _3216_ (.A1(_0665_),
    .A2(_0681_),
    .Y(_0682_),
    .B1(_0239_));
 sg13g2_or2_1 _3217_ (.X(_0003_),
    .B(_0682_),
    .A(_0680_));
 sg13g2_a22oi_1 _3218_ (.Y(_0683_),
    .B1(_0677_),
    .B2(_0649_),
    .A2(_0675_),
    .A1(_0666_));
 sg13g2_nor2_1 _3219_ (.A(_0239_),
    .B(_0658_),
    .Y(_0684_));
 sg13g2_a21o_1 _3220_ (.A2(_0684_),
    .A1(_0662_),
    .B1(_0683_),
    .X(_0004_));
 sg13g2_a21oi_1 _3221_ (.A1(_0641_),
    .A2(_0648_),
    .Y(_0685_),
    .B1(_0635_));
 sg13g2_xnor2_1 _3222_ (.Y(_0686_),
    .A(_0665_),
    .B(_0685_));
 sg13g2_a21o_1 _3223_ (.A2(_0686_),
    .A1(_0623_),
    .B1(_0680_),
    .X(_0005_));
 sg13g2_a21oi_1 _3224_ (.A1(_0668_),
    .A2(_0677_),
    .Y(_0687_),
    .B1(_0675_));
 sg13g2_nor3_1 _3225_ (.A(_0238_),
    .B(_0667_),
    .C(_0685_),
    .Y(_0688_));
 sg13g2_a21oi_1 _3226_ (.A1(_0238_),
    .A2(_0667_),
    .Y(_0689_),
    .B1(_0688_));
 sg13g2_a21o_1 _3227_ (.A2(_0689_),
    .A1(_0623_),
    .B1(_0687_),
    .X(_0006_));
 sg13g2_and3_1 _3228_ (.X(_0010_),
    .A(net682),
    .B(_1899_),
    .C(_0585_));
 sg13g2_xor2_1 _3229_ (.B(net440),
    .A(\dsp.digit ),
    .X(uo_out[5]));
 sg13g2_xor2_1 _3230_ (.B(\dsp.digit_sel_raw[1] ),
    .A(net440),
    .X(uo_out[6]));
 sg13g2_xor2_1 _3231_ (.B(\dsp.segments_raw[0] ),
    .A(net440),
    .X(uio_out[0]));
 sg13g2_xor2_1 _3232_ (.B(\dsp.segments_raw[1] ),
    .A(net440),
    .X(uio_out[1]));
 sg13g2_xor2_1 _3233_ (.B(\dsp.segments_raw[2] ),
    .A(net440),
    .X(uio_out[2]));
 sg13g2_xor2_1 _3234_ (.B(\dsp.segments_raw[3] ),
    .A(net440),
    .X(uio_out[3]));
 sg13g2_xor2_1 _3235_ (.B(\dsp.segments_raw[4] ),
    .A(net5),
    .X(uio_out[4]));
 sg13g2_xor2_1 _3236_ (.B(\dsp.segments_raw[5] ),
    .A(net440),
    .X(uio_out[5]));
 sg13g2_xor2_1 _3237_ (.B(\dsp.segments_raw[6] ),
    .A(net440),
    .X(uio_out[6]));
 sg13g2_nor2b_1 _3238_ (.A(net389),
    .B_N(\game.input_color[1] ),
    .Y(_0690_));
 sg13g2_a21oi_2 _3239_ (.B1(_0690_),
    .Y(_0691_),
    .A2(\game.slv.fsm_color[1] ),
    .A1(net389));
 sg13g2_xnor2_1 _3240_ (.Y(_0692_),
    .A(net354),
    .B(_0691_));
 sg13g2_nor2b_1 _3241_ (.A(net389),
    .B_N(\game.input_color[0] ),
    .Y(_0693_));
 sg13g2_a21oi_2 _3242_ (.B1(_0693_),
    .Y(_0694_),
    .A2(\game.slv.fsm_color[0] ),
    .A1(net389));
 sg13g2_a21o_1 _3243_ (.A2(\game.slv.fsm_color[0] ),
    .A1(net389),
    .B1(_0693_),
    .X(_0695_));
 sg13g2_nor3_2 _3244_ (.A(net396),
    .B(net397),
    .C(net401),
    .Y(_0696_));
 sg13g2_xnor2_1 _3245_ (.Y(_0697_),
    .A(net353),
    .B(_0694_));
 sg13g2_nor3_2 _3246_ (.A(_0692_),
    .B(_0696_),
    .C(_0697_),
    .Y(_0698_));
 sg13g2_nor2b_1 _3247_ (.A(\game.solver_active ),
    .B_N(\game.input_reset ),
    .Y(_0699_));
 sg13g2_a21oi_1 _3248_ (.A1(\game.solver_active ),
    .A2(\game.slv.fsm_reset ),
    .Y(_0700_),
    .B1(_0699_));
 sg13g2_a21o_1 _3249_ (.A2(\game.slv.fsm_reset ),
    .A1(\game.solver_active ),
    .B1(_0699_),
    .X(_0701_));
 sg13g2_or2_2 _3250_ (.X(_0702_),
    .B(_0499_),
    .A(_0064_));
 sg13g2_mux2_1 _3251_ (.A0(\game.input_update ),
    .A1(\game.slv.fsm_update ),
    .S(net389),
    .X(_0703_));
 sg13g2_and2_1 _3252_ (.A(_0702_),
    .B(_0703_),
    .X(_0704_));
 sg13g2_nand2_1 _3253_ (.Y(_0705_),
    .A(_0702_),
    .B(_0703_));
 sg13g2_nor2_1 _3254_ (.A(net355),
    .B(net348),
    .Y(_0706_));
 sg13g2_nand2_2 _3255_ (.Y(_0707_),
    .A(net365),
    .B(_0704_));
 sg13g2_nand2_1 _3256_ (.Y(_0708_),
    .A(_0698_),
    .B(net349));
 sg13g2_inv_1 _3257_ (.Y(_0709_),
    .A(_0708_));
 sg13g2_nor2_1 _3258_ (.A(net356),
    .B(_0708_),
    .Y(_0710_));
 sg13g2_nand2_2 _3259_ (.Y(_0711_),
    .A(_0698_),
    .B(net347));
 sg13g2_nor2_2 _3260_ (.A(net373),
    .B(_1945_),
    .Y(_0712_));
 sg13g2_or2_1 _3261_ (.X(_0713_),
    .B(_1945_),
    .A(_1911_));
 sg13g2_mux2_1 _3262_ (.A0(_0072_),
    .A1(_0073_),
    .S(net395),
    .X(_0714_));
 sg13g2_nand2_1 _3263_ (.Y(_0715_),
    .A(_0712_),
    .B(_0714_));
 sg13g2_xnor2_1 _3264_ (.Y(_0716_),
    .A(_0069_),
    .B(_1945_));
 sg13g2_xnor2_1 _3265_ (.Y(_0717_),
    .A(_1845_),
    .B(_1945_));
 sg13g2_a221oi_1 _3266_ (.B2(_0074_),
    .C1(_0716_),
    .B1(_1945_),
    .A1(_0075_),
    .Y(_0718_),
    .A2(net373));
 sg13g2_nand2_1 _3267_ (.Y(_0719_),
    .A(net394),
    .B(_0077_));
 sg13g2_o21ai_1 _3268_ (.B1(_0719_),
    .Y(_0720_),
    .A1(net394),
    .A2(_1856_));
 sg13g2_nor2_1 _3269_ (.A(_1845_),
    .B(\game.fsm.block_len[7][2] ),
    .Y(_0721_));
 sg13g2_a221oi_1 _3270_ (.B2(_0720_),
    .C1(_0721_),
    .B1(_0712_),
    .A1(_1829_),
    .Y(_0722_),
    .A2(net373));
 sg13g2_a22oi_1 _3271_ (.Y(_0723_),
    .B1(_0722_),
    .B2(_0716_),
    .A2(_0718_),
    .A1(_0715_));
 sg13g2_nand2_1 _3272_ (.Y(_0724_),
    .A(net395),
    .B(\game.fsm.block_len[0][1] ));
 sg13g2_o21ai_1 _3273_ (.B1(_0724_),
    .Y(_0725_),
    .A1(net395),
    .A2(_1849_));
 sg13g2_nand2_1 _3274_ (.Y(_0726_),
    .A(_0712_),
    .B(_0725_));
 sg13g2_a221oi_1 _3275_ (.B2(\game.fsm.block_len[3][1] ),
    .C1(_0716_),
    .B1(_1945_),
    .A1(\game.fsm.block_len[2][1] ),
    .Y(_0727_),
    .A2(_1911_));
 sg13g2_mux2_1 _3276_ (.A0(\game.fsm.block_len[5][1] ),
    .A1(\game.fsm.block_len[4][1] ),
    .S(net394),
    .X(_0728_));
 sg13g2_a21oi_1 _3277_ (.A1(\game.fsm.block_len[6][1] ),
    .A2(net373),
    .Y(_0729_),
    .B1(_0717_));
 sg13g2_a22oi_1 _3278_ (.Y(_0730_),
    .B1(_0712_),
    .B2(_0728_),
    .A2(\game.fsm.block_len[7][1] ),
    .A1(_0069_));
 sg13g2_a22oi_1 _3279_ (.Y(_0731_),
    .B1(_0729_),
    .B2(_0730_),
    .A2(_0727_),
    .A1(_0726_));
 sg13g2_mux2_1 _3280_ (.A0(_0065_),
    .A1(_0066_),
    .S(net395),
    .X(_0732_));
 sg13g2_a21oi_1 _3281_ (.A1(_0068_),
    .A2(_1911_),
    .Y(_0733_),
    .B1(_0716_));
 sg13g2_a22oi_1 _3282_ (.Y(_0734_),
    .B1(_0712_),
    .B2(_0732_),
    .A2(_1945_),
    .A1(_0067_));
 sg13g2_mux2_1 _3283_ (.A0(_0070_),
    .A1(_0071_),
    .S(net394),
    .X(_0735_));
 sg13g2_nand2_1 _3284_ (.Y(_0736_),
    .A(_1830_),
    .B(net373));
 sg13g2_a221oi_1 _3285_ (.B2(_0735_),
    .C1(_0717_),
    .B1(_0712_),
    .A1(_0069_),
    .Y(_0737_),
    .A2(_1848_));
 sg13g2_a22oi_1 _3286_ (.Y(_0738_),
    .B1(_0736_),
    .B2(_0737_),
    .A2(_0734_),
    .A1(_0733_));
 sg13g2_inv_2 _3287_ (.Y(_0739_),
    .A(_0738_));
 sg13g2_xnor2_1 _3288_ (.Y(_0740_),
    .A(_0731_),
    .B(_0738_));
 sg13g2_nand2_2 _3289_ (.Y(_0741_),
    .A(_0723_),
    .B(_0740_));
 sg13g2_nor2_2 _3290_ (.A(_0711_),
    .B(_0741_),
    .Y(_0742_));
 sg13g2_nor3_2 _3291_ (.A(net389),
    .B(_1858_),
    .C(_0696_),
    .Y(_0743_));
 sg13g2_nand2_2 _3292_ (.Y(_0744_),
    .A(_0705_),
    .B(_0743_));
 sg13g2_nor2_1 _3293_ (.A(net355),
    .B(_0744_),
    .Y(_0745_));
 sg13g2_nand3_1 _3294_ (.B(_0705_),
    .C(_0743_),
    .A(net368),
    .Y(_0746_));
 sg13g2_and2_1 _3295_ (.A(_0723_),
    .B(_0731_),
    .X(_0747_));
 sg13g2_inv_1 _3296_ (.Y(_0748_),
    .A(_0747_));
 sg13g2_nor2_2 _3297_ (.A(_0746_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_nor2_1 _3298_ (.A(_0742_),
    .B(_0749_),
    .Y(_0750_));
 sg13g2_o21ai_1 _3299_ (.B1(_0510_),
    .Y(_0751_),
    .A1(_0742_),
    .A2(_0749_));
 sg13g2_o21ai_1 _3300_ (.B1(_0520_),
    .Y(_0752_),
    .A1(_0742_),
    .A2(_0749_));
 sg13g2_nor2_1 _3301_ (.A(net352),
    .B(_0751_),
    .Y(_0753_));
 sg13g2_o21ai_1 _3302_ (.B1(net367),
    .Y(_0754_),
    .A1(net507),
    .A2(_0753_));
 sg13g2_a21oi_1 _3303_ (.A1(net507),
    .A2(_0753_),
    .Y(_0093_),
    .B1(_0754_));
 sg13g2_nor2_1 _3304_ (.A(net357),
    .B(_0753_),
    .Y(_0755_));
 sg13g2_mux4_1 _3305_ (.S0(net354),
    .A0(\game.fsm.len2_color_count[0][0] ),
    .A1(\game.fsm.len2_color_count[2][0] ),
    .A2(\game.fsm.len2_color_count[1][0] ),
    .A3(\game.fsm.len2_color_count[3][0] ),
    .S1(net352),
    .X(_0756_));
 sg13g2_mux4_1 _3306_ (.S0(_0509_),
    .A0(_0045_),
    .A1(_0047_),
    .A2(_0046_),
    .A3(_0048_),
    .S1(net352),
    .X(_0757_));
 sg13g2_xor2_1 _3307_ (.B(_0757_),
    .A(_0756_),
    .X(_0758_));
 sg13g2_nor2_2 _3308_ (.A(_0739_),
    .B(_0748_),
    .Y(_0759_));
 sg13g2_xnor2_1 _3309_ (.Y(_0760_),
    .A(_0758_),
    .B(_0759_));
 sg13g2_nand3_1 _3310_ (.B(_0749_),
    .C(_0758_),
    .A(_0738_),
    .Y(_0761_));
 sg13g2_nand2_1 _3311_ (.Y(_0762_),
    .A(_0739_),
    .B(_0749_));
 sg13g2_nand2_1 _3312_ (.Y(_0763_),
    .A(_0745_),
    .B(_0759_));
 sg13g2_o21ai_1 _3313_ (.B1(_0761_),
    .Y(_0764_),
    .A1(_0758_),
    .A2(_0762_));
 sg13g2_a21o_2 _3314_ (.A2(_0760_),
    .A1(_0742_),
    .B1(_0764_),
    .X(_0765_));
 sg13g2_mux2_1 _3315_ (.A0(_0765_),
    .A1(net599),
    .S(_0755_),
    .X(_0094_));
 sg13g2_xnor2_1 _3316_ (.Y(_0766_),
    .A(net458),
    .B(net627));
 sg13g2_nand2_1 _3317_ (.Y(_0095_),
    .A(net424),
    .B(_0766_));
 sg13g2_xnor2_1 _3318_ (.Y(_0767_),
    .A(net466),
    .B(net709));
 sg13g2_nand2_1 _3319_ (.Y(_0096_),
    .A(net422),
    .B(_0767_));
 sg13g2_nand2b_1 _3320_ (.Y(_0768_),
    .B(\game.slv.lfsr[18] ),
    .A_N(net605));
 sg13g2_nand2b_1 _3321_ (.Y(_0769_),
    .B(net605),
    .A_N(\game.slv.lfsr[18] ));
 sg13g2_nand3_1 _3322_ (.B(_0768_),
    .C(net606),
    .A(net422),
    .Y(_0097_));
 sg13g2_nand2b_1 _3323_ (.Y(_0098_),
    .B(net425),
    .A_N(net756));
 sg13g2_nand2b_1 _3324_ (.Y(_0099_),
    .B(net426),
    .A_N(net489));
 sg13g2_nand2b_1 _3325_ (.Y(_0100_),
    .B(net422),
    .A_N(net716));
 sg13g2_nand2b_1 _3326_ (.Y(_0101_),
    .B(net424),
    .A_N(net449));
 sg13g2_nand2b_1 _3327_ (.Y(_0102_),
    .B(net426),
    .A_N(net445));
 sg13g2_nand2b_1 _3328_ (.Y(_0103_),
    .B(net422),
    .A_N(net324));
 sg13g2_nand2b_1 _3329_ (.Y(_0104_),
    .B(net425),
    .A_N(net453));
 sg13g2_nand2b_1 _3330_ (.Y(_0105_),
    .B(net422),
    .A_N(net467));
 sg13g2_nand2b_1 _3331_ (.Y(_0106_),
    .B(net422),
    .A_N(net450));
 sg13g2_nand2b_1 _3332_ (.Y(_0107_),
    .B(net425),
    .A_N(net321));
 sg13g2_nand2b_1 _3333_ (.Y(_0108_),
    .B(net422),
    .A_N(net325));
 sg13g2_nand2b_1 _3334_ (.Y(_0109_),
    .B(net423),
    .A_N(net447));
 sg13g2_nand2b_1 _3335_ (.Y(_0110_),
    .B(net424),
    .A_N(net451));
 sg13g2_nand2b_1 _3336_ (.Y(_0111_),
    .B(net422),
    .A_N(net444));
 sg13g2_nand2b_1 _3337_ (.Y(_0112_),
    .B(net423),
    .A_N(net446));
 sg13g2_nand2b_1 _3338_ (.Y(_0113_),
    .B(net424),
    .A_N(net448));
 sg13g2_nand2b_1 _3339_ (.Y(_0114_),
    .B(net423),
    .A_N(net458));
 sg13g2_nand2b_1 _3340_ (.Y(_0115_),
    .B(net423),
    .A_N(net466));
 sg13g2_nor2_1 _3341_ (.A(_1832_),
    .B(\snd.counter[7] ),
    .Y(_0770_));
 sg13g2_nand2_1 _3342_ (.Y(_0771_),
    .A(_1836_),
    .B(\snd.counter[3] ));
 sg13g2_nor2_1 _3343_ (.A(_1839_),
    .B(\snd.counter[0] ),
    .Y(_0772_));
 sg13g2_o21ai_1 _3344_ (.B1(_0772_),
    .Y(_0773_),
    .A1(\snd.note_timing[1] ),
    .A2(_1889_));
 sg13g2_a22oi_1 _3345_ (.Y(_0774_),
    .B1(_1889_),
    .B2(\snd.note_timing[1] ),
    .A2(_1888_),
    .A1(\snd.note_timing[2] ));
 sg13g2_a22oi_1 _3346_ (.Y(_0775_),
    .B1(_0773_),
    .B2(_0774_),
    .A2(\snd.counter[2] ),
    .A1(_1837_));
 sg13g2_nor2_1 _3347_ (.A(_1836_),
    .B(\snd.counter[3] ),
    .Y(_0776_));
 sg13g2_a221oi_1 _3348_ (.B2(_0775_),
    .C1(_0776_),
    .B1(_0771_),
    .A1(\snd.note_timing[4] ),
    .Y(_0777_),
    .A2(_1887_));
 sg13g2_a221oi_1 _3349_ (.B2(_1835_),
    .C1(_0777_),
    .B1(\snd.counter[4] ),
    .A1(_1834_),
    .Y(_0778_),
    .A2(\snd.counter[5] ));
 sg13g2_a221oi_1 _3350_ (.B2(\snd.note_timing[5] ),
    .C1(_0778_),
    .B1(_1886_),
    .A1(\snd.note_timing[6] ),
    .Y(_0779_),
    .A2(_1885_));
 sg13g2_a21oi_1 _3351_ (.A1(_1833_),
    .A2(\snd.counter[6] ),
    .Y(_0780_),
    .B1(_0779_));
 sg13g2_a22oi_1 _3352_ (.Y(_0781_),
    .B1(\snd.counter[8] ),
    .B2(_1831_),
    .A2(\snd.counter[7] ),
    .A1(_1832_));
 sg13g2_o21ai_1 _3353_ (.B1(_0781_),
    .Y(_0782_),
    .A1(_0770_),
    .A2(_0780_));
 sg13g2_o21ai_1 _3354_ (.B1(_0782_),
    .Y(_0783_),
    .A1(_1831_),
    .A2(\snd.counter[8] ));
 sg13g2_o21ai_1 _3355_ (.B1(net437),
    .Y(_0784_),
    .A1(net476),
    .A2(net337));
 sg13g2_a21oi_1 _3356_ (.A1(_1841_),
    .A2(net337),
    .Y(_0116_),
    .B1(_0784_));
 sg13g2_o21ai_1 _3357_ (.B1(net437),
    .Y(_0785_),
    .A1(net564),
    .A2(net337));
 sg13g2_a21oi_1 _3358_ (.A1(_1840_),
    .A2(net337),
    .Y(_0117_),
    .B1(_0785_));
 sg13g2_nand2_1 _3359_ (.Y(_0786_),
    .A(_0501_),
    .B(net345));
 sg13g2_a22oi_1 _3360_ (.Y(_0787_),
    .B1(net345),
    .B2(_0501_),
    .A2(net347),
    .A1(_1859_));
 sg13g2_a22oi_1 _3361_ (.Y(_0788_),
    .B1(net345),
    .B2(_0504_),
    .A2(net347),
    .A1(_1820_));
 sg13g2_nor2_1 _3362_ (.A(net401),
    .B(_0707_),
    .Y(_0789_));
 sg13g2_a21oi_2 _3363_ (.B1(_0789_),
    .Y(_0790_),
    .A2(net345),
    .A1(net400));
 sg13g2_inv_1 _3364_ (.Y(_0791_),
    .A(_0790_));
 sg13g2_nand3_1 _3365_ (.B(_0788_),
    .C(_0791_),
    .A(_0787_),
    .Y(_0792_));
 sg13g2_nand3_1 _3366_ (.B(net363),
    .C(_0792_),
    .A(net717),
    .Y(_0793_));
 sg13g2_nand2_1 _3367_ (.Y(_0794_),
    .A(_0695_),
    .B(_0706_));
 sg13g2_o21ai_1 _3368_ (.B1(_0793_),
    .Y(_0118_),
    .A1(_0792_),
    .A2(net344));
 sg13g2_nand3_1 _3369_ (.B(net362),
    .C(_0792_),
    .A(net744),
    .Y(_0795_));
 sg13g2_nand2b_1 _3370_ (.Y(_0796_),
    .B(net347),
    .A_N(_0691_));
 sg13g2_o21ai_1 _3371_ (.B1(_0795_),
    .Y(_0119_),
    .A1(_0792_),
    .A2(net343));
 sg13g2_o21ai_1 _3372_ (.B1(net434),
    .Y(_0797_),
    .A1(\snd.next_note_timing[0] ),
    .A2(net335));
 sg13g2_a21oi_1 _3373_ (.A1(_1839_),
    .A2(net335),
    .Y(_0120_),
    .B1(_0797_));
 sg13g2_o21ai_1 _3374_ (.B1(net434),
    .Y(_0798_),
    .A1(net504),
    .A2(net335));
 sg13g2_a21oi_1 _3375_ (.A1(_1838_),
    .A2(net335),
    .Y(_0121_),
    .B1(_0798_));
 sg13g2_o21ai_1 _3376_ (.B1(net434),
    .Y(_0799_),
    .A1(net554),
    .A2(_0783_));
 sg13g2_a21oi_1 _3377_ (.A1(_1837_),
    .A2(net335),
    .Y(_0122_),
    .B1(_0799_));
 sg13g2_o21ai_1 _3378_ (.B1(net434),
    .Y(_0800_),
    .A1(net509),
    .A2(net335));
 sg13g2_a21oi_1 _3379_ (.A1(_1836_),
    .A2(net335),
    .Y(_0123_),
    .B1(_0800_));
 sg13g2_o21ai_1 _3380_ (.B1(net437),
    .Y(_0801_),
    .A1(net492),
    .A2(net336));
 sg13g2_a21oi_1 _3381_ (.A1(_1835_),
    .A2(net336),
    .Y(_0124_),
    .B1(_0801_));
 sg13g2_o21ai_1 _3382_ (.B1(net437),
    .Y(_0802_),
    .A1(net488),
    .A2(net336));
 sg13g2_a21oi_1 _3383_ (.A1(_1834_),
    .A2(net337),
    .Y(_0125_),
    .B1(_0802_));
 sg13g2_o21ai_1 _3384_ (.B1(net438),
    .Y(_0803_),
    .A1(\snd.next_note_timing[6] ),
    .A2(net336));
 sg13g2_a21oi_1 _3385_ (.A1(_1833_),
    .A2(net336),
    .Y(_0126_),
    .B1(_0803_));
 sg13g2_o21ai_1 _3386_ (.B1(net438),
    .Y(_0804_),
    .A1(net538),
    .A2(net337));
 sg13g2_a21oi_1 _3387_ (.A1(_1832_),
    .A2(net336),
    .Y(_0127_),
    .B1(_0804_));
 sg13g2_o21ai_1 _3388_ (.B1(net438),
    .Y(_0805_),
    .A1(net519),
    .A2(net337));
 sg13g2_a21oi_1 _3389_ (.A1(_1831_),
    .A2(net336),
    .Y(_0128_),
    .B1(_0805_));
 sg13g2_nor2_2 _3390_ (.A(net349),
    .B(_0743_),
    .Y(_0806_));
 sg13g2_nand2_2 _3391_ (.Y(_0807_),
    .A(net365),
    .B(_0806_));
 sg13g2_inv_1 _3392_ (.Y(_0808_),
    .A(_0807_));
 sg13g2_nand4_1 _3393_ (.B(_0788_),
    .C(_0790_),
    .A(_0787_),
    .Y(_0809_),
    .D(_0807_));
 sg13g2_nand2_1 _3394_ (.Y(_0810_),
    .A(net632),
    .B(_0809_));
 sg13g2_o21ai_1 _3395_ (.B1(_0810_),
    .Y(_0129_),
    .A1(net344),
    .A2(_0809_));
 sg13g2_nand2_1 _3396_ (.Y(_0811_),
    .A(net640),
    .B(_0809_));
 sg13g2_o21ai_1 _3397_ (.B1(_0811_),
    .Y(_0130_),
    .A1(net343),
    .A2(_0809_));
 sg13g2_nor2_1 _3398_ (.A(_0698_),
    .B(net348),
    .Y(_0812_));
 sg13g2_inv_1 _3399_ (.Y(_0813_),
    .A(_0812_));
 sg13g2_nor2_2 _3400_ (.A(_0698_),
    .B(_0707_),
    .Y(_0814_));
 sg13g2_nand2_2 _3401_ (.Y(_0815_),
    .A(_0711_),
    .B(_0746_));
 sg13g2_a22oi_1 _3402_ (.Y(_0816_),
    .B1(_0815_),
    .B2(_0713_),
    .A2(net341),
    .A1(\game.fsm.num_blocks[1] ));
 sg13g2_a22oi_1 _3403_ (.Y(_0817_),
    .B1(_0815_),
    .B2(_0717_),
    .A2(net341),
    .A1(_1818_));
 sg13g2_nand2_1 _3404_ (.Y(_0818_),
    .A(_0816_),
    .B(_0817_));
 sg13g2_mux2_2 _3405_ (.A0(net341),
    .A1(_0815_),
    .S(net394),
    .X(_0819_));
 sg13g2_nand2b_2 _3406_ (.Y(_0820_),
    .B(_0807_),
    .A_N(_0819_));
 sg13g2_nor2_2 _3407_ (.A(_0818_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_a21oi_2 _3408_ (.B1(net341),
    .Y(_0822_),
    .A2(_0815_),
    .A1(_0738_));
 sg13g2_a21o_1 _3409_ (.A2(_0815_),
    .A1(_0738_),
    .B1(net341),
    .X(_0823_));
 sg13g2_nor2_1 _3410_ (.A(net588),
    .B(_0821_),
    .Y(_0824_));
 sg13g2_a21oi_1 _3411_ (.A1(_0821_),
    .A2(_0822_),
    .Y(_0131_),
    .B1(_0824_));
 sg13g2_nor2_1 _3412_ (.A(net566),
    .B(_0821_),
    .Y(_0825_));
 sg13g2_xnor2_1 _3413_ (.Y(_0826_),
    .A(net349),
    .B(_0740_));
 sg13g2_nand2_2 _3414_ (.Y(_0827_),
    .A(_0815_),
    .B(_0826_));
 sg13g2_a21oi_1 _3415_ (.A1(_0821_),
    .A2(_0827_),
    .Y(_0132_),
    .B1(_0825_));
 sg13g2_nand2_2 _3416_ (.Y(_0828_),
    .A(_0710_),
    .B(_0747_));
 sg13g2_nor2_1 _3417_ (.A(_0738_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_nor3_1 _3418_ (.A(_0723_),
    .B(_0731_),
    .C(_0739_),
    .Y(_0830_));
 sg13g2_and2_1 _3419_ (.A(_0723_),
    .B(_0739_),
    .X(_0831_));
 sg13g2_nor4_1 _3420_ (.A(_0746_),
    .B(_0747_),
    .C(_0830_),
    .D(_0831_),
    .Y(_0832_));
 sg13g2_a21oi_1 _3421_ (.A1(_0731_),
    .A2(_0739_),
    .Y(_0833_),
    .B1(_0723_));
 sg13g2_nor2b_1 _3422_ (.A(_0711_),
    .B_N(_0833_),
    .Y(_0834_));
 sg13g2_nor3_2 _3423_ (.A(_0829_),
    .B(_0832_),
    .C(_0834_),
    .Y(_0835_));
 sg13g2_inv_1 _3424_ (.Y(_0836_),
    .A(_0835_));
 sg13g2_nor2_1 _3425_ (.A(net468),
    .B(_0821_),
    .Y(_0837_));
 sg13g2_a21oi_1 _3426_ (.A1(_0821_),
    .A2(_0835_),
    .Y(_0133_),
    .B1(_0837_));
 sg13g2_nand2b_1 _3427_ (.Y(_0838_),
    .B(_0817_),
    .A_N(_0816_));
 sg13g2_nand2b_2 _3428_ (.Y(_0839_),
    .B(_0819_),
    .A_N(_0838_));
 sg13g2_o21ai_1 _3429_ (.B1(net360),
    .Y(_0840_),
    .A1(_0823_),
    .A2(_0839_));
 sg13g2_a21oi_1 _3430_ (.A1(_1830_),
    .A2(_0839_),
    .Y(_0134_),
    .B1(_0840_));
 sg13g2_nor2b_1 _3431_ (.A(net677),
    .B_N(_0839_),
    .Y(_0841_));
 sg13g2_nor2b_1 _3432_ (.A(_0839_),
    .B_N(_0827_),
    .Y(_0842_));
 sg13g2_nor3_1 _3433_ (.A(net355),
    .B(_0841_),
    .C(_0842_),
    .Y(_0135_));
 sg13g2_o21ai_1 _3434_ (.B1(net360),
    .Y(_0843_),
    .A1(_0836_),
    .A2(_0839_));
 sg13g2_a21oi_1 _3435_ (.A1(_1829_),
    .A2(_0839_),
    .Y(_0136_),
    .B1(_0843_));
 sg13g2_a22oi_1 _3436_ (.Y(_0844_),
    .B1(net345),
    .B2(_0510_),
    .A2(net347),
    .A1(_0691_));
 sg13g2_a22oi_1 _3437_ (.Y(_0845_),
    .B1(net345),
    .B2(_0520_),
    .A2(net347),
    .A1(_0694_));
 sg13g2_nor2_2 _3438_ (.A(_0844_),
    .B(_0845_),
    .Y(_0846_));
 sg13g2_o21ai_1 _3439_ (.B1(net362),
    .Y(_0847_),
    .A1(net410),
    .A2(_0846_));
 sg13g2_a21oi_1 _3440_ (.A1(net410),
    .A2(_0846_),
    .Y(_0137_),
    .B1(_0847_));
 sg13g2_nand2_1 _3441_ (.Y(_0848_),
    .A(net353),
    .B(_0707_));
 sg13g2_and2_2 _3442_ (.A(_0794_),
    .B(_0848_),
    .X(_0849_));
 sg13g2_o21ai_1 _3443_ (.B1(_0796_),
    .Y(_0850_),
    .A1(_0510_),
    .A2(net347));
 sg13g2_mux4_1 _3444_ (.S0(_0849_),
    .A0(\game.fsm.color_count[1][0] ),
    .A1(net410),
    .A2(\game.fsm.color_count[3][0] ),
    .A3(\game.fsm.color_count[2][0] ),
    .S1(_0850_),
    .X(_0851_));
 sg13g2_mux4_1 _3445_ (.S0(_0849_),
    .A0(\game.fsm.color_count[1][1] ),
    .A1(net409),
    .A2(\game.fsm.color_count[3][1] ),
    .A3(\game.fsm.color_count[2][1] ),
    .S1(_0850_),
    .X(_0852_));
 sg13g2_nand2_1 _3446_ (.Y(_0853_),
    .A(_0851_),
    .B(_0852_));
 sg13g2_nor2_1 _3447_ (.A(_0851_),
    .B(_0852_),
    .Y(_0854_));
 sg13g2_xnor2_1 _3448_ (.Y(_0855_),
    .A(_0851_),
    .B(_0852_));
 sg13g2_o21ai_1 _3449_ (.B1(net362),
    .Y(_0856_),
    .A1(_0744_),
    .A2(_0855_));
 sg13g2_a21oi_2 _3450_ (.B1(_0856_),
    .Y(_0857_),
    .A2(_0855_),
    .A1(_0744_));
 sg13g2_nor2_1 _3451_ (.A(net355),
    .B(_0846_),
    .Y(_0858_));
 sg13g2_a22oi_1 _3452_ (.Y(_0859_),
    .B1(_0858_),
    .B2(net409),
    .A2(_0857_),
    .A1(_0846_));
 sg13g2_inv_1 _3453_ (.Y(_0138_),
    .A(_0859_));
 sg13g2_mux4_1 _3454_ (.S0(_0849_),
    .A0(\game.fsm.color_count[1][2] ),
    .A1(\game.fsm.color_count[0][2] ),
    .A2(_1868_),
    .A3(_1872_),
    .S1(_0850_),
    .X(_0860_));
 sg13g2_xnor2_1 _3455_ (.Y(_0861_),
    .A(_0853_),
    .B(_0860_));
 sg13g2_nand2_1 _3456_ (.Y(_0862_),
    .A(net347),
    .B(_0861_));
 sg13g2_xnor2_1 _3457_ (.Y(_0863_),
    .A(_0854_),
    .B(_0860_));
 sg13g2_o21ai_1 _3458_ (.B1(_0862_),
    .Y(_0864_),
    .A1(_0746_),
    .A2(_0863_));
 sg13g2_nor2_1 _3459_ (.A(_0858_),
    .B(_0864_),
    .Y(_0865_));
 sg13g2_a21oi_1 _3460_ (.A1(_1865_),
    .A2(_0858_),
    .Y(_0139_),
    .B1(_0865_));
 sg13g2_nand2b_2 _3461_ (.Y(_0866_),
    .B(_0819_),
    .A_N(_0818_));
 sg13g2_nand3_1 _3462_ (.B(net359),
    .C(_0866_),
    .A(net608),
    .Y(_0867_));
 sg13g2_o21ai_1 _3463_ (.B1(_0867_),
    .Y(_0140_),
    .A1(_0822_),
    .A2(_0866_));
 sg13g2_nand3_1 _3464_ (.B(net359),
    .C(_0866_),
    .A(net636),
    .Y(_0868_));
 sg13g2_o21ai_1 _3465_ (.B1(_0868_),
    .Y(_0141_),
    .A1(_0827_),
    .A2(_0866_));
 sg13g2_nand3_1 _3466_ (.B(net359),
    .C(_0866_),
    .A(net622),
    .Y(_0869_));
 sg13g2_o21ai_1 _3467_ (.B1(_0869_),
    .Y(_0142_),
    .A1(_0835_),
    .A2(_0866_));
 sg13g2_or2_1 _3468_ (.X(_0870_),
    .B(_0817_),
    .A(_0816_));
 sg13g2_or2_2 _3469_ (.X(_0871_),
    .B(_0870_),
    .A(_0820_));
 sg13g2_nand3_1 _3470_ (.B(net359),
    .C(_0871_),
    .A(net483),
    .Y(_0872_));
 sg13g2_o21ai_1 _3471_ (.B1(_0872_),
    .Y(_0143_),
    .A1(_0822_),
    .A2(_0871_));
 sg13g2_nand3_1 _3472_ (.B(net360),
    .C(_0871_),
    .A(net502),
    .Y(_0873_));
 sg13g2_o21ai_1 _3473_ (.B1(_0873_),
    .Y(_0144_),
    .A1(_0827_),
    .A2(_0871_));
 sg13g2_nand3_1 _3474_ (.B(net359),
    .C(_0871_),
    .A(net558),
    .Y(_0874_));
 sg13g2_o21ai_1 _3475_ (.B1(_0874_),
    .Y(_0145_),
    .A1(_0835_),
    .A2(_0871_));
 sg13g2_nand2b_2 _3476_ (.Y(_0875_),
    .B(_0819_),
    .A_N(_0870_));
 sg13g2_nand3_1 _3477_ (.B(net359),
    .C(_0875_),
    .A(net572),
    .Y(_0876_));
 sg13g2_o21ai_1 _3478_ (.B1(_0876_),
    .Y(_0146_),
    .A1(_0822_),
    .A2(_0875_));
 sg13g2_nand3_1 _3479_ (.B(net359),
    .C(_0875_),
    .A(net560),
    .Y(_0877_));
 sg13g2_o21ai_1 _3480_ (.B1(_0877_),
    .Y(_0147_),
    .A1(_0827_),
    .A2(_0875_));
 sg13g2_nand3_1 _3481_ (.B(net359),
    .C(_0875_),
    .A(net529),
    .Y(_0878_));
 sg13g2_o21ai_1 _3482_ (.B1(_0878_),
    .Y(_0148_),
    .A1(_0835_),
    .A2(_0875_));
 sg13g2_nand2b_1 _3483_ (.Y(_0879_),
    .B(_0816_),
    .A_N(_0817_));
 sg13g2_or2_2 _3484_ (.X(_0880_),
    .B(_0879_),
    .A(_0820_));
 sg13g2_nand3_1 _3485_ (.B(net361),
    .C(_0880_),
    .A(net459),
    .Y(_0881_));
 sg13g2_o21ai_1 _3486_ (.B1(_0881_),
    .Y(_0149_),
    .A1(_0822_),
    .A2(_0880_));
 sg13g2_nand3_1 _3487_ (.B(net365),
    .C(_0880_),
    .A(net594),
    .Y(_0882_));
 sg13g2_o21ai_1 _3488_ (.B1(_0882_),
    .Y(_0150_),
    .A1(_0827_),
    .A2(_0880_));
 sg13g2_nand3_1 _3489_ (.B(net361),
    .C(_0880_),
    .A(net641),
    .Y(_0883_));
 sg13g2_o21ai_1 _3490_ (.B1(_0883_),
    .Y(_0151_),
    .A1(_0835_),
    .A2(_0880_));
 sg13g2_nand2b_1 _3491_ (.Y(_0884_),
    .B(\snd.tune_counter[2] ),
    .A_N(_0081_));
 sg13g2_nor2_1 _3492_ (.A(\snd.tune_counter[1] ),
    .B(\snd.tune_counter[0] ),
    .Y(_0885_));
 sg13g2_nand2_1 _3493_ (.Y(_0886_),
    .A(\snd.tune_counter[5] ),
    .B(_0885_));
 sg13g2_nor4_2 _3494_ (.A(\snd.tune_counter[4] ),
    .B(\snd.tune_counter[3] ),
    .C(_0884_),
    .Y(_0887_),
    .D(_0886_));
 sg13g2_nand2b_2 _3495_ (.Y(_0888_),
    .B(\snd.sequencer_state[1] ),
    .A_N(\snd.sequencer_state[0] ));
 sg13g2_or2_2 _3496_ (.X(_0889_),
    .B(_0888_),
    .A(_0887_));
 sg13g2_nor2_2 _3497_ (.A(_0080_),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_nand2_2 _3498_ (.Y(_0891_),
    .A(_1776_),
    .B(\snd.sequencer_state[0] ));
 sg13g2_o21ai_1 _3499_ (.B1(_0891_),
    .Y(_0892_),
    .A1(net408),
    .A2(_0888_));
 sg13g2_nor2_1 _3500_ (.A(_0890_),
    .B(_0892_),
    .Y(_0893_));
 sg13g2_o21ai_1 _3501_ (.B1(net581),
    .Y(_0894_),
    .A1(_0890_),
    .A2(_0892_));
 sg13g2_nor2_2 _3502_ (.A(\snd.sequencer_state[1] ),
    .B(\snd.sequencer_state[0] ),
    .Y(_0895_));
 sg13g2_nand2_1 _3503_ (.Y(_0896_),
    .A(net684),
    .B(_0895_));
 sg13g2_mux2_1 _3504_ (.A0(_0079_),
    .A1(_1807_),
    .S(\game.sound_mode[0] ),
    .X(_0897_));
 sg13g2_nor2b_2 _3505_ (.A(_0896_),
    .B_N(_0897_),
    .Y(_0898_));
 sg13g2_nand2_1 _3506_ (.Y(_0899_),
    .A(net670),
    .B(_0895_));
 sg13g2_nor2b_1 _3507_ (.A(\game.sound_mode[1] ),
    .B_N(_0079_),
    .Y(_0900_));
 sg13g2_a21oi_1 _3508_ (.A1(_1807_),
    .A2(\game.sound_mode[1] ),
    .Y(_0901_),
    .B1(_0900_));
 sg13g2_nor2_2 _3509_ (.A(_0899_),
    .B(_0901_),
    .Y(_0902_));
 sg13g2_a22oi_1 _3510_ (.Y(_0903_),
    .B1(_0902_),
    .B2(\btn.button_state[3] ),
    .A2(_0898_),
    .A1(uo_out[3]));
 sg13g2_a21oi_1 _3511_ (.A1(_0894_),
    .A2(_0903_),
    .Y(_0152_),
    .B1(net419));
 sg13g2_nand2_1 _3512_ (.Y(_0904_),
    .A(net438),
    .B(net336));
 sg13g2_xnor2_1 _3513_ (.Y(_0905_),
    .A(net647),
    .B(\snd.counter[0] ));
 sg13g2_nor2_1 _3514_ (.A(net334),
    .B(net648),
    .Y(_0153_));
 sg13g2_and3_1 _3515_ (.X(_0906_),
    .A(net591),
    .B(net647),
    .C(net651));
 sg13g2_a21oi_1 _3516_ (.A1(\snd.counter[1] ),
    .A2(\snd.counter[0] ),
    .Y(_0907_),
    .B1(net591));
 sg13g2_nor3_1 _3517_ (.A(net334),
    .B(_0906_),
    .C(net592),
    .Y(_0154_));
 sg13g2_and2_1 _3518_ (.A(net658),
    .B(_0906_),
    .X(_0908_));
 sg13g2_nor2_1 _3519_ (.A(net658),
    .B(_0906_),
    .Y(_0909_));
 sg13g2_nor3_1 _3520_ (.A(net334),
    .B(_0908_),
    .C(_0909_),
    .Y(_0155_));
 sg13g2_and2_1 _3521_ (.A(net645),
    .B(_0908_),
    .X(_0910_));
 sg13g2_nor2_1 _3522_ (.A(net645),
    .B(_0908_),
    .Y(_0911_));
 sg13g2_nor3_1 _3523_ (.A(_0904_),
    .B(_0910_),
    .C(net646),
    .Y(_0156_));
 sg13g2_and2_1 _3524_ (.A(net653),
    .B(_0910_),
    .X(_0912_));
 sg13g2_nor2_1 _3525_ (.A(net653),
    .B(_0910_),
    .Y(_0913_));
 sg13g2_nor3_1 _3526_ (.A(net334),
    .B(_0912_),
    .C(_0913_),
    .Y(_0157_));
 sg13g2_and2_1 _3527_ (.A(net602),
    .B(_0912_),
    .X(_0914_));
 sg13g2_nor2_1 _3528_ (.A(net602),
    .B(_0912_),
    .Y(_0915_));
 sg13g2_nor3_1 _3529_ (.A(net334),
    .B(_0914_),
    .C(net603),
    .Y(_0158_));
 sg13g2_nand2_1 _3530_ (.Y(_0916_),
    .A(\snd.counter[7] ),
    .B(_0914_));
 sg13g2_xnor2_1 _3531_ (.Y(_0917_),
    .A(net703),
    .B(_0914_));
 sg13g2_nor2_1 _3532_ (.A(net334),
    .B(_0917_),
    .Y(_0159_));
 sg13g2_xor2_1 _3533_ (.B(_0916_),
    .A(net690),
    .X(_0918_));
 sg13g2_nor2_1 _3534_ (.A(net334),
    .B(net691),
    .Y(_0160_));
 sg13g2_nand4_1 _3535_ (.B(net534),
    .C(net530),
    .A(net544),
    .Y(_0919_),
    .D(net604));
 sg13g2_nand2_1 _3536_ (.Y(_0920_),
    .A(net696),
    .B(net494));
 sg13g2_nor4_1 _3537_ (.A(net620),
    .B(net460),
    .C(_0919_),
    .D(_0920_),
    .Y(_0921_));
 sg13g2_and2_1 _3538_ (.A(net430),
    .B(_0921_),
    .X(_0161_));
 sg13g2_nand2_1 _3539_ (.Y(_0922_),
    .A(net382),
    .B(_0589_));
 sg13g2_nor2_2 _3540_ (.A(_0590_),
    .B(_0610_),
    .Y(_0923_));
 sg13g2_nand3_1 _3541_ (.B(net383),
    .C(_0589_),
    .A(net381),
    .Y(_0924_));
 sg13g2_and3_1 _3542_ (.X(_0162_),
    .A(net465),
    .B(net421),
    .C(_0923_));
 sg13g2_or4_1 _3543_ (.A(_1878_),
    .B(net402),
    .C(net751),
    .D(_0582_),
    .X(_0925_));
 sg13g2_a21oi_1 _3544_ (.A1(_0584_),
    .A2(net752),
    .Y(_0926_),
    .B1(net720));
 sg13g2_nand2b_1 _3545_ (.Y(_0163_),
    .B(net427),
    .A_N(_0926_));
 sg13g2_nor2b_2 _3546_ (.A(net402),
    .B_N(net682),
    .Y(_0927_));
 sg13g2_and3_1 _3547_ (.X(_0164_),
    .A(_1899_),
    .B(_0586_),
    .C(_0927_));
 sg13g2_and2_1 _3548_ (.A(net756),
    .B(_0164_),
    .X(_0165_));
 sg13g2_and2_1 _3549_ (.A(net489),
    .B(_0164_),
    .X(_0166_));
 sg13g2_nand2_1 _3550_ (.Y(_0928_),
    .A(net484),
    .B(_1899_));
 sg13g2_nor2_1 _3551_ (.A(\game.slv.target[1] ),
    .B(\game.slv.target[0] ),
    .Y(_0929_));
 sg13g2_nand2b_1 _3552_ (.Y(_0930_),
    .B(\game.slv.target[1] ),
    .A_N(\game.slv.lfsr[0] ));
 sg13g2_nand3_1 _3553_ (.B(net427),
    .C(_0930_),
    .A(\game.slv.trigger ),
    .Y(_0931_));
 sg13g2_o21ai_1 _3554_ (.B1(net485),
    .Y(_0167_),
    .A1(_0929_),
    .A2(_0931_));
 sg13g2_and3_1 _3555_ (.X(_0932_),
    .A(_0083_),
    .B(_1879_),
    .C(net481));
 sg13g2_nor2_2 _3556_ (.A(\game.slv.state[1] ),
    .B(net403),
    .Y(_0933_));
 sg13g2_nand2_1 _3557_ (.Y(_0934_),
    .A(_0039_),
    .B(_0933_));
 sg13g2_nand2_1 _3558_ (.Y(_0935_),
    .A(_1898_),
    .B(_0934_));
 sg13g2_a21oi_1 _3559_ (.A1(_0582_),
    .A2(_0932_),
    .Y(_0936_),
    .B1(_0935_));
 sg13g2_a221oi_1 _3560_ (.B2(_0932_),
    .C1(_0935_),
    .B1(_0582_),
    .A1(\game.slv.state[1] ),
    .Y(_0937_),
    .A2(_1879_));
 sg13g2_and2_1 _3561_ (.A(net402),
    .B(\game.slv.lfsr[0] ),
    .X(_0938_));
 sg13g2_nor2_1 _3562_ (.A(net656),
    .B(net662),
    .Y(_0939_));
 sg13g2_nor3_2 _3563_ (.A(net735),
    .B(net656),
    .C(\game.slv.retries[0] ),
    .Y(_0940_));
 sg13g2_inv_1 _3564_ (.Y(_0941_),
    .A(_0940_));
 sg13g2_a21oi_1 _3565_ (.A1(\game.slv.length[2] ),
    .A2(\game.slv.length[1] ),
    .Y(_0942_),
    .B1(_0941_));
 sg13g2_xor2_1 _3566_ (.B(_0942_),
    .A(net713),
    .X(_0943_));
 sg13g2_a21oi_1 _3567_ (.A1(_1879_),
    .A2(_0943_),
    .Y(_0944_),
    .B1(_0938_));
 sg13g2_o21ai_1 _3568_ (.B1(net424),
    .Y(_0945_),
    .A1(net713),
    .A2(net333));
 sg13g2_a21oi_1 _3569_ (.A1(net333),
    .A2(_0944_),
    .Y(_0168_),
    .B1(_0945_));
 sg13g2_and2_1 _3570_ (.A(net402),
    .B(net489),
    .X(_0946_));
 sg13g2_a21oi_1 _3571_ (.A1(net796),
    .A2(_0940_),
    .Y(_0947_),
    .B1(net652));
 sg13g2_and2_1 _3572_ (.A(\game.slv.length[1] ),
    .B(\game.slv.length[0] ),
    .X(_0948_));
 sg13g2_a21oi_1 _3573_ (.A1(_0942_),
    .A2(_0948_),
    .Y(_0949_),
    .B1(_0947_));
 sg13g2_a21oi_1 _3574_ (.A1(_1879_),
    .A2(_0949_),
    .Y(_0950_),
    .B1(_0946_));
 sg13g2_o21ai_1 _3575_ (.B1(net424),
    .Y(_0951_),
    .A1(net652),
    .A2(net333));
 sg13g2_a21oi_1 _3576_ (.A1(net333),
    .A2(_0950_),
    .Y(_0169_),
    .B1(_0951_));
 sg13g2_a21oi_1 _3577_ (.A1(_0940_),
    .A2(_0948_),
    .Y(_0952_),
    .B1(net618));
 sg13g2_nor2_1 _3578_ (.A(net403),
    .B(_0952_),
    .Y(_0953_));
 sg13g2_or2_1 _3579_ (.X(_0954_),
    .B(_0953_),
    .A(_0927_));
 sg13g2_a21oi_1 _3580_ (.A1(net403),
    .A2(\game.slv.lfsr[2] ),
    .Y(_0955_),
    .B1(_0953_));
 sg13g2_o21ai_1 _3581_ (.B1(net424),
    .Y(_0956_),
    .A1(net618),
    .A2(net333));
 sg13g2_a21oi_1 _3582_ (.A1(net333),
    .A2(_0955_),
    .Y(_0170_),
    .B1(_0956_));
 sg13g2_nor2_1 _3583_ (.A(_0083_),
    .B(net402),
    .Y(_0957_));
 sg13g2_a221oi_1 _3584_ (.B2(_0585_),
    .C1(_0935_),
    .B1(_0957_),
    .A1(_0582_),
    .Y(_0958_),
    .A2(_0932_));
 sg13g2_a221oi_1 _3585_ (.B2(_0943_),
    .C1(_0938_),
    .B1(_0933_),
    .A1(net672),
    .Y(_0959_),
    .A2(_0927_));
 sg13g2_o21ai_1 _3586_ (.B1(net426),
    .Y(_0960_),
    .A1(\game.slv.pos[0] ),
    .A2(_0958_));
 sg13g2_a21oi_1 _3587_ (.A1(_0958_),
    .A2(_0959_),
    .Y(_0171_),
    .B1(_0960_));
 sg13g2_xnor2_1 _3588_ (.Y(_0961_),
    .A(\game.slv.pos[1] ),
    .B(\game.slv.pos[0] ));
 sg13g2_a221oi_1 _3589_ (.B2(_0927_),
    .C1(_0946_),
    .B1(_0961_),
    .A1(_0933_),
    .Y(_0962_),
    .A2(_0949_));
 sg13g2_o21ai_1 _3590_ (.B1(net426),
    .Y(_0963_),
    .A1(net726),
    .A2(_0958_));
 sg13g2_a21oi_1 _3591_ (.A1(_0958_),
    .A2(_0962_),
    .Y(_0172_),
    .B1(_0963_));
 sg13g2_o21ai_1 _3592_ (.B1(net680),
    .Y(_0964_),
    .A1(\game.slv.pos[1] ),
    .A2(\game.slv.pos[0] ));
 sg13g2_nand3_1 _3593_ (.B(_0586_),
    .C(_0964_),
    .A(\game.slv.state[1] ),
    .Y(_0965_));
 sg13g2_a22oi_1 _3594_ (.Y(_0966_),
    .B1(_0954_),
    .B2(_0965_),
    .A2(\game.slv.lfsr[2] ),
    .A1(net402));
 sg13g2_o21ai_1 _3595_ (.B1(net426),
    .Y(_0967_),
    .A1(net680),
    .A2(_0958_));
 sg13g2_a21oi_1 _3596_ (.A1(_0958_),
    .A2(_0966_),
    .Y(_0173_),
    .B1(_0967_));
 sg13g2_o21ai_1 _3597_ (.B1(_0937_),
    .Y(_0968_),
    .A1(_1827_),
    .A2(net403));
 sg13g2_nand2b_1 _3598_ (.Y(_0969_),
    .B(net662),
    .A_N(_0937_));
 sg13g2_a21oi_1 _3599_ (.A1(_0968_),
    .A2(_0969_),
    .Y(_0174_),
    .B1(net412));
 sg13g2_nor4_1 _3600_ (.A(_1826_),
    .B(\game.slv.retries[0] ),
    .C(\game.slv.state[1] ),
    .D(net403),
    .Y(_0970_));
 sg13g2_a221oi_1 _3601_ (.B2(_0936_),
    .C1(net412),
    .B1(_0970_),
    .A1(_1826_),
    .Y(_0175_),
    .A2(_0968_));
 sg13g2_a21o_1 _3602_ (.A2(_0939_),
    .A1(net333),
    .B1(_1825_),
    .X(_0971_));
 sg13g2_o21ai_1 _3603_ (.B1(net333),
    .Y(_0972_),
    .A1(net403),
    .A2(_0940_));
 sg13g2_a21oi_1 _3604_ (.A1(_0971_),
    .A2(_0972_),
    .Y(_0176_),
    .B1(net412));
 sg13g2_and4_1 _3605_ (.A(net481),
    .B(_1899_),
    .C(_0582_),
    .D(_0933_),
    .X(_0177_));
 sg13g2_nand2b_1 _3606_ (.Y(_0973_),
    .B(_0788_),
    .A_N(_0787_));
 sg13g2_or2_1 _3607_ (.X(_0974_),
    .B(_0973_),
    .A(_0790_));
 sg13g2_nand2_1 _3608_ (.Y(_0975_),
    .A(net364),
    .B(_0974_));
 sg13g2_a22oi_1 _3609_ (.Y(_0178_),
    .B1(_0975_),
    .B2(net344),
    .A2(_0974_),
    .A1(_1824_));
 sg13g2_a22oi_1 _3610_ (.Y(_0179_),
    .B1(_0975_),
    .B2(net343),
    .A2(_0974_),
    .A1(_1823_));
 sg13g2_nand2_1 _3611_ (.Y(_0976_),
    .A(net345),
    .B(_0830_));
 sg13g2_and3_1 _3612_ (.X(_0977_),
    .A(_0762_),
    .B(_0828_),
    .C(_0976_));
 sg13g2_nor2_2 _3613_ (.A(net354),
    .B(_0977_),
    .Y(_0978_));
 sg13g2_and2_1 _3614_ (.A(net367),
    .B(_0977_),
    .X(_0979_));
 sg13g2_nor2_1 _3615_ (.A(net352),
    .B(_0977_),
    .Y(_0980_));
 sg13g2_nor3_2 _3616_ (.A(_0978_),
    .B(_0979_),
    .C(_0980_),
    .Y(_0981_));
 sg13g2_mux4_1 _3617_ (.S0(net354),
    .A0(\game.fsm.len3_color_count[0][0] ),
    .A1(\game.fsm.len3_color_count[2][0] ),
    .A2(\game.fsm.len3_color_count[1][0] ),
    .A3(\game.fsm.len3_color_count[3][0] ),
    .S1(net352),
    .X(_0982_));
 sg13g2_nor2_1 _3618_ (.A(net357),
    .B(_0982_),
    .Y(_0983_));
 sg13g2_mux2_1 _3619_ (.A0(net539),
    .A1(_0983_),
    .S(_0981_),
    .X(_0180_));
 sg13g2_mux4_1 _3620_ (.S0(net354),
    .A0(_0041_),
    .A1(_0043_),
    .A2(_0042_),
    .A3(_0044_),
    .S1(net352),
    .X(_0984_));
 sg13g2_xor2_1 _3621_ (.B(_0984_),
    .A(_0982_),
    .X(_0985_));
 sg13g2_xnor2_1 _3622_ (.Y(_0986_),
    .A(_0738_),
    .B(_0985_));
 sg13g2_mux2_1 _3623_ (.A0(_0976_),
    .A1(_0762_),
    .S(_0985_),
    .X(_0987_));
 sg13g2_o21ai_1 _3624_ (.B1(_0987_),
    .Y(_0988_),
    .A1(_0828_),
    .A2(_0986_));
 sg13g2_mux2_1 _3625_ (.A0(net545),
    .A1(_0988_),
    .S(_0981_),
    .X(_0181_));
 sg13g2_nand2_1 _3626_ (.Y(_0989_),
    .A(_0844_),
    .B(_0845_));
 sg13g2_nand3_1 _3627_ (.B(_0844_),
    .C(_0845_),
    .A(_0807_),
    .Y(_0990_));
 sg13g2_a21oi_1 _3628_ (.A1(_1867_),
    .A2(net362),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_a21oi_1 _3629_ (.A1(_1867_),
    .A2(_0990_),
    .Y(_0182_),
    .B1(_0991_));
 sg13g2_mux2_1 _3630_ (.A0(_0857_),
    .A1(net404),
    .S(_0990_),
    .X(_0183_));
 sg13g2_nor2_1 _3631_ (.A(_0864_),
    .B(_0990_),
    .Y(_0992_));
 sg13g2_a21oi_1 _3632_ (.A1(_1866_),
    .A2(_0990_),
    .Y(_0184_),
    .B1(_0992_));
 sg13g2_nand2b_2 _3633_ (.Y(_0993_),
    .B(_0831_),
    .A_N(_0731_));
 sg13g2_nor2_2 _3634_ (.A(_0711_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_nor2_1 _3635_ (.A(_0814_),
    .B(_0994_),
    .Y(_0995_));
 sg13g2_o21ai_1 _3636_ (.B1(_0694_),
    .Y(_0996_),
    .A1(_0814_),
    .A2(_0994_));
 sg13g2_nor2_1 _3637_ (.A(_0741_),
    .B(_0746_),
    .Y(_0997_));
 sg13g2_inv_1 _3638_ (.Y(_0998_),
    .A(_0997_));
 sg13g2_o21ai_1 _3639_ (.B1(_0996_),
    .Y(_0999_),
    .A1(net353),
    .A2(_0998_));
 sg13g2_o21ai_1 _3640_ (.B1(_0691_),
    .Y(_1000_),
    .A1(net341),
    .A2(_0994_));
 sg13g2_o21ai_1 _3641_ (.B1(_1000_),
    .Y(_1001_),
    .A1(net354),
    .A2(_0998_));
 sg13g2_nand2b_1 _3642_ (.Y(_1002_),
    .B(_1001_),
    .A_N(_0999_));
 sg13g2_xor2_1 _3643_ (.B(_1002_),
    .A(net667),
    .X(_1003_));
 sg13g2_nor2_1 _3644_ (.A(net356),
    .B(_1003_),
    .Y(_0185_));
 sg13g2_and2_1 _3645_ (.A(net366),
    .B(_1002_),
    .X(_1004_));
 sg13g2_mux4_1 _3646_ (.S0(_0849_),
    .A0(_0050_),
    .A1(_0049_),
    .A2(_0052_),
    .A3(_0051_),
    .S1(_0850_),
    .X(_1005_));
 sg13g2_mux4_1 _3647_ (.S0(_0850_),
    .A0(\game.fsm.len1_color_count[1][0] ),
    .A1(\game.fsm.len1_color_count[3][0] ),
    .A2(\game.fsm.len1_color_count[0][0] ),
    .A3(\game.fsm.len1_color_count[2][0] ),
    .S1(_0849_),
    .X(_1006_));
 sg13g2_nand2b_1 _3648_ (.Y(_1007_),
    .B(_1006_),
    .A_N(_1005_));
 sg13g2_nor2b_1 _3649_ (.A(_1006_),
    .B_N(_1005_),
    .Y(_1008_));
 sg13g2_xor2_1 _3650_ (.B(_1006_),
    .A(_1005_),
    .X(_1009_));
 sg13g2_a21oi_1 _3651_ (.A1(_0738_),
    .A2(_0749_),
    .Y(_1010_),
    .B1(net341));
 sg13g2_nand3b_1 _3652_ (.B(_1009_),
    .C(_0815_),
    .Y(_1011_),
    .A_N(_0993_));
 sg13g2_o21ai_1 _3653_ (.B1(_1011_),
    .Y(_1012_),
    .A1(_1009_),
    .A2(_1010_));
 sg13g2_mux2_1 _3654_ (.A0(_1012_),
    .A1(net598),
    .S(_1004_),
    .X(_0186_));
 sg13g2_mux4_1 _3655_ (.S0(_0850_),
    .A0(_0036_),
    .A1(_0037_),
    .A2(_0035_),
    .A3(_0038_),
    .S1(_0849_),
    .X(_1013_));
 sg13g2_xnor2_1 _3656_ (.Y(_1014_),
    .A(_1007_),
    .B(_1013_));
 sg13g2_inv_1 _3657_ (.Y(_1015_),
    .A(_1014_));
 sg13g2_nand2_1 _3658_ (.Y(_1016_),
    .A(_0763_),
    .B(_1009_));
 sg13g2_xnor2_1 _3659_ (.Y(_1017_),
    .A(_1014_),
    .B(_1016_));
 sg13g2_xnor2_1 _3660_ (.Y(_1018_),
    .A(_1008_),
    .B(_1013_));
 sg13g2_a22oi_1 _3661_ (.Y(_1019_),
    .B1(_1018_),
    .B2(_0994_),
    .A2(_1015_),
    .A1(net341));
 sg13g2_o21ai_1 _3662_ (.B1(_1019_),
    .Y(_1020_),
    .A1(_0998_),
    .A2(_1017_));
 sg13g2_mux2_1 _3663_ (.A0(_1020_),
    .A1(net506),
    .S(_1004_),
    .X(_0187_));
 sg13g2_nand2b_1 _3664_ (.Y(_1021_),
    .B(_0999_),
    .A_N(_1001_));
 sg13g2_xor2_1 _3665_ (.B(_1021_),
    .A(net685),
    .X(_1022_));
 sg13g2_nor2_1 _3666_ (.A(net356),
    .B(_1022_),
    .Y(_0188_));
 sg13g2_and2_1 _3667_ (.A(net366),
    .B(_1021_),
    .X(_1023_));
 sg13g2_mux2_1 _3668_ (.A0(_1012_),
    .A1(net615),
    .S(_1023_),
    .X(_0189_));
 sg13g2_mux2_1 _3669_ (.A0(_1020_),
    .A1(net535),
    .S(_1023_),
    .X(_0190_));
 sg13g2_o21ai_1 _3670_ (.B1(net364),
    .Y(_1024_),
    .A1(net616),
    .A2(_0806_));
 sg13g2_a21oi_1 _3671_ (.A1(_1822_),
    .A2(_0806_),
    .Y(_0191_),
    .B1(_1024_));
 sg13g2_a22oi_1 _3672_ (.Y(_1025_),
    .B1(_0806_),
    .B2(net578),
    .A2(_0703_),
    .A1(_0500_));
 sg13g2_o21ai_1 _3673_ (.B1(_0786_),
    .Y(_0192_),
    .A1(net355),
    .A2(net579));
 sg13g2_a22oi_1 _3674_ (.Y(_1026_),
    .B1(_0808_),
    .B2(net396),
    .A2(net345),
    .A1(_0503_));
 sg13g2_o21ai_1 _3675_ (.B1(_1026_),
    .Y(_0193_),
    .A1(_0540_),
    .A2(_0707_));
 sg13g2_o21ai_1 _3676_ (.B1(_0813_),
    .Y(_1027_),
    .A1(_0744_),
    .A2(_0993_));
 sg13g2_nor2_1 _3677_ (.A(net395),
    .B(net338),
    .Y(_1028_));
 sg13g2_nor2b_1 _3678_ (.A(net330),
    .B_N(net338),
    .Y(_1029_));
 sg13g2_nor3_1 _3679_ (.A(net358),
    .B(_1028_),
    .C(_1029_),
    .Y(_0194_));
 sg13g2_nor2_1 _3680_ (.A(net348),
    .B(_0712_),
    .Y(_1030_));
 sg13g2_xnor2_1 _3681_ (.Y(_1031_),
    .A(net348),
    .B(_0712_));
 sg13g2_o21ai_1 _3682_ (.B1(net361),
    .Y(_1032_),
    .A1(net784),
    .A2(net338));
 sg13g2_a21oi_1 _3683_ (.A1(net338),
    .A2(_1031_),
    .Y(_0195_),
    .B1(_1032_));
 sg13g2_xnor2_1 _3684_ (.Y(_1033_),
    .A(_0716_),
    .B(_1030_));
 sg13g2_o21ai_1 _3685_ (.B1(net361),
    .Y(_1034_),
    .A1(net779),
    .A2(net338));
 sg13g2_a21oi_1 _3686_ (.A1(net338),
    .A2(_1033_),
    .Y(_0196_),
    .B1(_1034_));
 sg13g2_a221oi_1 _3687_ (.B2(_0709_),
    .C1(_0806_),
    .B1(_0993_),
    .A1(net348),
    .Y(_1035_),
    .A2(_0741_));
 sg13g2_o21ai_1 _3688_ (.B1(net366),
    .Y(_1036_),
    .A1(\game.fsm.len1_block_count[0] ),
    .A2(_1035_));
 sg13g2_a21oi_1 _3689_ (.A1(_1817_),
    .A2(_1035_),
    .Y(_0197_),
    .B1(_1036_));
 sg13g2_o21ai_1 _3690_ (.B1(_0708_),
    .Y(_1037_),
    .A1(net349),
    .A2(_0993_));
 sg13g2_and2_1 _3691_ (.A(\game.fsm.len1_block_count[1] ),
    .B(\game.fsm.len1_block_count[0] ),
    .X(_1038_));
 sg13g2_xor2_1 _3692_ (.B(\game.fsm.len1_block_count[0] ),
    .A(net746),
    .X(_1039_));
 sg13g2_xnor2_1 _3693_ (.Y(_1040_),
    .A(_1037_),
    .B(_1039_));
 sg13g2_o21ai_1 _3694_ (.B1(net366),
    .Y(_1041_),
    .A1(net746),
    .A2(_1035_));
 sg13g2_a21oi_1 _3695_ (.A1(_1035_),
    .A2(_1040_),
    .Y(_0198_),
    .B1(_1041_));
 sg13g2_o21ai_1 _3696_ (.B1(_1035_),
    .Y(_1042_),
    .A1(_1037_),
    .A2(_1038_));
 sg13g2_a21o_1 _3697_ (.A2(_1037_),
    .A1(_0489_),
    .B1(_1042_),
    .X(_1043_));
 sg13g2_xor2_1 _3698_ (.B(_1043_),
    .A(net674),
    .X(_1044_));
 sg13g2_nor2_1 _3699_ (.A(net356),
    .B(_1044_),
    .Y(_0199_));
 sg13g2_nor2b_1 _3700_ (.A(_0708_),
    .B_N(_0741_),
    .Y(_1045_));
 sg13g2_o21ai_1 _3701_ (.B1(_0723_),
    .Y(_1046_),
    .A1(net349),
    .A2(_0731_));
 sg13g2_nor4_2 _3702_ (.A(_0806_),
    .B(_0812_),
    .C(_1045_),
    .Y(_1047_),
    .D(_1046_));
 sg13g2_o21ai_1 _3703_ (.B1(net364),
    .Y(_1048_),
    .A1(\game.fsm.len2_block_count[0] ),
    .A2(_1047_));
 sg13g2_a21oi_1 _3704_ (.A1(_1816_),
    .A2(_1047_),
    .Y(_0200_),
    .B1(_1048_));
 sg13g2_nor2_1 _3705_ (.A(_2023_),
    .B(_0482_),
    .Y(_1049_));
 sg13g2_nor2_1 _3706_ (.A(net349),
    .B(_0759_),
    .Y(_1050_));
 sg13g2_o21ai_1 _3707_ (.B1(_0993_),
    .Y(_1051_),
    .A1(net349),
    .A2(_0759_));
 sg13g2_xnor2_1 _3708_ (.Y(_1052_),
    .A(_1049_),
    .B(_1051_));
 sg13g2_o21ai_1 _3709_ (.B1(net364),
    .Y(_1053_),
    .A1(net695),
    .A2(_1047_));
 sg13g2_a21oi_1 _3710_ (.A1(_1047_),
    .A2(_1052_),
    .Y(_0201_),
    .B1(_1053_));
 sg13g2_a21oi_1 _3711_ (.A1(net348),
    .A2(_0830_),
    .Y(_1054_),
    .B1(_0747_));
 sg13g2_a21oi_1 _3712_ (.A1(_0743_),
    .A2(_1050_),
    .Y(_1055_),
    .B1(_0709_));
 sg13g2_nor2_1 _3713_ (.A(_1054_),
    .B(_1055_),
    .Y(_1056_));
 sg13g2_o21ai_1 _3714_ (.B1(net366),
    .Y(_1057_),
    .A1(\game.fsm.len3_block_count[0] ),
    .A2(_1056_));
 sg13g2_a21oi_1 _3715_ (.A1(_1815_),
    .A2(_1056_),
    .Y(_0202_),
    .B1(_1057_));
 sg13g2_a21oi_1 _3716_ (.A1(net348),
    .A2(_0748_),
    .Y(_1058_),
    .B1(_0759_));
 sg13g2_xor2_1 _3717_ (.B(_1058_),
    .A(\game.fsm.len3_block_count[0] ),
    .X(_1059_));
 sg13g2_nand2_1 _3718_ (.Y(_1060_),
    .A(_1056_),
    .B(_1059_));
 sg13g2_xor2_1 _3719_ (.B(_1060_),
    .A(net628),
    .X(_1061_));
 sg13g2_nor2_1 _3720_ (.A(net355),
    .B(_1061_),
    .Y(_0203_));
 sg13g2_nand3_1 _3721_ (.B(net353),
    .C(net348),
    .A(_0510_),
    .Y(_1062_));
 sg13g2_nand3_1 _3722_ (.B(_0695_),
    .C(net349),
    .A(_0691_),
    .Y(_1063_));
 sg13g2_nand2_1 _3723_ (.Y(_1064_),
    .A(_1062_),
    .B(_1063_));
 sg13g2_a21oi_1 _3724_ (.A1(net339),
    .A2(_1064_),
    .Y(_1065_),
    .B1(net493));
 sg13g2_nand2_1 _3725_ (.Y(_1066_),
    .A(net493),
    .B(_1064_));
 sg13g2_nor2b_1 _3726_ (.A(_1066_),
    .B_N(net339),
    .Y(_1067_));
 sg13g2_nor3_1 _3727_ (.A(net356),
    .B(_1065_),
    .C(_1067_),
    .Y(_0204_));
 sg13g2_or2_1 _3728_ (.X(_1068_),
    .B(_1062_),
    .A(_1814_));
 sg13g2_xnor2_1 _3729_ (.Y(_1069_),
    .A(_1814_),
    .B(_1062_));
 sg13g2_xnor2_1 _3730_ (.Y(_1070_),
    .A(_1066_),
    .B(_1069_));
 sg13g2_o21ai_1 _3731_ (.B1(net368),
    .Y(_1071_),
    .A1(net540),
    .A2(net339));
 sg13g2_a21oi_1 _3732_ (.A1(net339),
    .A2(_1070_),
    .Y(_0205_),
    .B1(net541));
 sg13g2_o21ai_1 _3733_ (.B1(_1068_),
    .Y(_1072_),
    .A1(_1066_),
    .A2(_1069_));
 sg13g2_xnor2_1 _3734_ (.Y(_1073_),
    .A(net654),
    .B(_1062_));
 sg13g2_xnor2_1 _3735_ (.Y(_1074_),
    .A(_1072_),
    .B(_1073_));
 sg13g2_o21ai_1 _3736_ (.B1(net368),
    .Y(_1075_),
    .A1(net654),
    .A2(net338));
 sg13g2_a21oi_1 _3737_ (.A1(net338),
    .A2(_1074_),
    .Y(_0206_),
    .B1(net655));
 sg13g2_nor2_2 _3738_ (.A(\btn.input_event[0] ),
    .B(\btn.input_event[1] ),
    .Y(_1076_));
 sg13g2_inv_1 _3739_ (.Y(_1077_),
    .A(_1076_));
 sg13g2_and2_1 _3740_ (.A(_0040_),
    .B(_1076_),
    .X(_1078_));
 sg13g2_and3_2 _3741_ (.X(_1079_),
    .A(\btn.input_event[3] ),
    .B(\btn.input_event[2] ),
    .C(_1078_));
 sg13g2_nand3_1 _3742_ (.B(\btn.input_event[2] ),
    .C(_1078_),
    .A(\btn.input_event[3] ),
    .Y(_1080_));
 sg13g2_nor4_2 _3743_ (.A(_1881_),
    .B(\btn.input_event[3] ),
    .C(\btn.input_event[2] ),
    .Y(_1081_),
    .D(\btn.input_event[4] ));
 sg13g2_a21oi_2 _3744_ (.B1(_1079_),
    .Y(_1082_),
    .A2(_1081_),
    .A1(\btn.input_event[1] ));
 sg13g2_nand2_2 _3745_ (.Y(_1083_),
    .A(net372),
    .B(_1082_));
 sg13g2_o21ai_1 _3746_ (.B1(net346),
    .Y(_1084_),
    .A1(_1803_),
    .A2(_1083_));
 sg13g2_nor2_2 _3747_ (.A(_0600_),
    .B(_1084_),
    .Y(_1085_));
 sg13g2_nand2b_1 _3748_ (.Y(_1086_),
    .B(_0601_),
    .A_N(_1084_));
 sg13g2_nor3_2 _3749_ (.A(\game.challenge_num[2] ),
    .B(\game.challenge_num[1] ),
    .C(net393),
    .Y(_1087_));
 sg13g2_a21oi_2 _3750_ (.B1(_1079_),
    .Y(_1088_),
    .A2(_1087_),
    .A1(_1812_));
 sg13g2_nor2_1 _3751_ (.A(_0605_),
    .B(_1080_),
    .Y(_1089_));
 sg13g2_nor2_1 _3752_ (.A(_1803_),
    .B(net393),
    .Y(_1090_));
 sg13g2_o21ai_1 _3753_ (.B1(_1090_),
    .Y(_1091_),
    .A1(_1088_),
    .A2(_1089_));
 sg13g2_nand2b_1 _3754_ (.Y(_1092_),
    .B(_1091_),
    .A_N(_0637_));
 sg13g2_o21ai_1 _3755_ (.B1(net429),
    .Y(_1093_),
    .A1(_1086_),
    .A2(_1092_));
 sg13g2_a21oi_1 _3756_ (.A1(_1813_),
    .A2(_1086_),
    .Y(_0207_),
    .B1(_1093_));
 sg13g2_nor3_1 _3757_ (.A(_0605_),
    .B(_0644_),
    .C(_1080_),
    .Y(_1094_));
 sg13g2_a21o_1 _3758_ (.A2(_1080_),
    .A1(_0644_),
    .B1(net369),
    .X(_1095_));
 sg13g2_o21ai_1 _3759_ (.B1(_0645_),
    .Y(_1096_),
    .A1(_1094_),
    .A2(_1095_));
 sg13g2_o21ai_1 _3760_ (.B1(net429),
    .Y(_1097_),
    .A1(net765),
    .A2(_1085_));
 sg13g2_a21oi_1 _3761_ (.A1(_1085_),
    .A2(_1096_),
    .Y(_0208_),
    .B1(_1097_));
 sg13g2_nand2b_1 _3762_ (.Y(_1098_),
    .B(_0627_),
    .A_N(_0605_));
 sg13g2_xor2_1 _3763_ (.B(_0643_),
    .A(_0054_),
    .X(_1099_));
 sg13g2_a22oi_1 _3764_ (.Y(_1100_),
    .B1(_1099_),
    .B2(_1088_),
    .A2(_1098_),
    .A1(_1079_));
 sg13g2_nor2_1 _3765_ (.A(net369),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_o21ai_1 _3766_ (.B1(_1085_),
    .Y(_1102_),
    .A1(_0628_),
    .A2(_1101_));
 sg13g2_o21ai_1 _3767_ (.B1(_1102_),
    .Y(_1103_),
    .A1(net704),
    .A2(_1085_));
 sg13g2_nor2_1 _3768_ (.A(net418),
    .B(_1103_),
    .Y(_0209_));
 sg13g2_o21ai_1 _3769_ (.B1(_1079_),
    .Y(_1104_),
    .A1(_0605_),
    .A2(_0651_));
 sg13g2_xor2_1 _3770_ (.B(_1087_),
    .A(_0055_),
    .X(_1105_));
 sg13g2_a21oi_1 _3771_ (.A1(_1088_),
    .A2(_1105_),
    .Y(_1106_),
    .B1(net369));
 sg13g2_nand2_1 _3772_ (.Y(_1107_),
    .A(_1104_),
    .B(_1106_));
 sg13g2_a21oi_1 _3773_ (.A1(_0652_),
    .A2(_1107_),
    .Y(_1108_),
    .B1(_1084_));
 sg13g2_a21oi_1 _3774_ (.A1(net552),
    .A2(_1086_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_nor2_1 _3775_ (.A(net418),
    .B(_1109_),
    .Y(_0210_));
 sg13g2_nand2b_2 _3776_ (.Y(_1110_),
    .B(\btn.input_event[0] ),
    .A_N(\btn.input_event[1] ));
 sg13g2_nor2b_2 _3777_ (.A(\btn.input_event[2] ),
    .B_N(\btn.input_event[3] ),
    .Y(_1111_));
 sg13g2_nand2_1 _3778_ (.Y(_1112_),
    .A(_0040_),
    .B(_1111_));
 sg13g2_nor2_1 _3779_ (.A(_1110_),
    .B(_1112_),
    .Y(_1113_));
 sg13g2_o21ai_1 _3780_ (.B1(_0624_),
    .Y(_1114_),
    .A1(_1110_),
    .A2(_1112_));
 sg13g2_nand2b_1 _3781_ (.Y(_1115_),
    .B(_0608_),
    .A_N(_0605_));
 sg13g2_nand4_1 _3782_ (.B(_0616_),
    .C(_1114_),
    .A(_0601_),
    .Y(_1116_),
    .D(_1115_));
 sg13g2_o21ai_1 _3783_ (.B1(net429),
    .Y(_1117_),
    .A1(net351),
    .A2(_1116_));
 sg13g2_a21oi_1 _3784_ (.A1(_1811_),
    .A2(_1116_),
    .Y(_0211_),
    .B1(_1117_));
 sg13g2_nand3_1 _3785_ (.B(_1076_),
    .C(_1111_),
    .A(\btn.input_event[4] ),
    .Y(_1118_));
 sg13g2_nor3_2 _3786_ (.A(_0595_),
    .B(_0696_),
    .C(_1118_),
    .Y(_1119_));
 sg13g2_and2_1 _3787_ (.A(net421),
    .B(_1119_),
    .X(_0212_));
 sg13g2_nor2_2 _3788_ (.A(\btn.input_event[3] ),
    .B(_1882_),
    .Y(_1120_));
 sg13g2_or4_1 _3789_ (.A(\btn.input_event[3] ),
    .B(_1882_),
    .C(\btn.input_event[4] ),
    .D(_1110_),
    .X(_1121_));
 sg13g2_nand3_1 _3790_ (.B(_0596_),
    .C(_1111_),
    .A(_0040_),
    .Y(_1122_));
 sg13g2_nand3_1 _3791_ (.B(_1121_),
    .C(_1122_),
    .A(_0599_),
    .Y(_1123_));
 sg13g2_nor2_1 _3792_ (.A(net371),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_nand3_1 _3793_ (.B(_0612_),
    .C(net369),
    .A(_0609_),
    .Y(_1125_));
 sg13g2_or2_2 _3794_ (.X(_1126_),
    .B(_1125_),
    .A(_1124_));
 sg13g2_nor2_2 _3795_ (.A(_0615_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_o21ai_1 _3796_ (.B1(_0924_),
    .Y(_1128_),
    .A1(net465),
    .A2(_1127_));
 sg13g2_nor2_1 _3797_ (.A(net414),
    .B(_1128_),
    .Y(_0213_));
 sg13g2_o21ai_1 _3798_ (.B1(_1127_),
    .Y(_1129_),
    .A1(_0595_),
    .A2(_1122_));
 sg13g2_o21ai_1 _3799_ (.B1(_1129_),
    .Y(_1130_),
    .A1(net559),
    .A2(_1127_));
 sg13g2_nor2_1 _3800_ (.A(net411),
    .B(_1130_),
    .Y(_0214_));
 sg13g2_o21ai_1 _3801_ (.B1(net421),
    .Y(_1131_),
    .A1(net659),
    .A2(_1127_));
 sg13g2_a21oi_1 _3802_ (.A1(_0600_),
    .A2(_1127_),
    .Y(_0215_),
    .B1(_1131_));
 sg13g2_and4_1 _3803_ (.A(_0612_),
    .B(net369),
    .C(_1083_),
    .D(_1126_),
    .X(_1132_));
 sg13g2_nand4_1 _3804_ (.B(net369),
    .C(_1083_),
    .A(_0612_),
    .Y(_1133_),
    .D(_1126_));
 sg13g2_nor3_1 _3805_ (.A(\game.current_level[3] ),
    .B(net390),
    .C(_0481_),
    .Y(_1134_));
 sg13g2_inv_1 _3806_ (.Y(_1135_),
    .A(_1134_));
 sg13g2_a21o_1 _3807_ (.A2(_1134_),
    .A1(_0084_),
    .B1(net523),
    .X(_1136_));
 sg13g2_nand2_1 _3808_ (.Y(_1137_),
    .A(_0403_),
    .B(_0411_));
 sg13g2_nor2_2 _3809_ (.A(net371),
    .B(_1079_),
    .Y(_1138_));
 sg13g2_a22oi_1 _3810_ (.Y(_1139_),
    .B1(_1138_),
    .B2(_1136_),
    .A2(_1137_),
    .A1(net523));
 sg13g2_o21ai_1 _3811_ (.B1(net421),
    .Y(_1140_),
    .A1(net392),
    .A2(net340));
 sg13g2_a21oi_1 _3812_ (.A1(net340),
    .A2(net524),
    .Y(_0216_),
    .B1(_1140_));
 sg13g2_xor2_1 _3813_ (.B(_1138_),
    .A(_0642_),
    .X(_1141_));
 sg13g2_o21ai_1 _3814_ (.B1(net421),
    .Y(_1142_),
    .A1(net391),
    .A2(net340));
 sg13g2_a21oi_1 _3815_ (.A1(net340),
    .A2(_1141_),
    .Y(_0217_),
    .B1(_1142_));
 sg13g2_a21oi_2 _3816_ (.B1(_1138_),
    .Y(_1143_),
    .A2(_0411_),
    .A1(_0403_));
 sg13g2_xor2_1 _3817_ (.B(_0481_),
    .A(net390),
    .X(_1144_));
 sg13g2_a21oi_1 _3818_ (.A1(net787),
    .A2(_1134_),
    .Y(_1145_),
    .B1(_1144_));
 sg13g2_a22oi_1 _3819_ (.Y(_1146_),
    .B1(_1145_),
    .B2(_1138_),
    .A2(_1143_),
    .A1(_0631_));
 sg13g2_o21ai_1 _3820_ (.B1(net421),
    .Y(_1147_),
    .A1(net390),
    .A2(net340));
 sg13g2_a21oi_1 _3821_ (.A1(_1132_),
    .A2(net788),
    .Y(_0218_),
    .B1(_1147_));
 sg13g2_nor2_1 _3822_ (.A(_0084_),
    .B(_1135_),
    .Y(_1148_));
 sg13g2_o21ai_1 _3823_ (.B1(\game.current_level[3] ),
    .Y(_1149_),
    .A1(net390),
    .A2(_0481_));
 sg13g2_o21ai_1 _3824_ (.B1(_1149_),
    .Y(_1150_),
    .A1(_0084_),
    .A2(_1135_));
 sg13g2_a22oi_1 _3825_ (.Y(_1151_),
    .B1(_1150_),
    .B2(_1138_),
    .A2(_1143_),
    .A1(_0653_));
 sg13g2_o21ai_1 _3826_ (.B1(net429),
    .Y(_1152_),
    .A1(\game.current_level[3] ),
    .A2(net340));
 sg13g2_a21oi_1 _3827_ (.A1(net340),
    .A2(net774),
    .Y(_0219_),
    .B1(_1152_));
 sg13g2_a21oi_1 _3828_ (.A1(_1135_),
    .A2(_1138_),
    .Y(_1153_),
    .B1(_1133_));
 sg13g2_nand2_1 _3829_ (.Y(_1154_),
    .A(net766),
    .B(_1148_));
 sg13g2_a22oi_1 _3830_ (.Y(_1155_),
    .B1(_1154_),
    .B2(_1138_),
    .A2(_1143_),
    .A1(_0603_));
 sg13g2_o21ai_1 _3831_ (.B1(net429),
    .Y(_1156_),
    .A1(net766),
    .A2(_1153_));
 sg13g2_a21oi_1 _3832_ (.A1(net340),
    .A2(_1155_),
    .Y(_0220_),
    .B1(_1156_));
 sg13g2_nor2_2 _3833_ (.A(net383),
    .B(_0922_),
    .Y(_1157_));
 sg13g2_nand2_1 _3834_ (.Y(_1158_),
    .A(net408),
    .B(_1157_));
 sg13g2_nand2_1 _3835_ (.Y(_1159_),
    .A(\game.counter[6] ),
    .B(\game.counter[5] ));
 sg13g2_nor3_1 _3836_ (.A(\game.counter[4] ),
    .B(\game.counter[3] ),
    .C(\game.counter[2] ),
    .Y(_1160_));
 sg13g2_nor2_1 _3837_ (.A(_1159_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_nor2_1 _3838_ (.A(\game.counter[7] ),
    .B(_1161_),
    .Y(_1162_));
 sg13g2_nand2b_1 _3839_ (.Y(_1163_),
    .B(net397),
    .A_N(\game.fsm.read_pos[1] ));
 sg13g2_o21ai_1 _3840_ (.B1(_1163_),
    .Y(_1164_),
    .A1(\game.fsm.read_pos[0] ),
    .A2(_1822_));
 sg13g2_a22oi_1 _3841_ (.Y(_1165_),
    .B1(_1821_),
    .B2(\game.fsm.read_pos[1] ),
    .A2(_1820_),
    .A1(\game.fsm.read_pos[2] ));
 sg13g2_a22oi_1 _3842_ (.Y(_1166_),
    .B1(_1164_),
    .B2(_1165_),
    .A2(net396),
    .A1(_1808_));
 sg13g2_nor2_1 _3843_ (.A(_1162_),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_nor2_1 _3844_ (.A(_1158_),
    .B(_1167_),
    .Y(_1168_));
 sg13g2_nand2_2 _3845_ (.Y(_1169_),
    .A(net383),
    .B(_0592_));
 sg13g2_inv_1 _3846_ (.Y(_1170_),
    .A(_1169_));
 sg13g2_nor3_1 _3847_ (.A(\game.counter[7] ),
    .B(_1161_),
    .C(_1169_),
    .Y(_1171_));
 sg13g2_and2_1 _3848_ (.A(_0610_),
    .B(_0614_),
    .X(_1172_));
 sg13g2_nand2_1 _3849_ (.Y(_1173_),
    .A(_0610_),
    .B(_0614_));
 sg13g2_nor4_2 _3850_ (.A(_0080_),
    .B(_1168_),
    .C(_1171_),
    .Y(_1174_),
    .D(_1173_));
 sg13g2_inv_1 _3851_ (.Y(_1175_),
    .A(_1174_));
 sg13g2_a21oi_1 _3852_ (.A1(\game.state[1] ),
    .A2(_1174_),
    .Y(_1176_),
    .B1(net561));
 sg13g2_and2_1 _3853_ (.A(net561),
    .B(_1174_),
    .X(_1177_));
 sg13g2_nor3_1 _3854_ (.A(net411),
    .B(net562),
    .C(_1177_),
    .Y(_0221_));
 sg13g2_nand2_1 _3855_ (.Y(_1178_),
    .A(net722),
    .B(_1177_));
 sg13g2_o21ai_1 _3856_ (.B1(_1178_),
    .Y(_1179_),
    .A1(_1169_),
    .A2(_1175_));
 sg13g2_o21ai_1 _3857_ (.B1(net426),
    .Y(_1180_),
    .A1(net722),
    .A2(_1177_));
 sg13g2_nor2_1 _3858_ (.A(_1179_),
    .B(_1180_),
    .Y(_0222_));
 sg13g2_nand2_1 _3859_ (.Y(_1181_),
    .A(_1808_),
    .B(_1169_));
 sg13g2_a221oi_1 _3860_ (.B2(_1181_),
    .C1(net411),
    .B1(_1179_),
    .A1(_1808_),
    .Y(_0223_),
    .A2(_1178_));
 sg13g2_nand2_1 _3861_ (.Y(_1182_),
    .A(net389),
    .B(net428));
 sg13g2_a21oi_1 _3862_ (.A1(net778),
    .A2(_0923_),
    .Y(_1183_),
    .B1(_1182_));
 sg13g2_or2_1 _3863_ (.X(_0224_),
    .B(_1183_),
    .A(_0162_));
 sg13g2_nor2b_2 _3864_ (.A(\btn.input_event[1] ),
    .B_N(_1081_),
    .Y(_1184_));
 sg13g2_and3_1 _3865_ (.X(_1185_),
    .A(_0040_),
    .B(_0596_),
    .C(_0597_));
 sg13g2_nor2_1 _3866_ (.A(_1184_),
    .B(_1185_),
    .Y(_1186_));
 sg13g2_nand2_1 _3867_ (.Y(_1187_),
    .A(_1078_),
    .B(_1120_));
 sg13g2_o21ai_1 _3868_ (.B1(_1078_),
    .Y(_1188_),
    .A1(_1111_),
    .A2(_1120_));
 sg13g2_and2_2 _3869_ (.A(_1186_),
    .B(_1188_),
    .X(_1189_));
 sg13g2_nand2_1 _3870_ (.Y(_1190_),
    .A(net351),
    .B(_0702_));
 sg13g2_nor2_2 _3871_ (.A(_1189_),
    .B(_1190_),
    .Y(_1191_));
 sg13g2_nand2_1 _3872_ (.Y(_1192_),
    .A(net498),
    .B(net421));
 sg13g2_nor3_2 _3873_ (.A(net414),
    .B(_1189_),
    .C(_1190_),
    .Y(_0227_));
 sg13g2_nand3_1 _3874_ (.B(_1882_),
    .C(_0227_),
    .A(_1881_),
    .Y(_1193_));
 sg13g2_o21ai_1 _3875_ (.B1(_1193_),
    .Y(_0225_),
    .A1(_1191_),
    .A2(_1192_));
 sg13g2_o21ai_1 _3876_ (.B1(net421),
    .Y(_1194_),
    .A1(net612),
    .A2(_1191_));
 sg13g2_a21oi_1 _3877_ (.A1(_1077_),
    .A2(_1191_),
    .Y(_0226_),
    .B1(_1194_));
 sg13g2_o21ai_1 _3878_ (.B1(_1082_),
    .Y(_1195_),
    .A1(_0598_),
    .A2(_1110_));
 sg13g2_nand2_1 _3879_ (.Y(_1196_),
    .A(net350),
    .B(_1195_));
 sg13g2_nand2b_1 _3880_ (.Y(_0228_),
    .B(_1196_),
    .A_N(_1117_));
 sg13g2_and2_1 _3881_ (.A(net431),
    .B(net322),
    .X(_0229_));
 sg13g2_nand2_1 _3882_ (.Y(_1197_),
    .A(net431),
    .B(net781));
 sg13g2_inv_1 _3883_ (.Y(_0230_),
    .A(_1197_));
 sg13g2_nand3_1 _3884_ (.B(_1076_),
    .C(_1120_),
    .A(\btn.input_event[4] ),
    .Y(_1198_));
 sg13g2_nand2_2 _3885_ (.Y(_1199_),
    .A(_1187_),
    .B(_1198_));
 sg13g2_or4_1 _3886_ (.A(_1113_),
    .B(_1184_),
    .C(_1185_),
    .D(_1199_),
    .X(_1200_));
 sg13g2_nand2_1 _3887_ (.Y(_1201_),
    .A(_0597_),
    .B(_1078_));
 sg13g2_nand3_1 _3888_ (.B(_0596_),
    .C(_1120_),
    .A(_0040_),
    .Y(_1202_));
 sg13g2_nand3_1 _3889_ (.B(_1201_),
    .C(_1202_),
    .A(_1082_),
    .Y(_1203_));
 sg13g2_nor2_1 _3890_ (.A(_1200_),
    .B(_1203_),
    .Y(_1204_));
 sg13g2_o21ai_1 _3891_ (.B1(net370),
    .Y(_1205_),
    .A1(_0013_),
    .A2(_1204_));
 sg13g2_nor3_1 _3892_ (.A(_0013_),
    .B(_0607_),
    .C(_0610_),
    .Y(_1206_));
 sg13g2_and2_1 _3893_ (.A(_0895_),
    .B(_1206_),
    .X(_1207_));
 sg13g2_a21oi_1 _3894_ (.A1(net479),
    .A2(_1207_),
    .Y(_1208_),
    .B1(net372));
 sg13g2_nor2_1 _3895_ (.A(net351),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_nor3_1 _3896_ (.A(\game.state[2] ),
    .B(net382),
    .C(net383),
    .Y(_1210_));
 sg13g2_nor2_1 _3897_ (.A(_1802_),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_a21oi_1 _3898_ (.A1(_0080_),
    .A2(_1172_),
    .Y(_1212_),
    .B1(_1211_));
 sg13g2_nor2b_2 _3899_ (.A(_1157_),
    .B_N(net342),
    .Y(_1213_));
 sg13g2_inv_1 _3900_ (.Y(_1214_),
    .A(_1213_));
 sg13g2_a221oi_1 _3901_ (.B2(_1209_),
    .C1(_1214_),
    .B1(_1205_),
    .A1(net665),
    .Y(_1215_),
    .A2(net350));
 sg13g2_o21ai_1 _3902_ (.B1(net433),
    .Y(_1216_),
    .A1(net670),
    .A2(_1213_));
 sg13g2_nor2_1 _3903_ (.A(_1215_),
    .B(_1216_),
    .Y(_0231_));
 sg13g2_nand3b_1 _3904_ (.B(_0596_),
    .C(_1120_),
    .Y(_1217_),
    .A_N(\btn.input_event[4] ));
 sg13g2_nand3_1 _3905_ (.B(_1201_),
    .C(_1217_),
    .A(_1198_),
    .Y(_1218_));
 sg13g2_or2_1 _3906_ (.X(_1219_),
    .B(_1218_),
    .A(_1123_));
 sg13g2_nand3_1 _3907_ (.B(net350),
    .C(_1118_),
    .A(\game.sound_on ),
    .Y(_1220_));
 sg13g2_nor3_1 _3908_ (.A(_1195_),
    .B(_1219_),
    .C(_1220_),
    .Y(_1221_));
 sg13g2_o21ai_1 _3909_ (.B1(_1118_),
    .Y(_1222_),
    .A1(_0702_),
    .A2(_1189_));
 sg13g2_nor2_1 _3910_ (.A(_0696_),
    .B(_1118_),
    .Y(_1223_));
 sg13g2_nor3_1 _3911_ (.A(_0013_),
    .B(net371),
    .C(_1223_),
    .Y(_1224_));
 sg13g2_a22oi_1 _3912_ (.Y(_1225_),
    .B1(_1222_),
    .B2(_1224_),
    .A2(_1221_),
    .A1(_1189_));
 sg13g2_nand2_1 _3913_ (.Y(_1226_),
    .A(_1213_),
    .B(_1225_));
 sg13g2_a221oi_1 _3914_ (.B2(net469),
    .C1(_1226_),
    .B1(_1207_),
    .A1(net665),
    .Y(_1227_),
    .A2(_1170_));
 sg13g2_o21ai_1 _3915_ (.B1(net433),
    .Y(_1228_),
    .A1(net684),
    .A2(_1213_));
 sg13g2_nor2_1 _3916_ (.A(_1227_),
    .B(_1228_),
    .Y(_0232_));
 sg13g2_nand4_1 _3917_ (.B(net381),
    .C(net384),
    .A(net793),
    .Y(_1229_),
    .D(_0606_));
 sg13g2_inv_1 _3918_ (.Y(_1230_),
    .A(_1229_));
 sg13g2_nand2_1 _3919_ (.Y(_1231_),
    .A(_0895_),
    .B(_1230_));
 sg13g2_nor2b_1 _3920_ (.A(_1226_),
    .B_N(_1231_),
    .Y(_1232_));
 sg13g2_o21ai_1 _3921_ (.B1(net433),
    .Y(_1233_),
    .A1(net595),
    .A2(_1213_));
 sg13g2_nor2_1 _3922_ (.A(_1232_),
    .B(_1233_),
    .Y(_0233_));
 sg13g2_o21ai_1 _3923_ (.B1(net430),
    .Y(_1234_),
    .A1(net732),
    .A2(_0618_));
 sg13g2_nor2_1 _3924_ (.A(_0600_),
    .B(net733),
    .Y(_0234_));
 sg13g2_nand2b_1 _3925_ (.Y(_1235_),
    .B(net748),
    .A_N(net346));
 sg13g2_a21oi_1 _3926_ (.A1(_0633_),
    .A2(_1235_),
    .Y(_0237_),
    .B1(net417));
 sg13g2_nand3b_1 _3927_ (.B(net350),
    .C(_0581_),
    .Y(_1236_),
    .A_N(_0696_));
 sg13g2_nor2b_1 _3928_ (.A(_1166_),
    .B_N(_1157_),
    .Y(_1237_));
 sg13g2_nand2b_1 _3929_ (.Y(_1238_),
    .B(_0007_),
    .A_N(\game.fsm.seq[5][0] ));
 sg13g2_o21ai_1 _3930_ (.B1(_1238_),
    .Y(_1239_),
    .A1(\game.fsm.seq[4][0] ),
    .A2(_0007_));
 sg13g2_mux2_1 _3931_ (.A0(\game.fsm.seq[6][0] ),
    .A1(\game.fsm.seq[7][0] ),
    .S(_0007_),
    .X(_1240_));
 sg13g2_o21ai_1 _3932_ (.B1(_0009_),
    .Y(_1241_),
    .A1(_0008_),
    .A2(_1239_));
 sg13g2_a21oi_2 _3933_ (.B1(_1241_),
    .Y(_1242_),
    .A2(_1240_),
    .A1(_0008_));
 sg13g2_mux4_1 _3934_ (.S0(_0008_),
    .A0(\game.fsm.seq[0][0] ),
    .A1(\game.fsm.seq[2][0] ),
    .A2(\game.fsm.seq[1][0] ),
    .A3(\game.fsm.seq[3][0] ),
    .S1(_0007_),
    .X(_1243_));
 sg13g2_nor2_2 _3935_ (.A(_0009_),
    .B(_1243_),
    .Y(_1244_));
 sg13g2_nor2_1 _3936_ (.A(_1242_),
    .B(_1244_),
    .Y(_1245_));
 sg13g2_o21ai_1 _3937_ (.B1(_1237_),
    .Y(_1246_),
    .A1(_1242_),
    .A2(_1244_));
 sg13g2_nand2_1 _3938_ (.Y(_1247_),
    .A(net737),
    .B(\game.counter[0] ));
 sg13g2_nand4_1 _3939_ (.B(\game.counter[2] ),
    .C(\game.counter[1] ),
    .A(\game.counter[3] ),
    .Y(_1248_),
    .D(\game.counter[0] ));
 sg13g2_xnor2_1 _3940_ (.Y(_1249_),
    .A(net642),
    .B(_1248_));
 sg13g2_nor3_1 _3941_ (.A(_1801_),
    .B(\game.counter[2] ),
    .C(\game.counter[1] ),
    .Y(_1250_));
 sg13g2_nand4_1 _3942_ (.B(\game.counter[0] ),
    .C(_1162_),
    .A(\game.counter[3] ),
    .Y(_1251_),
    .D(_1250_));
 sg13g2_and2_1 _3943_ (.A(\game.counter[4] ),
    .B(\game.counter[3] ),
    .X(_1252_));
 sg13g2_o21ai_1 _3944_ (.B1(_1252_),
    .Y(_1253_),
    .A1(\game.counter[2] ),
    .A2(\game.counter[1] ));
 sg13g2_nor2_1 _3945_ (.A(\game.counter[6] ),
    .B(\game.counter[5] ),
    .Y(_1254_));
 sg13g2_and4_1 _3946_ (.A(_0058_),
    .B(_1251_),
    .C(_1253_),
    .D(_1254_),
    .X(_1255_));
 sg13g2_nand2b_1 _3947_ (.Y(_1256_),
    .B(_0007_),
    .A_N(\game.fsm.seq[5][1] ));
 sg13g2_o21ai_1 _3948_ (.B1(_1256_),
    .Y(_1257_),
    .A1(\game.fsm.seq[4][1] ),
    .A2(_0007_));
 sg13g2_mux2_1 _3949_ (.A0(\game.fsm.seq[6][1] ),
    .A1(\game.fsm.seq[7][1] ),
    .S(_0007_),
    .X(_1258_));
 sg13g2_o21ai_1 _3950_ (.B1(_0009_),
    .Y(_1259_),
    .A1(_0008_),
    .A2(_1257_));
 sg13g2_a21oi_1 _3951_ (.A1(_0008_),
    .A2(_1258_),
    .Y(_1260_),
    .B1(_1259_));
 sg13g2_mux4_1 _3952_ (.S0(_0008_),
    .A0(\game.fsm.seq[0][1] ),
    .A1(\game.fsm.seq[2][1] ),
    .A2(\game.fsm.seq[1][1] ),
    .A3(\game.fsm.seq[3][1] ),
    .S1(_0007_),
    .X(_1261_));
 sg13g2_nor2_1 _3953_ (.A(_0009_),
    .B(_1261_),
    .Y(_1262_));
 sg13g2_nor2_2 _3954_ (.A(_1260_),
    .B(_1262_),
    .Y(_1263_));
 sg13g2_or2_1 _3955_ (.X(_1264_),
    .B(_1263_),
    .A(_1255_));
 sg13g2_o21ai_1 _3956_ (.B1(_1236_),
    .Y(_1265_),
    .A1(_1246_),
    .A2(_1264_));
 sg13g2_inv_1 _3957_ (.Y(_1266_),
    .A(_1265_));
 sg13g2_o21ai_1 _3958_ (.B1(net433),
    .Y(_1267_),
    .A1(net783),
    .A2(net342));
 sg13g2_a21oi_1 _3959_ (.A1(net342),
    .A2(_1266_),
    .Y(_0240_),
    .B1(_1267_));
 sg13g2_nor3_1 _3960_ (.A(_0581_),
    .B(net371),
    .C(_0696_),
    .Y(_1268_));
 sg13g2_nand2_1 _3961_ (.Y(_1269_),
    .A(_1237_),
    .B(_1245_));
 sg13g2_o21ai_1 _3962_ (.B1(net342),
    .Y(_1270_),
    .A1(_1264_),
    .A2(_1269_));
 sg13g2_nor2_1 _3963_ (.A(_1268_),
    .B(_1270_),
    .Y(_1271_));
 sg13g2_o21ai_1 _3964_ (.B1(net433),
    .Y(_1272_),
    .A1(net754),
    .A2(net342));
 sg13g2_nor2_1 _3965_ (.A(_1271_),
    .B(_1272_),
    .Y(_0241_));
 sg13g2_nand2b_1 _3966_ (.Y(_1273_),
    .B(_1263_),
    .A_N(_1255_));
 sg13g2_nand2_1 _3967_ (.Y(_1274_),
    .A(net350),
    .B(_0696_));
 sg13g2_o21ai_1 _3968_ (.B1(_1274_),
    .Y(_1275_),
    .A1(_1246_),
    .A2(_1273_));
 sg13g2_a21oi_1 _3969_ (.A1(_1212_),
    .A2(_1275_),
    .Y(_1276_),
    .B1(net418));
 sg13g2_o21ai_1 _3970_ (.B1(_1276_),
    .Y(_0242_),
    .A1(_1805_),
    .A2(net342));
 sg13g2_nor2_1 _3971_ (.A(_0595_),
    .B(_0702_),
    .Y(_1277_));
 sg13g2_o21ai_1 _3972_ (.B1(net342),
    .Y(_1278_),
    .A1(_1269_),
    .A2(_1273_));
 sg13g2_nor2_1 _3973_ (.A(net734),
    .B(net342),
    .Y(_1279_));
 sg13g2_o21ai_1 _3974_ (.B1(net433),
    .Y(_1280_),
    .A1(_1277_),
    .A2(_1278_));
 sg13g2_nor2_1 _3975_ (.A(_1279_),
    .B(_1280_),
    .Y(_0243_));
 sg13g2_nand2_1 _3976_ (.Y(_1281_),
    .A(net354),
    .B(_0980_));
 sg13g2_xor2_1 _3977_ (.B(_1281_),
    .A(net706),
    .X(_1282_));
 sg13g2_nor2_1 _3978_ (.A(net357),
    .B(_1282_),
    .Y(_0244_));
 sg13g2_nand2_1 _3979_ (.Y(_1283_),
    .A(net366),
    .B(_1281_));
 sg13g2_mux2_1 _3980_ (.A0(net505),
    .A1(_0988_),
    .S(_1283_),
    .X(_0245_));
 sg13g2_nand2b_1 _3981_ (.Y(_1284_),
    .B(_0787_),
    .A_N(_0788_));
 sg13g2_or2_1 _3982_ (.X(_1285_),
    .B(_1284_),
    .A(_0790_));
 sg13g2_nand3_1 _3983_ (.B(net364),
    .C(_1285_),
    .A(net512),
    .Y(_1286_));
 sg13g2_o21ai_1 _3984_ (.B1(_1286_),
    .Y(_0246_),
    .A1(net344),
    .A2(_1285_));
 sg13g2_nand3_1 _3985_ (.B(net364),
    .C(_1285_),
    .A(net711),
    .Y(_1287_));
 sg13g2_o21ai_1 _3986_ (.B1(_1287_),
    .Y(_0247_),
    .A1(net343),
    .A2(_1285_));
 sg13g2_nand2_1 _3987_ (.Y(_1288_),
    .A(net352),
    .B(_0978_));
 sg13g2_xor2_1 _3988_ (.B(_1288_),
    .A(net668),
    .X(_1289_));
 sg13g2_nor2_1 _3989_ (.A(net357),
    .B(_1289_),
    .Y(_0248_));
 sg13g2_a21oi_1 _3990_ (.A1(net352),
    .A2(_0978_),
    .Y(_1290_),
    .B1(net357));
 sg13g2_mux2_1 _3991_ (.A0(_0988_),
    .A1(net587),
    .S(_1290_),
    .X(_0249_));
 sg13g2_nand2_1 _3992_ (.Y(_1291_),
    .A(net367),
    .B(_0750_));
 sg13g2_nand3_1 _3993_ (.B(_0752_),
    .C(_1291_),
    .A(_0751_),
    .Y(_1292_));
 sg13g2_nor3_1 _3994_ (.A(_0750_),
    .B(_0756_),
    .C(_1292_),
    .Y(_1293_));
 sg13g2_a21o_1 _3995_ (.A2(_1292_),
    .A1(net571),
    .B1(_1293_),
    .X(_0250_));
 sg13g2_mux2_1 _3996_ (.A0(_0765_),
    .A1(net614),
    .S(_1292_),
    .X(_0251_));
 sg13g2_nor2_2 _3997_ (.A(_0520_),
    .B(_0751_),
    .Y(_1294_));
 sg13g2_o21ai_1 _3998_ (.B1(net367),
    .Y(_1295_),
    .A1(net522),
    .A2(_1294_));
 sg13g2_a21oi_1 _3999_ (.A1(net522),
    .A2(_1294_),
    .Y(_0252_),
    .B1(_1295_));
 sg13g2_nor2_1 _4000_ (.A(net357),
    .B(_1294_),
    .Y(_1296_));
 sg13g2_mux2_1 _4001_ (.A0(_0765_),
    .A1(net623),
    .S(_1296_),
    .X(_0253_));
 sg13g2_nor2_2 _4002_ (.A(_0510_),
    .B(_0752_),
    .Y(_1297_));
 sg13g2_o21ai_1 _4003_ (.B1(net367),
    .Y(_1298_),
    .A1(net533),
    .A2(_1297_));
 sg13g2_a21oi_1 _4004_ (.A1(net533),
    .A2(_1297_),
    .Y(_0254_),
    .B1(_1298_));
 sg13g2_nor2_1 _4005_ (.A(net357),
    .B(_1297_),
    .Y(_1299_));
 sg13g2_mux2_1 _4006_ (.A0(_0765_),
    .A1(net633),
    .S(_1299_),
    .X(_0255_));
 sg13g2_nand2_1 _4007_ (.Y(_1300_),
    .A(_0520_),
    .B(_0978_));
 sg13g2_o21ai_1 _4008_ (.B1(net367),
    .Y(_1301_),
    .A1(_1876_),
    .A2(_1300_));
 sg13g2_a21oi_1 _4009_ (.A1(_1876_),
    .A2(_1300_),
    .Y(_0256_),
    .B1(_1301_));
 sg13g2_nand2_1 _4010_ (.Y(_1302_),
    .A(net366),
    .B(_1300_));
 sg13g2_mux2_1 _4011_ (.A0(net513),
    .A1(_0988_),
    .S(_1302_),
    .X(_0257_));
 sg13g2_nor2_1 _4012_ (.A(net356),
    .B(_0997_),
    .Y(_1303_));
 sg13g2_a21oi_2 _4013_ (.B1(_0989_),
    .Y(_1304_),
    .A2(_1303_),
    .A1(_0995_));
 sg13g2_nor2_1 _4014_ (.A(net356),
    .B(_1006_),
    .Y(_1305_));
 sg13g2_mux2_1 _4015_ (.A0(net600),
    .A1(_1305_),
    .S(_1304_),
    .X(_0258_));
 sg13g2_mux2_1 _4016_ (.A0(net511),
    .A1(_1012_),
    .S(_1304_),
    .X(_0259_));
 sg13g2_mux2_1 _4017_ (.A0(net480),
    .A1(_1020_),
    .S(_1304_),
    .X(_0260_));
 sg13g2_nand2b_2 _4018_ (.Y(_1306_),
    .B(_0819_),
    .A_N(_0879_));
 sg13g2_nand3_1 _4019_ (.B(net361),
    .C(_1306_),
    .A(net487),
    .Y(_1307_));
 sg13g2_o21ai_1 _4020_ (.B1(_1307_),
    .Y(_0261_),
    .A1(_0822_),
    .A2(_1306_));
 sg13g2_nand3_1 _4021_ (.B(net361),
    .C(_1306_),
    .A(net516),
    .Y(_1308_));
 sg13g2_o21ai_1 _4022_ (.B1(_1308_),
    .Y(_0262_),
    .A1(_0827_),
    .A2(_1306_));
 sg13g2_nand3_1 _4023_ (.B(net361),
    .C(_1306_),
    .A(net556),
    .Y(_1309_));
 sg13g2_o21ai_1 _4024_ (.B1(_1309_),
    .Y(_0263_),
    .A1(_0835_),
    .A2(_1306_));
 sg13g2_nand2b_1 _4025_ (.Y(_1310_),
    .B(_0790_),
    .A_N(_0973_));
 sg13g2_nand2_1 _4026_ (.Y(_1311_),
    .A(net590),
    .B(_1310_));
 sg13g2_o21ai_1 _4027_ (.B1(_1311_),
    .Y(_0264_),
    .A1(net344),
    .A2(_1310_));
 sg13g2_nand2_1 _4028_ (.Y(_1312_),
    .A(net584),
    .B(_1310_));
 sg13g2_o21ai_1 _4029_ (.B1(_1312_),
    .Y(_0265_),
    .A1(net343),
    .A2(_1310_));
 sg13g2_a22oi_1 _4030_ (.Y(_1313_),
    .B1(_1229_),
    .B2(net589),
    .A2(_0610_),
    .A1(_0606_));
 sg13g2_nand2_1 _4031_ (.Y(_1314_),
    .A(net370),
    .B(_1200_));
 sg13g2_mux2_1 _4032_ (.A0(_1184_),
    .A1(_1185_),
    .S(_0581_),
    .X(_1315_));
 sg13g2_nor3_1 _4033_ (.A(_1199_),
    .B(_1314_),
    .C(_1315_),
    .Y(_1316_));
 sg13g2_or3_1 _4034_ (.A(_0614_),
    .B(_1313_),
    .C(_1316_),
    .X(_1317_));
 sg13g2_nand2b_1 _4035_ (.Y(_1318_),
    .B(_1252_),
    .A_N(_1159_));
 sg13g2_o21ai_1 _4036_ (.B1(\game.counter[2] ),
    .Y(_1319_),
    .A1(\game.counter[1] ),
    .A2(\game.counter[0] ));
 sg13g2_o21ai_1 _4037_ (.B1(_1800_),
    .Y(_1320_),
    .A1(_1318_),
    .A2(_1319_));
 sg13g2_a21oi_1 _4038_ (.A1(_1166_),
    .A2(_1320_),
    .Y(_1321_),
    .B1(_1158_));
 sg13g2_nand2_1 _4039_ (.Y(_1322_),
    .A(net370),
    .B(_1203_));
 sg13g2_a21oi_1 _4040_ (.A1(_1860_),
    .A2(_1171_),
    .Y(_1323_),
    .B1(_1321_));
 sg13g2_nor3_1 _4041_ (.A(\game.solver_trigger_delayed ),
    .B(\game.slv.ready ),
    .C(_0924_),
    .Y(_1324_));
 sg13g2_a21o_1 _4042_ (.A2(_1210_),
    .A1(_0895_),
    .B1(_1802_),
    .X(_1325_));
 sg13g2_a21oi_2 _4043_ (.B1(net371),
    .Y(_1326_),
    .A2(_1202_),
    .A1(_1201_));
 sg13g2_a22oi_1 _4044_ (.Y(_1327_),
    .B1(_1172_),
    .B2(_0080_),
    .A2(_0923_),
    .A1(\game.solver_trigger_delayed ));
 sg13g2_nand3_1 _4045_ (.B(_1325_),
    .C(_1327_),
    .A(_1231_),
    .Y(_1328_));
 sg13g2_or2_1 _4046_ (.X(_1329_),
    .B(_1191_),
    .A(_1119_));
 sg13g2_nor4_1 _4047_ (.A(_1324_),
    .B(_1326_),
    .C(_1328_),
    .D(_1329_),
    .Y(_1330_));
 sg13g2_nand4_1 _4048_ (.B(_1322_),
    .C(_1323_),
    .A(_1196_),
    .Y(_1331_),
    .D(_1330_));
 sg13g2_inv_1 _4049_ (.Y(_1332_),
    .A(_1331_));
 sg13g2_nor3_1 _4050_ (.A(net350),
    .B(_0923_),
    .C(_1331_),
    .Y(_1333_));
 sg13g2_o21ai_1 _4051_ (.B1(net429),
    .Y(_1334_),
    .A1(net383),
    .A2(_1332_));
 sg13g2_a21oi_1 _4052_ (.A1(_1317_),
    .A2(_1333_),
    .Y(_0266_),
    .B1(_1334_));
 sg13g2_nand2_1 _4053_ (.Y(_1335_),
    .A(net586),
    .B(_1331_));
 sg13g2_nor2_1 _4054_ (.A(_0589_),
    .B(_1313_),
    .Y(_1336_));
 sg13g2_mux2_1 _4055_ (.A0(_1185_),
    .A1(_1184_),
    .S(_0581_),
    .X(_1337_));
 sg13g2_o21ai_1 _4056_ (.B1(_1336_),
    .Y(_1338_),
    .A1(_1314_),
    .A2(_1337_));
 sg13g2_o21ai_1 _4057_ (.B1(_1332_),
    .Y(_1339_),
    .A1(net371),
    .A2(_1198_));
 sg13g2_a21o_1 _4058_ (.A2(_1338_),
    .A1(_0593_),
    .B1(_1339_),
    .X(_1340_));
 sg13g2_a21oi_1 _4059_ (.A1(_1335_),
    .A2(_1340_),
    .Y(_0267_),
    .B1(net411));
 sg13g2_o21ai_1 _4060_ (.B1(net370),
    .Y(_1341_),
    .A1(_1113_),
    .A2(_1199_));
 sg13g2_nand2_1 _4061_ (.Y(_1342_),
    .A(net767),
    .B(_1229_));
 sg13g2_a22oi_1 _4062_ (.Y(_1343_),
    .B1(_0611_),
    .B2(_1342_),
    .A2(_0589_),
    .A1(net381));
 sg13g2_a22oi_1 _4063_ (.Y(_1344_),
    .B1(_1341_),
    .B2(_1343_),
    .A2(_1157_),
    .A1(net463));
 sg13g2_or2_1 _4064_ (.X(_1345_),
    .B(_1344_),
    .A(_0592_));
 sg13g2_a21oi_1 _4065_ (.A1(_1124_),
    .A2(_1198_),
    .Y(_1346_),
    .B1(_1331_));
 sg13g2_a221oi_1 _4066_ (.B2(_1346_),
    .C1(net411),
    .B1(_1345_),
    .A1(_1803_),
    .Y(_0268_),
    .A2(_1331_));
 sg13g2_o21ai_1 _4067_ (.B1(net432),
    .Y(_1347_),
    .A1(_1230_),
    .A2(_1331_));
 sg13g2_a21oi_1 _4068_ (.A1(_1802_),
    .A2(_1331_),
    .Y(_0269_),
    .B1(_1347_));
 sg13g2_a21o_1 _4069_ (.A2(_1199_),
    .A1(net372),
    .B1(_0589_),
    .X(_1348_));
 sg13g2_a22oi_1 _4070_ (.Y(_1349_),
    .B1(_1198_),
    .B2(net350),
    .A2(_0923_),
    .A1(_1883_));
 sg13g2_nand3_1 _4071_ (.B(_1348_),
    .C(_1349_),
    .A(_1327_),
    .Y(_1350_));
 sg13g2_a21oi_1 _4072_ (.A1(_1166_),
    .A2(_1169_),
    .Y(_1351_),
    .B1(_1162_));
 sg13g2_nor2_1 _4073_ (.A(_1173_),
    .B(_1351_),
    .Y(_1352_));
 sg13g2_o21ai_1 _4074_ (.B1(net427),
    .Y(_1353_),
    .A1(_1350_),
    .A2(_1352_));
 sg13g2_xor2_1 _4075_ (.B(_1350_),
    .A(net755),
    .X(_1354_));
 sg13g2_nor2b_2 _4076_ (.A(_1350_),
    .B_N(_1352_),
    .Y(_1355_));
 sg13g2_nor2_1 _4077_ (.A(_1353_),
    .B(_1354_),
    .Y(_0270_));
 sg13g2_a22oi_1 _4078_ (.Y(_1356_),
    .B1(_1355_),
    .B2(_1247_),
    .A2(_1350_),
    .A1(net737));
 sg13g2_o21ai_1 _4079_ (.B1(net427),
    .Y(_1357_),
    .A1(net737),
    .A2(\game.counter[0] ));
 sg13g2_nor2_1 _4080_ (.A(net738),
    .B(_1357_),
    .Y(_0271_));
 sg13g2_nor2_1 _4081_ (.A(_1247_),
    .B(_1350_),
    .Y(_1358_));
 sg13g2_nor2_1 _4082_ (.A(net729),
    .B(_1358_),
    .Y(_1359_));
 sg13g2_and2_1 _4083_ (.A(net729),
    .B(_1358_),
    .X(_1360_));
 sg13g2_nor3_1 _4084_ (.A(_1353_),
    .B(net730),
    .C(_1360_),
    .Y(_0272_));
 sg13g2_xnor2_1 _4085_ (.Y(_1361_),
    .A(net705),
    .B(_1360_));
 sg13g2_nor2_1 _4086_ (.A(_1353_),
    .B(_1361_),
    .Y(_0273_));
 sg13g2_a22oi_1 _4087_ (.Y(_1362_),
    .B1(_1355_),
    .B2(_1249_),
    .A2(_1350_),
    .A1(net642));
 sg13g2_nor2_1 _4088_ (.A(net412),
    .B(net643),
    .Y(_0274_));
 sg13g2_a21oi_1 _4089_ (.A1(_1252_),
    .A2(_1360_),
    .Y(_1363_),
    .B1(net546));
 sg13g2_and3_1 _4090_ (.X(_1364_),
    .A(net546),
    .B(_1252_),
    .C(_1360_));
 sg13g2_nor3_1 _4091_ (.A(_1353_),
    .B(net547),
    .C(_1364_),
    .Y(_0275_));
 sg13g2_xnor2_1 _4092_ (.Y(_1365_),
    .A(net611),
    .B(_1364_));
 sg13g2_nor2_1 _4093_ (.A(_1353_),
    .B(_1365_),
    .Y(_0276_));
 sg13g2_nor3_1 _4094_ (.A(_1801_),
    .B(_1159_),
    .C(_1248_),
    .Y(_1366_));
 sg13g2_xnor2_1 _4095_ (.Y(_1367_),
    .A(_0058_),
    .B(_1366_));
 sg13g2_a22oi_1 _4096_ (.Y(_1368_),
    .B1(_1355_),
    .B2(_1367_),
    .A2(_1350_),
    .A1(net536));
 sg13g2_nor2_1 _4097_ (.A(net411),
    .B(net537),
    .Y(_0277_));
 sg13g2_o21ai_1 _4098_ (.B1(net350),
    .Y(_1369_),
    .A1(_1195_),
    .A2(_1219_));
 sg13g2_nand4_1 _4099_ (.B(_1314_),
    .C(_1322_),
    .A(_0922_),
    .Y(_1370_),
    .D(_1369_));
 sg13g2_a21o_1 _4100_ (.A2(_0924_),
    .A1(_0611_),
    .B1(_1370_),
    .X(_1371_));
 sg13g2_nand3_1 _4101_ (.B(_0609_),
    .C(_0613_),
    .A(net432),
    .Y(_1372_));
 sg13g2_a21oi_1 _4102_ (.A1(_1799_),
    .A2(_1371_),
    .Y(_0278_),
    .B1(_1372_));
 sg13g2_o21ai_1 _4103_ (.B1(net432),
    .Y(_1373_),
    .A1(_1126_),
    .A2(_1371_));
 sg13g2_a21oi_1 _4104_ (.A1(_1798_),
    .A2(_1371_),
    .Y(_0279_),
    .B1(_1373_));
 sg13g2_a21oi_1 _4105_ (.A1(net651),
    .A2(net335),
    .Y(_0283_),
    .B1(net420));
 sg13g2_nand2b_2 _4106_ (.Y(_1374_),
    .B(net430),
    .A_N(_0921_));
 sg13g2_nor2_1 _4107_ (.A(_1893_),
    .B(_1374_),
    .Y(_0284_));
 sg13g2_xnor2_1 _4108_ (.Y(_1375_),
    .A(\clk_div_counter[0] ),
    .B(net620));
 sg13g2_nor2_1 _4109_ (.A(_1374_),
    .B(net621),
    .Y(_0285_));
 sg13g2_and3_1 _4110_ (.X(_1376_),
    .A(\clk_div_counter[0] ),
    .B(\clk_div_counter[1] ),
    .C(net460));
 sg13g2_a21oi_1 _4111_ (.A1(\clk_div_counter[0] ),
    .A2(\clk_div_counter[1] ),
    .Y(_1377_),
    .B1(net460));
 sg13g2_nor3_1 _4112_ (.A(_1374_),
    .B(_1376_),
    .C(net461),
    .Y(_0286_));
 sg13g2_and2_1 _4113_ (.A(net494),
    .B(_1376_),
    .X(_1378_));
 sg13g2_nor2_1 _4114_ (.A(net494),
    .B(_1376_),
    .Y(_1379_));
 sg13g2_nor3_1 _4115_ (.A(_1374_),
    .B(_1378_),
    .C(net495),
    .Y(_0287_));
 sg13g2_and2_1 _4116_ (.A(net534),
    .B(_1378_),
    .X(_1380_));
 sg13g2_nor2_1 _4117_ (.A(net534),
    .B(_1378_),
    .Y(_1381_));
 sg13g2_nor3_1 _4118_ (.A(_1374_),
    .B(_1380_),
    .C(_1381_),
    .Y(_0288_));
 sg13g2_nor2_1 _4119_ (.A(net544),
    .B(_1380_),
    .Y(_1382_));
 sg13g2_and2_1 _4120_ (.A(net544),
    .B(_1380_),
    .X(_1383_));
 sg13g2_nor3_1 _4121_ (.A(_1374_),
    .B(_1382_),
    .C(_1383_),
    .Y(_0289_));
 sg13g2_nor2_1 _4122_ (.A(net530),
    .B(_1383_),
    .Y(_1384_));
 sg13g2_and2_1 _4123_ (.A(net530),
    .B(_1383_),
    .X(_1385_));
 sg13g2_nor3_1 _4124_ (.A(_1374_),
    .B(net531),
    .C(_1385_),
    .Y(_0290_));
 sg13g2_a21oi_1 _4125_ (.A1(net604),
    .A2(_1385_),
    .Y(_1386_),
    .B1(_1374_));
 sg13g2_o21ai_1 _4126_ (.B1(_1386_),
    .Y(_1387_),
    .A1(net604),
    .A2(_1385_));
 sg13g2_inv_1 _4127_ (.Y(_0291_),
    .A(_1387_));
 sg13g2_nor4_1 _4128_ (.A(\game.state[3] ),
    .B(net381),
    .C(net384),
    .D(_1202_),
    .Y(_1388_));
 sg13g2_a21oi_1 _4129_ (.A1(_0013_),
    .A2(_1388_),
    .Y(_1389_),
    .B1(net418));
 sg13g2_o21ai_1 _4130_ (.B1(_1389_),
    .Y(_0292_),
    .A1(_1797_),
    .A2(_1388_));
 sg13g2_nand3_1 _4131_ (.B(\btn.sample_10ms[2] ),
    .C(\btn.sample_15ms[2] ),
    .A(net721),
    .Y(_1390_));
 sg13g2_xnor2_1 _4132_ (.Y(_1391_),
    .A(net557),
    .B(net3));
 sg13g2_nand3_1 _4133_ (.B(\btn.sample_10ms[0] ),
    .C(\btn.sample_15ms[0] ),
    .A(\btn.sample_5ms[0] ),
    .Y(_1392_));
 sg13g2_xor2_1 _4134_ (.B(net1),
    .A(net497),
    .X(_1393_));
 sg13g2_nand2b_1 _4135_ (.Y(_1394_),
    .B(_1393_),
    .A_N(_1392_));
 sg13g2_o21ai_1 _4136_ (.B1(_1394_),
    .Y(_1395_),
    .A1(_1390_),
    .A2(_1391_));
 sg13g2_nand3_1 _4137_ (.B(\btn.sample_10ms[3] ),
    .C(\btn.sample_15ms[3] ),
    .A(\btn.sample_5ms[3] ),
    .Y(_1396_));
 sg13g2_xnor2_1 _4138_ (.Y(_1397_),
    .A(\btn.button_state[3] ),
    .B(net4));
 sg13g2_nor2_1 _4139_ (.A(_1396_),
    .B(_1397_),
    .Y(_1398_));
 sg13g2_nand3_1 _4140_ (.B(\btn.sample_10ms[1] ),
    .C(\btn.sample_15ms[1] ),
    .A(\btn.sample_5ms[1] ),
    .Y(_1399_));
 sg13g2_xnor2_1 _4141_ (.Y(_1400_),
    .A(net477),
    .B(net2));
 sg13g2_nor2_1 _4142_ (.A(_1399_),
    .B(_1400_),
    .Y(_1401_));
 sg13g2_nor3_2 _4143_ (.A(_1395_),
    .B(_1398_),
    .C(_1401_),
    .Y(_1402_));
 sg13g2_nor2_1 _4144_ (.A(net3),
    .B(_1390_),
    .Y(_1403_));
 sg13g2_a21oi_1 _4145_ (.A1(_1784_),
    .A2(_1390_),
    .Y(_1404_),
    .B1(_1403_));
 sg13g2_or2_1 _4146_ (.X(_1405_),
    .B(_1404_),
    .A(_1402_));
 sg13g2_mux2_1 _4147_ (.A0(net2),
    .A1(\btn.button_state[1] ),
    .S(_1399_),
    .X(_1406_));
 sg13g2_nor2_1 _4148_ (.A(net376),
    .B(net478),
    .Y(_1407_));
 sg13g2_nor2_1 _4149_ (.A(net4),
    .B(_1396_),
    .Y(_1408_));
 sg13g2_a21oi_1 _4150_ (.A1(_1783_),
    .A2(_1396_),
    .Y(_1409_),
    .B1(_1408_));
 sg13g2_nor2_1 _4151_ (.A(net1),
    .B(_1392_),
    .Y(_1410_));
 sg13g2_a21oi_1 _4152_ (.A1(_1785_),
    .A2(_1392_),
    .Y(_1411_),
    .B1(_1410_));
 sg13g2_nor4_1 _4153_ (.A(net374),
    .B(_1406_),
    .C(_1409_),
    .D(_1411_),
    .Y(_1412_));
 sg13g2_nand2b_2 _4154_ (.Y(_1413_),
    .B(_1412_),
    .A_N(_1405_));
 sg13g2_nand2_2 _4155_ (.Y(_1414_),
    .A(net431),
    .B(_1413_));
 sg13g2_nor3_1 _4156_ (.A(\btn.button_state[3] ),
    .B(\btn.button_state[2] ),
    .C(\btn.button_state[1] ),
    .Y(_1415_));
 sg13g2_a21oi_2 _4157_ (.B1(net374),
    .Y(_1416_),
    .A2(_1415_),
    .A1(_1785_));
 sg13g2_nand2_2 _4158_ (.Y(_1417_),
    .A(_1402_),
    .B(_1416_));
 sg13g2_nand3_1 _4159_ (.B(\btn.change_timer[3] ),
    .C(\btn.change_timer[2] ),
    .A(\btn.change_timer[4] ),
    .Y(_1418_));
 sg13g2_nand2b_1 _4160_ (.Y(_1419_),
    .B(net576),
    .A_N(\btn.change_timer[6] ));
 sg13g2_nor4_2 _4161_ (.A(net514),
    .B(\btn.change_timer[0] ),
    .C(_1418_),
    .Y(_1420_),
    .D(_1419_));
 sg13g2_nand4_1 _4162_ (.B(_1402_),
    .C(_1416_),
    .A(net431),
    .Y(_1421_),
    .D(net515));
 sg13g2_o21ai_1 _4163_ (.B1(_1421_),
    .Y(_0293_),
    .A1(_1796_),
    .A2(_1414_));
 sg13g2_nand2b_1 _4164_ (.Y(_1422_),
    .B(net405),
    .A_N(_1402_));
 sg13g2_nand3_1 _4165_ (.B(_1416_),
    .C(_1420_),
    .A(net452),
    .Y(_1423_));
 sg13g2_nor2b_2 _4166_ (.A(_1416_),
    .B_N(_1422_),
    .Y(_1424_));
 sg13g2_nand2_1 _4167_ (.Y(_1425_),
    .A(_1422_),
    .B(_1423_));
 sg13g2_o21ai_1 _4168_ (.B1(_1425_),
    .Y(_1426_),
    .A1(_1402_),
    .A2(_1411_));
 sg13g2_a21oi_1 _4169_ (.A1(_1795_),
    .A2(_1426_),
    .Y(_0294_),
    .B1(_1414_));
 sg13g2_o21ai_1 _4170_ (.B1(_1425_),
    .Y(_1427_),
    .A1(_1402_),
    .A2(_1406_));
 sg13g2_a21oi_1 _4171_ (.A1(_1794_),
    .A2(_1427_),
    .Y(_0295_),
    .B1(_1414_));
 sg13g2_a21oi_1 _4172_ (.A1(_1405_),
    .A2(_1425_),
    .Y(_1428_),
    .B1(net332));
 sg13g2_nor2_1 _4173_ (.A(_1414_),
    .B(_1428_),
    .Y(_0296_));
 sg13g2_o21ai_1 _4174_ (.B1(_1425_),
    .Y(_1429_),
    .A1(_1402_),
    .A2(_1409_));
 sg13g2_a21oi_1 _4175_ (.A1(_1792_),
    .A2(_1429_),
    .Y(_0297_),
    .B1(_1414_));
 sg13g2_nand2_1 _4176_ (.Y(_1430_),
    .A(\btn.change_timer[1] ),
    .B(\btn.change_timer[0] ));
 sg13g2_nand3_1 _4177_ (.B(\btn.change_timer[1] ),
    .C(\btn.change_timer[0] ),
    .A(\btn.change_timer[2] ),
    .Y(_1431_));
 sg13g2_nor2_1 _4178_ (.A(_1791_),
    .B(_1431_),
    .Y(_1432_));
 sg13g2_nor2_1 _4179_ (.A(_1418_),
    .B(_1430_),
    .Y(_1433_));
 sg13g2_nand2_1 _4180_ (.Y(_1434_),
    .A(net576),
    .B(_1433_));
 sg13g2_nand3_1 _4181_ (.B(net686),
    .C(_1433_),
    .A(net634),
    .Y(_1435_));
 sg13g2_a21oi_1 _4182_ (.A1(net692),
    .A2(_1435_),
    .Y(_1436_),
    .B1(_1417_));
 sg13g2_a21oi_1 _4183_ (.A1(net692),
    .A2(_1424_),
    .Y(_1437_),
    .B1(_1436_));
 sg13g2_nor2_1 _4184_ (.A(net416),
    .B(_1437_),
    .Y(_0298_));
 sg13g2_xnor2_1 _4185_ (.Y(_1438_),
    .A(net514),
    .B(\btn.change_timer[0] ));
 sg13g2_a21oi_1 _4186_ (.A1(_1435_),
    .A2(_1438_),
    .Y(_1439_),
    .B1(_1417_));
 sg13g2_a21oi_1 _4187_ (.A1(net514),
    .A2(_1424_),
    .Y(_1440_),
    .B1(net687));
 sg13g2_nor2_1 _4188_ (.A(net416),
    .B(_1440_),
    .Y(_0299_));
 sg13g2_xor2_1 _4189_ (.B(_1430_),
    .A(net596),
    .X(_1441_));
 sg13g2_a21oi_1 _4190_ (.A1(_1435_),
    .A2(_1441_),
    .Y(_1442_),
    .B1(_1417_));
 sg13g2_a21oi_1 _4191_ (.A1(net596),
    .A2(_1424_),
    .Y(_1443_),
    .B1(_1442_));
 sg13g2_nor2_1 _4192_ (.A(net415),
    .B(net597),
    .Y(_0300_));
 sg13g2_xor2_1 _4193_ (.B(_1431_),
    .A(net638),
    .X(_1444_));
 sg13g2_a21oi_1 _4194_ (.A1(_1435_),
    .A2(_1444_),
    .Y(_1445_),
    .B1(_1417_));
 sg13g2_a21oi_1 _4195_ (.A1(net638),
    .A2(_1424_),
    .Y(_1446_),
    .B1(_1445_));
 sg13g2_nor2_1 _4196_ (.A(net415),
    .B(net639),
    .Y(_0301_));
 sg13g2_nor2_1 _4197_ (.A(_1417_),
    .B(_1433_),
    .Y(_1447_));
 sg13g2_o21ai_1 _4198_ (.B1(_1447_),
    .Y(_1448_),
    .A1(net697),
    .A2(_1432_));
 sg13g2_nor2_1 _4199_ (.A(_1417_),
    .B(_1435_),
    .Y(_1449_));
 sg13g2_a21oi_1 _4200_ (.A1(net697),
    .A2(_1424_),
    .Y(_1450_),
    .B1(_1449_));
 sg13g2_a21oi_1 _4201_ (.A1(_1448_),
    .A2(_1450_),
    .Y(_0302_),
    .B1(net415));
 sg13g2_o21ai_1 _4202_ (.B1(net576),
    .Y(_1451_),
    .A1(_1424_),
    .A2(_1447_));
 sg13g2_nand4_1 _4203_ (.B(_1416_),
    .C(_1419_),
    .A(_1402_),
    .Y(_1452_),
    .D(_1433_));
 sg13g2_a21oi_1 _4204_ (.A1(_1451_),
    .A2(_1452_),
    .Y(_0303_),
    .B1(net416));
 sg13g2_nor2_1 _4205_ (.A(_1424_),
    .B(_1434_),
    .Y(_1453_));
 sg13g2_o21ai_1 _4206_ (.B1(_1422_),
    .Y(_1454_),
    .A1(net634),
    .A2(_1453_));
 sg13g2_nor2_1 _4207_ (.A(net416),
    .B(_1454_),
    .Y(_0304_));
 sg13g2_o21ai_1 _4208_ (.B1(net437),
    .Y(_1455_),
    .A1(net406),
    .A2(\btn.sample_15ms[0] ));
 sg13g2_a21oi_1 _4209_ (.A1(net406),
    .A2(_1790_),
    .Y(_0305_),
    .B1(_1455_));
 sg13g2_o21ai_1 _4210_ (.B1(net436),
    .Y(_1456_),
    .A1(net407),
    .A2(\btn.sample_15ms[1] ));
 sg13g2_a21oi_1 _4211_ (.A1(net407),
    .A2(_1789_),
    .Y(_0306_),
    .B1(_1456_));
 sg13g2_o21ai_1 _4212_ (.B1(net436),
    .Y(_1457_),
    .A1(net406),
    .A2(\btn.sample_15ms[2] ));
 sg13g2_a21oi_1 _4213_ (.A1(net406),
    .A2(_1788_),
    .Y(_0307_),
    .B1(_1457_));
 sg13g2_o21ai_1 _4214_ (.B1(net435),
    .Y(_1458_),
    .A1(net405),
    .A2(net474));
 sg13g2_a21oi_1 _4215_ (.A1(net405),
    .A2(_1787_),
    .Y(_0308_),
    .B1(_1458_));
 sg13g2_o21ai_1 _4216_ (.B1(net437),
    .Y(_1459_),
    .A1(net405),
    .A2(net490));
 sg13g2_a21oi_1 _4217_ (.A1(net406),
    .A2(_1786_),
    .Y(_0309_),
    .B1(_1459_));
 sg13g2_o21ai_1 _4218_ (.B1(net436),
    .Y(_1460_),
    .A1(net376),
    .A2(net527));
 sg13g2_a21oi_1 _4219_ (.A1(net376),
    .A2(_1789_),
    .Y(_0310_),
    .B1(_1460_));
 sg13g2_o21ai_1 _4220_ (.B1(net436),
    .Y(_1461_),
    .A1(net375),
    .A2(net526));
 sg13g2_a21oi_1 _4221_ (.A1(net375),
    .A2(_1788_),
    .Y(_0311_),
    .B1(_1461_));
 sg13g2_o21ai_1 _4222_ (.B1(net435),
    .Y(_1462_),
    .A1(net375),
    .A2(\btn.sample_5ms[3] ));
 sg13g2_a21oi_1 _4223_ (.A1(net375),
    .A2(_1787_),
    .Y(_0312_),
    .B1(_1462_));
 sg13g2_o21ai_1 _4224_ (.B1(net435),
    .Y(_1463_),
    .A1(net375),
    .A2(_1393_));
 sg13g2_a21oi_1 _4225_ (.A1(net378),
    .A2(_1786_),
    .Y(_0313_),
    .B1(_1463_));
 sg13g2_o21ai_1 _4226_ (.B1(net436),
    .Y(_1464_),
    .A1(net407),
    .A2(net527));
 sg13g2_a21oi_1 _4227_ (.A1(net407),
    .A2(_1400_),
    .Y(_0314_),
    .B1(_1464_));
 sg13g2_o21ai_1 _4228_ (.B1(net435),
    .Y(_1465_),
    .A1(net405),
    .A2(net526));
 sg13g2_a21oi_1 _4229_ (.A1(net405),
    .A2(_1391_),
    .Y(_0315_),
    .B1(_1465_));
 sg13g2_o21ai_1 _4230_ (.B1(net435),
    .Y(_1466_),
    .A1(net405),
    .A2(net630));
 sg13g2_a21oi_1 _4231_ (.A1(net405),
    .A2(_1397_),
    .Y(_0316_),
    .B1(_1466_));
 sg13g2_o21ai_1 _4232_ (.B1(net435),
    .Y(_1467_),
    .A1(net374),
    .A2(_1411_));
 sg13g2_a21oi_1 _4233_ (.A1(net374),
    .A2(_1785_),
    .Y(_0317_),
    .B1(_1467_));
 sg13g2_o21ai_1 _4234_ (.B1(net436),
    .Y(_1468_),
    .A1(net407),
    .A2(net477));
 sg13g2_nor2_1 _4235_ (.A(_1407_),
    .B(_1468_),
    .Y(_0318_));
 sg13g2_o21ai_1 _4236_ (.B1(net435),
    .Y(_1469_),
    .A1(net374),
    .A2(_1404_));
 sg13g2_a21oi_1 _4237_ (.A1(net374),
    .A2(_1784_),
    .Y(_0319_),
    .B1(_1469_));
 sg13g2_o21ai_1 _4238_ (.B1(net435),
    .Y(_1470_),
    .A1(net374),
    .A2(_1409_));
 sg13g2_a21oi_1 _4239_ (.A1(net374),
    .A2(_1783_),
    .Y(_0320_),
    .B1(_1470_));
 sg13g2_nor2_1 _4240_ (.A(\display_value[4] ),
    .B(\display_value[2] ),
    .Y(_1471_));
 sg13g2_nand2_1 _4241_ (.Y(_1472_),
    .A(\display_value[1] ),
    .B(\display_value[0] ));
 sg13g2_nand2_1 _4242_ (.Y(_1473_),
    .A(_1471_),
    .B(_1472_));
 sg13g2_nand2_1 _4243_ (.Y(_1474_),
    .A(\display_value[1] ),
    .B(net760));
 sg13g2_nand2_1 _4244_ (.Y(_1475_),
    .A(net388),
    .B(_1474_));
 sg13g2_nor3_1 _4245_ (.A(net385),
    .B(_1473_),
    .C(_1475_),
    .Y(_1476_));
 sg13g2_nor2_2 _4246_ (.A(net417),
    .B(\dsp.digit ),
    .Y(_1477_));
 sg13g2_o21ai_1 _4247_ (.B1(_1477_),
    .Y(_1478_),
    .A1(display_graphical),
    .A2(net770));
 sg13g2_nor2_1 _4248_ (.A(net385),
    .B(_1806_),
    .Y(_1479_));
 sg13g2_nor2_1 _4249_ (.A(\display_value[1] ),
    .B(\display_value[0] ),
    .Y(_1480_));
 sg13g2_or2_1 _4250_ (.X(_1481_),
    .B(\display_value[0] ),
    .A(\display_value[1] ));
 sg13g2_nor2_1 _4251_ (.A(net387),
    .B(net760),
    .Y(_1482_));
 sg13g2_nand4_1 _4252_ (.B(_1479_),
    .C(_1480_),
    .A(_0230_),
    .Y(_1483_),
    .D(_1482_));
 sg13g2_and2_1 _4253_ (.A(net388),
    .B(_0230_),
    .X(_1484_));
 sg13g2_nand2_1 _4254_ (.Y(_1485_),
    .A(_1471_),
    .B(_1480_));
 sg13g2_o21ai_1 _4255_ (.B1(_1484_),
    .Y(_1486_),
    .A1(net386),
    .A2(_1485_));
 sg13g2_o21ai_1 _4256_ (.B1(_1486_),
    .Y(_1487_),
    .A1(_1476_),
    .A2(_1478_));
 sg13g2_nand2b_1 _4257_ (.Y(_0321_),
    .B(_1483_),
    .A_N(_1487_));
 sg13g2_o21ai_1 _4258_ (.B1(_1473_),
    .Y(_1488_),
    .A1(\display_value[4] ),
    .A2(net386));
 sg13g2_nor2_1 _4259_ (.A(\display_value[0] ),
    .B(_1474_),
    .Y(_1489_));
 sg13g2_nand3_1 _4260_ (.B(_1806_),
    .C(_1489_),
    .A(net385),
    .Y(_1490_));
 sg13g2_nand2_1 _4261_ (.Y(_1491_),
    .A(_1488_),
    .B(_1490_));
 sg13g2_a21oi_1 _4262_ (.A1(\display_value[2] ),
    .A2(_1481_),
    .Y(_1492_),
    .B1(net385));
 sg13g2_o21ai_1 _4263_ (.B1(_1491_),
    .Y(_1493_),
    .A1(net760),
    .A2(_1492_));
 sg13g2_nand3b_1 _4264_ (.B(_1479_),
    .C(_1480_),
    .Y(_1494_),
    .A_N(net760));
 sg13g2_o21ai_1 _4265_ (.B1(net387),
    .Y(_1495_),
    .A1(net385),
    .A2(\display_value[2] ));
 sg13g2_and3_1 _4266_ (.X(_1496_),
    .A(\dsp.digit ),
    .B(_1494_),
    .C(_1495_));
 sg13g2_o21ai_1 _4267_ (.B1(net387),
    .Y(_1497_),
    .A1(\display_value[4] ),
    .A2(net385));
 sg13g2_nand2_1 _4268_ (.Y(_1498_),
    .A(\display_value[2] ),
    .B(net387));
 sg13g2_o21ai_1 _4269_ (.B1(_1497_),
    .Y(_1499_),
    .A1(_1472_),
    .A2(_1498_));
 sg13g2_nand3_1 _4270_ (.B(_1479_),
    .C(_1489_),
    .A(net387),
    .Y(_1500_));
 sg13g2_nor2b_1 _4271_ (.A(net387),
    .B_N(_0015_),
    .Y(_1501_));
 sg13g2_nor3_1 _4272_ (.A(\dsp.digit ),
    .B(_1499_),
    .C(_1501_),
    .Y(_1502_));
 sg13g2_a221oi_1 _4273_ (.B2(_1502_),
    .C1(net417),
    .B1(_1500_),
    .A1(_1493_),
    .Y(_0322_),
    .A2(_1496_));
 sg13g2_nand2b_1 _4274_ (.Y(_1503_),
    .B(net749),
    .A_N(net387));
 sg13g2_o21ai_1 _4275_ (.B1(_1503_),
    .Y(_1504_),
    .A1(_1471_),
    .A2(_1497_));
 sg13g2_o21ai_1 _4276_ (.B1(_1482_),
    .Y(_1505_),
    .A1(net385),
    .A2(net748));
 sg13g2_a21oi_1 _4277_ (.A1(_1488_),
    .A2(_1490_),
    .Y(_1506_),
    .B1(_1197_));
 sg13g2_a22oi_1 _4278_ (.Y(_1507_),
    .B1(_1505_),
    .B2(_1506_),
    .A2(_1504_),
    .A1(_1477_));
 sg13g2_inv_1 _4279_ (.Y(_0323_),
    .A(net750));
 sg13g2_nor2b_1 _4280_ (.A(\display_value[4] ),
    .B_N(net387),
    .Y(_1508_));
 sg13g2_nand3_1 _4281_ (.B(_1472_),
    .C(_1474_),
    .A(_1891_),
    .Y(_1509_));
 sg13g2_nand4_1 _4282_ (.B(net748),
    .C(_1481_),
    .A(net385),
    .Y(_1510_),
    .D(_1509_));
 sg13g2_a21oi_1 _4283_ (.A1(_1891_),
    .A2(net762),
    .Y(_1511_),
    .B1(net388));
 sg13g2_o21ai_1 _4284_ (.B1(_1511_),
    .Y(_1512_),
    .A1(_1891_),
    .A2(_1494_));
 sg13g2_nand2_1 _4285_ (.Y(_1513_),
    .A(net431),
    .B(_1512_));
 sg13g2_a21oi_1 _4286_ (.A1(_1508_),
    .A2(_1510_),
    .Y(_0324_),
    .B1(_1513_));
 sg13g2_o21ai_1 _4287_ (.B1(_1477_),
    .Y(_1514_),
    .A1(net388),
    .A2(net780));
 sg13g2_a21o_1 _4288_ (.A2(_1488_),
    .A1(net388),
    .B1(_1514_),
    .X(_1515_));
 sg13g2_nor2_1 _4289_ (.A(_1197_),
    .B(_1497_),
    .Y(_1516_));
 sg13g2_nand2_1 _4290_ (.Y(_1517_),
    .A(_1485_),
    .B(_1516_));
 sg13g2_nand3_1 _4291_ (.B(_1515_),
    .C(_1517_),
    .A(_1483_),
    .Y(_0325_));
 sg13g2_nand2_1 _4292_ (.Y(_1518_),
    .A(_1492_),
    .B(_1508_));
 sg13g2_nand2_1 _4293_ (.Y(_1519_),
    .A(_1477_),
    .B(_1518_));
 sg13g2_o21ai_1 _4294_ (.B1(_1484_),
    .Y(_1520_),
    .A1(net386),
    .A2(_1473_));
 sg13g2_nor2_1 _4295_ (.A(net388),
    .B(net455),
    .Y(_1521_));
 sg13g2_a21oi_1 _4296_ (.A1(_1519_),
    .A2(_1520_),
    .Y(_0326_),
    .B1(_1521_));
 sg13g2_nand2_1 _4297_ (.Y(_1522_),
    .A(_0230_),
    .B(_1499_));
 sg13g2_o21ai_1 _4298_ (.B1(_1497_),
    .Y(_1523_),
    .A1(net388),
    .A2(_1892_));
 sg13g2_nand2_1 _4299_ (.Y(_1524_),
    .A(_1477_),
    .B(_1523_));
 sg13g2_nand3_1 _4300_ (.B(_1522_),
    .C(net769),
    .A(_1483_),
    .Y(_0327_));
 sg13g2_nor3_1 _4301_ (.A(_1795_),
    .B(net415),
    .C(_1413_),
    .Y(_0328_));
 sg13g2_nor3_1 _4302_ (.A(_1794_),
    .B(net415),
    .C(_1413_),
    .Y(_0329_));
 sg13g2_nor3_1 _4303_ (.A(_1793_),
    .B(net415),
    .C(_1413_),
    .Y(_0330_));
 sg13g2_nor3_1 _4304_ (.A(_1792_),
    .B(net415),
    .C(_1413_),
    .Y(_0331_));
 sg13g2_nor3_1 _4305_ (.A(_1796_),
    .B(net415),
    .C(_1413_),
    .Y(_0332_));
 sg13g2_and2_1 _4306_ (.A(_0999_),
    .B(_1001_),
    .X(_1525_));
 sg13g2_o21ai_1 _4307_ (.B1(net366),
    .Y(_1526_),
    .A1(net563),
    .A2(_1525_));
 sg13g2_a21oi_1 _4308_ (.A1(net563),
    .A2(_1525_),
    .Y(_0333_),
    .B1(_1526_));
 sg13g2_a21oi_1 _4309_ (.A1(_0999_),
    .A2(_1001_),
    .Y(_1527_),
    .B1(net356));
 sg13g2_mux2_1 _4310_ (.A0(_1012_),
    .A1(net629),
    .S(_1527_),
    .X(_0334_));
 sg13g2_mux2_1 _4311_ (.A0(_1020_),
    .A1(net548),
    .S(_1527_),
    .X(_0335_));
 sg13g2_nor2b_2 _4312_ (.A(_0845_),
    .B_N(_0844_),
    .Y(_1528_));
 sg13g2_o21ai_1 _4313_ (.B1(net362),
    .Y(_1529_),
    .A1(net759),
    .A2(_1528_));
 sg13g2_a21oi_1 _4314_ (.A1(net759),
    .A2(_1528_),
    .Y(_0336_),
    .B1(_1529_));
 sg13g2_nor2_1 _4315_ (.A(net355),
    .B(_1528_),
    .Y(_1530_));
 sg13g2_a22oi_1 _4316_ (.Y(_1531_),
    .B1(_1530_),
    .B2(net728),
    .A2(_1528_),
    .A1(_0857_));
 sg13g2_inv_1 _4317_ (.Y(_0337_),
    .A(_1531_));
 sg13g2_nor2_1 _4318_ (.A(_0864_),
    .B(_1530_),
    .Y(_1532_));
 sg13g2_a21oi_1 _4319_ (.A1(_1869_),
    .A2(_1530_),
    .Y(_0338_),
    .B1(_1532_));
 sg13g2_nor2b_1 _4320_ (.A(_0844_),
    .B_N(_0845_),
    .Y(_1533_));
 sg13g2_o21ai_1 _4321_ (.B1(net362),
    .Y(_1534_),
    .A1(net764),
    .A2(_1533_));
 sg13g2_a21oi_1 _4322_ (.A1(net764),
    .A2(_1533_),
    .Y(_0339_),
    .B1(_1534_));
 sg13g2_nor2_1 _4323_ (.A(net355),
    .B(_1533_),
    .Y(_1535_));
 sg13g2_a22oi_1 _4324_ (.Y(_1536_),
    .B1(_1535_),
    .B2(net741),
    .A2(_1533_),
    .A1(_0857_));
 sg13g2_inv_1 _4325_ (.Y(_0340_),
    .A(_1536_));
 sg13g2_nor2_1 _4326_ (.A(_0864_),
    .B(_1535_),
    .Y(_1537_));
 sg13g2_a21oi_1 _4327_ (.A1(_1861_),
    .A2(_1535_),
    .Y(_0341_),
    .B1(_1537_));
 sg13g2_or2_2 _4328_ (.X(_1538_),
    .B(_0838_),
    .A(_0820_));
 sg13g2_nor2_1 _4329_ (.A(_0823_),
    .B(_1538_),
    .Y(_1539_));
 sg13g2_a21oi_1 _4330_ (.A1(_1848_),
    .A2(_1538_),
    .Y(_0342_),
    .B1(_1539_));
 sg13g2_nand2_1 _4331_ (.Y(_1540_),
    .A(net472),
    .B(_1538_));
 sg13g2_o21ai_1 _4332_ (.B1(_1540_),
    .Y(_0343_),
    .A1(_0827_),
    .A2(_1538_));
 sg13g2_nand2_1 _4333_ (.Y(_1541_),
    .A(net475),
    .B(_1538_));
 sg13g2_o21ai_1 _4334_ (.B1(_1541_),
    .Y(_0344_),
    .A1(_0835_),
    .A2(_1538_));
 sg13g2_nand2_1 _4335_ (.Y(_1542_),
    .A(_1832_),
    .B(\snd.counter[6] ));
 sg13g2_nor2_1 _4336_ (.A(_1833_),
    .B(\snd.counter[5] ),
    .Y(_1543_));
 sg13g2_nor2_1 _4337_ (.A(_1838_),
    .B(\snd.counter[0] ),
    .Y(_1544_));
 sg13g2_o21ai_1 _4338_ (.B1(_1544_),
    .Y(_1545_),
    .A1(\snd.note_timing[2] ),
    .A2(_1889_));
 sg13g2_a22oi_1 _4339_ (.Y(_1546_),
    .B1(_1889_),
    .B2(\snd.note_timing[2] ),
    .A2(_1888_),
    .A1(\snd.note_timing[3] ));
 sg13g2_nand2_1 _4340_ (.Y(_1547_),
    .A(_1835_),
    .B(\snd.counter[3] ));
 sg13g2_a22oi_1 _4341_ (.Y(_1548_),
    .B1(_1545_),
    .B2(_1546_),
    .A2(\snd.counter[2] ),
    .A1(_1836_));
 sg13g2_nor2_1 _4342_ (.A(_1835_),
    .B(\snd.counter[3] ),
    .Y(_1549_));
 sg13g2_a221oi_1 _4343_ (.B2(_1548_),
    .C1(_1549_),
    .B1(_1547_),
    .A1(\snd.note_timing[5] ),
    .Y(_1550_),
    .A2(_1887_));
 sg13g2_a221oi_1 _4344_ (.B2(_1834_),
    .C1(_1550_),
    .B1(\snd.counter[4] ),
    .A1(_1833_),
    .Y(_1551_),
    .A2(\snd.counter[5] ));
 sg13g2_o21ai_1 _4345_ (.B1(_1542_),
    .Y(_1552_),
    .A1(_1543_),
    .A2(_1551_));
 sg13g2_a22oi_1 _4346_ (.Y(_1553_),
    .B1(_1885_),
    .B2(\snd.note_timing[7] ),
    .A2(_1884_),
    .A1(\snd.note_timing[8] ));
 sg13g2_nor2_1 _4347_ (.A(net568),
    .B(\snd.counter[8] ),
    .Y(_1554_));
 sg13g2_a22oi_1 _4348_ (.Y(_1555_),
    .B1(_1552_),
    .B2(_1553_),
    .A2(\snd.counter[7] ),
    .A1(_1831_));
 sg13g2_a21oi_1 _4349_ (.A1(net569),
    .A2(_1555_),
    .Y(_0345_),
    .B1(net334));
 sg13g2_nand2_1 _4350_ (.Y(_1556_),
    .A(_1840_),
    .B(\snd.note_sel[0] ));
 sg13g2_nor2_2 _4351_ (.A(\snd.chord[1][5] ),
    .B(\snd.chord[1][0] ),
    .Y(_1557_));
 sg13g2_nor2_1 _4352_ (.A(\snd.note_sel[1] ),
    .B(\snd.note_sel[0] ),
    .Y(_1558_));
 sg13g2_or4_1 _4353_ (.A(\snd.chord[0][3] ),
    .B(\snd.chord[0][2] ),
    .C(\snd.chord[0][1] ),
    .D(\snd.chord[0][0] ),
    .X(_1559_));
 sg13g2_nor3_2 _4354_ (.A(\snd.chord[0][5] ),
    .B(\snd.chord[0][4] ),
    .C(_1559_),
    .Y(_1560_));
 sg13g2_nand3_1 _4355_ (.B(\snd.note_sel[0] ),
    .C(_1560_),
    .A(\snd.note_sel[1] ),
    .Y(_1561_));
 sg13g2_nand2b_1 _4356_ (.Y(_1562_),
    .B(_1561_),
    .A_N(_1558_));
 sg13g2_nand2_1 _4357_ (.Y(_1563_),
    .A(_1557_),
    .B(_1562_));
 sg13g2_a22oi_1 _4358_ (.Y(_1564_),
    .B1(_1556_),
    .B2(_1563_),
    .A2(_1828_),
    .A1(_1780_));
 sg13g2_nand2_1 _4359_ (.Y(_1565_),
    .A(\snd.note_sel[1] ),
    .B(_1841_));
 sg13g2_nand3_1 _4360_ (.B(_1557_),
    .C(_1560_),
    .A(\snd.chord[2][2] ),
    .Y(_1566_));
 sg13g2_a21oi_1 _4361_ (.A1(net567),
    .A2(_1566_),
    .Y(_1567_),
    .B1(_1565_));
 sg13g2_nor2_2 _4362_ (.A(_1564_),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_inv_1 _4363_ (.Y(_1569_),
    .A(_1568_));
 sg13g2_o21ai_1 _4364_ (.B1(_1557_),
    .Y(_1570_),
    .A1(\snd.chord[2][2] ),
    .A2(_1828_));
 sg13g2_o21ai_1 _4365_ (.B1(_1565_),
    .Y(_1571_),
    .A1(\snd.chord[2][2] ),
    .A2(_1556_));
 sg13g2_nand2b_1 _4366_ (.Y(_1572_),
    .B(_1560_),
    .A_N(_1557_));
 sg13g2_o21ai_1 _4367_ (.B1(_1572_),
    .Y(_1573_),
    .A1(_0061_),
    .A2(_1558_));
 sg13g2_and2_1 _4368_ (.A(_1571_),
    .B(_1573_),
    .X(_1574_));
 sg13g2_a21o_2 _4369_ (.A2(_1570_),
    .A1(_1562_),
    .B1(_1574_),
    .X(_1575_));
 sg13g2_nor2_2 _4370_ (.A(_1569_),
    .B(_1575_),
    .Y(_1576_));
 sg13g2_nand2_2 _4371_ (.Y(_1577_),
    .A(\snd.chord[0][4] ),
    .B(_1576_));
 sg13g2_nand3_1 _4372_ (.B(_1569_),
    .C(_1575_),
    .A(\snd.chord[3][0] ),
    .Y(_1578_));
 sg13g2_inv_1 _4373_ (.Y(_1579_),
    .A(_1578_));
 sg13g2_mux4_1 _4374_ (.S0(_1568_),
    .A0(_1780_),
    .A1(_1778_),
    .A2(_1828_),
    .A3(_1779_),
    .S1(_1575_),
    .X(_1580_));
 sg13g2_a21oi_2 _4375_ (.B1(net379),
    .Y(_1581_),
    .A2(_1580_),
    .A1(_1577_));
 sg13g2_a21o_1 _4376_ (.A2(_1568_),
    .A1(\snd.chord[1][0] ),
    .B1(_1576_),
    .X(_1582_));
 sg13g2_mux4_1 _4377_ (.S0(_1568_),
    .A0(\snd.chord[2][2] ),
    .A1(\snd.chord[0][2] ),
    .A2(\snd.chord[3][0] ),
    .A3(\snd.chord[1][0] ),
    .S1(_1575_),
    .X(_1583_));
 sg13g2_nand2_2 _4378_ (.Y(_1584_),
    .A(\snd.chord[0][3] ),
    .B(_1576_));
 sg13g2_a21oi_2 _4379_ (.B1(_1579_),
    .Y(_1585_),
    .A2(_1576_),
    .A1(\snd.chord[0][1] ));
 sg13g2_nand2_1 _4380_ (.Y(_1586_),
    .A(_0059_),
    .B(_1576_));
 sg13g2_o21ai_1 _4381_ (.B1(_1586_),
    .Y(_1587_),
    .A1(_1579_),
    .A2(_1582_));
 sg13g2_nand2_2 _4382_ (.Y(_1588_),
    .A(_1585_),
    .B(_1587_));
 sg13g2_xnor2_1 _4383_ (.Y(_1589_),
    .A(_1584_),
    .B(_1588_));
 sg13g2_inv_1 _4384_ (.Y(_1590_),
    .A(_1589_));
 sg13g2_a21oi_2 _4385_ (.B1(_1580_),
    .Y(_1591_),
    .A2(_1576_),
    .A1(\snd.chord[0][4] ));
 sg13g2_o21ai_1 _4386_ (.B1(_1591_),
    .Y(_1592_),
    .A1(_1583_),
    .A2(_1590_));
 sg13g2_nor2_2 _4387_ (.A(_1778_),
    .B(_1577_),
    .Y(_1593_));
 sg13g2_nor2_1 _4388_ (.A(_1583_),
    .B(_1584_),
    .Y(_1594_));
 sg13g2_or2_1 _4389_ (.X(_1595_),
    .B(_1584_),
    .A(_1583_));
 sg13g2_nor2_1 _4390_ (.A(_1583_),
    .B(_1587_),
    .Y(_1596_));
 sg13g2_a21oi_2 _4391_ (.B1(_1596_),
    .Y(_1597_),
    .A2(_1594_),
    .A1(_1585_));
 sg13g2_nand2_1 _4392_ (.Y(_1598_),
    .A(_1593_),
    .B(_1597_));
 sg13g2_nand2_1 _4393_ (.Y(_1599_),
    .A(_1583_),
    .B(_1584_));
 sg13g2_o21ai_1 _4394_ (.B1(_1584_),
    .Y(_1600_),
    .A1(_1583_),
    .A2(_1588_));
 sg13g2_nand2_1 _4395_ (.Y(_1601_),
    .A(_1595_),
    .B(_1600_));
 sg13g2_nor2_1 _4396_ (.A(_1585_),
    .B(_1587_),
    .Y(_1602_));
 sg13g2_inv_1 _4397_ (.Y(_1603_),
    .A(_1602_));
 sg13g2_or2_1 _4398_ (.X(_1604_),
    .B(_1602_),
    .A(_1599_));
 sg13g2_inv_1 _4399_ (.Y(_1605_),
    .A(_1604_));
 sg13g2_nand2_1 _4400_ (.Y(_1606_),
    .A(_1588_),
    .B(_1605_));
 sg13g2_nand2_1 _4401_ (.Y(_1607_),
    .A(_1594_),
    .B(_1602_));
 sg13g2_nor2_2 _4402_ (.A(\snd.chord[0][5] ),
    .B(_1577_),
    .Y(_1608_));
 sg13g2_nand4_1 _4403_ (.B(_1606_),
    .C(_1607_),
    .A(_1601_),
    .Y(_1609_),
    .D(_1608_));
 sg13g2_nand3_1 _4404_ (.B(_1598_),
    .C(_1609_),
    .A(_1592_),
    .Y(_1610_));
 sg13g2_a22oi_1 _4405_ (.Y(_1611_),
    .B1(_1581_),
    .B2(_1610_),
    .A2(net508),
    .A1(net379));
 sg13g2_nor2_1 _4406_ (.A(net419),
    .B(_1611_),
    .Y(_0346_));
 sg13g2_o21ai_1 _4407_ (.B1(_1608_),
    .Y(_1612_),
    .A1(_1583_),
    .A2(_1590_));
 sg13g2_nor2_1 _4408_ (.A(_1583_),
    .B(_1585_),
    .Y(_1613_));
 sg13g2_o21ai_1 _4409_ (.B1(_1607_),
    .Y(_1614_),
    .A1(_1594_),
    .A2(_1613_));
 sg13g2_a22oi_1 _4410_ (.Y(_1615_),
    .B1(_1614_),
    .B2(_1593_),
    .A2(_1597_),
    .A1(_1591_));
 sg13g2_nand2_1 _4411_ (.Y(_1616_),
    .A(_1612_),
    .B(_1615_));
 sg13g2_a22oi_1 _4412_ (.Y(_1617_),
    .B1(_1581_),
    .B2(_1616_),
    .A2(net504),
    .A1(net379));
 sg13g2_nor2_1 _4413_ (.A(net419),
    .B(_1617_),
    .Y(_0347_));
 sg13g2_nand2b_1 _4414_ (.Y(_1618_),
    .B(_1587_),
    .A_N(_1599_));
 sg13g2_nand2b_1 _4415_ (.Y(_1619_),
    .B(_1618_),
    .A_N(_1596_));
 sg13g2_inv_1 _4416_ (.Y(_1620_),
    .A(_1619_));
 sg13g2_a22oi_1 _4417_ (.Y(_1621_),
    .B1(_1620_),
    .B2(_1593_),
    .A2(_1614_),
    .A1(_1591_));
 sg13g2_nand2b_1 _4418_ (.Y(_1622_),
    .B(_1581_),
    .A_N(_1621_));
 sg13g2_nor3_2 _4419_ (.A(\snd.chord[0][5] ),
    .B(net377),
    .C(_1577_),
    .Y(_1623_));
 sg13g2_nand2_1 _4420_ (.Y(_1624_),
    .A(net407),
    .B(_1608_));
 sg13g2_a22oi_1 _4421_ (.Y(_1625_),
    .B1(_1597_),
    .B2(_1623_),
    .A2(net554),
    .A1(net377));
 sg13g2_a21oi_1 _4422_ (.A1(_1622_),
    .A2(_1625_),
    .Y(_0348_),
    .B1(net419));
 sg13g2_a21oi_2 _4423_ (.B1(_1613_),
    .Y(_1626_),
    .A2(_1605_),
    .A1(_1588_));
 sg13g2_nand2_1 _4424_ (.Y(_1627_),
    .A(_1593_),
    .B(_1626_));
 sg13g2_a22oi_1 _4425_ (.Y(_1628_),
    .B1(_1620_),
    .B2(_1591_),
    .A2(_1614_),
    .A1(_1608_));
 sg13g2_nand2_1 _4426_ (.Y(_1629_),
    .A(_1627_),
    .B(_1628_));
 sg13g2_a22oi_1 _4427_ (.Y(_1630_),
    .B1(_1581_),
    .B2(_1629_),
    .A2(net509),
    .A1(net379));
 sg13g2_nor2_1 _4428_ (.A(net419),
    .B(_1630_),
    .Y(_0349_));
 sg13g2_nor3_1 _4429_ (.A(\snd.chord[0][5] ),
    .B(_1577_),
    .C(_1619_),
    .Y(_1631_));
 sg13g2_a221oi_1 _4430_ (.B2(_1591_),
    .C1(_1631_),
    .B1(_1626_),
    .A1(_1593_),
    .Y(_1632_),
    .A2(_1604_));
 sg13g2_inv_1 _4431_ (.Y(_1633_),
    .A(_1632_));
 sg13g2_a22oi_1 _4432_ (.Y(_1634_),
    .B1(_1581_),
    .B2(_1633_),
    .A2(net492),
    .A1(net377));
 sg13g2_nor2_1 _4433_ (.A(net420),
    .B(_1634_),
    .Y(_0350_));
 sg13g2_nand2_1 _4434_ (.Y(_1635_),
    .A(_1608_),
    .B(_1626_));
 sg13g2_o21ai_1 _4435_ (.B1(_1595_),
    .Y(_1636_),
    .A1(_1599_),
    .A2(_1603_));
 sg13g2_a22oi_1 _4436_ (.Y(_1637_),
    .B1(_1636_),
    .B2(_1593_),
    .A2(_1604_),
    .A1(_1591_));
 sg13g2_nand2_1 _4437_ (.Y(_1638_),
    .A(_1635_),
    .B(_1637_));
 sg13g2_a22oi_1 _4438_ (.Y(_1639_),
    .B1(_1581_),
    .B2(_1638_),
    .A2(net488),
    .A1(net377));
 sg13g2_nor2_1 _4439_ (.A(net420),
    .B(_1639_),
    .Y(_0351_));
 sg13g2_mux2_1 _4440_ (.A0(_1593_),
    .A1(_1591_),
    .S(_1636_),
    .X(_1640_));
 sg13g2_nand2_1 _4441_ (.Y(_1641_),
    .A(_1581_),
    .B(_1640_));
 sg13g2_a22oi_1 _4442_ (.Y(_1642_),
    .B1(_1604_),
    .B2(_1623_),
    .A2(net649),
    .A1(net377));
 sg13g2_a21oi_1 _4443_ (.A1(_1641_),
    .A2(_1642_),
    .Y(_0352_),
    .B1(net420));
 sg13g2_mux2_1 _4444_ (.A0(_1577_),
    .A1(_1608_),
    .S(_1636_),
    .X(_1643_));
 sg13g2_a22oi_1 _4445_ (.Y(_1644_),
    .B1(_1581_),
    .B2(_1643_),
    .A2(net538),
    .A1(net377));
 sg13g2_nor2_1 _4446_ (.A(net420),
    .B(_1644_),
    .Y(_0353_));
 sg13g2_nor2_1 _4447_ (.A(_1624_),
    .B(_1636_),
    .Y(_1645_));
 sg13g2_a21oi_1 _4448_ (.A1(net378),
    .A2(net519),
    .Y(_1646_),
    .B1(_1645_));
 sg13g2_nor2_1 _4449_ (.A(net420),
    .B(_1646_),
    .Y(_0354_));
 sg13g2_o21ai_1 _4450_ (.B1(net437),
    .Y(_1647_),
    .A1(net377),
    .A2(_1575_));
 sg13g2_a21oi_1 _4451_ (.A1(net377),
    .A2(_1782_),
    .Y(_0355_),
    .B1(_1647_));
 sg13g2_o21ai_1 _4452_ (.B1(net437),
    .Y(_1648_),
    .A1(net564),
    .A2(net407));
 sg13g2_a21oi_1 _4453_ (.A1(net407),
    .A2(_1568_),
    .Y(_0356_),
    .B1(_1648_));
 sg13g2_o21ai_1 _4454_ (.B1(net693),
    .Y(_1649_),
    .A1(_0890_),
    .A2(_0892_));
 sg13g2_a22oi_1 _4455_ (.Y(_1650_),
    .B1(_0902_),
    .B2(net557),
    .A2(_0898_),
    .A1(uo_out[2]));
 sg13g2_a21oi_1 _4456_ (.A1(_1649_),
    .A2(_1650_),
    .Y(_0357_),
    .B1(net419));
 sg13g2_nand2_1 _4457_ (.Y(_1651_),
    .A(\snd.active_tune[1] ),
    .B(\snd.active_tune[0] ));
 sg13g2_nor3_1 _4458_ (.A(\snd.tune_counter[6] ),
    .B(\snd.tune_counter[5] ),
    .C(\snd.tune_counter[4] ),
    .Y(_1652_));
 sg13g2_nor2_1 _4459_ (.A(\snd.tune_counter[3] ),
    .B(\snd.tune_counter[2] ),
    .Y(_1653_));
 sg13g2_nand3_1 _4460_ (.B(_1652_),
    .C(_1653_),
    .A(_0885_),
    .Y(_1654_));
 sg13g2_nor3_2 _4461_ (.A(_0080_),
    .B(_0888_),
    .C(_1654_),
    .Y(_1655_));
 sg13g2_nor2_1 _4462_ (.A(\snd.tune_pos[1] ),
    .B(\snd.tune_pos[0] ),
    .Y(_1656_));
 sg13g2_nand2b_1 _4463_ (.Y(_1657_),
    .B(_1656_),
    .A_N(\snd.tune_pos[2] ));
 sg13g2_nor2b_1 _4464_ (.A(_1651_),
    .B_N(_1657_),
    .Y(_1658_));
 sg13g2_nor3_1 _4465_ (.A(_0892_),
    .B(_1654_),
    .C(_1658_),
    .Y(_1659_));
 sg13g2_nor2_1 _4466_ (.A(_0893_),
    .B(_1659_),
    .Y(_1660_));
 sg13g2_a21oi_2 _4467_ (.B1(_1660_),
    .Y(_1661_),
    .A2(_1655_),
    .A1(_1651_));
 sg13g2_or2_1 _4468_ (.X(_1662_),
    .B(_1661_),
    .A(net785));
 sg13g2_nand2_1 _4469_ (.Y(_1663_),
    .A(_0889_),
    .B(_1661_));
 sg13g2_and3_1 _4470_ (.X(_0358_),
    .A(net433),
    .B(_1662_),
    .C(_1663_));
 sg13g2_a221oi_1 _4471_ (.B2(net477),
    .C1(_1663_),
    .B1(_0902_),
    .A1(uo_out[1]),
    .Y(_1664_),
    .A2(_0898_));
 sg13g2_o21ai_1 _4472_ (.B1(net433),
    .Y(_1665_),
    .A1(net724),
    .A2(_1661_));
 sg13g2_nor2_1 _4473_ (.A(_1664_),
    .B(_1665_),
    .Y(_0359_));
 sg13g2_nor4_1 _4474_ (.A(\game.state[3] ),
    .B(_1170_),
    .C(_1206_),
    .D(_1329_),
    .Y(_1666_));
 sg13g2_nor2b_2 _4475_ (.A(_1370_),
    .B_N(_1666_),
    .Y(_1667_));
 sg13g2_o21ai_1 _4476_ (.B1(net429),
    .Y(_1668_),
    .A1(net589),
    .A2(_1667_));
 sg13g2_a21oi_1 _4477_ (.A1(_1115_),
    .A2(_1667_),
    .Y(_0360_),
    .B1(_1668_));
 sg13g2_o21ai_1 _4478_ (.B1(net429),
    .Y(_1669_),
    .A1(net553),
    .A2(_1667_));
 sg13g2_a21oi_1 _4479_ (.A1(net369),
    .A2(_1667_),
    .Y(_0361_),
    .B1(_1669_));
 sg13g2_nand2b_1 _4480_ (.Y(_1670_),
    .B(\snd.tune_pos[0] ),
    .A_N(\snd.tune_pos[2] ));
 sg13g2_nor2b_1 _4481_ (.A(\snd.tune_pos[0] ),
    .B_N(\snd.tune_pos[1] ),
    .Y(_1671_));
 sg13g2_nor2_1 _4482_ (.A(\snd.tune_pos[1] ),
    .B(_0082_),
    .Y(_1672_));
 sg13g2_a21oi_1 _4483_ (.A1(_0082_),
    .A2(_1671_),
    .Y(_1673_),
    .B1(_1672_));
 sg13g2_nand2_1 _4484_ (.Y(_1674_),
    .A(_1670_),
    .B(_1673_));
 sg13g2_nor2b_1 _4485_ (.A(\snd.tune_pos[1] ),
    .B_N(\snd.tune_pos[0] ),
    .Y(_1675_));
 sg13g2_nand2_1 _4486_ (.Y(_1676_),
    .A(\snd.tune_pos[2] ),
    .B(_1675_));
 sg13g2_nand4_1 _4487_ (.B(_1670_),
    .C(_1673_),
    .A(_1657_),
    .Y(_1677_),
    .D(_1676_));
 sg13g2_nand2b_1 _4488_ (.Y(_1678_),
    .B(_1675_),
    .A_N(\snd.tune_pos[2] ));
 sg13g2_nor3_1 _4489_ (.A(\snd.active_tune[1] ),
    .B(\snd.tune_pos[2] ),
    .C(\snd.tune_pos[1] ),
    .Y(_1679_));
 sg13g2_o21ai_1 _4490_ (.B1(\snd.active_tune[1] ),
    .Y(_1680_),
    .A1(net380),
    .A2(_1677_));
 sg13g2_nand3b_1 _4491_ (.B(_1680_),
    .C(_1655_),
    .Y(_1681_),
    .A_N(_1679_));
 sg13g2_nor2_1 _4492_ (.A(_1777_),
    .B(net380),
    .Y(_1682_));
 sg13g2_nand2b_2 _4493_ (.Y(_1683_),
    .B(_1681_),
    .A_N(_1660_));
 sg13g2_inv_1 _4494_ (.Y(_1684_),
    .A(_1683_));
 sg13g2_nor3_1 _4495_ (.A(\snd.active_tune[1] ),
    .B(net380),
    .C(_1678_),
    .Y(_1685_));
 sg13g2_inv_1 _4496_ (.Y(_1686_),
    .A(_1685_));
 sg13g2_nor3_1 _4497_ (.A(_0889_),
    .B(_1683_),
    .C(_1685_),
    .Y(_1687_));
 sg13g2_a21oi_1 _4498_ (.A1(net380),
    .A2(_1678_),
    .Y(_1688_),
    .B1(net758));
 sg13g2_nor4_1 _4499_ (.A(_1777_),
    .B(net380),
    .C(\snd.tune_pos[0] ),
    .D(_1673_),
    .Y(_1689_));
 sg13g2_o21ai_1 _4500_ (.B1(_1687_),
    .Y(_1690_),
    .A1(_1688_),
    .A2(_1689_));
 sg13g2_and2_1 _4501_ (.A(\btn.button_state[0] ),
    .B(_0902_),
    .X(_1691_));
 sg13g2_a21o_1 _4502_ (.A2(_0898_),
    .A1(uo_out[0]),
    .B1(_1691_),
    .X(_1692_));
 sg13g2_a21oi_1 _4503_ (.A1(net635),
    .A2(_1683_),
    .Y(_1693_),
    .B1(_1692_));
 sg13g2_a21oi_1 _4504_ (.A1(_1690_),
    .A2(_1693_),
    .Y(_0362_),
    .B1(net419));
 sg13g2_or2_1 _4505_ (.X(_1694_),
    .B(_1675_),
    .A(_1671_));
 sg13g2_nor2_1 _4506_ (.A(net380),
    .B(_1694_),
    .Y(_1695_));
 sg13g2_a21oi_1 _4507_ (.A1(_1674_),
    .A2(_1695_),
    .Y(_1696_),
    .B1(_1777_));
 sg13g2_nor2_1 _4508_ (.A(_0889_),
    .B(_1696_),
    .Y(_1697_));
 sg13g2_nor3_1 _4509_ (.A(_1683_),
    .B(_1692_),
    .C(_1697_),
    .Y(_1698_));
 sg13g2_o21ai_1 _4510_ (.B1(net434),
    .Y(_1699_),
    .A1(net669),
    .A2(_1684_));
 sg13g2_nor2_1 _4511_ (.A(_1698_),
    .B(_1699_),
    .Y(_0363_));
 sg13g2_nand2_1 _4512_ (.Y(_1700_),
    .A(\snd.tune_pos[2] ),
    .B(_1656_));
 sg13g2_a21oi_1 _4513_ (.A1(_1678_),
    .A2(_1700_),
    .Y(_1701_),
    .B1(net380));
 sg13g2_o21ai_1 _4514_ (.B1(_1687_),
    .Y(_1702_),
    .A1(_1688_),
    .A2(_1701_));
 sg13g2_a21oi_1 _4515_ (.A1(net707),
    .A2(_1683_),
    .Y(_1703_),
    .B1(_1692_));
 sg13g2_a21oi_1 _4516_ (.A1(_1702_),
    .A2(_1703_),
    .Y(_0364_),
    .B1(net419));
 sg13g2_nand3_1 _4517_ (.B(_1671_),
    .C(_1682_),
    .A(_0082_),
    .Y(_1704_));
 sg13g2_o21ai_1 _4518_ (.B1(_1684_),
    .Y(_1705_),
    .A1(_0889_),
    .A2(_1704_));
 sg13g2_o21ai_1 _4519_ (.B1(net434),
    .Y(_1706_),
    .A1(net675),
    .A2(_1684_));
 sg13g2_nor2b_1 _4520_ (.A(_1706_),
    .B_N(_1705_),
    .Y(_0365_));
 sg13g2_nand2b_1 _4521_ (.Y(_1707_),
    .B(_1682_),
    .A_N(_1676_));
 sg13g2_a21oi_1 _4522_ (.A1(_1686_),
    .A2(_1707_),
    .Y(_1708_),
    .B1(_0889_));
 sg13g2_nor3_1 _4523_ (.A(_1683_),
    .B(_1692_),
    .C(_1708_),
    .Y(_1709_));
 sg13g2_o21ai_1 _4524_ (.B1(net434),
    .Y(_1710_),
    .A1(net757),
    .A2(_1684_));
 sg13g2_nor2_1 _4525_ (.A(_1709_),
    .B(_1710_),
    .Y(_0366_));
 sg13g2_a21oi_1 _4526_ (.A1(net664),
    .A2(_1683_),
    .Y(_1711_),
    .B1(_1687_));
 sg13g2_nor2_1 _4527_ (.A(net420),
    .B(_1711_),
    .Y(_0367_));
 sg13g2_a21oi_2 _4528_ (.B1(_0898_),
    .Y(_1712_),
    .A2(_0900_),
    .A1(_0895_));
 sg13g2_o21ai_1 _4529_ (.B1(_1860_),
    .Y(_1713_),
    .A1(net408),
    .A2(_0888_));
 sg13g2_nand2_1 _4530_ (.Y(_1714_),
    .A(_0892_),
    .B(_1713_));
 sg13g2_nand2_2 _4531_ (.Y(_1715_),
    .A(_1712_),
    .B(_1714_));
 sg13g2_inv_1 _4532_ (.Y(_1716_),
    .A(_1715_));
 sg13g2_nand2_1 _4533_ (.Y(_1717_),
    .A(_0889_),
    .B(_0891_));
 sg13g2_nand2_1 _4534_ (.Y(_1718_),
    .A(\snd.tune_counter[5] ),
    .B(\snd.tune_counter[4] ));
 sg13g2_nand3_1 _4535_ (.B(_0081_),
    .C(_1653_),
    .A(\snd.tune_counter[1] ),
    .Y(_1719_));
 sg13g2_nor3_1 _4536_ (.A(\snd.tune_counter[0] ),
    .B(_1718_),
    .C(_1719_),
    .Y(_1720_));
 sg13g2_nor2b_1 _4537_ (.A(_0891_),
    .B_N(_1720_),
    .Y(_1721_));
 sg13g2_a21oi_1 _4538_ (.A1(_0889_),
    .A2(_0891_),
    .Y(_1722_),
    .B1(_1721_));
 sg13g2_a21oi_1 _4539_ (.A1(_1716_),
    .A2(_1722_),
    .Y(_1723_),
    .B1(net637));
 sg13g2_a21oi_1 _4540_ (.A1(net637),
    .A2(_1716_),
    .Y(_1724_),
    .B1(net413));
 sg13g2_nor2b_1 _4541_ (.A(_1723_),
    .B_N(_1724_),
    .Y(_0368_));
 sg13g2_a21oi_1 _4542_ (.A1(\snd.tune_counter[0] ),
    .A2(_1716_),
    .Y(_1725_),
    .B1(net573));
 sg13g2_a21oi_1 _4543_ (.A1(_0888_),
    .A2(_0891_),
    .Y(_1726_),
    .B1(_1721_));
 sg13g2_o21ai_1 _4544_ (.B1(net428),
    .Y(_1727_),
    .A1(_1715_),
    .A2(_1726_));
 sg13g2_nand2_1 _4545_ (.Y(_1728_),
    .A(net573),
    .B(\snd.tune_counter[0] ));
 sg13g2_nor2_1 _4546_ (.A(_1715_),
    .B(_1728_),
    .Y(_1729_));
 sg13g2_nor3_1 _4547_ (.A(net574),
    .B(_1727_),
    .C(_1729_),
    .Y(_0369_));
 sg13g2_nor2_1 _4548_ (.A(net625),
    .B(_1729_),
    .Y(_1730_));
 sg13g2_o21ai_1 _4549_ (.B1(net427),
    .Y(_1731_),
    .A1(_1715_),
    .A2(_1717_));
 sg13g2_and2_1 _4550_ (.A(net625),
    .B(_1729_),
    .X(_1732_));
 sg13g2_nor3_1 _4551_ (.A(net626),
    .B(_1731_),
    .C(_1732_),
    .Y(_0370_));
 sg13g2_nor2_1 _4552_ (.A(net660),
    .B(_1732_),
    .Y(_1733_));
 sg13g2_nand2_1 _4553_ (.Y(_1734_),
    .A(\snd.tune_counter[3] ),
    .B(\snd.tune_counter[2] ));
 sg13g2_nor3_2 _4554_ (.A(_1715_),
    .B(_1728_),
    .C(_1734_),
    .Y(_1735_));
 sg13g2_and3_2 _4555_ (.X(_1736_),
    .A(_0888_),
    .B(_0891_),
    .C(_1712_));
 sg13g2_nor4_1 _4556_ (.A(net413),
    .B(_1733_),
    .C(_1735_),
    .D(_1736_),
    .Y(_0371_));
 sg13g2_xnor2_1 _4557_ (.Y(_1737_),
    .A(net718),
    .B(_1735_));
 sg13g2_nor2_1 _4558_ (.A(_1727_),
    .B(net719),
    .Y(_0372_));
 sg13g2_a21oi_1 _4559_ (.A1(\snd.tune_counter[4] ),
    .A2(_1735_),
    .Y(_1738_),
    .B1(net517));
 sg13g2_or3_1 _4560_ (.A(_1718_),
    .B(_1728_),
    .C(_1734_),
    .X(_1739_));
 sg13g2_a21oi_1 _4561_ (.A1(_1722_),
    .A2(_1739_),
    .Y(_1740_),
    .B1(_1715_));
 sg13g2_nor3_1 _4562_ (.A(net413),
    .B(net518),
    .C(_1740_),
    .Y(_0373_));
 sg13g2_xor2_1 _4563_ (.B(_1739_),
    .A(_0081_),
    .X(_1741_));
 sg13g2_nor2_1 _4564_ (.A(_1715_),
    .B(_1741_),
    .Y(_1742_));
 sg13g2_nor2_1 _4565_ (.A(net549),
    .B(_1716_),
    .Y(_1743_));
 sg13g2_nor3_1 _4566_ (.A(_1731_),
    .B(_1742_),
    .C(_1743_),
    .Y(_0374_));
 sg13g2_nand2_1 _4567_ (.Y(_1744_),
    .A(_0893_),
    .B(_1712_));
 sg13g2_inv_1 _4568_ (.Y(_1745_),
    .A(_1744_));
 sg13g2_nor2_1 _4569_ (.A(net379),
    .B(_0888_),
    .Y(_1746_));
 sg13g2_nor2b_2 _4570_ (.A(_0890_),
    .B_N(_1746_),
    .Y(_1747_));
 sg13g2_o21ai_1 _4571_ (.B1(net427),
    .Y(_1748_),
    .A1(net715),
    .A2(_1747_));
 sg13g2_a21oi_1 _4572_ (.A1(net715),
    .A2(_1745_),
    .Y(_0375_),
    .B1(_1748_));
 sg13g2_a22oi_1 _4573_ (.Y(_1749_),
    .B1(_1747_),
    .B2(_1694_),
    .A2(_1744_),
    .A1(net700));
 sg13g2_nor2_1 _4574_ (.A(net413),
    .B(_1749_),
    .Y(_0376_));
 sg13g2_nand2_1 _4575_ (.Y(_1750_),
    .A(\snd.tune_pos[1] ),
    .B(\snd.tune_pos[0] ));
 sg13g2_xor2_1 _4576_ (.B(_1750_),
    .A(_0082_),
    .X(_1751_));
 sg13g2_a22oi_1 _4577_ (.Y(_1752_),
    .B1(_1747_),
    .B2(_1751_),
    .A2(_1744_),
    .A1(net688));
 sg13g2_nor2_1 _4578_ (.A(net413),
    .B(net689),
    .Y(_0377_));
 sg13g2_nor2_1 _4579_ (.A(net380),
    .B(_1736_),
    .Y(_1753_));
 sg13g2_a21oi_1 _4580_ (.A1(_0899_),
    .A2(_1736_),
    .Y(_1754_),
    .B1(net412));
 sg13g2_nor2b_1 _4581_ (.A(_1753_),
    .B_N(_1754_),
    .Y(_0378_));
 sg13g2_nand2_1 _4582_ (.Y(_1755_),
    .A(_0896_),
    .B(_1736_));
 sg13g2_o21ai_1 _4583_ (.B1(_1755_),
    .Y(_1756_),
    .A1(net742),
    .A2(_1736_));
 sg13g2_nor2_1 _4584_ (.A(net412),
    .B(_1756_),
    .Y(_0379_));
 sg13g2_nor2_1 _4585_ (.A(_1654_),
    .B(_1679_),
    .Y(_1757_));
 sg13g2_o21ai_1 _4586_ (.B1(_1757_),
    .Y(_1758_),
    .A1(_1651_),
    .A2(_1657_));
 sg13g2_nand3_1 _4587_ (.B(_1677_),
    .C(_1682_),
    .A(_1655_),
    .Y(_1759_));
 sg13g2_nor3_1 _4588_ (.A(_0080_),
    .B(_0891_),
    .C(_1720_),
    .Y(_1760_));
 sg13g2_a221oi_1 _4589_ (.B2(_0890_),
    .C1(_1760_),
    .B1(_1758_),
    .A1(_0887_),
    .Y(_1761_),
    .A2(_1746_));
 sg13g2_and3_1 _4590_ (.X(_1762_),
    .A(_1716_),
    .B(_1759_),
    .C(_1761_));
 sg13g2_or2_1 _4591_ (.X(_1763_),
    .B(_1762_),
    .A(net790));
 sg13g2_nand2_1 _4592_ (.Y(_1764_),
    .A(net790),
    .B(_1762_));
 sg13g2_and3_1 _4593_ (.X(_0380_),
    .A(net427),
    .B(_1763_),
    .C(_1764_));
 sg13g2_o21ai_1 _4594_ (.B1(net427),
    .Y(_1765_),
    .A1(_1776_),
    .A2(_1764_));
 sg13g2_a21oi_1 _4595_ (.A1(_1776_),
    .A2(_1764_),
    .Y(_0381_),
    .B1(_1765_));
 sg13g2_nor2_1 _4596_ (.A(_0787_),
    .B(_0788_),
    .Y(_1766_));
 sg13g2_nand2_2 _4597_ (.Y(_1767_),
    .A(_0790_),
    .B(_1766_));
 sg13g2_nand3_1 _4598_ (.B(net363),
    .C(_1767_),
    .A(net699),
    .Y(_1768_));
 sg13g2_o21ai_1 _4599_ (.B1(_1768_),
    .Y(_0382_),
    .A1(net344),
    .A2(_1767_));
 sg13g2_nand3_1 _4600_ (.B(net363),
    .C(_1767_),
    .A(net740),
    .Y(_1769_));
 sg13g2_o21ai_1 _4601_ (.B1(_1769_),
    .Y(_0383_),
    .A1(net343),
    .A2(_1767_));
 sg13g2_nand2_2 _4602_ (.Y(_1770_),
    .A(_0791_),
    .B(_1766_));
 sg13g2_nand3_1 _4603_ (.B(net363),
    .C(_1770_),
    .A(net745),
    .Y(_1771_));
 sg13g2_o21ai_1 _4604_ (.B1(_1771_),
    .Y(_0384_),
    .A1(net344),
    .A2(_1770_));
 sg13g2_nand3_1 _4605_ (.B(net362),
    .C(_1770_),
    .A(net776),
    .Y(_1772_));
 sg13g2_o21ai_1 _4606_ (.B1(_1772_),
    .Y(_0385_),
    .A1(net343),
    .A2(_1770_));
 sg13g2_nand2b_1 _4607_ (.Y(_1773_),
    .B(_0790_),
    .A_N(_1284_));
 sg13g2_nand3_1 _4608_ (.B(net363),
    .C(_1773_),
    .A(net644),
    .Y(_1774_));
 sg13g2_o21ai_1 _4609_ (.B1(_1774_),
    .Y(_0386_),
    .A1(net344),
    .A2(_1773_));
 sg13g2_nand3_1 _4610_ (.B(net362),
    .C(_1773_),
    .A(net747),
    .Y(_1775_));
 sg13g2_o21ai_1 _4611_ (.B1(_1775_),
    .Y(_0387_),
    .A1(net343),
    .A2(_1773_));
 sg13g2_nor3_1 _4612_ (.A(net411),
    .B(net562),
    .C(_1177_),
    .Y(_0280_));
 sg13g2_nor2_1 _4613_ (.A(_1179_),
    .B(_1180_),
    .Y(_0281_));
 sg13g2_a221oi_1 _4614_ (.B2(_1181_),
    .C1(net411),
    .B1(_1179_),
    .A1(_1808_),
    .Y(_0282_),
    .A2(_1178_));
 sg13g2_dfrbp_1 _4615_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net100),
    .D(_0093_),
    .Q_N(_2300_),
    .Q(\game.fsm.len2_color_count[0][0] ));
 sg13g2_dfrbp_1 _4616_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net257),
    .D(_0094_),
    .Q_N(_0045_),
    .Q(\game.fsm.len2_color_count[0][1] ));
 sg13g2_dfrbp_1 _4617_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net255),
    .D(_0095_),
    .Q_N(_2299_),
    .Q(\game.slv.lfsr[0] ));
 sg13g2_dfrbp_1 _4618_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net254),
    .D(_0096_),
    .Q_N(_2298_),
    .Q(\game.slv.lfsr[1] ));
 sg13g2_dfrbp_1 _4619_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net253),
    .D(net607),
    .Q_N(_2297_),
    .Q(\game.slv.lfsr[2] ));
 sg13g2_dfrbp_1 _4620_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net252),
    .D(_0098_),
    .Q_N(_2296_),
    .Q(\game.slv.lfsr[3] ));
 sg13g2_dfrbp_1 _4621_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net251),
    .D(_0099_),
    .Q_N(_2295_),
    .Q(\game.slv.lfsr[4] ));
 sg13g2_dfrbp_1 _4622_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net250),
    .D(_0100_),
    .Q_N(_2294_),
    .Q(\game.slv.lfsr[5] ));
 sg13g2_dfrbp_1 _4623_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net249),
    .D(_0101_),
    .Q_N(_2293_),
    .Q(\game.slv.lfsr[6] ));
 sg13g2_dfrbp_1 _4624_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net248),
    .D(_0102_),
    .Q_N(_2292_),
    .Q(\game.slv.lfsr[7] ));
 sg13g2_dfrbp_1 _4625_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net247),
    .D(_0103_),
    .Q_N(_2291_),
    .Q(\game.slv.lfsr[8] ));
 sg13g2_dfrbp_1 _4626_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net246),
    .D(_0104_),
    .Q_N(_2290_),
    .Q(\game.slv.lfsr[9] ));
 sg13g2_dfrbp_1 _4627_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net245),
    .D(_0105_),
    .Q_N(_2289_),
    .Q(\game.slv.lfsr[10] ));
 sg13g2_dfrbp_1 _4628_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net244),
    .D(_0106_),
    .Q_N(_2288_),
    .Q(\game.slv.lfsr[11] ));
 sg13g2_dfrbp_1 _4629_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net243),
    .D(_0107_),
    .Q_N(_2287_),
    .Q(\game.slv.lfsr[12] ));
 sg13g2_dfrbp_1 _4630_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net242),
    .D(_0108_),
    .Q_N(_2286_),
    .Q(\game.slv.lfsr[13] ));
 sg13g2_dfrbp_1 _4631_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net241),
    .D(_0109_),
    .Q_N(_2285_),
    .Q(\game.slv.lfsr[14] ));
 sg13g2_dfrbp_1 _4632_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net240),
    .D(_0110_),
    .Q_N(_2284_),
    .Q(\game.slv.lfsr[15] ));
 sg13g2_dfrbp_1 _4633_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net239),
    .D(_0111_),
    .Q_N(_2283_),
    .Q(\game.slv.lfsr[16] ));
 sg13g2_dfrbp_1 _4634_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net238),
    .D(_0112_),
    .Q_N(_2282_),
    .Q(\game.slv.lfsr[17] ));
 sg13g2_dfrbp_1 _4635_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net237),
    .D(_0113_),
    .Q_N(_2281_),
    .Q(\game.slv.lfsr[18] ));
 sg13g2_dfrbp_1 _4636_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net236),
    .D(_0114_),
    .Q_N(_2280_),
    .Q(\game.slv.lfsr[19] ));
 sg13g2_dfrbp_1 _4637_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net235),
    .D(_0115_),
    .Q_N(_2279_),
    .Q(\game.slv.lfsr[20] ));
 sg13g2_dfrbp_1 _4638_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net234),
    .D(_0116_),
    .Q_N(_2278_),
    .Q(\snd.note_sel[0] ));
 sg13g2_dfrbp_1 _4639_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net232),
    .D(net565),
    .Q_N(_2277_),
    .Q(\snd.note_sel[1] ));
 sg13g2_dfrbp_1 _4640_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net230),
    .D(_0118_),
    .Q_N(_2276_),
    .Q(\game.fsm.seq[4][0] ));
 sg13g2_dfrbp_1 _4641_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net228),
    .D(_0119_),
    .Q_N(_2275_),
    .Q(\game.fsm.seq[4][1] ));
 sg13g2_dfrbp_1 _4642_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net226),
    .D(net471),
    .Q_N(_2274_),
    .Q(\snd.note_timing[0] ));
 sg13g2_dfrbp_1 _4643_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net224),
    .D(_0121_),
    .Q_N(_2273_),
    .Q(\snd.note_timing[1] ));
 sg13g2_dfrbp_1 _4644_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net222),
    .D(net555),
    .Q_N(_2272_),
    .Q(\snd.note_timing[2] ));
 sg13g2_dfrbp_1 _4645_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net220),
    .D(_0123_),
    .Q_N(_2271_),
    .Q(\snd.note_timing[3] ));
 sg13g2_dfrbp_1 _4646_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net218),
    .D(_0124_),
    .Q_N(_2270_),
    .Q(\snd.note_timing[4] ));
 sg13g2_dfrbp_1 _4647_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net216),
    .D(_0125_),
    .Q_N(_2269_),
    .Q(\snd.note_timing[5] ));
 sg13g2_dfrbp_1 _4648_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net214),
    .D(net610),
    .Q_N(_2268_),
    .Q(\snd.note_timing[6] ));
 sg13g2_dfrbp_1 _4649_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net212),
    .D(_0127_),
    .Q_N(_2267_),
    .Q(\snd.note_timing[7] ));
 sg13g2_dfrbp_1 _4650_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net210),
    .D(_0128_),
    .Q_N(_2266_),
    .Q(\snd.note_timing[8] ));
 sg13g2_dfrbp_1 _4651_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net208),
    .D(_0129_),
    .Q_N(_2265_),
    .Q(\game.fsm.seq[5][0] ));
 sg13g2_dfrbp_1 _4652_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net207),
    .D(_0130_),
    .Q_N(_2264_),
    .Q(\game.fsm.seq[5][1] ));
 sg13g2_dfrbp_1 _4653_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net206),
    .D(_0131_),
    .Q_N(_0070_),
    .Q(\game.fsm.block_len[5][0] ));
 sg13g2_dfrbp_1 _4654_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net205),
    .D(_0132_),
    .Q_N(_0027_),
    .Q(\game.fsm.block_len[5][1] ));
 sg13g2_dfrbp_1 _4655_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net204),
    .D(_0133_),
    .Q_N(_0076_),
    .Q(\game.fsm.block_len[5][2] ));
 sg13g2_dfrbp_1 _4656_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net203),
    .D(_0134_),
    .Q_N(_0026_),
    .Q(\game.fsm.block_len[6][0] ));
 sg13g2_dfrbp_1 _4657_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net201),
    .D(_0135_),
    .Q_N(_0034_),
    .Q(\game.fsm.block_len[6][1] ));
 sg13g2_dfrbp_1 _4658_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net199),
    .D(_0136_),
    .Q_N(_0029_),
    .Q(\game.fsm.block_len[6][2] ));
 sg13g2_dfrbp_1 _4659_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net197),
    .D(_0137_),
    .Q_N(_2263_),
    .Q(\game.fsm.color_count[0][0] ));
 sg13g2_dfrbp_1 _4660_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net195),
    .D(_0138_),
    .Q_N(_2262_),
    .Q(\game.fsm.color_count[0][1] ));
 sg13g2_dfrbp_1 _4661_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net193),
    .D(_0139_),
    .Q_N(_2261_),
    .Q(\game.fsm.color_count[0][2] ));
 sg13g2_dfrbp_1 _4662_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net191),
    .D(_0140_),
    .Q_N(_0071_),
    .Q(\game.fsm.block_len[4][0] ));
 sg13g2_dfrbp_1 _4663_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net189),
    .D(_0141_),
    .Q_N(_0028_),
    .Q(\game.fsm.block_len[4][1] ));
 sg13g2_dfrbp_1 _4664_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net187),
    .D(_0142_),
    .Q_N(_0077_),
    .Q(\game.fsm.block_len[4][2] ));
 sg13g2_dfrbp_1 _4665_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net185),
    .D(_0143_),
    .Q_N(_0067_),
    .Q(\game.fsm.block_len[3][0] ));
 sg13g2_dfrbp_1 _4666_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net183),
    .D(_0144_),
    .Q_N(_0032_),
    .Q(\game.fsm.block_len[3][1] ));
 sg13g2_dfrbp_1 _4667_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net181),
    .D(_0145_),
    .Q_N(_0074_),
    .Q(\game.fsm.block_len[3][2] ));
 sg13g2_dfrbp_1 _4668_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net179),
    .D(_0146_),
    .Q_N(_0068_),
    .Q(\game.fsm.block_len[2][0] ));
 sg13g2_dfrbp_1 _4669_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net177),
    .D(_0147_),
    .Q_N(_0033_),
    .Q(\game.fsm.block_len[2][1] ));
 sg13g2_dfrbp_1 _4670_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net175),
    .D(_0148_),
    .Q_N(_0075_),
    .Q(\game.fsm.block_len[2][2] ));
 sg13g2_dfrbp_1 _4671_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net173),
    .D(_0149_),
    .Q_N(_0065_),
    .Q(\game.fsm.block_len[1][0] ));
 sg13g2_dfrbp_1 _4672_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net171),
    .D(_0150_),
    .Q_N(_0030_),
    .Q(\game.fsm.block_len[1][1] ));
 sg13g2_dfrbp_1 _4673_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net169),
    .D(_0151_),
    .Q_N(_0072_),
    .Q(\game.fsm.block_len[1][2] ));
 sg13g2_dfrbp_1 _4674_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net167),
    .D(net582),
    .Q_N(_0061_),
    .Q(\snd.chord[3][0] ));
 sg13g2_dfrbp_1 _4675_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net165),
    .D(_0153_),
    .Q_N(_2260_),
    .Q(\snd.counter[1] ));
 sg13g2_dfrbp_1 _4676_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net164),
    .D(net593),
    .Q_N(_2259_),
    .Q(\snd.counter[2] ));
 sg13g2_dfrbp_1 _4677_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net163),
    .D(_0155_),
    .Q_N(_2258_),
    .Q(\snd.counter[3] ));
 sg13g2_dfrbp_1 _4678_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net162),
    .D(_0156_),
    .Q_N(_2257_),
    .Q(\snd.counter[4] ));
 sg13g2_dfrbp_1 _4679_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net161),
    .D(_0157_),
    .Q_N(_2256_),
    .Q(\snd.counter[5] ));
 sg13g2_dfrbp_1 _4680_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net160),
    .D(_0158_),
    .Q_N(_2255_),
    .Q(\snd.counter[6] ));
 sg13g2_dfrbp_1 _4681_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net159),
    .D(_0159_),
    .Q_N(_2254_),
    .Q(\snd.counter[7] ));
 sg13g2_dfrbp_1 _4682_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net158),
    .D(_0160_),
    .Q_N(_2253_),
    .Q(\snd.counter[8] ));
 sg13g2_dfrbp_1 _4683_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net157),
    .D(_0161_),
    .Q_N(_0080_),
    .Q(\btn.gate_200hz ));
 sg13g2_dfrbp_1 _4684_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net156),
    .D(_0162_),
    .Q_N(_2252_),
    .Q(\game.slv.trigger ));
 sg13g2_dfrbp_1 _4685_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net155),
    .D(_0163_),
    .Q_N(_2251_),
    .Q(\game.slv.fsm_reset ));
 sg13g2_dfrbp_1 _4686_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net154),
    .D(_0164_),
    .Q_N(_2250_),
    .Q(\game.slv.fsm_update ));
 sg13g2_dfrbp_1 _4687_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net153),
    .D(_0165_),
    .Q_N(_2249_),
    .Q(\game.slv.fsm_color[0] ));
 sg13g2_dfrbp_1 _4688_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net152),
    .D(_0166_),
    .Q_N(_2248_),
    .Q(\game.slv.fsm_color[1] ));
 sg13g2_dfrbp_1 _4689_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net151),
    .D(net486),
    .Q_N(_2247_),
    .Q(\game.slv.saved_target ));
 sg13g2_dfrbp_1 _4690_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net149),
    .D(net714),
    .Q_N(_2246_),
    .Q(\game.slv.length[0] ));
 sg13g2_dfrbp_1 _4691_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net147),
    .D(_0169_),
    .Q_N(_2245_),
    .Q(\game.slv.length[1] ));
 sg13g2_dfrbp_1 _4692_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net145),
    .D(net619),
    .Q_N(_2244_),
    .Q(\game.slv.length[2] ));
 sg13g2_dfrbp_1 _4693_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net143),
    .D(net673),
    .Q_N(_0056_),
    .Q(\game.slv.pos[0] ));
 sg13g2_dfrbp_1 _4694_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net141),
    .D(net727),
    .Q_N(_2243_),
    .Q(\game.slv.pos[1] ));
 sg13g2_dfrbp_1 _4695_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net139),
    .D(net681),
    .Q_N(_2242_),
    .Q(\game.slv.pos[2] ));
 sg13g2_dfrbp_1 _4696_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net137),
    .D(net663),
    .Q_N(_2241_),
    .Q(\game.slv.retries[0] ));
 sg13g2_dfrbp_1 _4697_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net135),
    .D(net657),
    .Q_N(_2240_),
    .Q(\game.slv.retries[1] ));
 sg13g2_dfrbp_1 _4698_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net133),
    .D(net736),
    .Q_N(_2239_),
    .Q(\game.slv.retries[2] ));
 sg13g2_dfrbp_1 _4699_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net131),
    .D(net482),
    .Q_N(_2238_),
    .Q(\game.slv.ready ));
 sg13g2_dfrbp_1 _4700_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net130),
    .D(_0178_),
    .Q_N(_2237_),
    .Q(\game.fsm.seq[6][0] ));
 sg13g2_dfrbp_1 _4701_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net128),
    .D(_0179_),
    .Q_N(_2236_),
    .Q(\game.fsm.seq[6][1] ));
 sg13g2_dfrbp_1 _4702_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net126),
    .D(_0180_),
    .Q_N(_2235_),
    .Q(\game.fsm.len3_color_count[3][0] ));
 sg13g2_dfrbp_1 _4703_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net125),
    .D(_0181_),
    .Q_N(_0044_),
    .Q(\game.fsm.len3_color_count[3][1] ));
 sg13g2_dfrbp_1 _4704_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net124),
    .D(_0182_),
    .Q_N(_2234_),
    .Q(\game.fsm.color_count[3][0] ));
 sg13g2_dfrbp_1 _4705_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net123),
    .D(_0183_),
    .Q_N(_2233_),
    .Q(\game.fsm.color_count[3][1] ));
 sg13g2_dfrbp_1 _4706_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net101),
    .D(_0184_),
    .Q_N(_0024_),
    .Q(\game.fsm.color_count[3][2] ));
 sg13g2_dfrbp_1 _4707_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net102),
    .D(_0011_),
    .Q_N(_0083_),
    .Q(\game.slv.state[1] ));
 sg13g2_dfrbp_1 _4708_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net103),
    .D(_0012_),
    .Q_N(_2301_),
    .Q(\game.slv.state[2] ));
 sg13g2_dfrbp_1 _4709_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net104),
    .D(net683),
    .Q_N(_0039_),
    .Q(\game.slv.state[3] ));
 sg13g2_dfrbp_1 _4710_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net105),
    .D(_0000_),
    .Q_N(_2302_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _4711_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net106),
    .D(_0001_),
    .Q_N(_2303_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _4712_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net107),
    .D(_0002_),
    .Q_N(_2304_),
    .Q(_0016_));
 sg13g2_dfrbp_1 _4713_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net108),
    .D(_0003_),
    .Q_N(_2305_),
    .Q(_0017_));
 sg13g2_dfrbp_1 _4714_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net109),
    .D(_0004_),
    .Q_N(_2306_),
    .Q(_0018_));
 sg13g2_dfrbp_1 _4715_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net68),
    .D(_0005_),
    .Q_N(_2307_),
    .Q(_0019_));
 sg13g2_dfrbp_1 _4716_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net122),
    .D(_0006_),
    .Q_N(_2232_),
    .Q(_0020_));
 sg13g2_dfrbp_1 _4717_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net121),
    .D(_0185_),
    .Q_N(_2231_),
    .Q(\game.fsm.len1_color_count[1][0] ));
 sg13g2_dfrbp_1 _4718_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net119),
    .D(_0186_),
    .Q_N(_0050_),
    .Q(\game.fsm.len1_color_count[1][1] ));
 sg13g2_dfrbp_1 _4719_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net117),
    .D(_0187_),
    .Q_N(_0036_),
    .Q(\game.fsm.len1_color_count[1][2] ));
 sg13g2_dfrbp_1 _4720_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net115),
    .D(_0188_),
    .Q_N(_2230_),
    .Q(\game.fsm.len1_color_count[2][0] ));
 sg13g2_dfrbp_1 _4721_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net113),
    .D(_0189_),
    .Q_N(_0051_),
    .Q(\game.fsm.len1_color_count[2][1] ));
 sg13g2_dfrbp_1 _4722_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net111),
    .D(_0190_),
    .Q_N(_0038_),
    .Q(\game.fsm.len1_color_count[2][2] ));
 sg13g2_dfrbp_1 _4723_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net99),
    .D(net617),
    .Q_N(_0092_),
    .Q(\game.fsm.length[0] ));
 sg13g2_dfrbp_1 _4724_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net97),
    .D(_0192_),
    .Q_N(_0078_),
    .Q(\game.fsm.length[1] ));
 sg13g2_dfrbp_1 _4725_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net95),
    .D(_0193_),
    .Q_N(_0064_),
    .Q(\game.fsm.length[2] ));
 sg13g2_dfrbp_1 _4726_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net93),
    .D(net331),
    .Q_N(_0091_),
    .Q(\game.fsm.num_blocks[0] ));
 sg13g2_dfrbp_1 _4727_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net91),
    .D(_0195_),
    .Q_N(_2229_),
    .Q(\game.fsm.num_blocks[1] ));
 sg13g2_dfrbp_1 _4728_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net89),
    .D(_0196_),
    .Q_N(_0069_),
    .Q(\game.fsm.num_blocks[2] ));
 sg13g2_dfrbp_1 _4729_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net87),
    .D(net327),
    .Q_N(_0090_),
    .Q(\game.fsm.len1_block_count[0] ));
 sg13g2_dfrbp_1 _4730_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net85),
    .D(_0198_),
    .Q_N(_2228_),
    .Q(\game.fsm.len1_block_count[1] ));
 sg13g2_dfrbp_1 _4731_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net83),
    .D(_0199_),
    .Q_N(_2227_),
    .Q(\game.fsm.len1_block_count[2] ));
 sg13g2_dfrbp_1 _4732_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net81),
    .D(net329),
    .Q_N(_0089_),
    .Q(\game.fsm.len2_block_count[0] ));
 sg13g2_dfrbp_1 _4733_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net79),
    .D(_0201_),
    .Q_N(_2226_),
    .Q(\game.fsm.len2_block_count[1] ));
 sg13g2_dfrbp_1 _4734_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net77),
    .D(net443),
    .Q_N(_0088_),
    .Q(\game.fsm.len3_block_count[0] ));
 sg13g2_dfrbp_1 _4735_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net75),
    .D(_0203_),
    .Q_N(_2225_),
    .Q(\game.fsm.len3_block_count[1] ));
 sg13g2_dfrbp_1 _4736_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net73),
    .D(_0204_),
    .Q_N(_2224_),
    .Q(\game.fsm.green_block_count[0] ));
 sg13g2_dfrbp_1 _4737_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net71),
    .D(_0205_),
    .Q_N(_2223_),
    .Q(\game.fsm.green_block_count[1] ));
 sg13g2_dfrbp_1 _4738_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net69),
    .D(_0206_),
    .Q_N(_2222_),
    .Q(\game.fsm.green_block_count[2] ));
 sg13g2_dfrbp_1 _4739_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net67),
    .D(_0207_),
    .Q_N(_2221_),
    .Q(\game.challenge_num[0] ));
 sg13g2_dfrbp_1 _4740_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net65),
    .D(_0208_),
    .Q_N(_0053_),
    .Q(\game.challenge_num[1] ));
 sg13g2_dfrbp_1 _4741_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net63),
    .D(_0209_),
    .Q_N(_0054_),
    .Q(\game.challenge_num[2] ));
 sg13g2_dfrbp_1 _4742_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net61),
    .D(_0210_),
    .Q_N(_0055_),
    .Q(\game.challenge_num[3] ));
 sg13g2_dfrbp_1 _4743_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net59),
    .D(net464),
    .Q_N(_2220_),
    .Q(\game.challenge_mode ));
 sg13g2_dfrbp_1 _4744_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net57),
    .D(_0212_),
    .Q_N(_2219_),
    .Q(\game.input_erase ));
 sg13g2_dfrbp_1 _4745_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net56),
    .D(_0213_),
    .Q_N(_2218_),
    .Q(\game.solver_trigger_delayed ));
 sg13g2_dfrbp_1 _4746_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net54),
    .D(_0214_),
    .Q_N(_2217_),
    .Q(\game.slv.target[0] ));
 sg13g2_dfrbp_1 _4747_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net52),
    .D(_0215_),
    .Q_N(_2216_),
    .Q(\game.slv.target[1] ));
 sg13g2_dfrbp_1 _4748_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net50),
    .D(net525),
    .Q_N(_0022_),
    .Q(\game.current_level[0] ));
 sg13g2_dfrbp_1 _4749_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net48),
    .D(_0217_),
    .Q_N(_2215_),
    .Q(\game.current_level[1] ));
 sg13g2_dfrbp_1 _4750_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net46),
    .D(net789),
    .Q_N(_0086_),
    .Q(\game.current_level[2] ));
 sg13g2_dfrbp_1 _4751_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net44),
    .D(net775),
    .Q_N(_0085_),
    .Q(\game.current_level[3] ));
 sg13g2_dfrbp_1 _4752_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net42),
    .D(_0220_),
    .Q_N(_0084_),
    .Q(\game.current_level[4] ));
 sg13g2_dfrbp_1 _4753_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net40),
    .D(_0221_),
    .Q_N(_2214_),
    .Q(\game.fsm.read_pos[0] ));
 sg13g2_dfrbp_1 _4754_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net38),
    .D(_0222_),
    .Q_N(_2213_),
    .Q(\game.fsm.read_pos[1] ));
 sg13g2_dfrbp_1 _4755_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net36),
    .D(net679),
    .Q_N(_2212_),
    .Q(\game.fsm.read_pos[2] ));
 sg13g2_dfrbp_1 _4756_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net34),
    .D(_0224_),
    .Q_N(_2211_),
    .Q(\game.solver_active ));
 sg13g2_dfrbp_1 _4757_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net32),
    .D(net499),
    .Q_N(_2210_),
    .Q(\game.input_color[0] ));
 sg13g2_dfrbp_1 _4758_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net30),
    .D(net613),
    .Q_N(_2209_),
    .Q(\game.input_color[1] ));
 sg13g2_dfrbp_1 _4759_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net28),
    .D(_0227_),
    .Q_N(_2208_),
    .Q(\game.input_update ));
 sg13g2_dfrbp_1 _4760_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net27),
    .D(_0228_),
    .Q_N(_2207_),
    .Q(\game.input_reset ));
 sg13g2_dfrbp_1 _4761_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net26),
    .D(_0229_),
    .Q_N(_0021_),
    .Q(\dsp.digit ));
 sg13g2_dfrbp_1 _4762_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net25),
    .D(_0230_),
    .Q_N(_2206_),
    .Q(\dsp.digit_sel_raw[1] ));
 sg13g2_dfrbp_1 _4763_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net24),
    .D(net671),
    .Q_N(_2205_),
    .Q(\game.sound_mode[0] ));
 sg13g2_dfrbp_1 _4764_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net22),
    .D(_0232_),
    .Q_N(_2204_),
    .Q(\game.sound_mode[1] ));
 sg13g2_dfrbp_1 _4765_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net20),
    .D(_0233_),
    .Q_N(_0079_),
    .Q(\game.sound_mode[2] ));
 sg13g2_dfrbp_1 _4766_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net18),
    .D(_0234_),
    .Q_N(_2203_),
    .Q(display_graphical));
 sg13g2_dfrbp_1 _4767_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net16),
    .D(_0235_),
    .Q_N(_2202_),
    .Q(\display_value[0] ));
 sg13g2_dfrbp_1 _4768_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net14),
    .D(_0236_),
    .Q_N(_2201_),
    .Q(\display_value[1] ));
 sg13g2_dfrbp_1 _4769_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net12),
    .D(_0237_),
    .Q_N(_0057_),
    .Q(\display_value[2] ));
 sg13g2_dfrbp_1 _4770_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net10),
    .D(_0238_),
    .Q_N(_2200_),
    .Q(\display_value[3] ));
 sg13g2_dfrbp_1 _4771_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net8),
    .D(_0239_),
    .Q_N(_0060_),
    .Q(\display_value[4] ));
 sg13g2_dfrbp_1 _4772_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net311),
    .D(_0240_),
    .Q_N(_2199_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _4773_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net309),
    .D(_0241_),
    .Q_N(_2198_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _4774_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net307),
    .D(_0242_),
    .Q_N(_2197_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _4775_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net305),
    .D(_0243_),
    .Q_N(_2196_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _4776_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net303),
    .D(_0244_),
    .Q_N(_2195_),
    .Q(\game.fsm.len3_color_count[2][0] ));
 sg13g2_dfrbp_1 _4777_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net301),
    .D(_0245_),
    .Q_N(_0043_),
    .Q(\game.fsm.len3_color_count[2][1] ));
 sg13g2_dfrbp_1 _4778_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net299),
    .D(_0246_),
    .Q_N(_0063_),
    .Q(\game.fsm.seq[0][0] ));
 sg13g2_dfrbp_1 _4779_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net297),
    .D(_0247_),
    .Q_N(_2194_),
    .Q(\game.fsm.seq[0][1] ));
 sg13g2_dfrbp_1 _4780_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net295),
    .D(_0248_),
    .Q_N(_2193_),
    .Q(\game.fsm.len3_color_count[1][0] ));
 sg13g2_dfrbp_1 _4781_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net293),
    .D(_0249_),
    .Q_N(_0042_),
    .Q(\game.fsm.len3_color_count[1][1] ));
 sg13g2_dfrbp_1 _4782_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net291),
    .D(_0250_),
    .Q_N(_2192_),
    .Q(\game.fsm.len2_color_count[3][0] ));
 sg13g2_dfrbp_1 _4783_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net290),
    .D(_0251_),
    .Q_N(_0048_),
    .Q(\game.fsm.len2_color_count[3][1] ));
 sg13g2_dfrbp_1 _4784_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net289),
    .D(_0252_),
    .Q_N(_2191_),
    .Q(\game.fsm.len2_color_count[1][0] ));
 sg13g2_dfrbp_1 _4785_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net287),
    .D(_0253_),
    .Q_N(_0046_),
    .Q(\game.fsm.len2_color_count[1][1] ));
 sg13g2_dfrbp_1 _4786_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net285),
    .D(_0254_),
    .Q_N(_2190_),
    .Q(\game.fsm.len2_color_count[2][0] ));
 sg13g2_dfrbp_1 _4787_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net283),
    .D(_0255_),
    .Q_N(_0047_),
    .Q(\game.fsm.len2_color_count[2][1] ));
 sg13g2_dfrbp_1 _4788_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net281),
    .D(_0256_),
    .Q_N(_2189_),
    .Q(\game.fsm.len3_color_count[0][0] ));
 sg13g2_dfrbp_1 _4789_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net279),
    .D(_0257_),
    .Q_N(_0041_),
    .Q(\game.fsm.len3_color_count[0][1] ));
 sg13g2_dfrbp_1 _4790_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net277),
    .D(_0258_),
    .Q_N(_2188_),
    .Q(\game.fsm.len1_color_count[3][0] ));
 sg13g2_dfrbp_1 _4791_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net276),
    .D(_0259_),
    .Q_N(_0052_),
    .Q(\game.fsm.len1_color_count[3][1] ));
 sg13g2_dfrbp_1 _4792_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net275),
    .D(_0260_),
    .Q_N(_0037_),
    .Q(\game.fsm.len1_color_count[3][2] ));
 sg13g2_dfrbp_1 _4793_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net274),
    .D(_0261_),
    .Q_N(_0066_),
    .Q(\game.fsm.block_len[0][0] ));
 sg13g2_dfrbp_1 _4794_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net272),
    .D(_0262_),
    .Q_N(_0031_),
    .Q(\game.fsm.block_len[0][1] ));
 sg13g2_dfrbp_1 _4795_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net270),
    .D(_0263_),
    .Q_N(_0073_),
    .Q(\game.fsm.block_len[0][2] ));
 sg13g2_dfrbp_1 _4796_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net268),
    .D(_0264_),
    .Q_N(_2187_),
    .Q(\game.fsm.seq[7][0] ));
 sg13g2_dfrbp_1 _4797_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net267),
    .D(_0265_),
    .Q_N(_2186_),
    .Q(\game.fsm.seq[7][1] ));
 sg13g2_dfrbp_1 _4798_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net266),
    .D(_0266_),
    .Q_N(_2185_),
    .Q(\game.state[0] ));
 sg13g2_dfrbp_1 _4799_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net264),
    .D(_0267_),
    .Q_N(_2184_),
    .Q(\game.state[1] ));
 sg13g2_dfrbp_1 _4800_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net262),
    .D(_0268_),
    .Q_N(_2183_),
    .Q(\game.state[2] ));
 sg13g2_dfrbp_1 _4801_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net260),
    .D(_0269_),
    .Q_N(_2182_),
    .Q(\game.state[3] ));
 sg13g2_dfrbp_1 _4802_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net258),
    .D(_0270_),
    .Q_N(_2181_),
    .Q(\game.counter[0] ));
 sg13g2_dfrbp_1 _4803_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net233),
    .D(net739),
    .Q_N(_2180_),
    .Q(\game.counter[1] ));
 sg13g2_dfrbp_1 _4804_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net229),
    .D(_0272_),
    .Q_N(_2179_),
    .Q(\game.counter[2] ));
 sg13g2_dfrbp_1 _4805_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net225),
    .D(_0273_),
    .Q_N(_2178_),
    .Q(\game.counter[3] ));
 sg13g2_dfrbp_1 _4806_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net221),
    .D(_0274_),
    .Q_N(_2177_),
    .Q(\game.counter[4] ));
 sg13g2_dfrbp_1 _4807_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net217),
    .D(_0275_),
    .Q_N(_2176_),
    .Q(\game.counter[5] ));
 sg13g2_dfrbp_1 _4808_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net213),
    .D(_0276_),
    .Q_N(_2175_),
    .Q(\game.counter[6] ));
 sg13g2_dfrbp_1 _4809_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net209),
    .D(_0277_),
    .Q_N(_0058_),
    .Q(\game.counter[7] ));
 sg13g2_dfrbp_1 _4810_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net200),
    .D(_0278_),
    .Q_N(_2174_),
    .Q(\game.tune[0] ));
 sg13g2_dfrbp_1 _4811_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net196),
    .D(_0279_),
    .Q_N(_2173_),
    .Q(\game.tune[1] ));
 sg13g2_dfrbp_1 _4812_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net192),
    .D(_0280_),
    .Q_N(_2172_),
    .Q(_0007_));
 sg13g2_dfrbp_1 _4813_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net190),
    .D(_0281_),
    .Q_N(_2171_),
    .Q(_0008_));
 sg13g2_dfrbp_1 _4814_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net188),
    .D(_0282_),
    .Q_N(_2170_),
    .Q(_0009_));
 sg13g2_dfrbp_1 _4815_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net186),
    .D(_0283_),
    .Q_N(_2169_),
    .Q(\snd.counter[0] ));
 sg13g2_dfrbp_1 _4816_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net184),
    .D(_0284_),
    .Q_N(_0087_),
    .Q(\clk_div_counter[0] ));
 sg13g2_dfrbp_1 _4817_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net182),
    .D(_0285_),
    .Q_N(_2168_),
    .Q(\clk_div_counter[1] ));
 sg13g2_dfrbp_1 _4818_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net180),
    .D(net462),
    .Q_N(_2167_),
    .Q(\clk_div_counter[2] ));
 sg13g2_dfrbp_1 _4819_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net178),
    .D(_0287_),
    .Q_N(_2166_),
    .Q(\clk_div_counter[3] ));
 sg13g2_dfrbp_1 _4820_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net176),
    .D(_0288_),
    .Q_N(_2165_),
    .Q(\clk_div_counter[4] ));
 sg13g2_dfrbp_1 _4821_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net174),
    .D(_0289_),
    .Q_N(_2164_),
    .Q(\clk_div_counter[5] ));
 sg13g2_dfrbp_1 _4822_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net172),
    .D(_0290_),
    .Q_N(_2163_),
    .Q(\clk_div_counter[6] ));
 sg13g2_dfrbp_1 _4823_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net170),
    .D(_0291_),
    .Q_N(_2162_),
    .Q(\clk_div_counter[7] ));
 sg13g2_dfrbp_1 _4824_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net168),
    .D(net666),
    .Q_N(_0013_),
    .Q(\game.sound_on ));
 sg13g2_dfrbp_1 _4825_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net150),
    .D(_0293_),
    .Q_N(_2161_),
    .Q(\btn.long_press ));
 sg13g2_dfrbp_1 _4826_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net146),
    .D(_0294_),
    .Q_N(_2160_),
    .Q(\btn.current_event[0] ));
 sg13g2_dfrbp_1 _4827_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net142),
    .D(_0295_),
    .Q_N(_2159_),
    .Q(\btn.current_event[1] ));
 sg13g2_dfrbp_1 _4828_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net138),
    .D(_0296_),
    .Q_N(_2158_),
    .Q(\btn.current_event[2] ));
 sg13g2_dfrbp_1 _4829_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net134),
    .D(_0297_),
    .Q_N(_2157_),
    .Q(\btn.current_event[3] ));
 sg13g2_dfrbp_1 _4830_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net129),
    .D(_0298_),
    .Q_N(_2156_),
    .Q(\btn.change_timer[0] ));
 sg13g2_dfrbp_1 _4831_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net120),
    .D(_0299_),
    .Q_N(_2155_),
    .Q(\btn.change_timer[1] ));
 sg13g2_dfrbp_1 _4832_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net116),
    .D(_0300_),
    .Q_N(_2154_),
    .Q(\btn.change_timer[2] ));
 sg13g2_dfrbp_1 _4833_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net112),
    .D(_0301_),
    .Q_N(_2153_),
    .Q(\btn.change_timer[3] ));
 sg13g2_dfrbp_1 _4834_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net98),
    .D(net698),
    .Q_N(_2152_),
    .Q(\btn.change_timer[4] ));
 sg13g2_dfrbp_1 _4835_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net94),
    .D(net577),
    .Q_N(_2151_),
    .Q(\btn.change_timer[5] ));
 sg13g2_dfrbp_1 _4836_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net90),
    .D(_0304_),
    .Q_N(_2150_),
    .Q(\btn.change_timer[6] ));
 sg13g2_dfrbp_1 _4837_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net86),
    .D(net491),
    .Q_N(_2149_),
    .Q(\btn.sample_15ms[0] ));
 sg13g2_dfrbp_1 _4838_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net82),
    .D(net543),
    .Q_N(_2148_),
    .Q(\btn.sample_15ms[1] ));
 sg13g2_dfrbp_1 _4839_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net78),
    .D(net521),
    .Q_N(_2147_),
    .Q(\btn.sample_15ms[2] ));
 sg13g2_dfrbp_1 _4840_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net74),
    .D(_0308_),
    .Q_N(_2146_),
    .Q(\btn.sample_15ms[3] ));
 sg13g2_dfrbp_1 _4841_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net70),
    .D(_0309_),
    .Q_N(_2145_),
    .Q(\btn.sample_10ms[0] ));
 sg13g2_dfrbp_1 _4842_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net66),
    .D(net528),
    .Q_N(_2144_),
    .Q(\btn.sample_10ms[1] ));
 sg13g2_dfrbp_1 _4843_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net62),
    .D(_0311_),
    .Q_N(_2143_),
    .Q(\btn.sample_10ms[2] ));
 sg13g2_dfrbp_1 _4844_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net58),
    .D(net501),
    .Q_N(_2142_),
    .Q(\btn.sample_10ms[3] ));
 sg13g2_dfrbp_1 _4845_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net53),
    .D(_0313_),
    .Q_N(_2141_),
    .Q(\btn.sample_5ms[0] ));
 sg13g2_dfrbp_1 _4846_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net49),
    .D(_0314_),
    .Q_N(_2140_),
    .Q(\btn.sample_5ms[1] ));
 sg13g2_dfrbp_1 _4847_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net45),
    .D(_0315_),
    .Q_N(_2139_),
    .Q(\btn.sample_5ms[2] ));
 sg13g2_dfrbp_1 _4848_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net41),
    .D(net631),
    .Q_N(_2138_),
    .Q(\btn.sample_5ms[3] ));
 sg13g2_dfrbp_1 _4849_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net37),
    .D(_0317_),
    .Q_N(_2137_),
    .Q(\btn.button_state[0] ));
 sg13g2_dfrbp_1 _4850_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net33),
    .D(_0318_),
    .Q_N(_2136_),
    .Q(\btn.button_state[1] ));
 sg13g2_dfrbp_1 _4851_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net29),
    .D(_0319_),
    .Q_N(_2135_),
    .Q(\btn.button_state[2] ));
 sg13g2_dfrbp_1 _4852_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net21),
    .D(_0320_),
    .Q_N(_2134_),
    .Q(\btn.button_state[3] ));
 sg13g2_dfrbp_1 _4853_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net17),
    .D(_0321_),
    .Q_N(_2133_),
    .Q(\dsp.segments_raw[0] ));
 sg13g2_dfrbp_1 _4854_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net15),
    .D(net761),
    .Q_N(_2132_),
    .Q(\dsp.segments_raw[1] ));
 sg13g2_dfrbp_1 _4855_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net13),
    .D(_0323_),
    .Q_N(_2131_),
    .Q(\dsp.segments_raw[2] ));
 sg13g2_dfrbp_1 _4856_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net11),
    .D(net763),
    .Q_N(_2130_),
    .Q(\dsp.segments_raw[3] ));
 sg13g2_dfrbp_1 _4857_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net9),
    .D(_0325_),
    .Q_N(_2129_),
    .Q(\dsp.segments_raw[4] ));
 sg13g2_dfrbp_1 _4858_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net312),
    .D(net456),
    .Q_N(_2128_),
    .Q(\dsp.segments_raw[5] ));
 sg13g2_dfrbp_1 _4859_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net310),
    .D(_0327_),
    .Q_N(_2127_),
    .Q(\dsp.segments_raw[6] ));
 sg13g2_dfrbp_1 _4860_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net308),
    .D(_0328_),
    .Q_N(_2126_),
    .Q(\btn.input_event[0] ));
 sg13g2_dfrbp_1 _4861_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net306),
    .D(_0329_),
    .Q_N(_2125_),
    .Q(\btn.input_event[1] ));
 sg13g2_dfrbp_1 _4862_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net304),
    .D(_0330_),
    .Q_N(_2124_),
    .Q(\btn.input_event[2] ));
 sg13g2_dfrbp_1 _4863_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net302),
    .D(_0331_),
    .Q_N(_2123_),
    .Q(\btn.input_event[3] ));
 sg13g2_dfrbp_1 _4864_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net300),
    .D(_0332_),
    .Q_N(_0040_),
    .Q(\btn.input_event[4] ));
 sg13g2_dfrbp_1 _4865_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net298),
    .D(_0333_),
    .Q_N(_2122_),
    .Q(\game.fsm.len1_color_count[0][0] ));
 sg13g2_dfrbp_1 _4866_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net294),
    .D(_0334_),
    .Q_N(_0049_),
    .Q(\game.fsm.len1_color_count[0][1] ));
 sg13g2_dfrbp_1 _4867_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net288),
    .D(_0335_),
    .Q_N(_0035_),
    .Q(\game.fsm.len1_color_count[0][2] ));
 sg13g2_dfrbp_1 _4868_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net284),
    .D(_0336_),
    .Q_N(_2121_),
    .Q(\game.fsm.color_count[2][0] ));
 sg13g2_dfrbp_1 _4869_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net280),
    .D(_0337_),
    .Q_N(_2120_),
    .Q(\game.fsm.color_count[2][1] ));
 sg13g2_dfrbp_1 _4870_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net273),
    .D(_0338_),
    .Q_N(_0025_),
    .Q(\game.fsm.color_count[2][2] ));
 sg13g2_dfrbp_1 _4871_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net269),
    .D(_0339_),
    .Q_N(_2119_),
    .Q(\game.fsm.color_count[1][0] ));
 sg13g2_dfrbp_1 _4872_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net263),
    .D(_0340_),
    .Q_N(_2118_),
    .Q(\game.fsm.color_count[1][1] ));
 sg13g2_dfrbp_1 _4873_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net259),
    .D(_0341_),
    .Q_N(_0023_),
    .Q(\game.fsm.color_count[1][2] ));
 sg13g2_dfrbp_1 _4874_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net231),
    .D(_0342_),
    .Q_N(_2117_),
    .Q(\game.fsm.block_len[7][0] ));
 sg13g2_dfrbp_1 _4875_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net227),
    .D(_0343_),
    .Q_N(_2116_),
    .Q(\game.fsm.block_len[7][1] ));
 sg13g2_dfrbp_1 _4876_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net223),
    .D(_0344_),
    .Q_N(_2115_),
    .Q(\game.fsm.block_len[7][2] ));
 sg13g2_dfrbp_1 _4877_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net219),
    .D(net570),
    .Q_N(_2114_),
    .Q(\snd.sound ));
 sg13g2_dfrbp_1 _4878_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net211),
    .D(_0346_),
    .Q_N(_2113_),
    .Q(\snd.next_note_timing[0] ));
 sg13g2_dfrbp_1 _4879_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net198),
    .D(_0347_),
    .Q_N(_2112_),
    .Q(\snd.next_note_timing[1] ));
 sg13g2_dfrbp_1 _4880_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net166),
    .D(_0348_),
    .Q_N(_2111_),
    .Q(\snd.next_note_timing[2] ));
 sg13g2_dfrbp_1 _4881_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net144),
    .D(_0349_),
    .Q_N(_2110_),
    .Q(\snd.next_note_timing[3] ));
 sg13g2_dfrbp_1 _4882_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net136),
    .D(_0350_),
    .Q_N(_2109_),
    .Q(\snd.next_note_timing[4] ));
 sg13g2_dfrbp_1 _4883_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net127),
    .D(_0351_),
    .Q_N(_2108_),
    .Q(\snd.next_note_timing[5] ));
 sg13g2_dfrbp_1 _4884_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net114),
    .D(_0352_),
    .Q_N(_2107_),
    .Q(\snd.next_note_timing[6] ));
 sg13g2_dfrbp_1 _4885_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net96),
    .D(_0353_),
    .Q_N(_2106_),
    .Q(\snd.next_note_timing[7] ));
 sg13g2_dfrbp_1 _4886_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net88),
    .D(_0354_),
    .Q_N(_2105_),
    .Q(\snd.next_note_timing[8] ));
 sg13g2_dfrbp_1 _4887_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net80),
    .D(_0355_),
    .Q_N(_2104_),
    .Q(\snd.next_note_sel[0] ));
 sg13g2_dfrbp_1 _4888_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net72),
    .D(_0356_),
    .Q_N(_2103_),
    .Q(\snd.next_note_sel[1] ));
 sg13g2_dfrbp_1 _4889_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net64),
    .D(net694),
    .Q_N(_2102_),
    .Q(\snd.chord[2][2] ));
 sg13g2_dfrbp_1 _4890_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net55),
    .D(_0358_),
    .Q_N(_2101_),
    .Q(\snd.chord[1][0] ));
 sg13g2_dfrbp_1 _4891_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net47),
    .D(net725),
    .Q_N(_2100_),
    .Q(\snd.chord[1][5] ));
 sg13g2_dfrbp_1 _4892_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net39),
    .D(_0360_),
    .Q_N(_2099_),
    .Q(\game.next_state[0] ));
 sg13g2_dfrbp_1 _4893_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net31),
    .D(_0361_),
    .Q_N(_2098_),
    .Q(\game.next_state[2] ));
 sg13g2_dfrbp_1 _4894_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net19),
    .D(_0362_),
    .Q_N(_0059_),
    .Q(\snd.chord[0][0] ));
 sg13g2_dfrbp_1 _4895_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net292),
    .D(_0363_),
    .Q_N(_2097_),
    .Q(\snd.chord[0][1] ));
 sg13g2_dfrbp_1 _4896_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net282),
    .D(_0364_),
    .Q_N(_2096_),
    .Q(\snd.chord[0][2] ));
 sg13g2_dfrbp_1 _4897_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net271),
    .D(net676),
    .Q_N(_2095_),
    .Q(\snd.chord[0][3] ));
 sg13g2_dfrbp_1 _4898_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net261),
    .D(_0366_),
    .Q_N(_2094_),
    .Q(\snd.chord[0][4] ));
 sg13g2_dfrbp_1 _4899_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net215),
    .D(_0367_),
    .Q_N(_2093_),
    .Q(\snd.chord[0][5] ));
 sg13g2_dfrbp_1 _4900_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net194),
    .D(_0368_),
    .Q_N(_2092_),
    .Q(\snd.tune_counter[0] ));
 sg13g2_dfrbp_1 _4901_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net140),
    .D(_0369_),
    .Q_N(_2091_),
    .Q(\snd.tune_counter[1] ));
 sg13g2_dfrbp_1 _4902_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net118),
    .D(_0370_),
    .Q_N(_2090_),
    .Q(\snd.tune_counter[2] ));
 sg13g2_dfrbp_1 _4903_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net92),
    .D(_0371_),
    .Q_N(_2089_),
    .Q(\snd.tune_counter[3] ));
 sg13g2_dfrbp_1 _4904_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net76),
    .D(_0372_),
    .Q_N(_2088_),
    .Q(\snd.tune_counter[4] ));
 sg13g2_dfrbp_1 _4905_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net60),
    .D(_0373_),
    .Q_N(_2087_),
    .Q(\snd.tune_counter[5] ));
 sg13g2_dfrbp_1 _4906_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net43),
    .D(net550),
    .Q_N(_0081_),
    .Q(\snd.tune_counter[6] ));
 sg13g2_dfrbp_1 _4907_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net23),
    .D(_0375_),
    .Q_N(_2086_),
    .Q(\snd.tune_pos[0] ));
 sg13g2_dfrbp_1 _4908_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net286),
    .D(_0376_),
    .Q_N(_2085_),
    .Q(\snd.tune_pos[1] ));
 sg13g2_dfrbp_1 _4909_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net265),
    .D(_0377_),
    .Q_N(_0082_),
    .Q(\snd.tune_pos[2] ));
 sg13g2_dfrbp_1 _4910_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net202),
    .D(_0378_),
    .Q_N(_2084_),
    .Q(\snd.active_tune[0] ));
 sg13g2_dfrbp_1 _4911_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net132),
    .D(_0379_),
    .Q_N(_2083_),
    .Q(\snd.active_tune[1] ));
 sg13g2_dfrbp_1 _4912_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net84),
    .D(_0380_),
    .Q_N(_2082_),
    .Q(\snd.sequencer_state[0] ));
 sg13g2_dfrbp_1 _4913_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net51),
    .D(net702),
    .Q_N(_2081_),
    .Q(\snd.sequencer_state[1] ));
 sg13g2_dfrbp_1 _4914_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net296),
    .D(_0382_),
    .Q_N(_2080_),
    .Q(\game.fsm.seq[3][0] ));
 sg13g2_dfrbp_1 _4915_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net256),
    .D(_0383_),
    .Q_N(_2079_),
    .Q(\game.fsm.seq[3][1] ));
 sg13g2_dfrbp_1 _4916_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net110),
    .D(_0384_),
    .Q_N(_2078_),
    .Q(\game.fsm.seq[2][0] ));
 sg13g2_dfrbp_1 _4917_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net35),
    .D(_0385_),
    .Q_N(_2077_),
    .Q(\game.fsm.seq[2][1] ));
 sg13g2_dfrbp_1 _4918_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net148),
    .D(_0386_),
    .Q_N(_0062_),
    .Q(\game.fsm.seq[1][0] ));
 sg13g2_dfrbp_1 _4919_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net278),
    .D(_0387_),
    .Q_N(_2076_),
    .Q(\game.fsm.seq[1][1] ));
 sg13g2_tiehi _4857__9 (.L_HI(net9));
 sg13g2_tiehi _4770__10 (.L_HI(net10));
 sg13g2_tiehi _4856__11 (.L_HI(net11));
 sg13g2_tiehi _4769__12 (.L_HI(net12));
 sg13g2_tiehi _4855__13 (.L_HI(net13));
 sg13g2_tiehi _4768__14 (.L_HI(net14));
 sg13g2_tiehi _4854__15 (.L_HI(net15));
 sg13g2_tiehi _4767__16 (.L_HI(net16));
 sg13g2_tiehi _4853__17 (.L_HI(net17));
 sg13g2_tiehi _4766__18 (.L_HI(net18));
 sg13g2_tiehi _4894__19 (.L_HI(net19));
 sg13g2_tiehi _4765__20 (.L_HI(net20));
 sg13g2_tiehi _4852__21 (.L_HI(net21));
 sg13g2_tiehi _4764__22 (.L_HI(net22));
 sg13g2_tiehi _4907__23 (.L_HI(net23));
 sg13g2_tiehi _4763__24 (.L_HI(net24));
 sg13g2_tiehi _4762__25 (.L_HI(net25));
 sg13g2_tiehi _4761__26 (.L_HI(net26));
 sg13g2_tiehi _4760__27 (.L_HI(net27));
 sg13g2_tiehi _4759__28 (.L_HI(net28));
 sg13g2_tiehi _4851__29 (.L_HI(net29));
 sg13g2_tiehi _4758__30 (.L_HI(net30));
 sg13g2_tiehi _4893__31 (.L_HI(net31));
 sg13g2_tiehi _4757__32 (.L_HI(net32));
 sg13g2_tiehi _4850__33 (.L_HI(net33));
 sg13g2_tiehi _4756__34 (.L_HI(net34));
 sg13g2_tiehi _4917__35 (.L_HI(net35));
 sg13g2_tiehi _4755__36 (.L_HI(net36));
 sg13g2_tiehi _4849__37 (.L_HI(net37));
 sg13g2_tiehi _4754__38 (.L_HI(net38));
 sg13g2_tiehi _4892__39 (.L_HI(net39));
 sg13g2_tiehi _4753__40 (.L_HI(net40));
 sg13g2_tiehi _4848__41 (.L_HI(net41));
 sg13g2_tiehi _4752__42 (.L_HI(net42));
 sg13g2_tiehi _4906__43 (.L_HI(net43));
 sg13g2_tiehi _4751__44 (.L_HI(net44));
 sg13g2_tiehi _4847__45 (.L_HI(net45));
 sg13g2_tiehi _4750__46 (.L_HI(net46));
 sg13g2_tiehi _4891__47 (.L_HI(net47));
 sg13g2_tiehi _4749__48 (.L_HI(net48));
 sg13g2_tiehi _4846__49 (.L_HI(net49));
 sg13g2_tiehi _4748__50 (.L_HI(net50));
 sg13g2_tiehi _4913__51 (.L_HI(net51));
 sg13g2_tiehi _4747__52 (.L_HI(net52));
 sg13g2_tiehi _4845__53 (.L_HI(net53));
 sg13g2_tiehi _4746__54 (.L_HI(net54));
 sg13g2_tiehi _4890__55 (.L_HI(net55));
 sg13g2_tiehi _4745__56 (.L_HI(net56));
 sg13g2_tiehi _4744__57 (.L_HI(net57));
 sg13g2_tiehi _4844__58 (.L_HI(net58));
 sg13g2_tiehi _4743__59 (.L_HI(net59));
 sg13g2_tiehi _4905__60 (.L_HI(net60));
 sg13g2_tiehi _4742__61 (.L_HI(net61));
 sg13g2_tiehi _4843__62 (.L_HI(net62));
 sg13g2_tiehi _4741__63 (.L_HI(net63));
 sg13g2_tiehi _4889__64 (.L_HI(net64));
 sg13g2_tiehi _4740__65 (.L_HI(net65));
 sg13g2_tiehi _4842__66 (.L_HI(net66));
 sg13g2_tiehi _4739__67 (.L_HI(net67));
 sg13g2_tiehi _4715__68 (.L_HI(net68));
 sg13g2_tiehi _4738__69 (.L_HI(net69));
 sg13g2_tiehi _4841__70 (.L_HI(net70));
 sg13g2_tiehi _4737__71 (.L_HI(net71));
 sg13g2_tiehi _4888__72 (.L_HI(net72));
 sg13g2_tiehi _4736__73 (.L_HI(net73));
 sg13g2_tiehi _4840__74 (.L_HI(net74));
 sg13g2_tiehi _4735__75 (.L_HI(net75));
 sg13g2_tiehi _4904__76 (.L_HI(net76));
 sg13g2_tiehi _4734__77 (.L_HI(net77));
 sg13g2_tiehi _4839__78 (.L_HI(net78));
 sg13g2_tiehi _4733__79 (.L_HI(net79));
 sg13g2_tiehi _4887__80 (.L_HI(net80));
 sg13g2_tiehi _4732__81 (.L_HI(net81));
 sg13g2_tiehi _4838__82 (.L_HI(net82));
 sg13g2_tiehi _4731__83 (.L_HI(net83));
 sg13g2_tiehi _4912__84 (.L_HI(net84));
 sg13g2_tiehi _4730__85 (.L_HI(net85));
 sg13g2_tiehi _4837__86 (.L_HI(net86));
 sg13g2_tiehi _4729__87 (.L_HI(net87));
 sg13g2_tiehi _4886__88 (.L_HI(net88));
 sg13g2_tiehi _4728__89 (.L_HI(net89));
 sg13g2_tiehi _4836__90 (.L_HI(net90));
 sg13g2_tiehi _4727__91 (.L_HI(net91));
 sg13g2_tiehi _4903__92 (.L_HI(net92));
 sg13g2_tiehi _4726__93 (.L_HI(net93));
 sg13g2_tiehi _4835__94 (.L_HI(net94));
 sg13g2_tiehi _4725__95 (.L_HI(net95));
 sg13g2_tiehi _4885__96 (.L_HI(net96));
 sg13g2_tiehi _4724__97 (.L_HI(net97));
 sg13g2_tiehi _4834__98 (.L_HI(net98));
 sg13g2_tiehi _4723__99 (.L_HI(net99));
 sg13g2_tiehi _4615__100 (.L_HI(net100));
 sg13g2_tiehi _4706__101 (.L_HI(net101));
 sg13g2_tiehi _4707__102 (.L_HI(net102));
 sg13g2_tiehi _4708__103 (.L_HI(net103));
 sg13g2_tiehi _4709__104 (.L_HI(net104));
 sg13g2_tiehi _4710__105 (.L_HI(net105));
 sg13g2_tiehi _4711__106 (.L_HI(net106));
 sg13g2_tiehi _4712__107 (.L_HI(net107));
 sg13g2_tiehi _4713__108 (.L_HI(net108));
 sg13g2_tiehi _4714__109 (.L_HI(net109));
 sg13g2_tiehi _4916__110 (.L_HI(net110));
 sg13g2_tiehi _4722__111 (.L_HI(net111));
 sg13g2_tiehi _4833__112 (.L_HI(net112));
 sg13g2_tiehi _4721__113 (.L_HI(net113));
 sg13g2_tiehi _4884__114 (.L_HI(net114));
 sg13g2_tiehi _4720__115 (.L_HI(net115));
 sg13g2_tiehi _4832__116 (.L_HI(net116));
 sg13g2_tiehi _4719__117 (.L_HI(net117));
 sg13g2_tiehi _4902__118 (.L_HI(net118));
 sg13g2_tiehi _4718__119 (.L_HI(net119));
 sg13g2_tiehi _4831__120 (.L_HI(net120));
 sg13g2_tiehi _4717__121 (.L_HI(net121));
 sg13g2_tiehi _4716__122 (.L_HI(net122));
 sg13g2_tiehi _4705__123 (.L_HI(net123));
 sg13g2_tiehi _4704__124 (.L_HI(net124));
 sg13g2_tiehi _4703__125 (.L_HI(net125));
 sg13g2_tiehi _4702__126 (.L_HI(net126));
 sg13g2_tiehi _4883__127 (.L_HI(net127));
 sg13g2_tiehi _4701__128 (.L_HI(net128));
 sg13g2_tiehi _4830__129 (.L_HI(net129));
 sg13g2_tiehi _4700__130 (.L_HI(net130));
 sg13g2_tiehi _4699__131 (.L_HI(net131));
 sg13g2_tiehi _4911__132 (.L_HI(net132));
 sg13g2_tiehi _4698__133 (.L_HI(net133));
 sg13g2_tiehi _4829__134 (.L_HI(net134));
 sg13g2_tiehi _4697__135 (.L_HI(net135));
 sg13g2_tiehi _4882__136 (.L_HI(net136));
 sg13g2_tiehi _4696__137 (.L_HI(net137));
 sg13g2_tiehi _4828__138 (.L_HI(net138));
 sg13g2_tiehi _4695__139 (.L_HI(net139));
 sg13g2_tiehi _4901__140 (.L_HI(net140));
 sg13g2_tiehi _4694__141 (.L_HI(net141));
 sg13g2_tiehi _4827__142 (.L_HI(net142));
 sg13g2_tiehi _4693__143 (.L_HI(net143));
 sg13g2_tiehi _4881__144 (.L_HI(net144));
 sg13g2_tiehi _4692__145 (.L_HI(net145));
 sg13g2_tiehi _4826__146 (.L_HI(net146));
 sg13g2_tiehi _4691__147 (.L_HI(net147));
 sg13g2_tiehi _4918__148 (.L_HI(net148));
 sg13g2_tiehi _4690__149 (.L_HI(net149));
 sg13g2_tiehi _4825__150 (.L_HI(net150));
 sg13g2_tiehi _4689__151 (.L_HI(net151));
 sg13g2_tiehi _4688__152 (.L_HI(net152));
 sg13g2_tiehi _4687__153 (.L_HI(net153));
 sg13g2_tiehi _4686__154 (.L_HI(net154));
 sg13g2_tiehi _4685__155 (.L_HI(net155));
 sg13g2_tiehi _4684__156 (.L_HI(net156));
 sg13g2_tiehi _4683__157 (.L_HI(net157));
 sg13g2_tiehi _4682__158 (.L_HI(net158));
 sg13g2_tiehi _4681__159 (.L_HI(net159));
 sg13g2_tiehi _4680__160 (.L_HI(net160));
 sg13g2_tiehi _4679__161 (.L_HI(net161));
 sg13g2_tiehi _4678__162 (.L_HI(net162));
 sg13g2_tiehi _4677__163 (.L_HI(net163));
 sg13g2_tiehi _4676__164 (.L_HI(net164));
 sg13g2_tiehi _4675__165 (.L_HI(net165));
 sg13g2_tiehi _4880__166 (.L_HI(net166));
 sg13g2_tiehi _4674__167 (.L_HI(net167));
 sg13g2_tiehi _4824__168 (.L_HI(net168));
 sg13g2_tiehi _4673__169 (.L_HI(net169));
 sg13g2_tiehi _4823__170 (.L_HI(net170));
 sg13g2_tiehi _4672__171 (.L_HI(net171));
 sg13g2_tiehi _4822__172 (.L_HI(net172));
 sg13g2_tiehi _4671__173 (.L_HI(net173));
 sg13g2_tiehi _4821__174 (.L_HI(net174));
 sg13g2_tiehi _4670__175 (.L_HI(net175));
 sg13g2_tiehi _4820__176 (.L_HI(net176));
 sg13g2_tiehi _4669__177 (.L_HI(net177));
 sg13g2_tiehi _4819__178 (.L_HI(net178));
 sg13g2_tiehi _4668__179 (.L_HI(net179));
 sg13g2_tiehi _4818__180 (.L_HI(net180));
 sg13g2_tiehi _4667__181 (.L_HI(net181));
 sg13g2_tiehi _4817__182 (.L_HI(net182));
 sg13g2_tiehi _4666__183 (.L_HI(net183));
 sg13g2_tiehi _4816__184 (.L_HI(net184));
 sg13g2_tiehi _4665__185 (.L_HI(net185));
 sg13g2_tiehi _4815__186 (.L_HI(net186));
 sg13g2_tiehi _4664__187 (.L_HI(net187));
 sg13g2_tiehi _4814__188 (.L_HI(net188));
 sg13g2_tiehi _4663__189 (.L_HI(net189));
 sg13g2_tiehi _4813__190 (.L_HI(net190));
 sg13g2_tiehi _4662__191 (.L_HI(net191));
 sg13g2_tiehi _4812__192 (.L_HI(net192));
 sg13g2_tiehi _4661__193 (.L_HI(net193));
 sg13g2_tiehi _4900__194 (.L_HI(net194));
 sg13g2_tiehi _4660__195 (.L_HI(net195));
 sg13g2_tiehi _4811__196 (.L_HI(net196));
 sg13g2_tiehi _4659__197 (.L_HI(net197));
 sg13g2_tiehi _4879__198 (.L_HI(net198));
 sg13g2_tiehi _4658__199 (.L_HI(net199));
 sg13g2_tiehi _4810__200 (.L_HI(net200));
 sg13g2_tiehi _4657__201 (.L_HI(net201));
 sg13g2_tiehi _4910__202 (.L_HI(net202));
 sg13g2_tiehi _4656__203 (.L_HI(net203));
 sg13g2_tiehi _4655__204 (.L_HI(net204));
 sg13g2_tiehi _4654__205 (.L_HI(net205));
 sg13g2_tiehi _4653__206 (.L_HI(net206));
 sg13g2_tiehi _4652__207 (.L_HI(net207));
 sg13g2_tiehi _4651__208 (.L_HI(net208));
 sg13g2_tiehi _4809__209 (.L_HI(net209));
 sg13g2_tiehi _4650__210 (.L_HI(net210));
 sg13g2_tiehi _4878__211 (.L_HI(net211));
 sg13g2_tiehi _4649__212 (.L_HI(net212));
 sg13g2_tiehi _4808__213 (.L_HI(net213));
 sg13g2_tiehi _4648__214 (.L_HI(net214));
 sg13g2_tiehi _4899__215 (.L_HI(net215));
 sg13g2_tiehi _4647__216 (.L_HI(net216));
 sg13g2_tiehi _4807__217 (.L_HI(net217));
 sg13g2_tiehi _4646__218 (.L_HI(net218));
 sg13g2_tiehi _4877__219 (.L_HI(net219));
 sg13g2_tiehi _4645__220 (.L_HI(net220));
 sg13g2_tiehi _4806__221 (.L_HI(net221));
 sg13g2_tiehi _4644__222 (.L_HI(net222));
 sg13g2_tiehi _4876__223 (.L_HI(net223));
 sg13g2_tiehi _4643__224 (.L_HI(net224));
 sg13g2_tiehi _4805__225 (.L_HI(net225));
 sg13g2_tiehi _4642__226 (.L_HI(net226));
 sg13g2_tiehi _4875__227 (.L_HI(net227));
 sg13g2_tiehi _4641__228 (.L_HI(net228));
 sg13g2_tiehi _4804__229 (.L_HI(net229));
 sg13g2_tiehi _4640__230 (.L_HI(net230));
 sg13g2_tiehi _4874__231 (.L_HI(net231));
 sg13g2_tiehi _4639__232 (.L_HI(net232));
 sg13g2_tiehi _4803__233 (.L_HI(net233));
 sg13g2_tiehi _4638__234 (.L_HI(net234));
 sg13g2_tiehi _4637__235 (.L_HI(net235));
 sg13g2_tiehi _4636__236 (.L_HI(net236));
 sg13g2_tiehi _4635__237 (.L_HI(net237));
 sg13g2_tiehi _4634__238 (.L_HI(net238));
 sg13g2_tiehi _4633__239 (.L_HI(net239));
 sg13g2_tiehi _4632__240 (.L_HI(net240));
 sg13g2_tiehi _4631__241 (.L_HI(net241));
 sg13g2_tiehi _4630__242 (.L_HI(net242));
 sg13g2_tiehi _4629__243 (.L_HI(net243));
 sg13g2_tiehi _4628__244 (.L_HI(net244));
 sg13g2_tiehi _4627__245 (.L_HI(net245));
 sg13g2_tiehi _4626__246 (.L_HI(net246));
 sg13g2_tiehi _4625__247 (.L_HI(net247));
 sg13g2_tiehi _4624__248 (.L_HI(net248));
 sg13g2_tiehi _4623__249 (.L_HI(net249));
 sg13g2_tiehi _4622__250 (.L_HI(net250));
 sg13g2_tiehi _4621__251 (.L_HI(net251));
 sg13g2_tiehi _4620__252 (.L_HI(net252));
 sg13g2_tiehi _4619__253 (.L_HI(net253));
 sg13g2_tiehi _4618__254 (.L_HI(net254));
 sg13g2_tiehi _4617__255 (.L_HI(net255));
 sg13g2_tiehi _4915__256 (.L_HI(net256));
 sg13g2_tiehi _4616__257 (.L_HI(net257));
 sg13g2_tiehi _4802__258 (.L_HI(net258));
 sg13g2_tiehi _4873__259 (.L_HI(net259));
 sg13g2_tiehi _4801__260 (.L_HI(net260));
 sg13g2_tiehi _4898__261 (.L_HI(net261));
 sg13g2_tiehi _4800__262 (.L_HI(net262));
 sg13g2_tiehi _4872__263 (.L_HI(net263));
 sg13g2_tiehi _4799__264 (.L_HI(net264));
 sg13g2_tiehi _4909__265 (.L_HI(net265));
 sg13g2_tiehi _4798__266 (.L_HI(net266));
 sg13g2_tiehi _4797__267 (.L_HI(net267));
 sg13g2_tiehi _4796__268 (.L_HI(net268));
 sg13g2_tiehi _4871__269 (.L_HI(net269));
 sg13g2_tiehi _4795__270 (.L_HI(net270));
 sg13g2_tiehi _4897__271 (.L_HI(net271));
 sg13g2_tiehi _4794__272 (.L_HI(net272));
 sg13g2_tiehi _4870__273 (.L_HI(net273));
 sg13g2_tiehi _4793__274 (.L_HI(net274));
 sg13g2_tiehi _4792__275 (.L_HI(net275));
 sg13g2_tiehi _4791__276 (.L_HI(net276));
 sg13g2_tiehi _4790__277 (.L_HI(net277));
 sg13g2_tiehi _4919__278 (.L_HI(net278));
 sg13g2_tiehi _4789__279 (.L_HI(net279));
 sg13g2_tiehi _4869__280 (.L_HI(net280));
 sg13g2_tiehi _4788__281 (.L_HI(net281));
 sg13g2_tiehi _4896__282 (.L_HI(net282));
 sg13g2_tiehi _4787__283 (.L_HI(net283));
 sg13g2_tiehi _4868__284 (.L_HI(net284));
 sg13g2_tiehi _4786__285 (.L_HI(net285));
 sg13g2_tiehi _4908__286 (.L_HI(net286));
 sg13g2_tiehi _4785__287 (.L_HI(net287));
 sg13g2_tiehi _4867__288 (.L_HI(net288));
 sg13g2_tiehi _4784__289 (.L_HI(net289));
 sg13g2_tiehi _4783__290 (.L_HI(net290));
 sg13g2_tiehi _4782__291 (.L_HI(net291));
 sg13g2_tiehi _4895__292 (.L_HI(net292));
 sg13g2_tiehi _4781__293 (.L_HI(net293));
 sg13g2_tiehi _4866__294 (.L_HI(net294));
 sg13g2_tiehi _4780__295 (.L_HI(net295));
 sg13g2_tiehi _4914__296 (.L_HI(net296));
 sg13g2_tiehi _4779__297 (.L_HI(net297));
 sg13g2_tiehi _4865__298 (.L_HI(net298));
 sg13g2_tiehi _4778__299 (.L_HI(net299));
 sg13g2_tiehi _4864__300 (.L_HI(net300));
 sg13g2_tiehi _4777__301 (.L_HI(net301));
 sg13g2_tiehi _4863__302 (.L_HI(net302));
 sg13g2_tiehi _4776__303 (.L_HI(net303));
 sg13g2_tiehi _4862__304 (.L_HI(net304));
 sg13g2_tiehi _4775__305 (.L_HI(net305));
 sg13g2_tiehi _4861__306 (.L_HI(net306));
 sg13g2_tiehi _4774__307 (.L_HI(net307));
 sg13g2_tiehi _4860__308 (.L_HI(net308));
 sg13g2_tiehi _4773__309 (.L_HI(net309));
 sg13g2_tiehi _4859__310 (.L_HI(net310));
 sg13g2_tiehi _4772__311 (.L_HI(net311));
 sg13g2_tiehi _4858__312 (.L_HI(net312));
 sg13g2_tiehi tt_um_htfab_caterpillar_313 (.L_HI(net313));
 sg13g2_tiehi tt_um_htfab_caterpillar_314 (.L_HI(net314));
 sg13g2_tiehi tt_um_htfab_caterpillar_315 (.L_HI(net315));
 sg13g2_tiehi tt_um_htfab_caterpillar_316 (.L_HI(net316));
 sg13g2_tiehi tt_um_htfab_caterpillar_317 (.L_HI(net317));
 sg13g2_tiehi tt_um_htfab_caterpillar_318 (.L_HI(net318));
 sg13g2_tiehi tt_um_htfab_caterpillar_319 (.L_HI(net319));
 sg13g2_tiehi tt_um_htfab_caterpillar_320 (.L_HI(net320));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_htfab_caterpillar_7 (.L_LO(net7));
 sg13g2_tiehi _4771__8 (.L_HI(net8));
 sg13g2_buf_1 _5235_ (.A(\snd.sound ),
    .X(uo_out[4]));
 sg13g2_buf_2 fanout333 (.A(_0937_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_0904_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_0783_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net337),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_0783_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_1027_),
    .X(net338));
 sg13g2_buf_1 fanout339 (.A(_1027_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_1132_),
    .X(net340));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_0814_));
 sg13g2_buf_2 fanout342 (.A(_1212_),
    .X(net342));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(_0796_));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_0794_));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(_0745_));
 sg13g2_buf_2 fanout346 (.A(_0617_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_0706_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_0705_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_0704_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_0594_),
    .X(net351));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net353));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(_0519_));
 sg13g2_buf_8 fanout354 (.A(_0509_),
    .X(net354));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(net358));
 sg13g2_buf_2 fanout356 (.A(net358),
    .X(net356));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(net358));
 sg13g2_buf_2 fanout358 (.A(_0701_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(net361),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(net365),
    .X(net361));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net364));
 sg13g2_buf_2 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(net365));
 sg13g2_buf_2 fanout365 (.A(_0700_),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(net368));
 sg13g2_buf_2 fanout367 (.A(net368),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_0700_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_0625_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_0624_),
    .X(net370));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(_0595_));
 sg13g2_buf_2 fanout372 (.A(_0618_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_1911_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_1 fanout376 (.A(net378),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(net378),
    .X(net377));
 sg13g2_buf_1 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(_1781_));
 sg13g2_buf_2 fanout380 (.A(net772),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(net382),
    .X(net381));
 sg13g2_buf_1 fanout382 (.A(\game.state[1] ),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(net708),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(net708),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(\display_value[3] ),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(display_graphical),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(\game.solver_active ),
    .X(net389));
 sg13g2_buf_4 fanout390 (.X(net390),
    .A(\game.current_level[2] ));
 sg13g2_buf_4 fanout391 (.X(net391),
    .A(net791));
 sg13g2_buf_4 fanout392 (.X(net392),
    .A(\game.current_level[0] ));
 sg13g2_buf_2 fanout393 (.A(\game.challenge_num[0] ),
    .X(net393));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(\game.fsm.num_blocks[0] ));
 sg13g2_buf_2 fanout395 (.A(\game.fsm.num_blocks[0] ),
    .X(net395));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(net792));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(\game.fsm.length[1] ));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(net400));
 sg13g2_buf_2 fanout399 (.A(net400),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(net401),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(\game.fsm.length[0] ),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(\game.slv.state[2] ),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(net794),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net408),
    .X(net405));
 sg13g2_buf_1 fanout406 (.A(net408),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_4 fanout408 (.X(net408),
    .A(\btn.gate_200hz ));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(net777));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(net771));
 sg13g2_buf_2 fanout411 (.A(net414),
    .X(net411));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(net414));
 sg13g2_buf_2 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_1880_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(net417),
    .X(net415));
 sg13g2_buf_1 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(net418),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_1880_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(_1880_));
 sg13g2_buf_2 fanout421 (.A(net428),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(net425),
    .X(net422));
 sg13g2_buf_1 fanout423 (.A(net425),
    .X(net423));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(net425));
 sg13g2_buf_2 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(net428),
    .X(net426));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(net428));
 sg13g2_buf_4 fanout428 (.X(net428),
    .A(rst_n));
 sg13g2_buf_4 fanout429 (.X(net429),
    .A(net432));
 sg13g2_buf_2 fanout430 (.A(net431),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(rst_n),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(net439),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(net439),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(net436),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(net439),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(net439),
    .X(net437));
 sg13g2_buf_1 fanout438 (.A(net439),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(rst_n),
    .X(net439));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(net5));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_tielo tt_um_htfab_caterpillar_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_41_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_43_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_2_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_3_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_38_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_33_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_36_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_37_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_8_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_10_clk));
 sg13g2_inv_8 clkload18 (.A(clknet_leaf_16_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_19_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\game.slv.lfsr[9] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0021_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0087_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold4 (.A(\game.slv.lfsr[5] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold5 (.A(\game.slv.lfsr[10] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0090_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0197_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0089_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0200_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0091_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0194_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold12 (.A(\btn.current_event[2] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold13 (.A(\btn.current_event[3] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0088_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0202_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold16 (.A(\game.slv.lfsr[13] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold17 (.A(\game.slv.lfsr[4] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold18 (.A(\game.slv.lfsr[14] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold19 (.A(\game.slv.lfsr[11] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold20 (.A(\game.slv.lfsr[15] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold21 (.A(\game.slv.lfsr[3] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold22 (.A(\game.slv.lfsr[8] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold23 (.A(\game.slv.lfsr[12] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold24 (.A(\btn.long_press ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold25 (.A(\game.slv.lfsr[6] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold26 (.A(\btn.current_event[0] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0019_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0326_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold29 (.A(\btn.current_event[1] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold30 (.A(\game.slv.lfsr[16] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold31 (.A(\game.fsm.block_len[1][0] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold32 (.A(\clk_div_counter[2] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold33 (.A(_1377_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0286_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold35 (.A(\game.challenge_mode ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0211_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold37 (.A(\game.solver_trigger_delayed ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold38 (.A(\game.slv.lfsr[17] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold39 (.A(\game.slv.lfsr[7] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold40 (.A(\game.fsm.block_len[5][2] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold41 (.A(\game.tune[1] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold42 (.A(\snd.note_timing[0] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0120_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold44 (.A(\game.fsm.block_len[7][1] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold45 (.A(\btn.sample_5ms[0] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold46 (.A(\btn.sample_15ms[3] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold47 (.A(\game.fsm.block_len[7][2] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold48 (.A(\snd.next_note_sel[0] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold49 (.A(\btn.button_state[1] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold50 (.A(_1406_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold51 (.A(\game.tune[0] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold52 (.A(\game.fsm.len1_color_count[3][2] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold53 (.A(\game.slv.state[3] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0177_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold55 (.A(\game.fsm.block_len[3][0] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold56 (.A(\game.slv.saved_target ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0928_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0167_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold59 (.A(\game.fsm.block_len[0][0] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold60 (.A(\snd.next_note_timing[5] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold61 (.A(\game.slv.lfsr[1] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold62 (.A(\btn.sample_10ms[0] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0305_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold64 (.A(\snd.next_note_timing[4] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold65 (.A(\game.fsm.green_block_count[0] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold66 (.A(\clk_div_counter[3] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold67 (.A(_1379_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold68 (.A(\game.challenge_num[0] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold69 (.A(\btn.button_state[0] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold70 (.A(\game.input_color[0] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0225_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold72 (.A(\btn.sample_10ms[3] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0312_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold74 (.A(\game.fsm.block_len[3][1] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold75 (.A(\game.fsm.block_len[7][0] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold76 (.A(\snd.next_note_timing[1] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold77 (.A(\game.fsm.len3_color_count[2][1] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold78 (.A(\game.fsm.len1_color_count[1][2] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold79 (.A(\game.fsm.len2_color_count[0][0] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold80 (.A(\snd.next_note_timing[0] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold81 (.A(\snd.next_note_timing[3] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold82 (.A(\snd.note_sel[0] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold83 (.A(\game.fsm.len1_color_count[3][1] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold84 (.A(\game.fsm.seq[0][0] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold85 (.A(\game.fsm.len3_color_count[0][1] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold86 (.A(\btn.change_timer[1] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold87 (.A(_1420_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold88 (.A(\game.fsm.block_len[0][1] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold89 (.A(\snd.tune_counter[5] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold90 (.A(_1738_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold91 (.A(\snd.next_note_timing[8] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold92 (.A(\btn.sample_10ms[2] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0307_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold94 (.A(\game.fsm.len2_color_count[1][0] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0022_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold96 (.A(_1139_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0216_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold98 (.A(\btn.sample_5ms[2] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold99 (.A(\btn.sample_5ms[1] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0310_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold101 (.A(\game.fsm.block_len[2][2] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold102 (.A(\clk_div_counter[6] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold103 (.A(_1384_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold104 (.A(\snd.note_timing[1] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold105 (.A(\game.fsm.len2_color_count[2][0] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold106 (.A(\clk_div_counter[4] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold107 (.A(\game.fsm.len1_color_count[2][2] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold108 (.A(\game.counter[7] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold109 (.A(_1368_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold110 (.A(\snd.next_note_timing[7] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold111 (.A(\game.fsm.len3_color_count[3][0] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold112 (.A(\game.fsm.green_block_count[1] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold113 (.A(_1071_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold114 (.A(\btn.sample_10ms[1] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0306_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold116 (.A(\clk_div_counter[5] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold117 (.A(\game.fsm.len3_color_count[3][1] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold118 (.A(\game.counter[5] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold119 (.A(_1363_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold120 (.A(\game.fsm.len1_color_count[0][2] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold121 (.A(\snd.tune_counter[6] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0374_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold123 (.A(\snd.note_timing[3] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold124 (.A(\game.challenge_num[3] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold125 (.A(\game.next_state[2] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold126 (.A(\snd.next_note_timing[2] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0122_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold128 (.A(\game.fsm.block_len[0][2] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold129 (.A(\btn.button_state[2] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold130 (.A(\game.fsm.block_len[3][2] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold131 (.A(\game.slv.target[0] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold132 (.A(\game.fsm.block_len[2][1] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold133 (.A(\game.fsm.read_pos[0] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold134 (.A(_1176_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold135 (.A(\game.fsm.len1_color_count[0][0] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold136 (.A(\snd.next_note_sel[1] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0117_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold138 (.A(\game.fsm.block_len[5][1] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0061_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold140 (.A(\snd.sound ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold141 (.A(_1554_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0345_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold143 (.A(\game.fsm.len2_color_count[3][0] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold144 (.A(\game.fsm.block_len[2][0] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold145 (.A(\snd.tune_counter[1] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold146 (.A(_1725_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold147 (.A(\snd.note_timing[7] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold148 (.A(\btn.change_timer[5] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0303_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold150 (.A(\game.fsm.length[1] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold151 (.A(_1025_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold152 (.A(\snd.note_timing[5] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold153 (.A(\snd.chord[3][0] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0152_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold155 (.A(\snd.note_timing[8] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold156 (.A(\game.fsm.seq[7][1] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold157 (.A(\game.fsm.block_len[6][0] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold158 (.A(\game.state[1] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold159 (.A(\game.fsm.len3_color_count[1][1] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold160 (.A(\game.fsm.block_len[5][0] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold161 (.A(\game.next_state[0] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold162 (.A(\game.fsm.seq[7][0] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold163 (.A(\snd.counter[2] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0907_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0154_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold166 (.A(\game.fsm.block_len[1][1] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold167 (.A(\game.sound_mode[2] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold168 (.A(\btn.change_timer[2] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold169 (.A(_1443_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold170 (.A(\game.fsm.len1_color_count[1][1] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold171 (.A(\game.fsm.len2_color_count[0][1] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold172 (.A(\game.fsm.len1_color_count[3][0] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold173 (.A(\game.fsm.len3_color_count[0][0] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold174 (.A(\snd.counter[6] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0915_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold176 (.A(\clk_div_counter[7] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold177 (.A(\game.slv.lfsr[20] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0769_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0097_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold180 (.A(\game.fsm.block_len[4][0] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold181 (.A(\snd.note_timing[6] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0126_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold183 (.A(\game.counter[6] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold184 (.A(\game.input_color[1] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0226_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold186 (.A(\game.fsm.len2_color_count[3][1] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold187 (.A(\game.fsm.len1_color_count[2][1] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0092_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0191_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold190 (.A(\game.slv.length[2] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0170_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold192 (.A(\clk_div_counter[1] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold193 (.A(_1375_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold194 (.A(\game.fsm.block_len[4][2] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold195 (.A(\game.fsm.len2_color_count[1][1] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold196 (.A(\game.fsm.block_len[6][2] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold197 (.A(\snd.tune_counter[2] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold198 (.A(_1730_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold199 (.A(\game.slv.lfsr[18] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold200 (.A(\game.fsm.len3_block_count[1] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold201 (.A(\game.fsm.len1_color_count[0][1] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold202 (.A(\btn.sample_5ms[3] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0316_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold204 (.A(\game.fsm.seq[5][0] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold205 (.A(\game.fsm.len2_color_count[2][1] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold206 (.A(\btn.change_timer[6] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold207 (.A(\snd.chord[0][0] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold208 (.A(\game.fsm.block_len[4][1] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold209 (.A(\snd.tune_counter[0] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold210 (.A(\btn.change_timer[3] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold211 (.A(_1446_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold212 (.A(\game.fsm.seq[5][1] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold213 (.A(\game.fsm.block_len[1][2] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold214 (.A(\game.counter[4] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold215 (.A(_1362_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold216 (.A(\game.fsm.seq[1][0] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold217 (.A(\snd.counter[4] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0911_),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold219 (.A(\snd.counter[1] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0905_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold221 (.A(\snd.next_note_timing[6] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold222 (.A(\snd.note_timing[4] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold223 (.A(\snd.counter[0] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold224 (.A(\game.slv.length[1] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold225 (.A(\snd.counter[5] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold226 (.A(\game.fsm.green_block_count[2] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold227 (.A(_1075_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold228 (.A(\game.slv.retries[1] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0175_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold230 (.A(\snd.counter[3] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold231 (.A(\game.slv.target[1] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold232 (.A(\snd.tune_counter[3] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold233 (.A(\game.fsm.seq[6][0] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold234 (.A(\game.slv.retries[0] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0174_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold236 (.A(\snd.chord[0][5] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold237 (.A(\game.sound_on ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0292_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold239 (.A(\game.fsm.len1_color_count[1][0] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold240 (.A(\game.fsm.len3_color_count[1][0] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold241 (.A(\snd.chord[0][1] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold242 (.A(\game.sound_mode[0] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0231_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0056_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0171_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold246 (.A(\game.fsm.len1_block_count[2] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold247 (.A(\snd.chord[0][3] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0365_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold249 (.A(\game.fsm.block_len[6][1] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold250 (.A(\game.fsm.read_pos[2] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0223_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold252 (.A(\game.slv.pos[2] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0173_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold254 (.A(\game.slv.state[1] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0010_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold256 (.A(\game.sound_mode[1] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold257 (.A(\game.fsm.len1_color_count[2][0] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold258 (.A(\btn.change_timer[5] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold259 (.A(_1439_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold260 (.A(\snd.tune_pos[2] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold261 (.A(_1752_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold262 (.A(\snd.counter[8] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0918_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold264 (.A(\btn.change_timer[0] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold265 (.A(\snd.chord[2][2] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0357_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold267 (.A(\game.fsm.len2_block_count[1] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold268 (.A(\clk_div_counter[0] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold269 (.A(\btn.change_timer[4] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0302_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold271 (.A(\game.fsm.seq[3][0] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold272 (.A(\snd.tune_pos[1] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold273 (.A(\snd.sequencer_state[1] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0381_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold275 (.A(\snd.counter[7] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold276 (.A(\game.challenge_num[2] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold277 (.A(\game.counter[3] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold278 (.A(\game.fsm.len3_color_count[2][0] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold279 (.A(\snd.chord[0][2] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold280 (.A(\game.state[0] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold281 (.A(\game.slv.lfsr[19] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold282 (.A(uo_out[2]),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold283 (.A(\game.fsm.seq[0][1] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold284 (.A(\btn.button_state[3] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold285 (.A(\game.slv.length[0] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0168_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold287 (.A(\snd.tune_pos[0] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold288 (.A(\game.slv.lfsr[2] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold289 (.A(\game.fsm.seq[4][0] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold290 (.A(\snd.tune_counter[4] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold291 (.A(_1737_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold292 (.A(\game.slv.trigger ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold293 (.A(\btn.sample_5ms[2] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold294 (.A(\game.fsm.read_pos[1] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold295 (.A(\game.fsm.color_count[3][2] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold296 (.A(\snd.chord[1][5] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0359_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold298 (.A(\game.slv.pos[1] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0172_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold300 (.A(\game.fsm.color_count[2][1] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold301 (.A(\game.counter[2] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold302 (.A(_1359_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold303 (.A(\game.fsm.color_count[2][2] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold304 (.A(display_graphical),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold305 (.A(_1234_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold306 (.A(uo_out[3]),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold307 (.A(\game.slv.retries[2] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0176_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold309 (.A(\game.counter[1] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold310 (.A(_1356_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0271_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold312 (.A(\game.fsm.seq[3][1] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold313 (.A(\game.fsm.color_count[1][1] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold314 (.A(\snd.active_tune[1] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold315 (.A(\game.fsm.seq[6][1] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold316 (.A(\game.fsm.seq[4][1] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold317 (.A(\game.fsm.seq[2][0] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold318 (.A(\game.fsm.len1_block_count[1] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold319 (.A(\game.fsm.seq[1][1] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold320 (.A(\display_value[2] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0016_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold322 (.A(_1507_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0039_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0925_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold325 (.A(\game.fsm.color_count[1][2] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold326 (.A(uo_out[1]),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold327 (.A(\game.counter[0] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold328 (.A(\game.slv.lfsr[0] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold329 (.A(\snd.chord[0][4] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold330 (.A(\snd.active_tune[1] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold331 (.A(\game.fsm.color_count[2][0] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0060_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0322_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0017_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0324_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold336 (.A(\game.fsm.color_count[1][0] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold337 (.A(\game.challenge_num[1] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold338 (.A(\game.current_level[4] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold339 (.A(\game.next_state[2] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0020_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold341 (.A(_1524_),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0014_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold343 (.A(\game.fsm.color_count[0][0] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold344 (.A(\snd.active_tune[0] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0085_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold346 (.A(_1151_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0219_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold348 (.A(\game.fsm.seq[2][1] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold349 (.A(\game.fsm.color_count[0][1] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold350 (.A(\game.slv.ready ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold351 (.A(\game.fsm.num_blocks[2] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0018_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold353 (.A(\dsp.digit ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold354 (.A(\game.state[3] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold355 (.A(uo_out[0]),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold356 (.A(\game.fsm.num_blocks[1] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold357 (.A(\snd.chord[1][0] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold358 (.A(\game.fsm.color_count[3][0] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0084_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold360 (.A(_1146_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0218_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold362 (.A(\snd.sequencer_state[0] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold363 (.A(\game.current_level[1] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold364 (.A(\game.fsm.length[2] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold365 (.A(\game.sound_on ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold366 (.A(\game.fsm.color_count[3][1] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold367 (.A(\game.fsm.color_count[0][2] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold368 (.A(\game.slv.length[0] ),
    .X(net796));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_fill_1 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_46 ();
 sg13g2_fill_2 FILLER_0_53 ();
 sg13g2_fill_1 FILLER_0_55 ();
 sg13g2_decap_4 FILLER_0_82 ();
 sg13g2_fill_2 FILLER_0_86 ();
 sg13g2_decap_8 FILLER_0_92 ();
 sg13g2_decap_8 FILLER_0_99 ();
 sg13g2_decap_4 FILLER_0_106 ();
 sg13g2_fill_2 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_116 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_decap_4 FILLER_0_130 ();
 sg13g2_fill_1 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_142 ();
 sg13g2_decap_4 FILLER_0_149 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_4 FILLER_0_164 ();
 sg13g2_fill_1 FILLER_0_168 ();
 sg13g2_decap_4 FILLER_0_174 ();
 sg13g2_fill_1 FILLER_0_178 ();
 sg13g2_fill_2 FILLER_0_184 ();
 sg13g2_fill_1 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_191 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_219 ();
 sg13g2_decap_8 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_240 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_4 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_25 ();
 sg13g2_decap_4 FILLER_1_53 ();
 sg13g2_fill_1 FILLER_1_66 ();
 sg13g2_fill_1 FILLER_1_71 ();
 sg13g2_fill_2 FILLER_1_101 ();
 sg13g2_fill_2 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_227 ();
 sg13g2_decap_8 FILLER_1_234 ();
 sg13g2_decap_8 FILLER_1_241 ();
 sg13g2_decap_8 FILLER_1_248 ();
 sg13g2_decap_8 FILLER_1_255 ();
 sg13g2_decap_8 FILLER_1_262 ();
 sg13g2_decap_8 FILLER_1_269 ();
 sg13g2_decap_8 FILLER_1_276 ();
 sg13g2_decap_8 FILLER_1_283 ();
 sg13g2_decap_8 FILLER_1_290 ();
 sg13g2_decap_8 FILLER_1_297 ();
 sg13g2_decap_8 FILLER_1_304 ();
 sg13g2_decap_8 FILLER_1_311 ();
 sg13g2_decap_8 FILLER_1_318 ();
 sg13g2_decap_8 FILLER_1_325 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_4 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_35 ();
 sg13g2_fill_2 FILLER_2_72 ();
 sg13g2_fill_1 FILLER_2_74 ();
 sg13g2_fill_1 FILLER_2_98 ();
 sg13g2_fill_2 FILLER_2_108 ();
 sg13g2_fill_1 FILLER_2_110 ();
 sg13g2_fill_2 FILLER_2_199 ();
 sg13g2_decap_8 FILLER_2_227 ();
 sg13g2_decap_8 FILLER_2_234 ();
 sg13g2_decap_8 FILLER_2_241 ();
 sg13g2_decap_8 FILLER_2_248 ();
 sg13g2_decap_8 FILLER_2_255 ();
 sg13g2_decap_8 FILLER_2_262 ();
 sg13g2_decap_8 FILLER_2_269 ();
 sg13g2_decap_8 FILLER_2_276 ();
 sg13g2_decap_8 FILLER_2_283 ();
 sg13g2_decap_8 FILLER_2_290 ();
 sg13g2_decap_8 FILLER_2_297 ();
 sg13g2_decap_8 FILLER_2_304 ();
 sg13g2_decap_8 FILLER_2_311 ();
 sg13g2_decap_8 FILLER_2_318 ();
 sg13g2_decap_8 FILLER_2_325 ();
 sg13g2_decap_8 FILLER_2_332 ();
 sg13g2_decap_8 FILLER_2_339 ();
 sg13g2_decap_8 FILLER_2_346 ();
 sg13g2_decap_8 FILLER_2_353 ();
 sg13g2_decap_8 FILLER_2_360 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_21 ();
 sg13g2_fill_1 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_233 ();
 sg13g2_decap_8 FILLER_3_240 ();
 sg13g2_decap_8 FILLER_3_247 ();
 sg13g2_decap_8 FILLER_3_254 ();
 sg13g2_decap_8 FILLER_3_261 ();
 sg13g2_decap_8 FILLER_3_268 ();
 sg13g2_decap_8 FILLER_3_275 ();
 sg13g2_decap_8 FILLER_3_282 ();
 sg13g2_decap_8 FILLER_3_289 ();
 sg13g2_decap_8 FILLER_3_296 ();
 sg13g2_decap_8 FILLER_3_303 ();
 sg13g2_decap_8 FILLER_3_310 ();
 sg13g2_decap_8 FILLER_3_317 ();
 sg13g2_decap_8 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_331 ();
 sg13g2_decap_8 FILLER_3_338 ();
 sg13g2_decap_8 FILLER_3_345 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_28 ();
 sg13g2_fill_2 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_37 ();
 sg13g2_fill_2 FILLER_4_46 ();
 sg13g2_fill_1 FILLER_4_48 ();
 sg13g2_fill_1 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_86 ();
 sg13g2_fill_2 FILLER_4_132 ();
 sg13g2_fill_1 FILLER_4_134 ();
 sg13g2_decap_4 FILLER_4_180 ();
 sg13g2_fill_1 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_decap_8 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_240 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_decap_8 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_2 FILLER_5_53 ();
 sg13g2_fill_1 FILLER_5_55 ();
 sg13g2_fill_2 FILLER_5_61 ();
 sg13g2_fill_1 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_103 ();
 sg13g2_fill_2 FILLER_5_110 ();
 sg13g2_fill_1 FILLER_5_112 ();
 sg13g2_fill_2 FILLER_5_127 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_fill_1 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_148 ();
 sg13g2_fill_1 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_288 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_59 ();
 sg13g2_fill_1 FILLER_6_61 ();
 sg13g2_fill_1 FILLER_6_75 ();
 sg13g2_fill_1 FILLER_6_103 ();
 sg13g2_decap_8 FILLER_6_114 ();
 sg13g2_decap_4 FILLER_6_121 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_2 FILLER_6_198 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_decap_8 FILLER_6_261 ();
 sg13g2_decap_8 FILLER_6_268 ();
 sg13g2_decap_8 FILLER_6_275 ();
 sg13g2_decap_8 FILLER_6_282 ();
 sg13g2_decap_8 FILLER_6_289 ();
 sg13g2_decap_8 FILLER_6_296 ();
 sg13g2_decap_8 FILLER_6_303 ();
 sg13g2_decap_8 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_317 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_fill_1 FILLER_7_15 ();
 sg13g2_decap_4 FILLER_7_46 ();
 sg13g2_decap_4 FILLER_7_64 ();
 sg13g2_fill_1 FILLER_7_72 ();
 sg13g2_fill_2 FILLER_7_81 ();
 sg13g2_fill_1 FILLER_7_83 ();
 sg13g2_fill_1 FILLER_7_91 ();
 sg13g2_fill_2 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_151 ();
 sg13g2_fill_2 FILLER_7_158 ();
 sg13g2_fill_1 FILLER_7_160 ();
 sg13g2_fill_1 FILLER_7_174 ();
 sg13g2_fill_1 FILLER_7_186 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_255 ();
 sg13g2_decap_8 FILLER_7_262 ();
 sg13g2_decap_8 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_276 ();
 sg13g2_decap_8 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_decap_4 FILLER_8_175 ();
 sg13g2_fill_2 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_209 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_decap_8 FILLER_8_257 ();
 sg13g2_decap_8 FILLER_8_264 ();
 sg13g2_decap_8 FILLER_8_271 ();
 sg13g2_decap_8 FILLER_8_278 ();
 sg13g2_decap_8 FILLER_8_285 ();
 sg13g2_decap_8 FILLER_8_292 ();
 sg13g2_decap_8 FILLER_8_299 ();
 sg13g2_decap_8 FILLER_8_306 ();
 sg13g2_decap_8 FILLER_8_313 ();
 sg13g2_decap_8 FILLER_8_320 ();
 sg13g2_decap_8 FILLER_8_327 ();
 sg13g2_decap_8 FILLER_8_334 ();
 sg13g2_decap_8 FILLER_8_341 ();
 sg13g2_decap_8 FILLER_8_348 ();
 sg13g2_decap_8 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_362 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_114 ();
 sg13g2_fill_2 FILLER_9_153 ();
 sg13g2_fill_2 FILLER_9_159 ();
 sg13g2_decap_4 FILLER_9_173 ();
 sg13g2_fill_1 FILLER_9_177 ();
 sg13g2_decap_8 FILLER_9_187 ();
 sg13g2_fill_2 FILLER_9_194 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_fill_1 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_250 ();
 sg13g2_decap_8 FILLER_9_257 ();
 sg13g2_decap_8 FILLER_9_264 ();
 sg13g2_decap_8 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_278 ();
 sg13g2_decap_8 FILLER_9_285 ();
 sg13g2_decap_8 FILLER_9_292 ();
 sg13g2_decap_8 FILLER_9_299 ();
 sg13g2_decap_8 FILLER_9_306 ();
 sg13g2_decap_8 FILLER_9_313 ();
 sg13g2_decap_8 FILLER_9_320 ();
 sg13g2_decap_8 FILLER_9_327 ();
 sg13g2_decap_8 FILLER_9_334 ();
 sg13g2_decap_8 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_348 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_2 FILLER_10_30 ();
 sg13g2_decap_8 FILLER_10_106 ();
 sg13g2_decap_8 FILLER_10_113 ();
 sg13g2_decap_8 FILLER_10_120 ();
 sg13g2_fill_2 FILLER_10_130 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_decap_8 FILLER_10_164 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_fill_1 FILLER_10_173 ();
 sg13g2_fill_2 FILLER_10_210 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_219 ();
 sg13g2_decap_8 FILLER_10_226 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_decap_8 FILLER_10_247 ();
 sg13g2_decap_8 FILLER_10_254 ();
 sg13g2_decap_8 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_268 ();
 sg13g2_decap_8 FILLER_10_275 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_25 ();
 sg13g2_decap_8 FILLER_11_37 ();
 sg13g2_decap_8 FILLER_11_47 ();
 sg13g2_fill_1 FILLER_11_54 ();
 sg13g2_decap_8 FILLER_11_78 ();
 sg13g2_fill_1 FILLER_11_85 ();
 sg13g2_fill_1 FILLER_11_94 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_decap_4 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_251 ();
 sg13g2_decap_8 FILLER_11_258 ();
 sg13g2_decap_8 FILLER_11_265 ();
 sg13g2_decap_8 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_279 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_decap_8 FILLER_11_293 ();
 sg13g2_decap_8 FILLER_11_300 ();
 sg13g2_decap_8 FILLER_11_307 ();
 sg13g2_decap_4 FILLER_11_314 ();
 sg13g2_fill_2 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_335 ();
 sg13g2_decap_8 FILLER_11_342 ();
 sg13g2_decap_8 FILLER_11_349 ();
 sg13g2_decap_8 FILLER_11_356 ();
 sg13g2_decap_8 FILLER_11_363 ();
 sg13g2_decap_8 FILLER_11_370 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_decap_4 FILLER_12_31 ();
 sg13g2_decap_8 FILLER_12_54 ();
 sg13g2_decap_8 FILLER_12_61 ();
 sg13g2_fill_2 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_76 ();
 sg13g2_fill_1 FILLER_12_78 ();
 sg13g2_fill_2 FILLER_12_104 ();
 sg13g2_fill_1 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_125 ();
 sg13g2_fill_2 FILLER_12_134 ();
 sg13g2_fill_1 FILLER_12_142 ();
 sg13g2_decap_4 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_308 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_fill_2 FILLER_12_325 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_39 ();
 sg13g2_decap_4 FILLER_13_48 ();
 sg13g2_fill_1 FILLER_13_52 ();
 sg13g2_fill_2 FILLER_13_70 ();
 sg13g2_fill_2 FILLER_13_77 ();
 sg13g2_fill_1 FILLER_13_79 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_fill_1 FILLER_13_141 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_decap_4 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_fill_1 FILLER_13_179 ();
 sg13g2_fill_2 FILLER_13_189 ();
 sg13g2_fill_2 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_212 ();
 sg13g2_decap_4 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_255 ();
 sg13g2_decap_8 FILLER_13_262 ();
 sg13g2_decap_8 FILLER_13_269 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_decap_8 FILLER_13_282 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_1 FILLER_14_40 ();
 sg13g2_fill_1 FILLER_14_54 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_fill_2 FILLER_14_95 ();
 sg13g2_fill_1 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_102 ();
 sg13g2_fill_1 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_164 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_4 FILLER_14_202 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_decap_4 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_239 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_1 FILLER_15_12 ();
 sg13g2_fill_2 FILLER_15_57 ();
 sg13g2_fill_2 FILLER_15_64 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_decap_8 FILLER_15_83 ();
 sg13g2_decap_8 FILLER_15_90 ();
 sg13g2_decap_8 FILLER_15_97 ();
 sg13g2_decap_8 FILLER_15_104 ();
 sg13g2_fill_2 FILLER_15_111 ();
 sg13g2_fill_1 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_decap_8 FILLER_15_145 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_173 ();
 sg13g2_fill_1 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_180 ();
 sg13g2_fill_2 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_230 ();
 sg13g2_fill_2 FILLER_15_261 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_275 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_fill_2 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_fill_2 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_fill_2 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_58 ();
 sg13g2_decap_8 FILLER_16_78 ();
 sg13g2_decap_8 FILLER_16_85 ();
 sg13g2_decap_8 FILLER_16_107 ();
 sg13g2_decap_8 FILLER_16_114 ();
 sg13g2_decap_4 FILLER_16_142 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_decap_4 FILLER_16_158 ();
 sg13g2_fill_2 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_250 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_fill_1 FILLER_16_318 ();
 sg13g2_fill_2 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_31 ();
 sg13g2_decap_8 FILLER_17_57 ();
 sg13g2_decap_8 FILLER_17_64 ();
 sg13g2_decap_4 FILLER_17_71 ();
 sg13g2_fill_2 FILLER_17_75 ();
 sg13g2_fill_2 FILLER_17_93 ();
 sg13g2_decap_8 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_159 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_fill_1 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_299 ();
 sg13g2_fill_2 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_307 ();
 sg13g2_fill_1 FILLER_17_313 ();
 sg13g2_fill_1 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_fill_1 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_53 ();
 sg13g2_fill_1 FILLER_18_98 ();
 sg13g2_fill_1 FILLER_18_107 ();
 sg13g2_fill_2 FILLER_18_168 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_195 ();
 sg13g2_fill_1 FILLER_18_197 ();
 sg13g2_decap_4 FILLER_18_202 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_fill_1 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_decap_4 FILLER_18_261 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_fill_2 FILLER_19_26 ();
 sg13g2_fill_2 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_decap_8 FILLER_19_107 ();
 sg13g2_decap_4 FILLER_19_114 ();
 sg13g2_decap_4 FILLER_19_159 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_fill_2 FILLER_19_297 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_55 ();
 sg13g2_fill_1 FILLER_20_57 ();
 sg13g2_decap_4 FILLER_20_78 ();
 sg13g2_fill_1 FILLER_20_92 ();
 sg13g2_fill_2 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_104 ();
 sg13g2_decap_8 FILLER_20_111 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_decap_4 FILLER_20_146 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_170 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_decap_8 FILLER_20_198 ();
 sg13g2_decap_4 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_263 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_fill_2 FILLER_21_9 ();
 sg13g2_decap_8 FILLER_21_20 ();
 sg13g2_decap_4 FILLER_21_27 ();
 sg13g2_fill_1 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_57 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_decap_8 FILLER_21_113 ();
 sg13g2_decap_4 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_fill_2 FILLER_21_164 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_179 ();
 sg13g2_decap_4 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_fill_2 FILLER_21_286 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_114 ();
 sg13g2_decap_8 FILLER_22_124 ();
 sg13g2_decap_8 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_138 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_4 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_235 ();
 sg13g2_fill_1 FILLER_22_237 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_259 ();
 sg13g2_fill_1 FILLER_22_261 ();
 sg13g2_fill_2 FILLER_22_299 ();
 sg13g2_fill_2 FILLER_22_309 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_fill_1 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_51 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_fill_2 FILLER_23_73 ();
 sg13g2_fill_1 FILLER_23_80 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_decap_8 FILLER_23_138 ();
 sg13g2_decap_4 FILLER_23_145 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_231 ();
 sg13g2_fill_1 FILLER_23_233 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_1 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_52 ();
 sg13g2_fill_1 FILLER_24_54 ();
 sg13g2_fill_1 FILLER_24_69 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_decap_4 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_decap_4 FILLER_24_129 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_fill_2 FILLER_24_176 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_decap_4 FILLER_24_268 ();
 sg13g2_fill_2 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_36 ();
 sg13g2_decap_8 FILLER_25_69 ();
 sg13g2_fill_2 FILLER_25_76 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_decap_8 FILLER_25_89 ();
 sg13g2_decap_8 FILLER_25_96 ();
 sg13g2_decap_8 FILLER_25_103 ();
 sg13g2_fill_1 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_decap_8 FILLER_25_142 ();
 sg13g2_decap_4 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_fill_1 FILLER_25_232 ();
 sg13g2_decap_4 FILLER_25_273 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_fill_2 FILLER_26_13 ();
 sg13g2_fill_1 FILLER_26_15 ();
 sg13g2_fill_1 FILLER_26_64 ();
 sg13g2_decap_8 FILLER_26_73 ();
 sg13g2_decap_8 FILLER_26_80 ();
 sg13g2_decap_8 FILLER_26_87 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_2 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_fill_2 FILLER_27_26 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_38 ();
 sg13g2_fill_2 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_64 ();
 sg13g2_decap_8 FILLER_27_71 ();
 sg13g2_decap_8 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_85 ();
 sg13g2_fill_2 FILLER_27_138 ();
 sg13g2_decap_4 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_337 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_58 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_fill_2 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_53 ();
 sg13g2_fill_1 FILLER_29_55 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_fill_1 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_decap_4 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_74 ();
 sg13g2_fill_1 FILLER_30_76 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_171 ();
 sg13g2_decap_4 FILLER_30_178 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_194 ();
 sg13g2_decap_4 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_decap_8 FILLER_30_355 ();
 sg13g2_decap_8 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_369 ();
 sg13g2_decap_8 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_18 ();
 sg13g2_fill_2 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_31 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_68 ();
 sg13g2_decap_4 FILLER_31_81 ();
 sg13g2_fill_1 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_114 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_decap_8 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_decap_4 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_178 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_decap_8 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_206 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_4 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_17 ();
 sg13g2_decap_8 FILLER_32_24 ();
 sg13g2_decap_4 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_fill_2 FILLER_32_97 ();
 sg13g2_decap_8 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_131 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_267 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_26 ();
 sg13g2_decap_8 FILLER_33_33 ();
 sg13g2_fill_2 FILLER_33_40 ();
 sg13g2_fill_2 FILLER_33_46 ();
 sg13g2_fill_1 FILLER_33_48 ();
 sg13g2_fill_1 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_120 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_162 ();
 sg13g2_decap_4 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_37 ();
 sg13g2_fill_1 FILLER_34_69 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_fill_2 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_2 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_decap_4 FILLER_34_324 ();
 sg13g2_fill_2 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_4 FILLER_35_44 ();
 sg13g2_decap_4 FILLER_35_76 ();
 sg13g2_fill_2 FILLER_35_80 ();
 sg13g2_fill_2 FILLER_35_85 ();
 sg13g2_decap_4 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_decap_4 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_decap_4 FILLER_35_194 ();
 sg13g2_fill_2 FILLER_35_202 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_18 ();
 sg13g2_fill_1 FILLER_36_20 ();
 sg13g2_decap_4 FILLER_36_49 ();
 sg13g2_fill_1 FILLER_36_53 ();
 sg13g2_decap_4 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_76 ();
 sg13g2_decap_8 FILLER_36_99 ();
 sg13g2_decap_8 FILLER_36_106 ();
 sg13g2_decap_4 FILLER_36_113 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_fill_2 FILLER_36_123 ();
 sg13g2_fill_2 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_4 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_198 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_decap_4 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_330 ();
 sg13g2_decap_8 FILLER_36_356 ();
 sg13g2_decap_8 FILLER_36_363 ();
 sg13g2_decap_8 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_11 ();
 sg13g2_fill_1 FILLER_37_13 ();
 sg13g2_fill_2 FILLER_37_29 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_decap_4 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_171 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_183 ();
 sg13g2_decap_4 FILLER_37_211 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_decap_4 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_236 ();
 sg13g2_fill_1 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_370 ();
 sg13g2_decap_8 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_18 ();
 sg13g2_fill_1 FILLER_38_25 ();
 sg13g2_fill_1 FILLER_38_52 ();
 sg13g2_fill_2 FILLER_38_80 ();
 sg13g2_fill_1 FILLER_38_82 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_fill_1 FILLER_38_187 ();
 sg13g2_fill_1 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_fill_2 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_253 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_1 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_59 ();
 sg13g2_fill_1 FILLER_39_78 ();
 sg13g2_decap_8 FILLER_39_83 ();
 sg13g2_fill_2 FILLER_39_90 ();
 sg13g2_fill_2 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_160 ();
 sg13g2_decap_4 FILLER_39_167 ();
 sg13g2_fill_1 FILLER_39_171 ();
 sg13g2_fill_1 FILLER_39_176 ();
 sg13g2_decap_8 FILLER_39_181 ();
 sg13g2_fill_2 FILLER_39_188 ();
 sg13g2_fill_1 FILLER_39_190 ();
 sg13g2_fill_1 FILLER_39_199 ();
 sg13g2_fill_1 FILLER_39_213 ();
 sg13g2_decap_4 FILLER_39_240 ();
 sg13g2_fill_1 FILLER_39_248 ();
 sg13g2_decap_8 FILLER_39_362 ();
 sg13g2_decap_8 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_39_376 ();
 sg13g2_decap_8 FILLER_39_383 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_fill_1 FILLER_40_38 ();
 sg13g2_decap_8 FILLER_40_65 ();
 sg13g2_decap_8 FILLER_40_72 ();
 sg13g2_decap_8 FILLER_40_79 ();
 sg13g2_fill_2 FILLER_40_86 ();
 sg13g2_fill_2 FILLER_40_100 ();
 sg13g2_decap_8 FILLER_40_110 ();
 sg13g2_decap_8 FILLER_40_117 ();
 sg13g2_decap_8 FILLER_40_124 ();
 sg13g2_fill_1 FILLER_40_131 ();
 sg13g2_fill_1 FILLER_40_136 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_198 ();
 sg13g2_decap_8 FILLER_40_214 ();
 sg13g2_fill_2 FILLER_40_221 ();
 sg13g2_fill_1 FILLER_40_223 ();
 sg13g2_fill_1 FILLER_40_289 ();
 sg13g2_fill_1 FILLER_40_298 ();
 sg13g2_fill_2 FILLER_40_305 ();
 sg13g2_fill_2 FILLER_40_320 ();
 sg13g2_decap_8 FILLER_40_359 ();
 sg13g2_decap_8 FILLER_40_366 ();
 sg13g2_decap_8 FILLER_40_373 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_41_18 ();
 sg13g2_fill_1 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_54 ();
 sg13g2_decap_4 FILLER_41_61 ();
 sg13g2_fill_2 FILLER_41_65 ();
 sg13g2_fill_2 FILLER_41_72 ();
 sg13g2_fill_1 FILLER_41_74 ();
 sg13g2_fill_2 FILLER_41_131 ();
 sg13g2_fill_2 FILLER_41_139 ();
 sg13g2_fill_1 FILLER_41_141 ();
 sg13g2_decap_4 FILLER_41_148 ();
 sg13g2_fill_1 FILLER_41_196 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_decap_4 FILLER_41_300 ();
 sg13g2_fill_2 FILLER_41_304 ();
 sg13g2_decap_4 FILLER_41_311 ();
 sg13g2_fill_1 FILLER_41_315 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_decap_8 FILLER_41_365 ();
 sg13g2_decap_8 FILLER_41_372 ();
 sg13g2_decap_8 FILLER_41_379 ();
 sg13g2_decap_8 FILLER_41_386 ();
 sg13g2_decap_8 FILLER_41_393 ();
 sg13g2_decap_8 FILLER_41_400 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_fill_1 FILLER_42_20 ();
 sg13g2_decap_8 FILLER_42_47 ();
 sg13g2_decap_8 FILLER_42_54 ();
 sg13g2_fill_1 FILLER_42_92 ();
 sg13g2_fill_2 FILLER_42_141 ();
 sg13g2_fill_2 FILLER_42_204 ();
 sg13g2_fill_1 FILLER_42_206 ();
 sg13g2_decap_8 FILLER_42_211 ();
 sg13g2_fill_2 FILLER_42_218 ();
 sg13g2_decap_8 FILLER_42_228 ();
 sg13g2_fill_1 FILLER_42_235 ();
 sg13g2_fill_2 FILLER_42_257 ();
 sg13g2_fill_2 FILLER_42_303 ();
 sg13g2_fill_1 FILLER_42_305 ();
 sg13g2_fill_2 FILLER_42_311 ();
 sg13g2_decap_8 FILLER_42_366 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_4 ();
 sg13g2_fill_2 FILLER_43_35 ();
 sg13g2_decap_4 FILLER_43_47 ();
 sg13g2_fill_2 FILLER_43_55 ();
 sg13g2_fill_2 FILLER_43_60 ();
 sg13g2_fill_1 FILLER_43_62 ();
 sg13g2_fill_1 FILLER_43_76 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_93 ();
 sg13g2_decap_4 FILLER_43_98 ();
 sg13g2_fill_2 FILLER_43_107 ();
 sg13g2_fill_1 FILLER_43_109 ();
 sg13g2_fill_2 FILLER_43_150 ();
 sg13g2_fill_1 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_196 ();
 sg13g2_decap_4 FILLER_43_205 ();
 sg13g2_decap_4 FILLER_43_214 ();
 sg13g2_fill_1 FILLER_43_218 ();
 sg13g2_decap_8 FILLER_43_222 ();
 sg13g2_fill_1 FILLER_43_233 ();
 sg13g2_fill_2 FILLER_43_300 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_340 ();
 sg13g2_decap_8 FILLER_43_372 ();
 sg13g2_decap_8 FILLER_43_379 ();
 sg13g2_decap_8 FILLER_43_386 ();
 sg13g2_decap_8 FILLER_43_393 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_fill_2 FILLER_44_26 ();
 sg13g2_fill_2 FILLER_44_68 ();
 sg13g2_fill_1 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_80 ();
 sg13g2_decap_8 FILLER_44_87 ();
 sg13g2_fill_2 FILLER_44_94 ();
 sg13g2_fill_2 FILLER_44_134 ();
 sg13g2_fill_1 FILLER_44_136 ();
 sg13g2_fill_1 FILLER_44_170 ();
 sg13g2_fill_2 FILLER_44_179 ();
 sg13g2_fill_1 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_189 ();
 sg13g2_fill_2 FILLER_44_204 ();
 sg13g2_fill_1 FILLER_44_206 ();
 sg13g2_fill_1 FILLER_44_218 ();
 sg13g2_fill_2 FILLER_44_240 ();
 sg13g2_fill_1 FILLER_44_242 ();
 sg13g2_fill_2 FILLER_44_248 ();
 sg13g2_fill_2 FILLER_44_257 ();
 sg13g2_fill_1 FILLER_44_259 ();
 sg13g2_fill_1 FILLER_44_299 ();
 sg13g2_fill_2 FILLER_44_307 ();
 sg13g2_fill_1 FILLER_44_309 ();
 sg13g2_fill_1 FILLER_44_323 ();
 sg13g2_fill_2 FILLER_44_347 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_4 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_fill_1 FILLER_45_35 ();
 sg13g2_fill_2 FILLER_45_67 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_4 FILLER_45_116 ();
 sg13g2_decap_4 FILLER_45_158 ();
 sg13g2_fill_2 FILLER_45_202 ();
 sg13g2_fill_2 FILLER_45_210 ();
 sg13g2_fill_1 FILLER_45_212 ();
 sg13g2_fill_1 FILLER_45_225 ();
 sg13g2_fill_2 FILLER_45_248 ();
 sg13g2_fill_2 FILLER_45_255 ();
 sg13g2_decap_4 FILLER_45_309 ();
 sg13g2_fill_1 FILLER_45_313 ();
 sg13g2_decap_8 FILLER_45_318 ();
 sg13g2_fill_1 FILLER_45_325 ();
 sg13g2_decap_8 FILLER_45_367 ();
 sg13g2_decap_8 FILLER_45_374 ();
 sg13g2_decap_8 FILLER_45_381 ();
 sg13g2_decap_8 FILLER_45_388 ();
 sg13g2_decap_8 FILLER_45_395 ();
 sg13g2_decap_8 FILLER_45_402 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_15 ();
 sg13g2_fill_2 FILLER_46_37 ();
 sg13g2_fill_1 FILLER_46_66 ();
 sg13g2_decap_4 FILLER_46_96 ();
 sg13g2_decap_8 FILLER_46_108 ();
 sg13g2_fill_2 FILLER_46_115 ();
 sg13g2_decap_4 FILLER_46_121 ();
 sg13g2_fill_1 FILLER_46_159 ();
 sg13g2_fill_2 FILLER_46_201 ();
 sg13g2_fill_1 FILLER_46_203 ();
 sg13g2_fill_1 FILLER_46_241 ();
 sg13g2_decap_8 FILLER_46_255 ();
 sg13g2_decap_8 FILLER_46_283 ();
 sg13g2_decap_8 FILLER_46_290 ();
 sg13g2_decap_4 FILLER_46_297 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_fill_1 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_363 ();
 sg13g2_decap_8 FILLER_46_370 ();
 sg13g2_decap_8 FILLER_46_377 ();
 sg13g2_decap_8 FILLER_46_384 ();
 sg13g2_decap_8 FILLER_46_391 ();
 sg13g2_decap_8 FILLER_46_398 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_4 ();
 sg13g2_fill_2 FILLER_47_21 ();
 sg13g2_fill_1 FILLER_47_23 ();
 sg13g2_fill_1 FILLER_47_36 ();
 sg13g2_fill_2 FILLER_47_45 ();
 sg13g2_fill_1 FILLER_47_47 ();
 sg13g2_fill_1 FILLER_47_80 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_fill_2 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_157 ();
 sg13g2_decap_4 FILLER_47_193 ();
 sg13g2_fill_1 FILLER_47_214 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_fill_2 FILLER_47_238 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_decap_4 FILLER_47_245 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_decap_8 FILLER_47_260 ();
 sg13g2_decap_8 FILLER_47_267 ();
 sg13g2_decap_8 FILLER_47_274 ();
 sg13g2_fill_1 FILLER_47_281 ();
 sg13g2_fill_1 FILLER_47_290 ();
 sg13g2_fill_2 FILLER_47_324 ();
 sg13g2_fill_1 FILLER_47_333 ();
 sg13g2_fill_2 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_362 ();
 sg13g2_decap_8 FILLER_47_369 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_decap_8 FILLER_47_383 ();
 sg13g2_decap_8 FILLER_47_390 ();
 sg13g2_decap_8 FILLER_47_397 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_57 ();
 sg13g2_fill_2 FILLER_48_72 ();
 sg13g2_fill_1 FILLER_48_74 ();
 sg13g2_decap_8 FILLER_48_90 ();
 sg13g2_fill_2 FILLER_48_101 ();
 sg13g2_fill_1 FILLER_48_103 ();
 sg13g2_decap_4 FILLER_48_109 ();
 sg13g2_fill_2 FILLER_48_113 ();
 sg13g2_fill_2 FILLER_48_137 ();
 sg13g2_fill_1 FILLER_48_171 ();
 sg13g2_fill_2 FILLER_48_177 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_fill_1 FILLER_48_227 ();
 sg13g2_decap_4 FILLER_48_257 ();
 sg13g2_fill_2 FILLER_48_269 ();
 sg13g2_fill_2 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_299 ();
 sg13g2_fill_1 FILLER_48_317 ();
 sg13g2_decap_8 FILLER_48_349 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_decap_8 FILLER_48_370 ();
 sg13g2_decap_8 FILLER_48_377 ();
 sg13g2_decap_8 FILLER_48_384 ();
 sg13g2_decap_8 FILLER_48_391 ();
 sg13g2_decap_8 FILLER_48_398 ();
 sg13g2_decap_4 FILLER_48_405 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_39 ();
 sg13g2_fill_1 FILLER_49_43 ();
 sg13g2_fill_2 FILLER_49_69 ();
 sg13g2_fill_1 FILLER_49_71 ();
 sg13g2_fill_2 FILLER_49_120 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_decap_4 FILLER_49_200 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_268 ();
 sg13g2_fill_2 FILLER_49_289 ();
 sg13g2_fill_2 FILLER_49_315 ();
 sg13g2_fill_2 FILLER_49_322 ();
 sg13g2_fill_1 FILLER_49_324 ();
 sg13g2_fill_1 FILLER_49_339 ();
 sg13g2_decap_8 FILLER_49_353 ();
 sg13g2_decap_8 FILLER_49_360 ();
 sg13g2_decap_8 FILLER_49_367 ();
 sg13g2_decap_8 FILLER_49_374 ();
 sg13g2_decap_8 FILLER_49_381 ();
 sg13g2_decap_8 FILLER_49_388 ();
 sg13g2_decap_8 FILLER_49_395 ();
 sg13g2_decap_8 FILLER_49_402 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_23 ();
 sg13g2_fill_1 FILLER_50_27 ();
 sg13g2_fill_1 FILLER_50_38 ();
 sg13g2_fill_2 FILLER_50_47 ();
 sg13g2_decap_8 FILLER_50_57 ();
 sg13g2_decap_4 FILLER_50_64 ();
 sg13g2_fill_2 FILLER_50_68 ();
 sg13g2_fill_2 FILLER_50_110 ();
 sg13g2_fill_1 FILLER_50_112 ();
 sg13g2_fill_2 FILLER_50_139 ();
 sg13g2_fill_2 FILLER_50_169 ();
 sg13g2_fill_2 FILLER_50_176 ();
 sg13g2_fill_2 FILLER_50_196 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_fill_1 FILLER_50_218 ();
 sg13g2_fill_2 FILLER_50_224 ();
 sg13g2_fill_2 FILLER_50_231 ();
 sg13g2_fill_2 FILLER_50_247 ();
 sg13g2_fill_1 FILLER_50_249 ();
 sg13g2_fill_2 FILLER_50_310 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_decap_8 FILLER_50_359 ();
 sg13g2_decap_8 FILLER_50_366 ();
 sg13g2_decap_8 FILLER_50_373 ();
 sg13g2_decap_8 FILLER_50_380 ();
 sg13g2_decap_8 FILLER_50_387 ();
 sg13g2_decap_8 FILLER_50_394 ();
 sg13g2_decap_8 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_26 ();
 sg13g2_fill_1 FILLER_51_33 ();
 sg13g2_fill_2 FILLER_51_44 ();
 sg13g2_fill_2 FILLER_51_59 ();
 sg13g2_fill_1 FILLER_51_61 ();
 sg13g2_fill_1 FILLER_51_86 ();
 sg13g2_fill_2 FILLER_51_109 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_fill_1 FILLER_51_138 ();
 sg13g2_fill_2 FILLER_51_145 ();
 sg13g2_fill_1 FILLER_51_147 ();
 sg13g2_fill_2 FILLER_51_185 ();
 sg13g2_fill_2 FILLER_51_192 ();
 sg13g2_decap_8 FILLER_51_226 ();
 sg13g2_decap_8 FILLER_51_233 ();
 sg13g2_decap_4 FILLER_51_240 ();
 sg13g2_fill_1 FILLER_51_248 ();
 sg13g2_fill_2 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_265 ();
 sg13g2_fill_2 FILLER_51_272 ();
 sg13g2_fill_1 FILLER_51_274 ();
 sg13g2_fill_2 FILLER_51_279 ();
 sg13g2_decap_8 FILLER_51_356 ();
 sg13g2_decap_8 FILLER_51_363 ();
 sg13g2_decap_8 FILLER_51_370 ();
 sg13g2_decap_8 FILLER_51_377 ();
 sg13g2_decap_8 FILLER_51_384 ();
 sg13g2_decap_8 FILLER_51_391 ();
 sg13g2_decap_8 FILLER_51_398 ();
 sg13g2_decap_4 FILLER_51_405 ();
 sg13g2_decap_4 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_4 ();
 sg13g2_fill_2 FILLER_52_81 ();
 sg13g2_fill_1 FILLER_52_83 ();
 sg13g2_fill_1 FILLER_52_121 ();
 sg13g2_fill_1 FILLER_52_131 ();
 sg13g2_fill_2 FILLER_52_141 ();
 sg13g2_decap_8 FILLER_52_152 ();
 sg13g2_fill_2 FILLER_52_159 ();
 sg13g2_fill_1 FILLER_52_161 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_241 ();
 sg13g2_decap_8 FILLER_52_254 ();
 sg13g2_decap_8 FILLER_52_261 ();
 sg13g2_fill_2 FILLER_52_279 ();
 sg13g2_fill_1 FILLER_52_281 ();
 sg13g2_fill_1 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_325 ();
 sg13g2_decap_8 FILLER_52_347 ();
 sg13g2_decap_4 FILLER_52_354 ();
 sg13g2_decap_8 FILLER_52_363 ();
 sg13g2_decap_8 FILLER_52_370 ();
 sg13g2_decap_8 FILLER_52_377 ();
 sg13g2_decap_8 FILLER_52_384 ();
 sg13g2_decap_8 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_398 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_65 ();
 sg13g2_fill_1 FILLER_53_92 ();
 sg13g2_fill_2 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_126 ();
 sg13g2_fill_2 FILLER_53_135 ();
 sg13g2_fill_1 FILLER_53_137 ();
 sg13g2_decap_4 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_159 ();
 sg13g2_fill_2 FILLER_53_166 ();
 sg13g2_fill_1 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_191 ();
 sg13g2_fill_2 FILLER_53_246 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_fill_2 FILLER_53_275 ();
 sg13g2_fill_2 FILLER_53_290 ();
 sg13g2_fill_1 FILLER_53_292 ();
 sg13g2_decap_8 FILLER_53_336 ();
 sg13g2_decap_4 FILLER_53_343 ();
 sg13g2_fill_2 FILLER_53_347 ();
 sg13g2_decap_8 FILLER_53_358 ();
 sg13g2_decap_8 FILLER_53_365 ();
 sg13g2_decap_8 FILLER_53_372 ();
 sg13g2_decap_8 FILLER_53_379 ();
 sg13g2_decap_8 FILLER_53_386 ();
 sg13g2_decap_8 FILLER_53_393 ();
 sg13g2_decap_8 FILLER_53_400 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_fill_2 FILLER_54_37 ();
 sg13g2_fill_2 FILLER_54_70 ();
 sg13g2_fill_1 FILLER_54_72 ();
 sg13g2_fill_2 FILLER_54_88 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_2 FILLER_54_159 ();
 sg13g2_decap_4 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_206 ();
 sg13g2_decap_8 FILLER_54_213 ();
 sg13g2_decap_8 FILLER_54_220 ();
 sg13g2_fill_1 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_fill_1 FILLER_54_303 ();
 sg13g2_fill_1 FILLER_54_321 ();
 sg13g2_decap_8 FILLER_54_331 ();
 sg13g2_fill_1 FILLER_54_338 ();
 sg13g2_decap_8 FILLER_54_391 ();
 sg13g2_decap_8 FILLER_54_398 ();
 sg13g2_decap_4 FILLER_54_405 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_9 ();
 sg13g2_fill_1 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_101 ();
 sg13g2_fill_1 FILLER_55_123 ();
 sg13g2_fill_2 FILLER_55_155 ();
 sg13g2_fill_1 FILLER_55_169 ();
 sg13g2_decap_8 FILLER_55_180 ();
 sg13g2_decap_8 FILLER_55_187 ();
 sg13g2_decap_8 FILLER_55_208 ();
 sg13g2_fill_2 FILLER_55_215 ();
 sg13g2_decap_4 FILLER_55_234 ();
 sg13g2_decap_4 FILLER_55_241 ();
 sg13g2_fill_2 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_251 ();
 sg13g2_fill_1 FILLER_55_262 ();
 sg13g2_decap_8 FILLER_55_292 ();
 sg13g2_fill_1 FILLER_55_299 ();
 sg13g2_decap_4 FILLER_55_303 ();
 sg13g2_fill_1 FILLER_55_307 ();
 sg13g2_fill_1 FILLER_55_343 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_37 ();
 sg13g2_fill_1 FILLER_56_39 ();
 sg13g2_fill_1 FILLER_56_50 ();
 sg13g2_decap_4 FILLER_56_120 ();
 sg13g2_fill_1 FILLER_56_124 ();
 sg13g2_fill_2 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_150 ();
 sg13g2_decap_4 FILLER_56_169 ();
 sg13g2_fill_2 FILLER_56_173 ();
 sg13g2_fill_2 FILLER_56_188 ();
 sg13g2_fill_1 FILLER_56_242 ();
 sg13g2_fill_2 FILLER_56_281 ();
 sg13g2_fill_1 FILLER_56_299 ();
 sg13g2_decap_4 FILLER_56_304 ();
 sg13g2_decap_4 FILLER_56_311 ();
 sg13g2_fill_2 FILLER_56_330 ();
 sg13g2_fill_1 FILLER_56_332 ();
 sg13g2_fill_2 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_400 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_21 ();
 sg13g2_fill_1 FILLER_57_52 ();
 sg13g2_fill_2 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_fill_1 FILLER_57_147 ();
 sg13g2_fill_2 FILLER_57_168 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_fill_1 FILLER_57_188 ();
 sg13g2_fill_1 FILLER_57_200 ();
 sg13g2_fill_1 FILLER_57_214 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_fill_2 FILLER_57_313 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_2 FILLER_57_348 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_fill_2 FILLER_57_390 ();
 sg13g2_decap_8 FILLER_57_395 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_4 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_18 ();
 sg13g2_fill_1 FILLER_58_55 ();
 sg13g2_decap_4 FILLER_58_117 ();
 sg13g2_fill_1 FILLER_58_121 ();
 sg13g2_fill_2 FILLER_58_130 ();
 sg13g2_decap_4 FILLER_58_160 ();
 sg13g2_fill_2 FILLER_58_164 ();
 sg13g2_fill_2 FILLER_58_208 ();
 sg13g2_fill_2 FILLER_58_215 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_fill_1 FILLER_58_253 ();
 sg13g2_decap_8 FILLER_58_268 ();
 sg13g2_fill_2 FILLER_58_288 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_1 FILLER_58_303 ();
 sg13g2_fill_1 FILLER_58_318 ();
 sg13g2_fill_2 FILLER_58_328 ();
 sg13g2_fill_2 FILLER_58_353 ();
 sg13g2_fill_2 FILLER_58_369 ();
 sg13g2_fill_2 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_397 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_4 FILLER_59_21 ();
 sg13g2_fill_1 FILLER_59_65 ();
 sg13g2_fill_1 FILLER_59_71 ();
 sg13g2_fill_1 FILLER_59_81 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_decap_8 FILLER_59_100 ();
 sg13g2_decap_4 FILLER_59_107 ();
 sg13g2_decap_8 FILLER_59_124 ();
 sg13g2_fill_2 FILLER_59_131 ();
 sg13g2_fill_2 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_153 ();
 sg13g2_fill_2 FILLER_59_163 ();
 sg13g2_fill_1 FILLER_59_165 ();
 sg13g2_fill_1 FILLER_59_172 ();
 sg13g2_fill_2 FILLER_59_180 ();
 sg13g2_fill_2 FILLER_59_202 ();
 sg13g2_fill_1 FILLER_59_204 ();
 sg13g2_decap_8 FILLER_59_211 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_fill_1 FILLER_59_235 ();
 sg13g2_fill_2 FILLER_59_245 ();
 sg13g2_fill_2 FILLER_59_256 ();
 sg13g2_fill_2 FILLER_59_263 ();
 sg13g2_fill_2 FILLER_59_398 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_fill_2 FILLER_60_11 ();
 sg13g2_decap_8 FILLER_60_16 ();
 sg13g2_fill_2 FILLER_60_23 ();
 sg13g2_fill_1 FILLER_60_25 ();
 sg13g2_fill_1 FILLER_60_61 ();
 sg13g2_decap_4 FILLER_60_66 ();
 sg13g2_fill_1 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_75 ();
 sg13g2_decap_8 FILLER_60_82 ();
 sg13g2_decap_8 FILLER_60_89 ();
 sg13g2_decap_8 FILLER_60_96 ();
 sg13g2_fill_2 FILLER_60_103 ();
 sg13g2_fill_1 FILLER_60_105 ();
 sg13g2_fill_2 FILLER_60_120 ();
 sg13g2_fill_1 FILLER_60_137 ();
 sg13g2_fill_1 FILLER_60_154 ();
 sg13g2_fill_1 FILLER_60_169 ();
 sg13g2_fill_2 FILLER_60_175 ();
 sg13g2_fill_1 FILLER_60_186 ();
 sg13g2_decap_8 FILLER_60_195 ();
 sg13g2_decap_4 FILLER_60_237 ();
 sg13g2_fill_2 FILLER_60_241 ();
 sg13g2_fill_2 FILLER_60_304 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_27 ();
 sg13g2_fill_2 FILLER_61_34 ();
 sg13g2_fill_1 FILLER_61_36 ();
 sg13g2_decap_8 FILLER_61_45 ();
 sg13g2_decap_4 FILLER_61_52 ();
 sg13g2_fill_2 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_61 ();
 sg13g2_decap_8 FILLER_61_68 ();
 sg13g2_decap_8 FILLER_61_75 ();
 sg13g2_decap_4 FILLER_61_82 ();
 sg13g2_fill_1 FILLER_61_86 ();
 sg13g2_fill_2 FILLER_61_162 ();
 sg13g2_fill_2 FILLER_61_169 ();
 sg13g2_fill_2 FILLER_61_178 ();
 sg13g2_fill_1 FILLER_61_221 ();
 sg13g2_decap_4 FILLER_61_226 ();
 sg13g2_decap_8 FILLER_61_239 ();
 sg13g2_decap_8 FILLER_61_246 ();
 sg13g2_fill_1 FILLER_61_253 ();
 sg13g2_fill_2 FILLER_61_258 ();
 sg13g2_fill_1 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_311 ();
 sg13g2_fill_2 FILLER_61_321 ();
 sg13g2_fill_1 FILLER_61_327 ();
 sg13g2_decap_4 FILLER_61_332 ();
 sg13g2_fill_1 FILLER_61_336 ();
 sg13g2_fill_2 FILLER_61_340 ();
 sg13g2_fill_1 FILLER_61_342 ();
 sg13g2_fill_1 FILLER_61_357 ();
 sg13g2_decap_4 FILLER_61_379 ();
 sg13g2_fill_2 FILLER_62_43 ();
 sg13g2_fill_1 FILLER_62_45 ();
 sg13g2_fill_2 FILLER_62_110 ();
 sg13g2_fill_2 FILLER_62_148 ();
 sg13g2_decap_4 FILLER_62_167 ();
 sg13g2_fill_1 FILLER_62_171 ();
 sg13g2_fill_2 FILLER_62_192 ();
 sg13g2_fill_1 FILLER_62_194 ();
 sg13g2_fill_2 FILLER_62_268 ();
 sg13g2_fill_1 FILLER_62_309 ();
 sg13g2_fill_1 FILLER_62_319 ();
 sg13g2_fill_2 FILLER_62_326 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_fill_2 FILLER_62_349 ();
 sg13g2_fill_1 FILLER_62_351 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_53 ();
 sg13g2_fill_2 FILLER_63_59 ();
 sg13g2_fill_1 FILLER_63_61 ();
 sg13g2_fill_2 FILLER_63_88 ();
 sg13g2_fill_1 FILLER_63_90 ();
 sg13g2_fill_1 FILLER_63_101 ();
 sg13g2_fill_2 FILLER_63_116 ();
 sg13g2_decap_8 FILLER_63_160 ();
 sg13g2_decap_4 FILLER_63_167 ();
 sg13g2_fill_2 FILLER_63_171 ();
 sg13g2_fill_1 FILLER_63_177 ();
 sg13g2_fill_2 FILLER_63_182 ();
 sg13g2_fill_1 FILLER_63_184 ();
 sg13g2_decap_8 FILLER_63_198 ();
 sg13g2_decap_8 FILLER_63_205 ();
 sg13g2_decap_4 FILLER_63_212 ();
 sg13g2_fill_2 FILLER_63_216 ();
 sg13g2_fill_1 FILLER_63_222 ();
 sg13g2_fill_2 FILLER_63_236 ();
 sg13g2_fill_1 FILLER_63_238 ();
 sg13g2_fill_2 FILLER_63_323 ();
 sg13g2_fill_2 FILLER_63_361 ();
 sg13g2_fill_1 FILLER_63_377 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_20 ();
 sg13g2_fill_1 FILLER_64_39 ();
 sg13g2_fill_1 FILLER_64_72 ();
 sg13g2_fill_2 FILLER_64_81 ();
 sg13g2_decap_4 FILLER_64_88 ();
 sg13g2_fill_2 FILLER_64_109 ();
 sg13g2_decap_8 FILLER_64_116 ();
 sg13g2_fill_2 FILLER_64_123 ();
 sg13g2_fill_1 FILLER_64_125 ();
 sg13g2_decap_4 FILLER_64_139 ();
 sg13g2_fill_1 FILLER_64_161 ();
 sg13g2_decap_4 FILLER_64_240 ();
 sg13g2_fill_2 FILLER_64_253 ();
 sg13g2_fill_1 FILLER_64_255 ();
 sg13g2_fill_2 FILLER_64_268 ();
 sg13g2_fill_1 FILLER_64_310 ();
 sg13g2_fill_2 FILLER_64_332 ();
 sg13g2_fill_2 FILLER_64_353 ();
 sg13g2_fill_1 FILLER_64_386 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_fill_2 FILLER_65_42 ();
 sg13g2_fill_1 FILLER_65_58 ();
 sg13g2_decap_8 FILLER_65_89 ();
 sg13g2_decap_8 FILLER_65_96 ();
 sg13g2_decap_4 FILLER_65_107 ();
 sg13g2_fill_2 FILLER_65_111 ();
 sg13g2_decap_8 FILLER_65_127 ();
 sg13g2_decap_8 FILLER_65_134 ();
 sg13g2_fill_2 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_143 ();
 sg13g2_fill_2 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_65_190 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_fill_1 FILLER_65_252 ();
 sg13g2_decap_4 FILLER_65_261 ();
 sg13g2_fill_2 FILLER_65_344 ();
 sg13g2_fill_2 FILLER_65_380 ();
 sg13g2_fill_2 FILLER_65_398 ();
 sg13g2_fill_2 FILLER_66_31 ();
 sg13g2_fill_2 FILLER_66_56 ();
 sg13g2_fill_2 FILLER_66_84 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_decap_4 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_95 ();
 sg13g2_fill_1 FILLER_66_100 ();
 sg13g2_fill_2 FILLER_66_131 ();
 sg13g2_fill_1 FILLER_66_133 ();
 sg13g2_fill_1 FILLER_66_160 ();
 sg13g2_decap_8 FILLER_66_187 ();
 sg13g2_decap_4 FILLER_66_194 ();
 sg13g2_decap_8 FILLER_66_206 ();
 sg13g2_decap_4 FILLER_66_213 ();
 sg13g2_fill_2 FILLER_66_217 ();
 sg13g2_fill_2 FILLER_66_224 ();
 sg13g2_fill_1 FILLER_66_226 ();
 sg13g2_decap_4 FILLER_66_253 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_decap_8 FILLER_66_262 ();
 sg13g2_decap_4 FILLER_66_269 ();
 sg13g2_fill_1 FILLER_66_273 ();
 sg13g2_fill_1 FILLER_66_324 ();
 sg13g2_fill_2 FILLER_66_355 ();
 sg13g2_fill_1 FILLER_66_357 ();
 sg13g2_fill_2 FILLER_66_366 ();
 sg13g2_fill_1 FILLER_66_368 ();
 sg13g2_fill_2 FILLER_66_381 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_33 ();
 sg13g2_decap_8 FILLER_67_60 ();
 sg13g2_fill_2 FILLER_67_67 ();
 sg13g2_decap_8 FILLER_67_73 ();
 sg13g2_fill_1 FILLER_67_106 ();
 sg13g2_decap_8 FILLER_67_138 ();
 sg13g2_decap_8 FILLER_67_145 ();
 sg13g2_decap_8 FILLER_67_152 ();
 sg13g2_decap_4 FILLER_67_159 ();
 sg13g2_fill_1 FILLER_67_163 ();
 sg13g2_fill_2 FILLER_67_169 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_fill_2 FILLER_67_210 ();
 sg13g2_fill_2 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_fill_1 FILLER_67_293 ();
 sg13g2_fill_1 FILLER_67_300 ();
 sg13g2_fill_2 FILLER_67_314 ();
 sg13g2_decap_4 FILLER_67_329 ();
 sg13g2_decap_4 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_344 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_11 ();
 sg13g2_fill_2 FILLER_68_64 ();
 sg13g2_fill_2 FILLER_68_138 ();
 sg13g2_fill_1 FILLER_68_140 ();
 sg13g2_fill_1 FILLER_68_181 ();
 sg13g2_fill_2 FILLER_68_218 ();
 sg13g2_fill_2 FILLER_68_262 ();
 sg13g2_fill_2 FILLER_68_295 ();
 sg13g2_fill_1 FILLER_68_297 ();
 sg13g2_decap_4 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_328 ();
 sg13g2_fill_1 FILLER_68_330 ();
 sg13g2_decap_8 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_350 ();
 sg13g2_decap_8 FILLER_68_357 ();
 sg13g2_fill_1 FILLER_68_372 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_fill_2 FILLER_69_35 ();
 sg13g2_fill_1 FILLER_69_37 ();
 sg13g2_fill_2 FILLER_69_56 ();
 sg13g2_fill_1 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_97 ();
 sg13g2_fill_2 FILLER_69_129 ();
 sg13g2_fill_1 FILLER_69_131 ();
 sg13g2_decap_4 FILLER_69_157 ();
 sg13g2_fill_2 FILLER_69_161 ();
 sg13g2_fill_2 FILLER_69_173 ();
 sg13g2_fill_2 FILLER_69_199 ();
 sg13g2_decap_4 FILLER_69_209 ();
 sg13g2_fill_2 FILLER_69_222 ();
 sg13g2_fill_2 FILLER_69_237 ();
 sg13g2_fill_1 FILLER_69_261 ();
 sg13g2_decap_4 FILLER_69_288 ();
 sg13g2_fill_1 FILLER_69_292 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_decap_4 FILLER_69_349 ();
 sg13g2_fill_1 FILLER_69_353 ();
 sg13g2_fill_2 FILLER_69_398 ();
 sg13g2_fill_2 FILLER_70_13 ();
 sg13g2_fill_1 FILLER_70_15 ();
 sg13g2_fill_2 FILLER_70_26 ();
 sg13g2_fill_1 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_33 ();
 sg13g2_fill_2 FILLER_70_66 ();
 sg13g2_fill_1 FILLER_70_127 ();
 sg13g2_decap_8 FILLER_70_132 ();
 sg13g2_decap_8 FILLER_70_139 ();
 sg13g2_decap_8 FILLER_70_146 ();
 sg13g2_decap_8 FILLER_70_153 ();
 sg13g2_decap_8 FILLER_70_160 ();
 sg13g2_fill_1 FILLER_70_167 ();
 sg13g2_fill_1 FILLER_70_205 ();
 sg13g2_fill_1 FILLER_70_214 ();
 sg13g2_fill_2 FILLER_70_220 ();
 sg13g2_decap_8 FILLER_70_311 ();
 sg13g2_fill_2 FILLER_70_318 ();
 sg13g2_fill_1 FILLER_70_320 ();
 sg13g2_fill_1 FILLER_70_327 ();
 sg13g2_fill_2 FILLER_70_369 ();
 sg13g2_fill_1 FILLER_71_40 ();
 sg13g2_fill_2 FILLER_71_66 ();
 sg13g2_fill_2 FILLER_71_75 ();
 sg13g2_fill_1 FILLER_71_114 ();
 sg13g2_fill_2 FILLER_71_120 ();
 sg13g2_decap_4 FILLER_71_126 ();
 sg13g2_fill_1 FILLER_71_130 ();
 sg13g2_fill_2 FILLER_71_139 ();
 sg13g2_decap_4 FILLER_71_145 ();
 sg13g2_fill_1 FILLER_71_149 ();
 sg13g2_fill_2 FILLER_71_154 ();
 sg13g2_fill_1 FILLER_71_156 ();
 sg13g2_fill_2 FILLER_71_218 ();
 sg13g2_fill_1 FILLER_71_220 ();
 sg13g2_fill_1 FILLER_71_284 ();
 sg13g2_decap_4 FILLER_71_319 ();
 sg13g2_fill_1 FILLER_71_340 ();
 sg13g2_fill_1 FILLER_71_347 ();
 sg13g2_fill_1 FILLER_71_391 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_44 ();
 sg13g2_decap_8 FILLER_72_51 ();
 sg13g2_fill_2 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_109 ();
 sg13g2_fill_2 FILLER_72_137 ();
 sg13g2_fill_1 FILLER_72_169 ();
 sg13g2_fill_1 FILLER_72_209 ();
 sg13g2_fill_1 FILLER_72_216 ();
 sg13g2_fill_2 FILLER_72_254 ();
 sg13g2_fill_1 FILLER_72_266 ();
 sg13g2_fill_1 FILLER_72_290 ();
 sg13g2_fill_2 FILLER_72_309 ();
 sg13g2_fill_2 FILLER_72_353 ();
 sg13g2_fill_2 FILLER_72_381 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_1 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_11 ();
 sg13g2_fill_1 FILLER_73_52 ();
 sg13g2_fill_2 FILLER_73_135 ();
 sg13g2_fill_1 FILLER_73_137 ();
 sg13g2_fill_2 FILLER_73_172 ();
 sg13g2_fill_1 FILLER_73_193 ();
 sg13g2_decap_8 FILLER_73_202 ();
 sg13g2_fill_2 FILLER_73_214 ();
 sg13g2_decap_4 FILLER_73_282 ();
 sg13g2_fill_1 FILLER_73_286 ();
 sg13g2_fill_2 FILLER_73_302 ();
 sg13g2_fill_1 FILLER_73_304 ();
 sg13g2_decap_4 FILLER_73_315 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_fill_2 FILLER_73_332 ();
 sg13g2_fill_1 FILLER_73_340 ();
 sg13g2_fill_1 FILLER_73_363 ();
 sg13g2_fill_1 FILLER_73_387 ();
 sg13g2_fill_2 FILLER_73_393 ();
 sg13g2_fill_2 FILLER_74_39 ();
 sg13g2_fill_1 FILLER_74_107 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_decap_8 FILLER_74_194 ();
 sg13g2_decap_8 FILLER_74_201 ();
 sg13g2_decap_8 FILLER_74_208 ();
 sg13g2_decap_4 FILLER_74_215 ();
 sg13g2_fill_2 FILLER_74_223 ();
 sg13g2_decap_4 FILLER_74_229 ();
 sg13g2_fill_1 FILLER_74_233 ();
 sg13g2_fill_2 FILLER_74_238 ();
 sg13g2_fill_2 FILLER_74_268 ();
 sg13g2_fill_1 FILLER_74_270 ();
 sg13g2_fill_1 FILLER_74_274 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_15 ();
 sg13g2_decap_8 FILLER_75_22 ();
 sg13g2_decap_8 FILLER_75_29 ();
 sg13g2_decap_8 FILLER_75_36 ();
 sg13g2_decap_4 FILLER_75_43 ();
 sg13g2_fill_2 FILLER_75_67 ();
 sg13g2_fill_2 FILLER_75_78 ();
 sg13g2_fill_2 FILLER_75_100 ();
 sg13g2_fill_2 FILLER_75_115 ();
 sg13g2_fill_2 FILLER_75_137 ();
 sg13g2_fill_2 FILLER_75_198 ();
 sg13g2_decap_4 FILLER_75_205 ();
 sg13g2_fill_1 FILLER_75_209 ();
 sg13g2_fill_2 FILLER_75_232 ();
 sg13g2_fill_1 FILLER_75_234 ();
 sg13g2_decap_8 FILLER_75_239 ();
 sg13g2_decap_4 FILLER_75_246 ();
 sg13g2_fill_2 FILLER_75_250 ();
 sg13g2_fill_2 FILLER_75_275 ();
 sg13g2_fill_2 FILLER_75_290 ();
 sg13g2_fill_1 FILLER_75_292 ();
 sg13g2_fill_1 FILLER_75_322 ();
 sg13g2_fill_1 FILLER_75_339 ();
 sg13g2_fill_1 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_fill_1 FILLER_76_75 ();
 sg13g2_fill_1 FILLER_76_91 ();
 sg13g2_decap_4 FILLER_76_115 ();
 sg13g2_fill_2 FILLER_76_119 ();
 sg13g2_fill_1 FILLER_76_133 ();
 sg13g2_fill_1 FILLER_76_161 ();
 sg13g2_fill_2 FILLER_76_286 ();
 sg13g2_fill_1 FILLER_76_288 ();
 sg13g2_fill_2 FILLER_76_330 ();
 sg13g2_fill_2 FILLER_76_347 ();
 sg13g2_fill_1 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_4 FILLER_77_49 ();
 sg13g2_fill_1 FILLER_77_53 ();
 sg13g2_fill_1 FILLER_77_80 ();
 sg13g2_fill_2 FILLER_77_97 ();
 sg13g2_fill_2 FILLER_77_130 ();
 sg13g2_fill_1 FILLER_77_132 ();
 sg13g2_fill_1 FILLER_77_261 ();
 sg13g2_fill_1 FILLER_77_310 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_4 FILLER_78_49 ();
 sg13g2_fill_1 FILLER_78_53 ();
 sg13g2_fill_2 FILLER_78_103 ();
 sg13g2_fill_1 FILLER_78_105 ();
 sg13g2_fill_1 FILLER_78_176 ();
 sg13g2_fill_1 FILLER_78_198 ();
 sg13g2_fill_2 FILLER_78_275 ();
 sg13g2_fill_1 FILLER_78_277 ();
 sg13g2_fill_1 FILLER_78_287 ();
 sg13g2_fill_1 FILLER_78_297 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_4 FILLER_79_56 ();
 sg13g2_fill_1 FILLER_79_64 ();
 sg13g2_fill_2 FILLER_79_73 ();
 sg13g2_fill_1 FILLER_79_75 ();
 sg13g2_fill_1 FILLER_79_115 ();
 sg13g2_fill_2 FILLER_79_136 ();
 sg13g2_fill_1 FILLER_79_138 ();
 sg13g2_fill_1 FILLER_79_170 ();
 sg13g2_fill_1 FILLER_79_202 ();
 sg13g2_fill_1 FILLER_79_354 ();
 sg13g2_fill_1 FILLER_79_381 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_68 ();
 sg13g2_fill_1 FILLER_80_70 ();
 sg13g2_fill_2 FILLER_80_93 ();
 sg13g2_fill_1 FILLER_80_95 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_fill_2 FILLER_80_162 ();
 sg13g2_fill_1 FILLER_80_169 ();
 sg13g2_fill_2 FILLER_80_184 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_fill_1 FILLER_80_213 ();
 sg13g2_fill_2 FILLER_80_227 ();
 sg13g2_fill_1 FILLER_80_229 ();
 sg13g2_fill_2 FILLER_80_322 ();
 assign uio_oe[0] = net313;
 assign uio_oe[1] = net314;
 assign uio_oe[2] = net315;
 assign uio_oe[3] = net316;
 assign uio_oe[4] = net317;
 assign uio_oe[5] = net318;
 assign uio_oe[6] = net319;
 assign uio_oe[7] = net320;
 assign uio_out[7] = net6;
 assign uo_out[7] = net7;
endmodule

module tt_um_rejunity_z80 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire clknet_leaf_0_clk;
 wire \addr_bus[0] ;
 wire \addr_bus[10] ;
 wire \addr_bus[11] ;
 wire \addr_bus[12] ;
 wire \addr_bus[13] ;
 wire \addr_bus[14] ;
 wire \addr_bus[15] ;
 wire \addr_bus[1] ;
 wire \addr_bus[2] ;
 wire \addr_bus[3] ;
 wire \addr_bus[4] ;
 wire \addr_bus[5] ;
 wire \addr_bus[6] ;
 wire \addr_bus[7] ;
 wire \addr_bus[8] ;
 wire \addr_bus[9] ;
 wire doe;
 wire \z80.iorq_n ;
 wire \z80.m1_n ;
 wire \z80.mreq_n ;
 wire \z80.rd_n ;
 wire \z80.rfsh_n ;
 wire \z80.tv80s.di_reg[0] ;
 wire \z80.tv80s.di_reg[1] ;
 wire \z80.tv80s.di_reg[2] ;
 wire \z80.tv80s.di_reg[3] ;
 wire \z80.tv80s.di_reg[4] ;
 wire \z80.tv80s.di_reg[5] ;
 wire \z80.tv80s.di_reg[6] ;
 wire \z80.tv80s.di_reg[7] ;
 wire \z80.tv80s.i_tv80_core.ACC[0] ;
 wire \z80.tv80s.i_tv80_core.ACC[1] ;
 wire \z80.tv80s.i_tv80_core.ACC[2] ;
 wire \z80.tv80s.i_tv80_core.ACC[3] ;
 wire \z80.tv80s.i_tv80_core.ACC[4] ;
 wire \z80.tv80s.i_tv80_core.ACC[5] ;
 wire \z80.tv80s.i_tv80_core.ACC[6] ;
 wire \z80.tv80s.i_tv80_core.ACC[7] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[0] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[1] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[2] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[3] ;
 wire \z80.tv80s.i_tv80_core.Alternate ;
 wire \z80.tv80s.i_tv80_core.Ap[0] ;
 wire \z80.tv80s.i_tv80_core.Ap[1] ;
 wire \z80.tv80s.i_tv80_core.Ap[2] ;
 wire \z80.tv80s.i_tv80_core.Ap[3] ;
 wire \z80.tv80s.i_tv80_core.Ap[4] ;
 wire \z80.tv80s.i_tv80_core.Ap[5] ;
 wire \z80.tv80s.i_tv80_core.Ap[6] ;
 wire \z80.tv80s.i_tv80_core.Ap[7] ;
 wire \z80.tv80s.i_tv80_core.Arith16_r ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t1 ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t2 ;
 wire \z80.tv80s.i_tv80_core.BTR_r ;
 wire \z80.tv80s.i_tv80_core.BusA[0] ;
 wire \z80.tv80s.i_tv80_core.BusA[1] ;
 wire \z80.tv80s.i_tv80_core.BusA[2] ;
 wire \z80.tv80s.i_tv80_core.BusA[3] ;
 wire \z80.tv80s.i_tv80_core.BusA[4] ;
 wire \z80.tv80s.i_tv80_core.BusA[5] ;
 wire \z80.tv80s.i_tv80_core.BusA[6] ;
 wire \z80.tv80s.i_tv80_core.BusA[7] ;
 wire \z80.tv80s.i_tv80_core.BusAck ;
 wire \z80.tv80s.i_tv80_core.BusB[0] ;
 wire \z80.tv80s.i_tv80_core.BusB[1] ;
 wire \z80.tv80s.i_tv80_core.BusB[2] ;
 wire \z80.tv80s.i_tv80_core.BusB[3] ;
 wire \z80.tv80s.i_tv80_core.BusB[4] ;
 wire \z80.tv80s.i_tv80_core.BusB[5] ;
 wire \z80.tv80s.i_tv80_core.BusB[6] ;
 wire \z80.tv80s.i_tv80_core.BusB[7] ;
 wire \z80.tv80s.i_tv80_core.BusReq_s ;
 wire \z80.tv80s.i_tv80_core.F[0] ;
 wire \z80.tv80s.i_tv80_core.F[1] ;
 wire \z80.tv80s.i_tv80_core.F[2] ;
 wire \z80.tv80s.i_tv80_core.F[3] ;
 wire \z80.tv80s.i_tv80_core.F[4] ;
 wire \z80.tv80s.i_tv80_core.F[5] ;
 wire \z80.tv80s.i_tv80_core.F[6] ;
 wire \z80.tv80s.i_tv80_core.F[7] ;
 wire \z80.tv80s.i_tv80_core.Fp[0] ;
 wire \z80.tv80s.i_tv80_core.Fp[1] ;
 wire \z80.tv80s.i_tv80_core.Fp[2] ;
 wire \z80.tv80s.i_tv80_core.Fp[3] ;
 wire \z80.tv80s.i_tv80_core.Fp[4] ;
 wire \z80.tv80s.i_tv80_core.Fp[5] ;
 wire \z80.tv80s.i_tv80_core.Fp[6] ;
 wire \z80.tv80s.i_tv80_core.Fp[7] ;
 wire \z80.tv80s.i_tv80_core.Halt_FF ;
 wire \z80.tv80s.i_tv80_core.INT_s ;
 wire \z80.tv80s.i_tv80_core.IR[0] ;
 wire \z80.tv80s.i_tv80_core.IR[1] ;
 wire \z80.tv80s.i_tv80_core.IR[2] ;
 wire \z80.tv80s.i_tv80_core.IR[3] ;
 wire \z80.tv80s.i_tv80_core.IR[4] ;
 wire \z80.tv80s.i_tv80_core.IR[5] ;
 wire \z80.tv80s.i_tv80_core.IR[6] ;
 wire \z80.tv80s.i_tv80_core.IR[7] ;
 wire \z80.tv80s.i_tv80_core.ISet[0] ;
 wire \z80.tv80s.i_tv80_core.ISet[1] ;
 wire \z80.tv80s.i_tv80_core.ISet[2] ;
 wire \z80.tv80s.i_tv80_core.ISet[3] ;
 wire \z80.tv80s.i_tv80_core.IStatus[1] ;
 wire \z80.tv80s.i_tv80_core.IStatus[2] ;
 wire \z80.tv80s.i_tv80_core.I[0] ;
 wire \z80.tv80s.i_tv80_core.I[1] ;
 wire \z80.tv80s.i_tv80_core.I[2] ;
 wire \z80.tv80s.i_tv80_core.I[3] ;
 wire \z80.tv80s.i_tv80_core.I[4] ;
 wire \z80.tv80s.i_tv80_core.I[5] ;
 wire \z80.tv80s.i_tv80_core.I[6] ;
 wire \z80.tv80s.i_tv80_core.I[7] ;
 wire \z80.tv80s.i_tv80_core.IncDecZ ;
 wire \z80.tv80s.i_tv80_core.IntCycle ;
 wire \z80.tv80s.i_tv80_core.IntE ;
 wire \z80.tv80s.i_tv80_core.IntE_FF2 ;
 wire \z80.tv80s.i_tv80_core.NMICycle ;
 wire \z80.tv80s.i_tv80_core.NMI_s ;
 wire \z80.tv80s.i_tv80_core.No_BTR ;
 wire \z80.tv80s.i_tv80_core.Oldnmi_n ;
 wire \z80.tv80s.i_tv80_core.PC[0] ;
 wire \z80.tv80s.i_tv80_core.PC[10] ;
 wire \z80.tv80s.i_tv80_core.PC[11] ;
 wire \z80.tv80s.i_tv80_core.PC[12] ;
 wire \z80.tv80s.i_tv80_core.PC[13] ;
 wire \z80.tv80s.i_tv80_core.PC[14] ;
 wire \z80.tv80s.i_tv80_core.PC[15] ;
 wire \z80.tv80s.i_tv80_core.PC[1] ;
 wire \z80.tv80s.i_tv80_core.PC[2] ;
 wire \z80.tv80s.i_tv80_core.PC[3] ;
 wire \z80.tv80s.i_tv80_core.PC[4] ;
 wire \z80.tv80s.i_tv80_core.PC[5] ;
 wire \z80.tv80s.i_tv80_core.PC[6] ;
 wire \z80.tv80s.i_tv80_core.PC[7] ;
 wire \z80.tv80s.i_tv80_core.PC[8] ;
 wire \z80.tv80s.i_tv80_core.PC[9] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ;
 wire \z80.tv80s.i_tv80_core.PreserveC_r ;
 wire \z80.tv80s.i_tv80_core.R[0] ;
 wire \z80.tv80s.i_tv80_core.R[1] ;
 wire \z80.tv80s.i_tv80_core.R[2] ;
 wire \z80.tv80s.i_tv80_core.R[3] ;
 wire \z80.tv80s.i_tv80_core.R[4] ;
 wire \z80.tv80s.i_tv80_core.R[5] ;
 wire \z80.tv80s.i_tv80_core.R[6] ;
 wire \z80.tv80s.i_tv80_core.R[7] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[10] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[11] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[12] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[13] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[14] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[15] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[3] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[5] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[6] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[7] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[8] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[9] ;
 wire \z80.tv80s.i_tv80_core.SP[0] ;
 wire \z80.tv80s.i_tv80_core.SP[10] ;
 wire \z80.tv80s.i_tv80_core.SP[11] ;
 wire \z80.tv80s.i_tv80_core.SP[12] ;
 wire \z80.tv80s.i_tv80_core.SP[13] ;
 wire \z80.tv80s.i_tv80_core.SP[14] ;
 wire \z80.tv80s.i_tv80_core.SP[15] ;
 wire \z80.tv80s.i_tv80_core.SP[1] ;
 wire \z80.tv80s.i_tv80_core.SP[2] ;
 wire \z80.tv80s.i_tv80_core.SP[3] ;
 wire \z80.tv80s.i_tv80_core.SP[4] ;
 wire \z80.tv80s.i_tv80_core.SP[5] ;
 wire \z80.tv80s.i_tv80_core.SP[6] ;
 wire \z80.tv80s.i_tv80_core.SP[7] ;
 wire \z80.tv80s.i_tv80_core.SP[8] ;
 wire \z80.tv80s.i_tv80_core.SP[9] ;
 wire \z80.tv80s.i_tv80_core.Save_ALU_r ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[0] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[10] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[11] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[12] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[13] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[14] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[15] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[1] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[2] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[3] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[4] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[5] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[6] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[7] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[8] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[9] ;
 wire \z80.tv80s.i_tv80_core.XY_Ind ;
 wire \z80.tv80s.i_tv80_core.XY_State[0] ;
 wire \z80.tv80s.i_tv80_core.XY_State[1] ;
 wire \z80.tv80s.i_tv80_core.Z16_r ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ;
 wire \z80.tv80s.i_tv80_core.mcycles[1] ;
 wire \z80.tv80s.i_tv80_core.mcycles[2] ;
 wire \z80.tv80s.i_tv80_core.mcycles[4] ;
 wire \z80.tv80s.i_tv80_core.mcycles[5] ;
 wire \z80.tv80s.i_tv80_core.ts[0] ;
 wire \z80.tv80s.i_tv80_core.ts[1] ;
 wire \z80.tv80s.i_tv80_core.ts[2] ;
 wire \z80.tv80s.i_tv80_core.ts[3] ;
 wire \z80.tv80s.i_tv80_core.ts[4] ;
 wire \z80.tv80s.i_tv80_core.ts[5] ;
 wire \z80.tv80s.i_tv80_core.ts[6] ;
 wire \z80.tv80s.wr_n ;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;

 sg13g2_inv_1 _4803_ (.Y(_0654_),
    .A(net333));
 sg13g2_inv_1 _4804_ (.Y(_0655_),
    .A(_0293_));
 sg13g2_inv_1 _4805_ (.Y(_0656_),
    .A(net323));
 sg13g2_inv_1 _4806_ (.Y(_0657_),
    .A(net309));
 sg13g2_inv_1 _4807_ (.Y(_0658_),
    .A(net338));
 sg13g2_inv_1 _4808_ (.Y(_0659_),
    .A(net229));
 sg13g2_inv_1 _4809_ (.Y(_0660_),
    .A(net341));
 sg13g2_inv_2 _4810_ (.Y(_0661_),
    .A(\z80.tv80s.i_tv80_core.F[7] ));
 sg13g2_inv_2 _4811_ (.Y(_0662_),
    .A(\z80.tv80s.i_tv80_core.F[6] ));
 sg13g2_inv_1 _4812_ (.Y(_0663_),
    .A(\z80.tv80s.i_tv80_core.F[3] ));
 sg13g2_inv_1 _4813_ (.Y(_0664_),
    .A(net2148));
 sg13g2_inv_4 _4814_ (.A(net2151),
    .Y(_0665_));
 sg13g2_inv_1 _4815_ (.Y(_0666_),
    .A(net248));
 sg13g2_inv_1 _4816_ (.Y(_0667_),
    .A(net342));
 sg13g2_inv_1 _4817_ (.Y(_0668_),
    .A(net2103));
 sg13g2_inv_2 _4818_ (.Y(_0669_),
    .A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sg13g2_inv_1 _4819_ (.Y(_0670_),
    .A(net2099));
 sg13g2_inv_4 _4820_ (.A(net2092),
    .Y(_0671_));
 sg13g2_inv_1 _4821_ (.Y(_0672_),
    .A(net2077));
 sg13g2_inv_2 _4822_ (.Y(_0673_),
    .A(net2072));
 sg13g2_inv_1 _4823_ (.Y(_0674_),
    .A(net2123));
 sg13g2_inv_1 _4824_ (.Y(_0675_),
    .A(net2166));
 sg13g2_inv_2 _4825_ (.Y(_0676_),
    .A(net2172));
 sg13g2_inv_2 _4826_ (.Y(_0677_),
    .A(net2113));
 sg13g2_inv_1 _4827_ (.Y(_0678_),
    .A(net2060));
 sg13g2_inv_1 _4828_ (.Y(_0679_),
    .A(net2110));
 sg13g2_inv_2 _4829_ (.Y(_0680_),
    .A(_0022_));
 sg13g2_inv_2 _4830_ (.Y(_0681_),
    .A(\z80.tv80s.i_tv80_core.NMICycle ));
 sg13g2_inv_1 _4831_ (.Y(_0682_),
    .A(net2138));
 sg13g2_inv_1 _4832_ (.Y(_0683_),
    .A(\z80.tv80s.i_tv80_core.ts[1] ));
 sg13g2_inv_1 _4833_ (.Y(_0684_),
    .A(_0021_));
 sg13g2_inv_1 _4834_ (.Y(_0685_),
    .A(net2227));
 sg13g2_inv_1 _4835_ (.Y(_0686_),
    .A(net469));
 sg13g2_inv_1 _4836_ (.Y(_0687_),
    .A(net219));
 sg13g2_inv_1 _4837_ (.Y(_0688_),
    .A(_0031_));
 sg13g2_inv_1 _4838_ (.Y(_0689_),
    .A(net2052));
 sg13g2_inv_2 _4839_ (.Y(_0690_),
    .A(net2032));
 sg13g2_inv_1 _4840_ (.Y(_0691_),
    .A(net225));
 sg13g2_inv_1 _4841_ (.Y(_0692_),
    .A(_0016_));
 sg13g2_inv_1 _4842_ (.Y(_0693_),
    .A(\z80.tv80s.i_tv80_core.Halt_FF ));
 sg13g2_inv_1 _4843_ (.Y(_0694_),
    .A(net446));
 sg13g2_inv_1 _4844_ (.Y(_0695_),
    .A(_0040_));
 sg13g2_inv_2 _4845_ (.Y(_0696_),
    .A(_0039_));
 sg13g2_inv_1 _4846_ (.Y(_0697_),
    .A(_0048_));
 sg13g2_inv_1 _4847_ (.Y(_0698_),
    .A(_0052_));
 sg13g2_inv_1 _4848_ (.Y(_0699_),
    .A(net387));
 sg13g2_inv_1 _4849_ (.Y(_0700_),
    .A(net450));
 sg13g2_inv_1 _4850_ (.Y(_0701_),
    .A(\z80.tv80s.i_tv80_core.SP[10] ));
 sg13g2_inv_1 _4851_ (.Y(_0702_),
    .A(_0059_));
 sg13g2_inv_1 _4852_ (.Y(_0703_),
    .A(_0068_));
 sg13g2_inv_1 _4853_ (.Y(_0704_),
    .A(_0067_));
 sg13g2_inv_1 _4854_ (.Y(_0705_),
    .A(net2048));
 sg13g2_inv_1 _4855_ (.Y(_0706_),
    .A(_0070_));
 sg13g2_inv_1 _4856_ (.Y(_0707_),
    .A(_0074_));
 sg13g2_inv_1 _4857_ (.Y(_0708_),
    .A(_0082_));
 sg13g2_inv_1 _4858_ (.Y(_0709_),
    .A(_0084_));
 sg13g2_inv_1 _4859_ (.Y(_0710_),
    .A(\z80.tv80s.i_tv80_core.SP[12] ));
 sg13g2_inv_1 _4860_ (.Y(_0711_),
    .A(_0092_));
 sg13g2_inv_1 _4861_ (.Y(_0712_),
    .A(_0096_));
 sg13g2_inv_1 _4862_ (.Y(_0713_),
    .A(_0100_));
 sg13g2_inv_1 _4863_ (.Y(_0714_),
    .A(_0107_));
 sg13g2_inv_1 _4864_ (.Y(_0715_),
    .A(_0114_));
 sg13g2_inv_1 _4865_ (.Y(_0716_),
    .A(_0116_));
 sg13g2_inv_1 _4866_ (.Y(_0717_),
    .A(_0115_));
 sg13g2_inv_1 _4867_ (.Y(_0718_),
    .A(\z80.tv80s.i_tv80_core.SP[14] ));
 sg13g2_inv_2 _4868_ (.Y(_0719_),
    .A(net2045));
 sg13g2_inv_1 _4869_ (.Y(_0720_),
    .A(_0124_));
 sg13g2_inv_1 _4870_ (.Y(_0721_),
    .A(_0130_));
 sg13g2_inv_1 _4871_ (.Y(_0722_),
    .A(_0132_));
 sg13g2_inv_1 _4872_ (.Y(_0723_),
    .A(_0131_));
 sg13g2_inv_1 _4873_ (.Y(_0724_),
    .A(\z80.tv80s.i_tv80_core.SP[15] ));
 sg13g2_inv_1 _4874_ (.Y(_0725_),
    .A(\z80.tv80s.i_tv80_core.SP[7] ));
 sg13g2_inv_1 _4875_ (.Y(_0726_),
    .A(_0138_));
 sg13g2_inv_1 _4876_ (.Y(_0727_),
    .A(_0139_));
 sg13g2_inv_1 _4877_ (.Y(_0728_),
    .A(_0144_));
 sg13g2_inv_1 _4878_ (.Y(_0729_),
    .A(_0143_));
 sg13g2_inv_1 _4879_ (.Y(_0730_),
    .A(_0146_));
 sg13g2_inv_1 _4880_ (.Y(_0731_),
    .A(_0148_));
 sg13g2_inv_1 _4881_ (.Y(_0732_),
    .A(_0147_));
 sg13g2_inv_1 _4882_ (.Y(_0733_),
    .A(_0149_));
 sg13g2_inv_1 _4883_ (.Y(_0734_),
    .A(net619));
 sg13g2_inv_1 _4884_ (.Y(_0735_),
    .A(net518));
 sg13g2_inv_1 _4885_ (.Y(_0736_),
    .A(net2165));
 sg13g2_inv_1 _4886_ (.Y(_0737_),
    .A(_0156_));
 sg13g2_inv_1 _4887_ (.Y(_0738_),
    .A(_0158_));
 sg13g2_inv_1 _4888_ (.Y(_0739_),
    .A(_0157_));
 sg13g2_inv_2 _4889_ (.Y(_0740_),
    .A(net560));
 sg13g2_inv_1 _4890_ (.Y(_0741_),
    .A(\z80.tv80s.i_tv80_core.PC[1] ));
 sg13g2_inv_1 _4891_ (.Y(_0742_),
    .A(_0161_));
 sg13g2_inv_1 _4892_ (.Y(_0743_),
    .A(_0165_));
 sg13g2_inv_1 _4893_ (.Y(_0744_),
    .A(net622));
 sg13g2_inv_2 _4894_ (.Y(_0745_),
    .A(net583));
 sg13g2_inv_1 _4895_ (.Y(_0746_),
    .A(\z80.tv80s.i_tv80_core.PC[12] ));
 sg13g2_inv_2 _4896_ (.Y(_0747_),
    .A(\z80.tv80s.i_tv80_core.PC[13] ));
 sg13g2_inv_1 _4897_ (.Y(_0748_),
    .A(\z80.tv80s.i_tv80_core.PC[14] ));
 sg13g2_inv_1 _4898_ (.Y(_0749_),
    .A(net632));
 sg13g2_inv_2 _4899_ (.Y(_0750_),
    .A(net590));
 sg13g2_inv_1 _4900_ (.Y(_0751_),
    .A(net628));
 sg13g2_inv_2 _4901_ (.Y(_0752_),
    .A(net481));
 sg13g2_inv_1 _4902_ (.Y(_0753_),
    .A(\z80.mreq_n ));
 sg13g2_inv_1 _4903_ (.Y(_0754_),
    .A(\z80.iorq_n ));
 sg13g2_inv_1 _4904_ (.Y(_0755_),
    .A(\z80.rd_n ));
 sg13g2_inv_1 _4905_ (.Y(_0756_),
    .A(\z80.tv80s.wr_n ));
 sg13g2_inv_1 _4906_ (.Y(_0757_),
    .A(\z80.rfsh_n ));
 sg13g2_inv_2 _4907_ (.Y(_0758_),
    .A(net500));
 sg13g2_inv_1 _4908_ (.Y(_0759_),
    .A(_0168_));
 sg13g2_inv_1 _4909_ (.Y(_0760_),
    .A(net2179));
 sg13g2_inv_2 _4910_ (.Y(_0761_),
    .A(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sg13g2_inv_1 _4911_ (.Y(_0762_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sg13g2_inv_1 _4912_ (.Y(_0763_),
    .A(net2134));
 sg13g2_inv_1 _4913_ (.Y(_0764_),
    .A(_0175_));
 sg13g2_inv_1 _4914_ (.Y(_0765_),
    .A(_0177_));
 sg13g2_inv_1 _4915_ (.Y(_0766_),
    .A(_0180_));
 sg13g2_inv_1 _4916_ (.Y(_0767_),
    .A(_0186_));
 sg13g2_inv_1 _4917_ (.Y(_0768_),
    .A(net507));
 sg13g2_inv_1 _4918_ (.Y(_0769_),
    .A(_0192_));
 sg13g2_inv_1 _4919_ (.Y(_0770_),
    .A(_0194_));
 sg13g2_inv_1 _4920_ (.Y(_0771_),
    .A(_0196_));
 sg13g2_inv_1 _4921_ (.Y(_0772_),
    .A(net540));
 sg13g2_inv_1 _4922_ (.Y(_0773_),
    .A(_0200_));
 sg13g2_inv_1 _4923_ (.Y(_0774_),
    .A(net537));
 sg13g2_inv_1 _4924_ (.Y(_0775_),
    .A(net550));
 sg13g2_inv_1 _4925_ (.Y(_0776_),
    .A(_0205_));
 sg13g2_inv_1 _4926_ (.Y(_0777_),
    .A(_0207_));
 sg13g2_inv_2 _4927_ (.Y(_0778_),
    .A(net2035));
 sg13g2_inv_2 _4928_ (.Y(_0779_),
    .A(net2036));
 sg13g2_inv_2 _4929_ (.Y(_0780_),
    .A(net2038));
 sg13g2_inv_4 _4930_ (.A(_0210_),
    .Y(_0781_));
 sg13g2_inv_2 _4931_ (.Y(_0782_),
    .A(net592));
 sg13g2_inv_2 _4932_ (.Y(_0783_),
    .A(\z80.tv80s.i_tv80_core.BusA[3] ));
 sg13g2_inv_1 _4933_ (.Y(_0784_),
    .A(\z80.tv80s.i_tv80_core.BusB[2] ));
 sg13g2_inv_1 _4934_ (.Y(_0785_),
    .A(\z80.tv80s.i_tv80_core.BusB[4] ));
 sg13g2_inv_1 _4935_ (.Y(_0786_),
    .A(\z80.tv80s.i_tv80_core.BusB[5] ));
 sg13g2_inv_1 _4936_ (.Y(_0787_),
    .A(\z80.tv80s.i_tv80_core.BusB[6] ));
 sg13g2_inv_1 _4937_ (.Y(_0788_),
    .A(\z80.tv80s.i_tv80_core.BusB[7] ));
 sg13g2_inv_1 _4938_ (.Y(_0789_),
    .A(_0225_));
 sg13g2_inv_1 _4939_ (.Y(_0790_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ));
 sg13g2_inv_1 _4940_ (.Y(_0791_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ));
 sg13g2_inv_1 _4941_ (.Y(_0792_),
    .A(net465));
 sg13g2_inv_1 _4942_ (.Y(_0793_),
    .A(net475));
 sg13g2_inv_1 _4943_ (.Y(_0794_),
    .A(net12));
 sg13g2_inv_1 _4944_ (.Y(_0795_),
    .A(net505));
 sg13g2_inv_1 _4945_ (.Y(_0796_),
    .A(net495));
 sg13g2_inv_1 _4946_ (.Y(_0797_),
    .A(net498));
 sg13g2_inv_1 _4947_ (.Y(_0798_),
    .A(_0229_));
 sg13g2_inv_1 _4948_ (.Y(_0799_),
    .A(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sg13g2_inv_2 _4949_ (.Y(_0800_),
    .A(net530));
 sg13g2_inv_1 _4950_ (.Y(_0801_),
    .A(\z80.tv80s.i_tv80_core.Fp[4] ));
 sg13g2_inv_1 _4951_ (.Y(_0802_),
    .A(\z80.tv80s.i_tv80_core.Fp[7] ));
 sg13g2_inv_1 _4952_ (.Y(_0803_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[9] ));
 sg13g2_inv_1 _4953_ (.Y(_0804_),
    .A(_0236_));
 sg13g2_inv_1 _4954_ (.Y(_0805_),
    .A(_0238_));
 sg13g2_inv_1 _4955_ (.Y(_0806_),
    .A(net478));
 sg13g2_nor2_2 _4956_ (.A(\z80.tv80s.i_tv80_core.ts[1] ),
    .B(\z80.tv80s.i_tv80_core.ts[2] ),
    .Y(_0807_));
 sg13g2_a21oi_2 _4957_ (.B1(net2020),
    .Y(_0808_),
    .A2(_0807_),
    .A1(_0023_));
 sg13g2_a21o_1 _4958_ (.A2(_0807_),
    .A1(_0023_),
    .B1(net2020),
    .X(_0809_));
 sg13g2_nand2_2 _4959_ (.Y(_0810_),
    .A(net2094),
    .B(net2098));
 sg13g2_nor2b_1 _4960_ (.A(net2089),
    .B_N(net2086),
    .Y(_0811_));
 sg13g2_nand2b_1 _4961_ (.Y(_0812_),
    .B(net2084),
    .A_N(net2090));
 sg13g2_and2_1 _4962_ (.A(net2055),
    .B(net2058),
    .X(_0813_));
 sg13g2_nand2_1 _4963_ (.Y(_0814_),
    .A(net2055),
    .B(net2058));
 sg13g2_nor2_2 _4964_ (.A(net2071),
    .B(net2062),
    .Y(_0815_));
 sg13g2_or2_2 _4965_ (.X(_0816_),
    .B(net2065),
    .A(net2073));
 sg13g2_nor2_1 _4966_ (.A(net1998),
    .B(_0816_),
    .Y(_0817_));
 sg13g2_nor4_2 _4967_ (.A(net2005),
    .B(net2003),
    .C(net1999),
    .Y(_0818_),
    .D(_0816_));
 sg13g2_a21o_1 _4968_ (.A2(_0818_),
    .A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B1(net1913),
    .X(_0819_));
 sg13g2_and2_2 _4969_ (.A(\z80.tv80s.i_tv80_core.ts[2] ),
    .B(net1),
    .X(_0820_));
 sg13g2_nand2_2 _4970_ (.Y(_0821_),
    .A(\z80.tv80s.i_tv80_core.ts[2] ),
    .B(net1));
 sg13g2_nor2_2 _4971_ (.A(net2182),
    .B(\z80.tv80s.i_tv80_core.BusAck ),
    .Y(_0822_));
 sg13g2_nand2b_2 _4972_ (.Y(_0823_),
    .B(net2227),
    .A_N(\z80.tv80s.i_tv80_core.BusAck ));
 sg13g2_nand2_1 _4973_ (.Y(_0824_),
    .A(net2229),
    .B(_0820_));
 sg13g2_nand2_1 _4974_ (.Y(_0825_),
    .A(net1901),
    .B(net1995));
 sg13g2_a21oi_2 _4975_ (.B1(net1981),
    .Y(_0826_),
    .A2(_0821_),
    .A1(net1913));
 sg13g2_nor2b_1 _4976_ (.A(net2094),
    .B_N(net2090),
    .Y(_0827_));
 sg13g2_and4_2 _4977_ (.A(net2098),
    .B(net2084),
    .C(net2002),
    .D(_0827_),
    .X(_0828_));
 sg13g2_nand2b_1 _4978_ (.Y(_0829_),
    .B(net2099),
    .A_N(net2095));
 sg13g2_nand2_2 _4979_ (.Y(_0830_),
    .A(net2090),
    .B(net2084));
 sg13g2_nand2_2 _4980_ (.Y(_0831_),
    .A(net2074),
    .B(_0828_));
 sg13g2_nand3_1 _4981_ (.B(_0826_),
    .C(_0831_),
    .A(_0819_),
    .Y(_0832_));
 sg13g2_nor2_2 _4982_ (.A(net2020),
    .B(net1997),
    .Y(_0833_));
 sg13g2_nor3_2 _4983_ (.A(net2020),
    .B(net1997),
    .C(net1980),
    .Y(_0834_));
 sg13g2_nand2_2 _4984_ (.Y(_0835_),
    .A(net1995),
    .B(_0833_));
 sg13g2_nand2b_1 _4985_ (.Y(_0836_),
    .B(_0831_),
    .A_N(_0818_));
 sg13g2_nand2_1 _4986_ (.Y(_0837_),
    .A(net2168),
    .B(_0836_));
 sg13g2_nor2b_2 _4987_ (.A(net2070),
    .B_N(net2062),
    .Y(_0838_));
 sg13g2_nand2b_1 _4988_ (.Y(_0839_),
    .B(net2064),
    .A_N(net2074));
 sg13g2_nor2_2 _4989_ (.A(net1998),
    .B(net1956),
    .Y(_0840_));
 sg13g2_nor4_2 _4990_ (.A(net2000),
    .B(_0815_),
    .C(net1958),
    .Y(_0841_),
    .D(_0830_));
 sg13g2_nand2_1 _4991_ (.Y(_0842_),
    .A(net2168),
    .B(_0841_));
 sg13g2_o21ai_1 _4992_ (.B1(net2168),
    .Y(_0843_),
    .A1(_0836_),
    .A2(_0841_));
 sg13g2_or4_1 _4993_ (.A(net2166),
    .B(net526),
    .C(net258),
    .D(_0843_),
    .X(_0844_));
 sg13g2_a22oi_1 _4994_ (.Y(_0296_),
    .B1(_0834_),
    .B2(_0844_),
    .A2(_0832_),
    .A1(net2172));
 sg13g2_nor2_1 _4995_ (.A(net2166),
    .B(net2168),
    .Y(_0845_));
 sg13g2_nand2_1 _4996_ (.Y(_0846_),
    .A(_0675_),
    .B(net2015));
 sg13g2_nor2b_1 _4997_ (.A(net2056),
    .B_N(net2059),
    .Y(_0847_));
 sg13g2_nand2b_1 _4998_ (.Y(_0848_),
    .B(net2059),
    .A_N(net2056));
 sg13g2_and3_2 _4999_ (.X(_0849_),
    .A(net2096),
    .B(net2100),
    .C(net2089));
 sg13g2_nand3_1 _5000_ (.B(net2098),
    .C(net2090),
    .A(net2094),
    .Y(_0850_));
 sg13g2_nand2_2 _5001_ (.Y(_0851_),
    .A(net1951),
    .B(_0849_));
 sg13g2_nor2_2 _5002_ (.A(net2104),
    .B(net2125),
    .Y(_0852_));
 sg13g2_nand2_1 _5003_ (.Y(_0853_),
    .A(net2026),
    .B(net2018));
 sg13g2_o21ai_1 _5004_ (.B1(_0852_),
    .Y(_0854_),
    .A1(net2068),
    .A2(_0851_));
 sg13g2_nor2b_2 _5005_ (.A(net2098),
    .B_N(net2095),
    .Y(_0855_));
 sg13g2_nand2b_2 _5006_ (.Y(_0856_),
    .B(net2095),
    .A_N(net2099));
 sg13g2_nor2_2 _5007_ (.A(net2091),
    .B(net1948),
    .Y(_0857_));
 sg13g2_nand2_2 _5008_ (.Y(_0858_),
    .A(_0671_),
    .B(_0855_));
 sg13g2_nor2_2 _5009_ (.A(net1949),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_nand2_2 _5010_ (.Y(_0860_),
    .A(net1951),
    .B(_0857_));
 sg13g2_nor2_2 _5011_ (.A(net2117),
    .B(net2124),
    .Y(_0861_));
 sg13g2_or2_1 _5012_ (.X(_0862_),
    .B(net2126),
    .A(net2115));
 sg13g2_nor2b_2 _5013_ (.A(net2059),
    .B_N(net2056),
    .Y(_0863_));
 sg13g2_nand2b_2 _5014_ (.Y(_0864_),
    .B(net2056),
    .A_N(net2059));
 sg13g2_and2_2 _5015_ (.A(net2066),
    .B(_0863_),
    .X(_0865_));
 sg13g2_nand2_1 _5016_ (.Y(_0866_),
    .A(net2065),
    .B(_0863_));
 sg13g2_nand3b_1 _5017_ (.B(net2098),
    .C(net2094),
    .Y(_0867_),
    .A_N(net2090));
 sg13g2_nor2_2 _5018_ (.A(net1890),
    .B(net1945),
    .Y(_0868_));
 sg13g2_nor2_1 _5019_ (.A(net2122),
    .B(net2110),
    .Y(_0869_));
 sg13g2_or2_2 _5020_ (.X(_0870_),
    .B(net2109),
    .A(net2114));
 sg13g2_nand2_1 _5021_ (.Y(_0871_),
    .A(net2014),
    .B(net2108));
 sg13g2_nand2_2 _5022_ (.Y(_0872_),
    .A(net2107),
    .B(net1942));
 sg13g2_inv_2 _5023_ (.Y(_0873_),
    .A(_0872_));
 sg13g2_nor2_1 _5024_ (.A(net2126),
    .B(_0873_),
    .Y(_0874_));
 sg13g2_o21ai_1 _5025_ (.B1(_0868_),
    .Y(_0875_),
    .A1(net2124),
    .A2(_0873_));
 sg13g2_o21ai_1 _5026_ (.B1(_0875_),
    .Y(_0876_),
    .A1(_0860_),
    .A2(_0861_));
 sg13g2_nor2_2 _5027_ (.A(_0858_),
    .B(net1890),
    .Y(_0877_));
 sg13g2_nor2_1 _5028_ (.A(net2097),
    .B(net2093),
    .Y(_0878_));
 sg13g2_and2_2 _5029_ (.A(_0865_),
    .B(_0878_),
    .X(_0879_));
 sg13g2_nor2_2 _5030_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .B(net2108),
    .Y(_0880_));
 sg13g2_nor2_1 _5031_ (.A(net2119),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_o21ai_1 _5032_ (.B1(net2018),
    .Y(_0882_),
    .A1(net2116),
    .A2(_0880_));
 sg13g2_o21ai_1 _5033_ (.B1(_0882_),
    .Y(_0883_),
    .A1(_0877_),
    .A2(_0879_));
 sg13g2_nor2_2 _5034_ (.A(net1956),
    .B(_0851_),
    .Y(_0884_));
 sg13g2_nand3_1 _5035_ (.B(_0847_),
    .C(_0849_),
    .A(_0838_),
    .Y(_0885_));
 sg13g2_nor2_1 _5036_ (.A(net2121),
    .B(net2014),
    .Y(_0886_));
 sg13g2_nand2b_2 _5037_ (.Y(_0887_),
    .B(net2109),
    .A_N(net2120));
 sg13g2_nor2_2 _5038_ (.A(net2128),
    .B(net1889),
    .Y(_0888_));
 sg13g2_nor2_1 _5039_ (.A(_0885_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_nor3_1 _5040_ (.A(_0854_),
    .B(_0876_),
    .C(_0889_),
    .Y(_0890_));
 sg13g2_a22oi_1 _5041_ (.Y(_0891_),
    .B1(_0883_),
    .B2(_0890_),
    .A2(net1892),
    .A1(net2025));
 sg13g2_nor2_1 _5042_ (.A(net2055),
    .B(net2058),
    .Y(_0892_));
 sg13g2_or2_1 _5043_ (.X(_0893_),
    .B(net2059),
    .A(net2056));
 sg13g2_nor4_2 _5044_ (.A(net2074),
    .B(net2064),
    .C(net2055),
    .Y(_0894_),
    .D(net2058));
 sg13g2_or4_2 _5045_ (.A(net2073),
    .B(net2065),
    .C(net2055),
    .D(net2058),
    .X(_0895_));
 sg13g2_nand3_1 _5046_ (.B(_0855_),
    .C(_0894_),
    .A(_0671_),
    .Y(_0896_));
 sg13g2_and2_1 _5047_ (.A(net2071),
    .B(net2063),
    .X(_0897_));
 sg13g2_nand2_1 _5048_ (.Y(_0898_),
    .A(net2073),
    .B(net2065));
 sg13g2_and2_2 _5049_ (.A(net2064),
    .B(net1940),
    .X(_0899_));
 sg13g2_nor2_2 _5050_ (.A(net1939),
    .B(net1934),
    .Y(_0900_));
 sg13g2_nor2_1 _5051_ (.A(net2004),
    .B(net1948),
    .Y(_0901_));
 sg13g2_and2_1 _5052_ (.A(_0900_),
    .B(_0901_),
    .X(_0902_));
 sg13g2_nand4_1 _5053_ (.B(_0855_),
    .C(net1940),
    .A(_0811_),
    .Y(_0903_),
    .D(net1935));
 sg13g2_nor2b_2 _5054_ (.A(net2064),
    .B_N(net2074),
    .Y(_0904_));
 sg13g2_nand2b_1 _5055_ (.Y(_0905_),
    .B(net2073),
    .A_N(net2067));
 sg13g2_nor2_2 _5056_ (.A(net1938),
    .B(net1931),
    .Y(_0906_));
 sg13g2_nand2_1 _5057_ (.Y(_0907_),
    .A(net1941),
    .B(_0904_));
 sg13g2_nand4_1 _5058_ (.B(_0855_),
    .C(net1940),
    .A(_0811_),
    .Y(_0908_),
    .D(_0904_));
 sg13g2_and2_1 _5059_ (.A(_0903_),
    .B(_0908_),
    .X(_0909_));
 sg13g2_and3_1 _5060_ (.X(_0910_),
    .A(_0896_),
    .B(_0903_),
    .C(_0908_));
 sg13g2_nand3_1 _5061_ (.B(_0903_),
    .C(_0908_),
    .A(_0896_),
    .Y(_0911_));
 sg13g2_nor2_1 _5062_ (.A(net2089),
    .B(net2086),
    .Y(_0912_));
 sg13g2_or2_2 _5063_ (.X(_0913_),
    .B(net2085),
    .A(net2091));
 sg13g2_nor2_1 _5064_ (.A(net1948),
    .B(_0913_),
    .Y(_0914_));
 sg13g2_nor4_2 _5065_ (.A(_0856_),
    .B(net1939),
    .C(net1933),
    .Y(_0915_),
    .D(_0913_));
 sg13g2_nand4_1 _5066_ (.B(net1940),
    .C(net1935),
    .A(_0855_),
    .Y(_0916_),
    .D(_0912_));
 sg13g2_nand4_1 _5067_ (.B(net1940),
    .C(_0904_),
    .A(_0855_),
    .Y(_0917_),
    .D(_0912_));
 sg13g2_nor2_1 _5068_ (.A(net1957),
    .B(_0913_),
    .Y(_0918_));
 sg13g2_nand2_1 _5069_ (.Y(_0919_),
    .A(_0899_),
    .B(_0918_));
 sg13g2_a221oi_1 _5070_ (.B2(_0899_),
    .C1(_0915_),
    .B1(_0918_),
    .A1(_0906_),
    .Y(_0920_),
    .A2(_0914_));
 sg13g2_nand3_1 _5071_ (.B(_0917_),
    .C(_0919_),
    .A(_0916_),
    .Y(_0921_));
 sg13g2_nor2_1 _5072_ (.A(_0911_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_nor4_2 _5073_ (.A(net2064),
    .B(net1957),
    .C(net1938),
    .Y(_0923_),
    .D(_0913_));
 sg13g2_nand2_2 _5074_ (.Y(_0924_),
    .A(_0857_),
    .B(_0899_));
 sg13g2_nor2_2 _5075_ (.A(net1955),
    .B(net1938),
    .Y(_0925_));
 sg13g2_nor4_2 _5076_ (.A(net2091),
    .B(net1955),
    .C(net1948),
    .Y(_0926_),
    .D(net1937));
 sg13g2_nand2_2 _5077_ (.Y(_0927_),
    .A(_0857_),
    .B(_0925_));
 sg13g2_nor2_2 _5078_ (.A(_0923_),
    .B(_0926_),
    .Y(_0928_));
 sg13g2_nand3b_1 _5079_ (.B(_0233_),
    .C(net2089),
    .Y(_0929_),
    .A_N(net2058));
 sg13g2_nor2_2 _5080_ (.A(net1948),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_or2_2 _5081_ (.X(_0931_),
    .B(_0929_),
    .A(net1948));
 sg13g2_nor4_2 _5082_ (.A(_0810_),
    .B(net2003),
    .C(net1998),
    .Y(_0932_),
    .D(net1955));
 sg13g2_nor3_2 _5083_ (.A(net2000),
    .B(_0829_),
    .C(_0913_),
    .Y(_0933_));
 sg13g2_nand2_2 _5084_ (.Y(_0934_),
    .A(net2002),
    .B(net1888));
 sg13g2_nor4_1 _5085_ (.A(net1951),
    .B(_0930_),
    .C(_0932_),
    .D(_0933_),
    .Y(_0935_));
 sg13g2_nand4_1 _5086_ (.B(_0916_),
    .C(_0917_),
    .A(net1950),
    .Y(_0936_),
    .D(_0931_));
 sg13g2_nand4_1 _5087_ (.B(_0920_),
    .C(_0928_),
    .A(_0910_),
    .Y(_0937_),
    .D(_0935_));
 sg13g2_nand2b_1 _5088_ (.Y(_0938_),
    .B(net2090),
    .A_N(net2083));
 sg13g2_nor2_2 _5089_ (.A(_0810_),
    .B(net1930),
    .Y(_0939_));
 sg13g2_or2_1 _5090_ (.X(_0940_),
    .B(net1930),
    .A(net2005));
 sg13g2_nor4_2 _5091_ (.A(net2005),
    .B(net1937),
    .C(net1931),
    .Y(_0941_),
    .D(net1929));
 sg13g2_and4_2 _5092_ (.A(net2094),
    .B(net2098),
    .C(net2090),
    .D(net2083),
    .X(_0942_));
 sg13g2_nand4_1 _5093_ (.B(net2098),
    .C(net2090),
    .A(net2094),
    .Y(_0943_),
    .D(net2084));
 sg13g2_nor2_1 _5094_ (.A(_0895_),
    .B(_0943_),
    .Y(_0944_));
 sg13g2_nor3_2 _5095_ (.A(net2005),
    .B(_0895_),
    .C(net1929),
    .Y(_0945_));
 sg13g2_a22oi_1 _5096_ (.Y(_0946_),
    .B1(_0940_),
    .B2(_0943_),
    .A2(_0907_),
    .A1(_0895_));
 sg13g2_nor3_2 _5097_ (.A(_0850_),
    .B(net1937),
    .C(net1933),
    .Y(_0947_));
 sg13g2_nor2_1 _5098_ (.A(net1999),
    .B(net1933),
    .Y(_0948_));
 sg13g2_nand4_1 _5099_ (.B(net2064),
    .C(net2055),
    .A(net2073),
    .Y(_0949_),
    .D(net2058));
 sg13g2_nor2_2 _5100_ (.A(net1944),
    .B(_0949_),
    .Y(_0950_));
 sg13g2_nor2_1 _5101_ (.A(_0947_),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_or2_1 _5102_ (.X(_0952_),
    .B(_0950_),
    .A(_0947_));
 sg13g2_nor2_1 _5103_ (.A(_0946_),
    .B(_0952_),
    .Y(_0953_));
 sg13g2_nor2_1 _5104_ (.A(_0671_),
    .B(net1948),
    .Y(_0954_));
 sg13g2_nand2_2 _5105_ (.Y(_0955_),
    .A(net2091),
    .B(_0855_));
 sg13g2_nand2_1 _5106_ (.Y(_0956_),
    .A(net2057),
    .B(net1886));
 sg13g2_a21oi_1 _5107_ (.A1(net2055),
    .A2(net1887),
    .Y(_0957_),
    .B1(_0863_));
 sg13g2_nor2_1 _5108_ (.A(net2000),
    .B(net1932),
    .Y(_0958_));
 sg13g2_nor3_2 _5109_ (.A(net2001),
    .B(net1944),
    .C(net1932),
    .Y(_0959_));
 sg13g2_nor2_1 _5110_ (.A(net2004),
    .B(net1957),
    .Y(_0960_));
 sg13g2_nor4_2 _5111_ (.A(net2003),
    .B(net1999),
    .C(net1958),
    .Y(_0961_),
    .D(net1931));
 sg13g2_nor2_1 _5112_ (.A(net2096),
    .B(net2100),
    .Y(_0962_));
 sg13g2_or2_2 _5113_ (.X(_0963_),
    .B(net2098),
    .A(net2094));
 sg13g2_nor3_2 _5114_ (.A(net2003),
    .B(_0895_),
    .C(_0963_),
    .Y(_0964_));
 sg13g2_nor2_1 _5115_ (.A(_0961_),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_or2_1 _5116_ (.X(_0966_),
    .B(_0964_),
    .A(_0961_));
 sg13g2_nor2_2 _5117_ (.A(net2082),
    .B(net1944),
    .Y(_0967_));
 sg13g2_nor4_2 _5118_ (.A(net2082),
    .B(net2001),
    .C(_0816_),
    .Y(_0968_),
    .D(net1944));
 sg13g2_nand2_2 _5119_ (.Y(_0969_),
    .A(_0817_),
    .B(_0967_));
 sg13g2_nor3_2 _5120_ (.A(net2089),
    .B(net2001),
    .C(net1948),
    .Y(_0970_));
 sg13g2_or2_2 _5121_ (.X(_0971_),
    .B(_0970_),
    .A(_0968_));
 sg13g2_nor4_2 _5122_ (.A(net2003),
    .B(net1999),
    .C(net1958),
    .Y(_0972_),
    .D(net1955));
 sg13g2_nor2_1 _5123_ (.A(_0841_),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_nor3_2 _5124_ (.A(net1955),
    .B(_0850_),
    .C(net1937),
    .Y(_0974_));
 sg13g2_nand2_1 _5125_ (.Y(_0975_),
    .A(_0849_),
    .B(_0925_));
 sg13g2_nor3_2 _5126_ (.A(_0818_),
    .B(_0947_),
    .C(_0974_),
    .Y(_0976_));
 sg13g2_nand4_1 _5127_ (.B(_0965_),
    .C(_0973_),
    .A(_0957_),
    .Y(_0977_),
    .D(_0976_));
 sg13g2_or4_2 _5128_ (.A(_0946_),
    .B(_0952_),
    .C(_0959_),
    .D(_0971_),
    .X(_0978_));
 sg13g2_nor2_1 _5129_ (.A(net2094),
    .B(net1930),
    .Y(_0979_));
 sg13g2_nor2_1 _5130_ (.A(net1957),
    .B(net1929),
    .Y(_0980_));
 sg13g2_nor3_2 _5131_ (.A(net2000),
    .B(net1958),
    .C(net1930),
    .Y(_0981_));
 sg13g2_nor2_2 _5132_ (.A(net1999),
    .B(_0850_),
    .Y(_0982_));
 sg13g2_nand2_2 _5133_ (.Y(_0983_),
    .A(net2002),
    .B(_0849_));
 sg13g2_nand2b_2 _5134_ (.Y(_0984_),
    .B(_0983_),
    .A_N(_0981_));
 sg13g2_nor3_2 _5135_ (.A(net2096),
    .B(net2099),
    .C(net2091),
    .Y(_0985_));
 sg13g2_or3_2 _5136_ (.A(net2095),
    .B(net2099),
    .C(net2092),
    .X(_0986_));
 sg13g2_nand2_1 _5137_ (.Y(_0987_),
    .A(net2002),
    .B(_0985_));
 sg13g2_nor2_1 _5138_ (.A(net2065),
    .B(net2000),
    .Y(_0988_));
 sg13g2_nor4_2 _5139_ (.A(net2004),
    .B(net2000),
    .C(_0816_),
    .Y(_0989_),
    .D(net1958));
 sg13g2_nor2_2 _5140_ (.A(net2083),
    .B(_0986_),
    .Y(_0990_));
 sg13g2_a221oi_1 _5141_ (.B2(_0840_),
    .C1(_0989_),
    .B1(_0990_),
    .A1(_0985_),
    .Y(_0991_),
    .A2(_0988_));
 sg13g2_nor3_2 _5142_ (.A(net2003),
    .B(_0949_),
    .C(_0963_),
    .Y(_0992_));
 sg13g2_nor4_2 _5143_ (.A(net2003),
    .B(net1998),
    .C(net1955),
    .Y(_0993_),
    .D(_0963_));
 sg13g2_nor3_1 _5144_ (.A(net2083),
    .B(_0949_),
    .C(_0986_),
    .Y(_0994_));
 sg13g2_nor2_1 _5145_ (.A(_0993_),
    .B(_0994_),
    .Y(_0995_));
 sg13g2_nor3_2 _5146_ (.A(_0992_),
    .B(_0993_),
    .C(_0994_),
    .Y(_0996_));
 sg13g2_nand2_1 _5147_ (.Y(_0997_),
    .A(_0991_),
    .B(_0995_));
 sg13g2_and2_2 _5148_ (.A(_0991_),
    .B(_0996_),
    .X(_0998_));
 sg13g2_nand3b_1 _5149_ (.B(_0991_),
    .C(_0996_),
    .Y(_0999_),
    .A_N(_0984_));
 sg13g2_nor4_2 _5150_ (.A(_0937_),
    .B(_0977_),
    .C(_0978_),
    .Y(_1000_),
    .D(_0999_));
 sg13g2_nor3_2 _5151_ (.A(net2083),
    .B(_0895_),
    .C(_0986_),
    .Y(_1001_));
 sg13g2_nand2_2 _5152_ (.Y(_1002_),
    .A(_0894_),
    .B(_0990_));
 sg13g2_nor4_2 _5153_ (.A(net2000),
    .B(_0816_),
    .C(net1958),
    .Y(_1003_),
    .D(_0830_));
 sg13g2_nand2_2 _5154_ (.Y(_1004_),
    .A(_0815_),
    .B(_0828_));
 sg13g2_nor3_2 _5155_ (.A(_0671_),
    .B(net2001),
    .C(net1928),
    .Y(_1005_));
 sg13g2_nand3_1 _5156_ (.B(net2002),
    .C(_0962_),
    .A(net2089),
    .Y(_1006_));
 sg13g2_nand3_1 _5157_ (.B(_1004_),
    .C(_1006_),
    .A(_1002_),
    .Y(_1007_));
 sg13g2_nor2_2 _5158_ (.A(net2096),
    .B(_0929_),
    .Y(_1008_));
 sg13g2_or2_1 _5159_ (.X(_1009_),
    .B(_0929_),
    .A(net2097));
 sg13g2_nand4_1 _5160_ (.B(_1004_),
    .C(_1006_),
    .A(_1002_),
    .Y(_1010_),
    .D(_1009_));
 sg13g2_nor4_2 _5161_ (.A(net2083),
    .B(net1939),
    .C(net1932),
    .Y(_1011_),
    .D(_0986_));
 sg13g2_nand2_2 _5162_ (.Y(_1012_),
    .A(_0906_),
    .B(_0990_));
 sg13g2_nor3_2 _5163_ (.A(net2004),
    .B(net1957),
    .C(net1939),
    .Y(_1013_));
 sg13g2_nand2_2 _5164_ (.Y(_1014_),
    .A(net1941),
    .B(_0960_));
 sg13g2_nor2_2 _5165_ (.A(_1011_),
    .B(net1882),
    .Y(_1015_));
 sg13g2_nand2_1 _5166_ (.Y(_1016_),
    .A(_1012_),
    .B(_1014_));
 sg13g2_nor4_2 _5167_ (.A(net2004),
    .B(net1937),
    .C(net1931),
    .Y(_1017_),
    .D(net1928));
 sg13g2_and3_2 _5168_ (.X(_1018_),
    .A(net2066),
    .B(net1940),
    .C(_0985_));
 sg13g2_or2_2 _5169_ (.X(_1019_),
    .B(_1018_),
    .A(_1017_));
 sg13g2_nor2_1 _5170_ (.A(net1945),
    .B(net1937),
    .Y(_1020_));
 sg13g2_nor3_2 _5171_ (.A(net2003),
    .B(net1958),
    .C(_0949_),
    .Y(_1021_));
 sg13g2_nor2_2 _5172_ (.A(net1881),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_nand2_1 _5173_ (.Y(_1023_),
    .A(_1015_),
    .B(_1022_));
 sg13g2_nor3_2 _5174_ (.A(_1010_),
    .B(_1019_),
    .C(_1023_),
    .Y(_1024_));
 sg13g2_nor4_1 _5175_ (.A(_0937_),
    .B(_0977_),
    .C(_0978_),
    .D(_1019_),
    .Y(_1025_));
 sg13g2_and2_2 _5176_ (.A(_1000_),
    .B(_1024_),
    .X(_1026_));
 sg13g2_nand2_1 _5177_ (.Y(_1027_),
    .A(_0888_),
    .B(_1026_));
 sg13g2_nand2b_1 _5178_ (.Y(_1028_),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .A_N(net2108));
 sg13g2_nor2_1 _5179_ (.A(net2114),
    .B(_1028_),
    .Y(_1029_));
 sg13g2_nor2_1 _5180_ (.A(_1027_),
    .B(_1029_),
    .Y(_1030_));
 sg13g2_nor2_1 _5181_ (.A(net2128),
    .B(_1000_),
    .Y(_1031_));
 sg13g2_nand2_1 _5182_ (.Y(_1032_),
    .A(_0888_),
    .B(_1003_));
 sg13g2_nor2_1 _5183_ (.A(net2081),
    .B(net2021),
    .Y(_1033_));
 sg13g2_nand2b_2 _5184_ (.Y(_1034_),
    .B(net2070),
    .A_N(net2078));
 sg13g2_nand3b_1 _5185_ (.B(net2071),
    .C(net2060),
    .Y(_1035_),
    .A_N(net2077));
 sg13g2_nor2_1 _5186_ (.A(net2151),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_nor2_1 _5187_ (.A(net2024),
    .B(net2070),
    .Y(_1037_));
 sg13g2_nand2b_2 _5188_ (.Y(_1038_),
    .B(net2078),
    .A_N(net2070));
 sg13g2_nor3_1 _5189_ (.A(_0662_),
    .B(net2062),
    .C(_1038_),
    .Y(_1039_));
 sg13g2_nor2_1 _5190_ (.A(net2024),
    .B(net2021),
    .Y(_1040_));
 sg13g2_nand2_2 _5191_ (.Y(_1041_),
    .A(net2078),
    .B(net2070));
 sg13g2_nand2_1 _5192_ (.Y(_1042_),
    .A(net2060),
    .B(net1878));
 sg13g2_nor3_1 _5193_ (.A(_0665_),
    .B(_0678_),
    .C(_1041_),
    .Y(_1043_));
 sg13g2_nand2_2 _5194_ (.Y(_1044_),
    .A(net2077),
    .B(_0838_));
 sg13g2_and3_1 _5195_ (.X(_1045_),
    .A(net2147),
    .B(net2077),
    .C(_0838_));
 sg13g2_nor2_1 _5196_ (.A(net2061),
    .B(_1034_),
    .Y(_1046_));
 sg13g2_nand2_2 _5197_ (.Y(_1047_),
    .A(_0678_),
    .B(net1879));
 sg13g2_nor3_1 _5198_ (.A(\z80.tv80s.i_tv80_core.F[7] ),
    .B(net2060),
    .C(_1034_),
    .Y(_1048_));
 sg13g2_nor3_1 _5199_ (.A(_0661_),
    .B(net2060),
    .C(_1041_),
    .Y(_1049_));
 sg13g2_nor2_2 _5200_ (.A(net2077),
    .B(net2070),
    .Y(_1050_));
 sg13g2_or2_2 _5201_ (.X(_1051_),
    .B(net2070),
    .A(net2077));
 sg13g2_nor2_1 _5202_ (.A(_0678_),
    .B(_1051_),
    .Y(_1052_));
 sg13g2_nor4_1 _5203_ (.A(_1043_),
    .B(_1045_),
    .C(_1049_),
    .D(_1052_),
    .Y(_1053_));
 sg13g2_nand2_1 _5204_ (.Y(_1054_),
    .A(_0678_),
    .B(_1050_));
 sg13g2_nor3_1 _5205_ (.A(net2147),
    .B(net2060),
    .C(_1051_),
    .Y(_1055_));
 sg13g2_nor4_1 _5206_ (.A(_1036_),
    .B(_1039_),
    .C(_1048_),
    .D(_1055_),
    .Y(_1056_));
 sg13g2_a22oi_1 _5207_ (.Y(_1057_),
    .B1(_1053_),
    .B2(_1056_),
    .A2(_1052_),
    .A1(\z80.tv80s.i_tv80_core.F[6] ));
 sg13g2_nand2_1 _5208_ (.Y(_1058_),
    .A(net1889),
    .B(_1057_));
 sg13g2_nand3_1 _5209_ (.B(net1884),
    .C(_1058_),
    .A(net2019),
    .Y(_1059_));
 sg13g2_nand2_1 _5210_ (.Y(_1060_),
    .A(_1032_),
    .B(_1059_));
 sg13g2_nor2_1 _5211_ (.A(_1011_),
    .B(_1017_),
    .Y(_1061_));
 sg13g2_nor3_2 _5212_ (.A(_1011_),
    .B(_1017_),
    .C(_1018_),
    .Y(_1062_));
 sg13g2_nand2b_1 _5213_ (.Y(_1063_),
    .B(_0888_),
    .A_N(_1062_));
 sg13g2_nor2_2 _5214_ (.A(\z80.tv80s.i_tv80_core.IntCycle ),
    .B(\z80.tv80s.i_tv80_core.NMICycle ),
    .Y(_1064_));
 sg13g2_a21oi_1 _5215_ (.A1(net2127),
    .A2(_1064_),
    .Y(_1065_),
    .B1(_1002_));
 sg13g2_nor2_1 _5216_ (.A(net2128),
    .B(_0870_),
    .Y(_1066_));
 sg13g2_o21ai_1 _5217_ (.B1(_1065_),
    .Y(_1067_),
    .A1(_1064_),
    .A2(_1066_));
 sg13g2_a21oi_1 _5218_ (.A1(net2119),
    .A2(net1875),
    .Y(_1068_),
    .B1(net2127));
 sg13g2_nand2b_1 _5219_ (.Y(_1069_),
    .B(net1882),
    .A_N(net2120));
 sg13g2_nor2_1 _5220_ (.A(net2129),
    .B(_1069_),
    .Y(_1070_));
 sg13g2_a21oi_1 _5221_ (.A1(_1008_),
    .A2(_1068_),
    .Y(_1071_),
    .B1(_1070_));
 sg13g2_nand4_1 _5222_ (.B(_1063_),
    .C(_1067_),
    .A(_1022_),
    .Y(_1072_),
    .D(_1071_));
 sg13g2_or4_1 _5223_ (.A(_1030_),
    .B(_1031_),
    .C(_1060_),
    .D(_1072_),
    .X(_1073_));
 sg13g2_nor2b_2 _5224_ (.A(net2104),
    .B_N(net2116),
    .Y(_1074_));
 sg13g2_o21ai_1 _5225_ (.B1(_1074_),
    .Y(_1075_),
    .A1(_0233_),
    .A2(net1939));
 sg13g2_o21ai_1 _5226_ (.B1(net2018),
    .Y(_1076_),
    .A1(_0955_),
    .A2(_1075_));
 sg13g2_or2_1 _5227_ (.X(_1077_),
    .B(_1076_),
    .A(_0675_));
 sg13g2_a21oi_1 _5228_ (.A1(net2168),
    .A2(_1073_),
    .Y(_1078_),
    .B1(net1952));
 sg13g2_a21oi_2 _5229_ (.B1(_0891_),
    .Y(_1079_),
    .A2(_1078_),
    .A1(_1077_));
 sg13g2_nand2_1 _5230_ (.Y(_1080_),
    .A(_1000_),
    .B(_1006_));
 sg13g2_nor2_1 _5231_ (.A(_1006_),
    .B(_1058_),
    .Y(_1081_));
 sg13g2_a21oi_1 _5232_ (.A1(_1004_),
    .A2(_1062_),
    .Y(_1082_),
    .B1(_0888_));
 sg13g2_nand2_1 _5233_ (.Y(_1083_),
    .A(net2113),
    .B(_0679_));
 sg13g2_a21oi_1 _5234_ (.A1(net2111),
    .A2(net2014),
    .Y(_1084_),
    .B1(_1064_));
 sg13g2_o21ai_1 _5235_ (.B1(_1001_),
    .Y(_1085_),
    .A1(net2128),
    .A2(_1084_));
 sg13g2_o21ai_1 _5236_ (.B1(_1085_),
    .Y(_1086_),
    .A1(net1883),
    .A2(_1068_));
 sg13g2_o21ai_1 _5237_ (.B1(_1022_),
    .Y(_1087_),
    .A1(_0861_),
    .A2(_1014_));
 sg13g2_o21ai_1 _5238_ (.B1(_1080_),
    .Y(_1088_),
    .A1(net2128),
    .A2(_1081_));
 sg13g2_nor4_1 _5239_ (.A(_1026_),
    .B(_1082_),
    .C(_1086_),
    .D(_1087_),
    .Y(_1089_));
 sg13g2_nand2_1 _5240_ (.Y(_1090_),
    .A(_1088_),
    .B(_1089_));
 sg13g2_nor2_1 _5241_ (.A(net2015),
    .B(_1030_),
    .Y(_1091_));
 sg13g2_a221oi_1 _5242_ (.B2(_1091_),
    .C1(_0891_),
    .B1(_1090_),
    .A1(net2167),
    .Y(_1092_),
    .A2(_1076_));
 sg13g2_nand2_1 _5243_ (.Y(_1093_),
    .A(_1079_),
    .B(_1092_));
 sg13g2_nor2_1 _5244_ (.A(net2127),
    .B(net1943),
    .Y(_1094_));
 sg13g2_nand2_2 _5245_ (.Y(_1095_),
    .A(net2019),
    .B(_0870_));
 sg13g2_o21ai_1 _5246_ (.B1(_1065_),
    .Y(_1096_),
    .A1(_1064_),
    .A2(_1095_));
 sg13g2_nand2_1 _5247_ (.Y(_1097_),
    .A(net1889),
    .B(_1019_));
 sg13g2_nand4_1 _5248_ (.B(_1071_),
    .C(_1096_),
    .A(_1012_),
    .Y(_1098_),
    .D(_1097_));
 sg13g2_nor3_1 _5249_ (.A(_0999_),
    .B(_1060_),
    .C(_1098_),
    .Y(_1099_));
 sg13g2_o21ai_1 _5250_ (.B1(_1099_),
    .Y(_1100_),
    .A1(net2127),
    .A2(_1025_));
 sg13g2_nand2b_1 _5251_ (.Y(_1101_),
    .B(_1027_),
    .A_N(_1100_));
 sg13g2_or2_1 _5252_ (.X(_1102_),
    .B(_0021_),
    .A(net2116));
 sg13g2_a21oi_1 _5253_ (.A1(_0877_),
    .A2(_1102_),
    .Y(_1103_),
    .B1(_0879_));
 sg13g2_nor2_2 _5254_ (.A(_0866_),
    .B(_0986_),
    .Y(_1104_));
 sg13g2_nand2_1 _5255_ (.Y(_1105_),
    .A(_0865_),
    .B(_0985_));
 sg13g2_nor2_2 _5256_ (.A(_0868_),
    .B(_0877_),
    .Y(_1106_));
 sg13g2_a21oi_2 _5257_ (.B1(net1890),
    .Y(_1107_),
    .A2(net1945),
    .A1(_0858_));
 sg13g2_nand2_1 _5258_ (.Y(_1108_),
    .A(_1105_),
    .B(_1106_));
 sg13g2_and2_1 _5259_ (.A(net2102),
    .B(_0879_),
    .X(_1109_));
 sg13g2_nand2_2 _5260_ (.Y(_1110_),
    .A(net2102),
    .B(_0879_));
 sg13g2_o21ai_1 _5261_ (.B1(_0885_),
    .Y(_1111_),
    .A1(net2093),
    .A2(net1890));
 sg13g2_nand2b_1 _5262_ (.Y(_1112_),
    .B(_0860_),
    .A_N(_1111_));
 sg13g2_a21oi_1 _5263_ (.A1(_1103_),
    .A2(_1112_),
    .Y(_1113_),
    .B1(net2124));
 sg13g2_a221oi_1 _5264_ (.B2(_0888_),
    .C1(_0868_),
    .B1(_0884_),
    .A1(_0859_),
    .Y(_1114_),
    .A2(_0861_));
 sg13g2_nand2b_1 _5265_ (.Y(_1115_),
    .B(_1114_),
    .A_N(_1113_));
 sg13g2_nor3_2 _5266_ (.A(net2069),
    .B(net1891),
    .C(_0851_),
    .Y(_1116_));
 sg13g2_nand3b_1 _5267_ (.B(_0230_),
    .C(_1077_),
    .Y(_1117_),
    .A_N(_1116_));
 sg13g2_a221oi_1 _5268_ (.B2(net1953),
    .C1(_1117_),
    .B1(_1115_),
    .A1(net2168),
    .Y(_1118_),
    .A2(_1101_));
 sg13g2_or2_1 _5269_ (.X(_1119_),
    .B(_1118_),
    .A(_1079_));
 sg13g2_nand2b_1 _5270_ (.Y(_1120_),
    .B(_1118_),
    .A_N(_1092_));
 sg13g2_nand3_1 _5271_ (.B(_1119_),
    .C(_1120_),
    .A(_1093_),
    .Y(_1121_));
 sg13g2_or2_1 _5272_ (.X(_1122_),
    .B(_1079_),
    .A(\z80.tv80s.i_tv80_core.ts[4] ));
 sg13g2_a21oi_1 _5273_ (.A1(_0029_),
    .A2(_1079_),
    .Y(_1123_),
    .B1(_1120_));
 sg13g2_nand2_1 _5274_ (.Y(_1124_),
    .A(_0031_),
    .B(_1118_));
 sg13g2_o21ai_1 _5275_ (.B1(_1124_),
    .Y(_1125_),
    .A1(net2142),
    .A2(_1118_));
 sg13g2_mux2_1 _5276_ (.A0(_0030_),
    .A1(_0032_),
    .S(_1092_),
    .X(_1126_));
 sg13g2_nor2_1 _5277_ (.A(_1119_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_a21oi_1 _5278_ (.A1(_1122_),
    .A2(_1123_),
    .Y(_1128_),
    .B1(_1127_));
 sg13g2_o21ai_1 _5279_ (.B1(_1128_),
    .Y(_1129_),
    .A1(_1093_),
    .A2(_1125_));
 sg13g2_mux2_1 _5280_ (.A0(\z80.tv80s.i_tv80_core.ts[0] ),
    .A1(_1129_),
    .S(_1121_),
    .X(_1130_));
 sg13g2_inv_4 _5281_ (.A(net1689),
    .Y(_1131_));
 sg13g2_nor2_1 _5282_ (.A(\z80.tv80s.i_tv80_core.BusReq_s ),
    .B(_1131_),
    .Y(_1132_));
 sg13g2_nand2b_2 _5283_ (.Y(_1133_),
    .B(\z80.tv80s.i_tv80_core.ts[2] ),
    .A_N(net1));
 sg13g2_and2_2 _5284_ (.A(net2227),
    .B(_1133_),
    .X(_1134_));
 sg13g2_and2_2 _5285_ (.A(_1132_),
    .B(_1134_),
    .X(_1135_));
 sg13g2_nor3_2 _5286_ (.A(_0856_),
    .B(net1933),
    .C(net1929),
    .Y(_1136_));
 sg13g2_nand3_1 _5287_ (.B(net1936),
    .C(net1887),
    .A(net2023),
    .Y(_1137_));
 sg13g2_nand2_2 _5288_ (.Y(_1138_),
    .A(net1940),
    .B(_1136_));
 sg13g2_nor2_1 _5289_ (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .B(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .Y(_1139_));
 sg13g2_or2_2 _5290_ (.X(_1140_),
    .B(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .A(\z80.tv80s.i_tv80_core.XY_State[1] ));
 sg13g2_nor2_2 _5291_ (.A(net2052),
    .B(net1924),
    .Y(_1141_));
 sg13g2_nor3_1 _5292_ (.A(net2172),
    .B(\z80.tv80s.i_tv80_core.ISet[1] ),
    .C(\z80.tv80s.i_tv80_core.ISet[3] ),
    .Y(_1142_));
 sg13g2_nand2b_2 _5293_ (.Y(_1143_),
    .B(net2105),
    .A_N(_1142_));
 sg13g2_nand2b_2 _5294_ (.Y(_1144_),
    .B(_1138_),
    .A_N(_0818_));
 sg13g2_a21oi_2 _5295_ (.B1(net2167),
    .Y(_1145_),
    .A2(_1144_),
    .A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sg13g2_a22oi_1 _5296_ (.Y(_1146_),
    .B1(_0948_),
    .B2(_0939_),
    .A2(_0942_),
    .A1(_0840_));
 sg13g2_a221oi_1 _5297_ (.B2(net1936),
    .C1(_0972_),
    .B1(_0982_),
    .A1(_0840_),
    .Y(_1147_),
    .A2(_0942_));
 sg13g2_nor4_2 _5298_ (.A(net2024),
    .B(net2001),
    .C(net1944),
    .Y(_1148_),
    .D(net1932));
 sg13g2_nand2_1 _5299_ (.Y(_1149_),
    .A(net2088),
    .B(_0959_));
 sg13g2_nand2_2 _5300_ (.Y(_1150_),
    .A(_0969_),
    .B(_1149_));
 sg13g2_and2_2 _5301_ (.A(net2005),
    .B(_0912_),
    .X(_1151_));
 sg13g2_nand2_1 _5302_ (.Y(_1152_),
    .A(net1928),
    .B(_1151_));
 sg13g2_nor3_1 _5303_ (.A(net1998),
    .B(net1931),
    .C(_1152_),
    .Y(_1153_));
 sg13g2_nor4_1 _5304_ (.A(_0992_),
    .B(_1003_),
    .C(_1150_),
    .D(_1153_),
    .Y(_1154_));
 sg13g2_nor2_1 _5305_ (.A(net2095),
    .B(_0830_),
    .Y(_1155_));
 sg13g2_nor3_1 _5306_ (.A(_0857_),
    .B(net1888),
    .C(_0979_),
    .Y(_1156_));
 sg13g2_o21ai_1 _5307_ (.B1(_1156_),
    .Y(_1157_),
    .A1(_0830_),
    .A2(net1928));
 sg13g2_nand2_1 _5308_ (.Y(_1158_),
    .A(_0817_),
    .B(_1157_));
 sg13g2_nand3_1 _5309_ (.B(_1154_),
    .C(_1158_),
    .A(_1147_),
    .Y(_1159_));
 sg13g2_nor2_2 _5310_ (.A(_0818_),
    .B(_1021_),
    .Y(_1160_));
 sg13g2_or2_1 _5311_ (.X(_1161_),
    .B(_1021_),
    .A(_0818_));
 sg13g2_nor2_2 _5312_ (.A(_0974_),
    .B(_1161_),
    .Y(_1162_));
 sg13g2_nand2_1 _5313_ (.Y(_1163_),
    .A(_0975_),
    .B(_1160_));
 sg13g2_nor4_2 _5314_ (.A(net2086),
    .B(net2001),
    .C(net1955),
    .Y(_1164_),
    .D(net1944));
 sg13g2_nand2_2 _5315_ (.Y(_1165_),
    .A(_0840_),
    .B(_0967_));
 sg13g2_nand4_1 _5316_ (.B(_0953_),
    .C(_1162_),
    .A(_0928_),
    .Y(_1166_),
    .D(_1165_));
 sg13g2_nor3_1 _5317_ (.A(net1998),
    .B(net1931),
    .C(_0943_),
    .Y(_1167_));
 sg13g2_a21o_2 _5318_ (.A2(_0939_),
    .A1(_0840_),
    .B1(_1167_),
    .X(_1168_));
 sg13g2_inv_1 _5319_ (.Y(_1169_),
    .A(_1168_));
 sg13g2_nor3_1 _5320_ (.A(net1998),
    .B(_0816_),
    .C(_0850_),
    .Y(_1170_));
 sg13g2_nor4_1 _5321_ (.A(net2005),
    .B(net1999),
    .C(net1931),
    .D(net1929),
    .Y(_1171_));
 sg13g2_or3_2 _5322_ (.A(_0841_),
    .B(_1170_),
    .C(_1171_),
    .X(_1172_));
 sg13g2_or2_1 _5323_ (.X(_1173_),
    .B(_1172_),
    .A(_1168_));
 sg13g2_nor4_2 _5324_ (.A(net2082),
    .B(net1998),
    .C(net1944),
    .Y(_1174_),
    .D(net1931));
 sg13g2_nand2_1 _5325_ (.Y(_1175_),
    .A(net2023),
    .B(_0959_));
 sg13g2_nor2_2 _5326_ (.A(_1001_),
    .B(_1174_),
    .Y(_1176_));
 sg13g2_nor2_2 _5327_ (.A(_0932_),
    .B(_0966_),
    .Y(_1177_));
 sg13g2_nand4_1 _5328_ (.B(_0995_),
    .C(_1176_),
    .A(_0922_),
    .Y(_1178_),
    .D(_1177_));
 sg13g2_nor4_2 _5329_ (.A(_1159_),
    .B(_1166_),
    .C(_1173_),
    .Y(_1179_),
    .D(_1178_));
 sg13g2_nand2_2 _5330_ (.Y(_1180_),
    .A(_0931_),
    .B(_0956_));
 sg13g2_nand2_1 _5331_ (.Y(_1181_),
    .A(net2121),
    .B(_1180_));
 sg13g2_a22oi_1 _5332_ (.Y(_1182_),
    .B1(_1181_),
    .B2(_0852_),
    .A2(_1144_),
    .A1(net2106));
 sg13g2_nor2_1 _5333_ (.A(_0864_),
    .B(net1932),
    .Y(_1183_));
 sg13g2_nor2_2 _5334_ (.A(_0816_),
    .B(_0864_),
    .Y(_1184_));
 sg13g2_nand4_1 _5335_ (.B(net1885),
    .C(_0986_),
    .A(net2085),
    .Y(_1185_),
    .D(_1184_));
 sg13g2_o21ai_1 _5336_ (.B1(_1185_),
    .Y(_1186_),
    .A1(net2092),
    .A2(net1890));
 sg13g2_a21oi_1 _5337_ (.A1(_1151_),
    .A2(_1183_),
    .Y(_1187_),
    .B1(_1186_));
 sg13g2_nor3_2 _5338_ (.A(_0671_),
    .B(net1957),
    .C(net1950),
    .Y(_1188_));
 sg13g2_or3_2 _5339_ (.A(_0671_),
    .B(net1957),
    .C(net1949),
    .X(_1189_));
 sg13g2_nor2_2 _5340_ (.A(net2024),
    .B(_0860_),
    .Y(_1190_));
 sg13g2_and2_1 _5341_ (.A(net1951),
    .B(_0878_),
    .X(_1191_));
 sg13g2_and2_2 _5342_ (.A(net2102),
    .B(_1191_),
    .X(_1192_));
 sg13g2_nand2_1 _5343_ (.Y(_1193_),
    .A(_0815_),
    .B(_1192_));
 sg13g2_o21ai_1 _5344_ (.B1(_1193_),
    .Y(_1194_),
    .A1(_0838_),
    .A2(_0851_));
 sg13g2_a221oi_1 _5345_ (.B2(net2065),
    .C1(_1194_),
    .B1(_1190_),
    .A1(net1935),
    .Y(_1195_),
    .A2(_1188_));
 sg13g2_a21oi_1 _5346_ (.A1(net2086),
    .A2(net2065),
    .Y(_1196_),
    .B1(_0858_));
 sg13g2_o21ai_1 _5347_ (.B1(net1951),
    .Y(_1197_),
    .A1(_0962_),
    .A2(_1196_));
 sg13g2_a22oi_1 _5348_ (.Y(_1198_),
    .B1(_1192_),
    .B2(_0816_),
    .A2(_1188_),
    .A1(net1933));
 sg13g2_nor2_2 _5349_ (.A(net1949),
    .B(net1945),
    .Y(_1199_));
 sg13g2_or2_2 _5350_ (.X(_1200_),
    .B(net1945),
    .A(net1949));
 sg13g2_and4_1 _5351_ (.A(_0885_),
    .B(_1197_),
    .C(_1198_),
    .D(_1200_),
    .X(_1201_));
 sg13g2_or3_1 _5352_ (.A(_0939_),
    .B(_0960_),
    .C(_0985_),
    .X(_1202_));
 sg13g2_nor2_1 _5353_ (.A(net1886),
    .B(_1151_),
    .Y(_1203_));
 sg13g2_nor2_1 _5354_ (.A(net1929),
    .B(net1928),
    .Y(_1204_));
 sg13g2_nand2_1 _5355_ (.Y(_1205_),
    .A(_0670_),
    .B(_0979_));
 sg13g2_o21ai_1 _5356_ (.B1(_0850_),
    .Y(_1206_),
    .A1(net2095),
    .A2(net1929));
 sg13g2_nor3_1 _5357_ (.A(net2073),
    .B(net1890),
    .C(_1205_),
    .Y(_1207_));
 sg13g2_a22oi_1 _5358_ (.Y(_1208_),
    .B1(_1206_),
    .B2(_0865_),
    .A2(_1203_),
    .A1(_1183_));
 sg13g2_nand2_1 _5359_ (.Y(_1209_),
    .A(_0958_),
    .B(_1204_));
 sg13g2_a21oi_1 _5360_ (.A1(net2095),
    .A2(net2091),
    .Y(_1210_),
    .B1(net2085));
 sg13g2_a22oi_1 _5361_ (.Y(_1211_),
    .B1(_1184_),
    .B2(_1210_),
    .A2(_1155_),
    .A1(_0865_));
 sg13g2_nand3_1 _5362_ (.B(_1209_),
    .C(_1211_),
    .A(_1208_),
    .Y(_1212_));
 sg13g2_a21oi_1 _5363_ (.A1(_1184_),
    .A2(_1202_),
    .Y(_1213_),
    .B1(_1212_));
 sg13g2_and2_1 _5364_ (.A(_1201_),
    .B(_1213_),
    .X(_1214_));
 sg13g2_nand4_1 _5365_ (.B(_1187_),
    .C(_1195_),
    .A(_1182_),
    .Y(_1215_),
    .D(_1214_));
 sg13g2_nor3_1 _5366_ (.A(net2064),
    .B(_0827_),
    .C(_0967_),
    .Y(_1216_));
 sg13g2_o21ai_1 _5367_ (.B1(_1216_),
    .Y(_1217_),
    .A1(_0670_),
    .A2(net2004));
 sg13g2_a21o_1 _5368_ (.A2(net2091),
    .A1(net2096),
    .B1(_0855_),
    .X(_1218_));
 sg13g2_o21ai_1 _5369_ (.B1(net2064),
    .Y(_1219_),
    .A1(net1888),
    .A2(_1218_));
 sg13g2_nand3_1 _5370_ (.B(_1217_),
    .C(_1219_),
    .A(net1941),
    .Y(_1220_));
 sg13g2_nand3_1 _5371_ (.B(_1061_),
    .C(_1220_),
    .A(_0991_),
    .Y(_1221_));
 sg13g2_nor2_1 _5372_ (.A(_0901_),
    .B(_0980_),
    .Y(_1222_));
 sg13g2_o21ai_1 _5373_ (.B1(_1222_),
    .Y(_1223_),
    .A1(_0830_),
    .A2(net1928));
 sg13g2_nand3_1 _5374_ (.B(_0813_),
    .C(_1223_),
    .A(net2073),
    .Y(_1224_));
 sg13g2_a21oi_1 _5375_ (.A1(_1152_),
    .A2(_1205_),
    .Y(_1225_),
    .B1(_0949_));
 sg13g2_a221oi_1 _5376_ (.B2(_0958_),
    .C1(_1225_),
    .B1(_1204_),
    .A1(_0840_),
    .Y(_1226_),
    .A2(_1157_));
 sg13g2_nand2_2 _5377_ (.Y(_1227_),
    .A(_1224_),
    .B(_1226_));
 sg13g2_nor3_2 _5378_ (.A(_1215_),
    .B(_1221_),
    .C(_1227_),
    .Y(_1228_));
 sg13g2_nand3_1 _5379_ (.B(_0847_),
    .C(_0962_),
    .A(net2089),
    .Y(_1229_));
 sg13g2_nand2_2 _5380_ (.Y(_1230_),
    .A(net1951),
    .B(_0985_));
 sg13g2_a21oi_1 _5381_ (.A1(_1179_),
    .A2(_1228_),
    .Y(_1231_),
    .B1(_1145_));
 sg13g2_nand2b_1 _5382_ (.Y(_1232_),
    .B(_0934_),
    .A_N(_0999_));
 sg13g2_o21ai_1 _5383_ (.B1(_0857_),
    .Y(_1233_),
    .A1(_0894_),
    .A2(_0906_));
 sg13g2_nor2_2 _5384_ (.A(_0863_),
    .B(_1164_),
    .Y(_1234_));
 sg13g2_a21oi_1 _5385_ (.A1(_0857_),
    .A2(_0899_),
    .Y(_1235_),
    .B1(_0930_));
 sg13g2_nor2b_1 _5386_ (.A(_1010_),
    .B_N(_1235_),
    .Y(_1236_));
 sg13g2_nand3_1 _5387_ (.B(_1234_),
    .C(_1236_),
    .A(_1233_),
    .Y(_1237_));
 sg13g2_nand2_2 _5388_ (.Y(_1238_),
    .A(net1885),
    .B(_1047_));
 sg13g2_nand3_1 _5389_ (.B(_1137_),
    .C(_1238_),
    .A(net2126),
    .Y(_1239_));
 sg13g2_or2_2 _5390_ (.X(_1240_),
    .B(_1020_),
    .A(_0946_));
 sg13g2_nor2_2 _5391_ (.A(_0952_),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_nand2_2 _5392_ (.Y(_1242_),
    .A(_1162_),
    .B(_1241_));
 sg13g2_nand2_2 _5393_ (.Y(_1243_),
    .A(net1941),
    .B(net1888));
 sg13g2_nor3_2 _5394_ (.A(net1957),
    .B(net1939),
    .C(_0913_),
    .Y(_1244_));
 sg13g2_nand2_2 _5395_ (.Y(_1245_),
    .A(net2002),
    .B(net1886));
 sg13g2_nor2_1 _5396_ (.A(_0968_),
    .B(net1882),
    .Y(_1246_));
 sg13g2_nand3_1 _5397_ (.B(_1245_),
    .C(_1246_),
    .A(_1177_),
    .Y(_1247_));
 sg13g2_nor3_1 _5398_ (.A(_0841_),
    .B(_0970_),
    .C(_0972_),
    .Y(_1248_));
 sg13g2_nand2_1 _5399_ (.Y(_1249_),
    .A(_1062_),
    .B(_1248_));
 sg13g2_or4_1 _5400_ (.A(_1242_),
    .B(_1244_),
    .C(_1247_),
    .D(_1249_),
    .X(_1250_));
 sg13g2_nand2_1 _5401_ (.Y(_1251_),
    .A(_0998_),
    .B(_1012_));
 sg13g2_nor2_1 _5402_ (.A(_0970_),
    .B(_1003_),
    .Y(_1252_));
 sg13g2_nand3_1 _5403_ (.B(_0996_),
    .C(_1062_),
    .A(_0991_),
    .Y(_1253_));
 sg13g2_nor4_2 _5404_ (.A(_0970_),
    .B(_1003_),
    .C(_1150_),
    .Y(_1254_),
    .D(_1253_));
 sg13g2_nor4_2 _5405_ (.A(net2083),
    .B(net1955),
    .C(_0850_),
    .Y(_1255_),
    .D(net1937));
 sg13g2_nor2_1 _5406_ (.A(_0946_),
    .B(_1255_),
    .Y(_1256_));
 sg13g2_or2_2 _5407_ (.X(_1257_),
    .B(_1255_),
    .A(_0946_));
 sg13g2_nand2b_1 _5408_ (.Y(_1258_),
    .B(net2005),
    .A_N(_0929_));
 sg13g2_and3_2 _5409_ (.X(_1259_),
    .A(net2067),
    .B(net1940),
    .C(_0942_));
 sg13g2_nand2_2 _5410_ (.Y(_1260_),
    .A(_0899_),
    .B(_0942_));
 sg13g2_nor2_2 _5411_ (.A(net2073),
    .B(_1260_),
    .Y(_1261_));
 sg13g2_nor3_1 _5412_ (.A(net1881),
    .B(_1161_),
    .C(_1261_),
    .Y(_1262_));
 sg13g2_nor2_2 _5413_ (.A(_0972_),
    .B(_1005_),
    .Y(_1263_));
 sg13g2_nor2_1 _5414_ (.A(net2088),
    .B(_1233_),
    .Y(_1264_));
 sg13g2_o21ai_1 _5415_ (.B1(_0909_),
    .Y(_1265_),
    .A1(net2082),
    .A2(_1233_));
 sg13g2_nor2_1 _5416_ (.A(_0932_),
    .B(_0981_),
    .Y(_1266_));
 sg13g2_or4_1 _5417_ (.A(_0959_),
    .B(_1232_),
    .C(_1237_),
    .D(_1250_),
    .X(_1267_));
 sg13g2_inv_2 _5418_ (.Y(_1268_),
    .A(net1843));
 sg13g2_o21ai_1 _5419_ (.B1(net2168),
    .Y(_1269_),
    .A1(_1239_),
    .A2(net1843));
 sg13g2_or2_1 _5420_ (.X(_1270_),
    .B(_1233_),
    .A(net2130));
 sg13g2_a21oi_1 _5421_ (.A1(net2131),
    .A2(net1886),
    .Y(_1271_),
    .B1(_1234_));
 sg13g2_a21oi_1 _5422_ (.A1(net1947),
    .A2(net1875),
    .Y(_1272_),
    .B1(_1009_));
 sg13g2_a21oi_1 _5423_ (.A1(net2118),
    .A2(net1875),
    .Y(_1273_),
    .B1(_0931_));
 sg13g2_nor4_1 _5424_ (.A(_1007_),
    .B(_1271_),
    .C(_1272_),
    .D(_1273_),
    .Y(_1274_));
 sg13g2_nand4_1 _5425_ (.B(_1237_),
    .C(_1270_),
    .A(_0924_),
    .Y(_1275_),
    .D(_1274_));
 sg13g2_nand2b_1 _5426_ (.Y(_1276_),
    .B(_1275_),
    .A_N(_1269_));
 sg13g2_nor2_1 _5427_ (.A(net1891),
    .B(_1200_),
    .Y(_1277_));
 sg13g2_nand2_2 _5428_ (.Y(_1278_),
    .A(net1953),
    .B(_1199_));
 sg13g2_or4_1 _5429_ (.A(_1111_),
    .B(_1188_),
    .C(_1191_),
    .D(_1199_),
    .X(_1279_));
 sg13g2_nand2_1 _5430_ (.Y(_1280_),
    .A(net1942),
    .B(_0884_));
 sg13g2_nor2_1 _5431_ (.A(net2129),
    .B(_1110_),
    .Y(_1281_));
 sg13g2_a21oi_1 _5432_ (.A1(net2018),
    .A2(_1191_),
    .Y(_1282_),
    .B1(_1188_));
 sg13g2_a21oi_1 _5433_ (.A1(_0861_),
    .A2(_1107_),
    .Y(_1283_),
    .B1(_1281_));
 sg13g2_and4_1 _5434_ (.A(_1279_),
    .B(_1280_),
    .C(_1282_),
    .D(_1283_),
    .X(_1284_));
 sg13g2_o21ai_1 _5435_ (.B1(_1284_),
    .Y(_1285_),
    .A1(net1946),
    .A2(_1105_));
 sg13g2_a21oi_1 _5436_ (.A1(net1953),
    .A2(_1285_),
    .Y(_1286_),
    .B1(_1231_));
 sg13g2_nand3_1 _5437_ (.B(_1278_),
    .C(_1286_),
    .A(_1276_),
    .Y(_1287_));
 sg13g2_and2_1 _5438_ (.A(_1143_),
    .B(_1287_),
    .X(_1288_));
 sg13g2_mux2_1 _5439_ (.A0(_0680_),
    .A1(_1057_),
    .S(net2109),
    .X(_1289_));
 sg13g2_a21oi_1 _5440_ (.A1(net2113),
    .A2(_1289_),
    .Y(_1290_),
    .B1(_1006_));
 sg13g2_nand2_1 _5441_ (.Y(_1291_),
    .A(net2019),
    .B(net2112));
 sg13g2_inv_1 _5442_ (.Y(_1292_),
    .A(_1291_));
 sg13g2_nand2b_1 _5443_ (.Y(_1293_),
    .B(net2131),
    .A_N(_1057_));
 sg13g2_a21oi_1 _5444_ (.A1(_1291_),
    .A2(_1293_),
    .Y(_1294_),
    .B1(_0987_));
 sg13g2_nor2_1 _5445_ (.A(_0677_),
    .B(_0880_),
    .Y(_1295_));
 sg13g2_o21ai_1 _5446_ (.B1(net2113),
    .Y(_1296_),
    .A1(net2109),
    .A2(net2108));
 sg13g2_nor2_1 _5447_ (.A(net2127),
    .B(_1165_),
    .Y(_1297_));
 sg13g2_nand2_1 _5448_ (.Y(_1298_),
    .A(net2019),
    .B(_1164_));
 sg13g2_a21oi_1 _5449_ (.A1(net2111),
    .A2(_1297_),
    .Y(_1299_),
    .B1(_1003_));
 sg13g2_nor2_1 _5450_ (.A(_1295_),
    .B(_1299_),
    .Y(_1300_));
 sg13g2_nor3_2 _5451_ (.A(net2083),
    .B(net1999),
    .C(net1958),
    .Y(_1301_));
 sg13g2_nor3_1 _5452_ (.A(_0982_),
    .B(_0989_),
    .C(_1301_),
    .Y(_1302_));
 sg13g2_o21ai_1 _5453_ (.B1(_0864_),
    .Y(_1303_),
    .A1(net2096),
    .A2(_0929_));
 sg13g2_or2_1 _5454_ (.X(_1304_),
    .B(_1303_),
    .A(net2017));
 sg13g2_a21oi_1 _5455_ (.A1(_1002_),
    .A2(_1302_),
    .Y(_1305_),
    .B1(net1947));
 sg13g2_a21oi_1 _5456_ (.A1(_1001_),
    .A2(_1064_),
    .Y(_1306_),
    .B1(_1304_));
 sg13g2_nand3_1 _5457_ (.B(_1270_),
    .C(_1306_),
    .A(_1235_),
    .Y(_1307_));
 sg13g2_nor4_1 _5458_ (.A(_1294_),
    .B(_1300_),
    .C(_1305_),
    .D(_1307_),
    .Y(_1308_));
 sg13g2_a21oi_1 _5459_ (.A1(net2111),
    .A2(_0959_),
    .Y(_1309_),
    .B1(_1250_));
 sg13g2_and2_1 _5460_ (.A(net1844),
    .B(_1309_),
    .X(_1310_));
 sg13g2_nand2_1 _5461_ (.Y(_1311_),
    .A(_1308_),
    .B(_1310_));
 sg13g2_nor2b_1 _5462_ (.A(net2126),
    .B_N(net2114),
    .Y(_1312_));
 sg13g2_nand2_2 _5463_ (.Y(_1313_),
    .A(net2120),
    .B(net2018));
 sg13g2_o21ai_1 _5464_ (.B1(_1313_),
    .Y(_1314_),
    .A1(_0868_),
    .A2(_1104_));
 sg13g2_nor4_1 _5465_ (.A(net2169),
    .B(_0884_),
    .C(_1109_),
    .D(_1199_),
    .Y(_1315_));
 sg13g2_nor2_1 _5466_ (.A(_0877_),
    .B(_1191_),
    .Y(_1316_));
 sg13g2_o21ai_1 _5467_ (.B1(_1316_),
    .Y(_1317_),
    .A1(net2116),
    .A2(_1189_));
 sg13g2_nand2_1 _5468_ (.Y(_1318_),
    .A(net2018),
    .B(_1317_));
 sg13g2_nand4_1 _5469_ (.B(_1314_),
    .C(_1315_),
    .A(_1279_),
    .Y(_1319_),
    .D(_1318_));
 sg13g2_o21ai_1 _5470_ (.B1(_1319_),
    .Y(_1320_),
    .A1(_1290_),
    .A2(_1311_));
 sg13g2_nand3_1 _5471_ (.B(_1145_),
    .C(_1320_),
    .A(_1143_),
    .Y(_1321_));
 sg13g2_nand2b_1 _5472_ (.Y(_1322_),
    .B(net2019),
    .A_N(_0896_));
 sg13g2_o21ai_1 _5473_ (.B1(_0916_),
    .Y(_1323_),
    .A1(net2109),
    .A2(_0903_));
 sg13g2_nand2_1 _5474_ (.Y(_1324_),
    .A(_0887_),
    .B(_1323_));
 sg13g2_a22oi_1 _5475_ (.Y(_1325_),
    .B1(_0926_),
    .B2(_1296_),
    .A2(_0906_),
    .A1(_0857_));
 sg13g2_nand2_1 _5476_ (.Y(_1326_),
    .A(_1274_),
    .B(_1325_));
 sg13g2_nand3_1 _5477_ (.B(_1322_),
    .C(_1324_),
    .A(_1310_),
    .Y(_1327_));
 sg13g2_nor3_1 _5478_ (.A(_1232_),
    .B(_1326_),
    .C(_1327_),
    .Y(_1328_));
 sg13g2_a22oi_1 _5479_ (.Y(_1329_),
    .B1(_1199_),
    .B2(_1296_),
    .A2(_1104_),
    .A1(net2019));
 sg13g2_a21oi_1 _5480_ (.A1(_1284_),
    .A2(_1329_),
    .Y(_1330_),
    .B1(net1893));
 sg13g2_nor2_1 _5481_ (.A(_1231_),
    .B(_1330_),
    .Y(_1331_));
 sg13g2_o21ai_1 _5482_ (.B1(_1331_),
    .Y(_1332_),
    .A1(_1269_),
    .A2(_1328_));
 sg13g2_and2_2 _5483_ (.A(_1143_),
    .B(_1332_),
    .X(_1333_));
 sg13g2_inv_1 _5484_ (.Y(_1334_),
    .A(_1333_));
 sg13g2_nand3b_1 _5485_ (.B(_1321_),
    .C(_1334_),
    .Y(_1335_),
    .A_N(_1288_));
 sg13g2_inv_1 _5486_ (.Y(_1336_),
    .A(net1701));
 sg13g2_a21oi_1 _5487_ (.A1(net2128),
    .A2(_1144_),
    .Y(_1337_),
    .B1(_1336_));
 sg13g2_nor2b_2 _5488_ (.A(_1337_),
    .B_N(_1141_),
    .Y(_1338_));
 sg13g2_nand3_1 _5489_ (.B(_1138_),
    .C(_1338_),
    .A(_1135_),
    .Y(_1339_));
 sg13g2_nand2_1 _5490_ (.Y(_1340_),
    .A(net2026),
    .B(net2107));
 sg13g2_nor2_1 _5491_ (.A(net2106),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .Y(_1341_));
 sg13g2_nand3_1 _5492_ (.B(net2107),
    .C(_1341_),
    .A(net2026),
    .Y(_1342_));
 sg13g2_nand2_1 _5493_ (.Y(_1343_),
    .A(_1132_),
    .B(_1338_));
 sg13g2_nand2_2 _5494_ (.Y(_1344_),
    .A(\z80.tv80s.i_tv80_core.BusAck ),
    .B(\z80.tv80s.i_tv80_core.BusReq_s ));
 sg13g2_nand2_1 _5495_ (.Y(_1345_),
    .A(_1133_),
    .B(_1344_));
 sg13g2_nand2_1 _5496_ (.Y(_1346_),
    .A(_1134_),
    .B(_1344_));
 sg13g2_or2_2 _5497_ (.X(_1347_),
    .B(_1346_),
    .A(_1343_));
 sg13g2_nand2_1 _5498_ (.Y(_1348_),
    .A(net344),
    .B(_1347_));
 sg13g2_o21ai_1 _5499_ (.B1(_1348_),
    .Y(_0005_),
    .A1(_1339_),
    .A2(_1342_));
 sg13g2_nand3_1 _5500_ (.B(_1074_),
    .C(_1341_),
    .A(_0880_),
    .Y(_1349_));
 sg13g2_nand2_1 _5501_ (.Y(_1350_),
    .A(_1138_),
    .B(_1349_));
 sg13g2_nor2_2 _5502_ (.A(net2107),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .Y(_1351_));
 sg13g2_and4_1 _5503_ (.A(_0669_),
    .B(net2109),
    .C(_0230_),
    .D(_1351_),
    .X(_1352_));
 sg13g2_nand2_1 _5504_ (.Y(_1353_),
    .A(net2026),
    .B(net2106));
 sg13g2_and2_1 _5505_ (.A(_0230_),
    .B(_1353_),
    .X(_1354_));
 sg13g2_nand3_1 _5506_ (.B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .C(_0230_),
    .A(_0669_),
    .Y(_1355_));
 sg13g2_nand4_1 _5507_ (.B(_1342_),
    .C(_1354_),
    .A(_1134_),
    .Y(_1356_),
    .D(_1355_));
 sg13g2_nor4_1 _5508_ (.A(_1343_),
    .B(_1350_),
    .C(_1352_),
    .D(_1356_),
    .Y(_1357_));
 sg13g2_a21o_1 _5509_ (.A2(_1347_),
    .A1(net408),
    .B1(_1357_),
    .X(_0008_));
 sg13g2_nand2_1 _5510_ (.Y(_1358_),
    .A(net488),
    .B(_1347_));
 sg13g2_o21ai_1 _5511_ (.B1(_1358_),
    .Y(_0009_),
    .A1(_1339_),
    .A2(_1355_));
 sg13g2_nor2b_1 _5512_ (.A(_1339_),
    .B_N(_1352_),
    .Y(_1359_));
 sg13g2_a21o_1 _5513_ (.A2(_1347_),
    .A1(net463),
    .B1(_1359_),
    .X(_0010_));
 sg13g2_nand2_1 _5514_ (.Y(_1360_),
    .A(net525),
    .B(_1347_));
 sg13g2_o21ai_1 _5515_ (.B1(_1360_),
    .Y(_0011_),
    .A1(net2025),
    .A2(_1339_));
 sg13g2_nand2_1 _5516_ (.Y(_1361_),
    .A(net260),
    .B(_1347_));
 sg13g2_nand3_1 _5517_ (.B(_1338_),
    .C(_1350_),
    .A(_1135_),
    .Y(_1362_));
 sg13g2_nand2_1 _5518_ (.Y(_0006_),
    .A(_1361_),
    .B(_1362_));
 sg13g2_nor2_1 _5519_ (.A(_1339_),
    .B(_1353_),
    .Y(_1363_));
 sg13g2_a21oi_1 _5520_ (.A1(net443),
    .A2(_1347_),
    .Y(_1364_),
    .B1(_1363_));
 sg13g2_inv_1 _5521_ (.Y(_0007_),
    .A(_1364_));
 sg13g2_or4_1 _5522_ (.A(_0010_),
    .B(_0011_),
    .C(_0006_),
    .D(_0007_),
    .X(_0018_));
 sg13g2_nor2_2 _5523_ (.A(net1981),
    .B(net1892),
    .Y(_1365_));
 sg13g2_nor2_2 _5524_ (.A(net2015),
    .B(net1980),
    .Y(_1366_));
 sg13g2_nand3_1 _5525_ (.B(_0900_),
    .C(_1366_),
    .A(_0857_),
    .Y(_1367_));
 sg13g2_a22oi_1 _5526_ (.Y(_1368_),
    .B1(_1111_),
    .B2(_1365_),
    .A2(net1981),
    .A1(net509));
 sg13g2_nand2_1 _5527_ (.Y(_0012_),
    .A(_1367_),
    .B(_1368_));
 sg13g2_or4_1 _5528_ (.A(_0008_),
    .B(_0009_),
    .C(_0010_),
    .D(_0011_),
    .X(_0017_));
 sg13g2_nor2_2 _5529_ (.A(net1887),
    .B(_1047_),
    .Y(_1369_));
 sg13g2_and3_1 _5530_ (.X(_1370_),
    .A(\z80.tv80s.i_tv80_core.F[0] ),
    .B(net2114),
    .C(net1880));
 sg13g2_a22oi_1 _5531_ (.Y(_1371_),
    .B1(_1370_),
    .B2(_1018_),
    .A2(_1369_),
    .A1(net1951));
 sg13g2_nor2_2 _5532_ (.A(net1949),
    .B(net1885),
    .Y(_1372_));
 sg13g2_nor2_1 _5533_ (.A(_0931_),
    .B(net1875),
    .Y(_1373_));
 sg13g2_a21oi_1 _5534_ (.A1(_1137_),
    .A2(_1372_),
    .Y(_1374_),
    .B1(_1373_));
 sg13g2_nand4_1 _5535_ (.B(_1233_),
    .C(_1371_),
    .A(_0956_),
    .Y(_1375_),
    .D(_1374_));
 sg13g2_nand2_1 _5536_ (.Y(_1376_),
    .A(_1366_),
    .B(_1375_));
 sg13g2_nor4_1 _5537_ (.A(_0033_),
    .B(net1980),
    .C(net1949),
    .D(net1885),
    .Y(_1377_));
 sg13g2_a221oi_1 _5538_ (.B2(_1365_),
    .C1(_1377_),
    .B1(_1191_),
    .A1(net576),
    .Y(_1378_),
    .A2(net1981));
 sg13g2_a22oi_1 _5539_ (.Y(_1379_),
    .B1(_1050_),
    .B2(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(net1878),
    .A1(_0665_));
 sg13g2_o21ai_1 _5540_ (.B1(_1379_),
    .Y(_1380_),
    .A1(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(_1038_));
 sg13g2_nand3_1 _5541_ (.B(_1018_),
    .C(_1366_),
    .A(net2114),
    .Y(_1381_));
 sg13g2_nand2b_1 _5542_ (.Y(_1382_),
    .B(_1380_),
    .A_N(_1381_));
 sg13g2_nand3_1 _5543_ (.B(_1378_),
    .C(_1382_),
    .A(_1376_),
    .Y(_0013_));
 sg13g2_or4_1 _5544_ (.A(_0005_),
    .B(_0009_),
    .C(_0011_),
    .D(_0007_),
    .X(_0019_));
 sg13g2_nor2b_1 _5545_ (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .B_N(\z80.tv80s.i_tv80_core.IntCycle ),
    .Y(_1383_));
 sg13g2_a21o_1 _5546_ (.A2(_0021_),
    .A1(net2113),
    .B1(net2119),
    .X(_1384_));
 sg13g2_a22oi_1 _5547_ (.Y(_1385_),
    .B1(_1384_),
    .B2(net1884),
    .A2(_1383_),
    .A1(_1001_));
 sg13g2_nand4_1 _5548_ (.B(_1004_),
    .C(_1165_),
    .A(_0927_),
    .Y(_1386_),
    .D(_1385_));
 sg13g2_o21ai_1 _5549_ (.B1(_1366_),
    .Y(_1387_),
    .A1(_1081_),
    .A2(_1386_));
 sg13g2_a22oi_1 _5550_ (.Y(_1388_),
    .B1(_1199_),
    .B2(_1365_),
    .A2(net1980),
    .A1(net512));
 sg13g2_nand2_1 _5551_ (.Y(_0014_),
    .A(_1387_),
    .B(_1388_));
 sg13g2_nand2b_1 _5552_ (.Y(_1389_),
    .B(_1293_),
    .A_N(_0987_));
 sg13g2_nor2_1 _5553_ (.A(net2119),
    .B(_1006_),
    .Y(_1390_));
 sg13g2_nor4_1 _5554_ (.A(net2119),
    .B(net2014),
    .C(_1006_),
    .D(_1057_),
    .Y(_1391_));
 sg13g2_nor2_1 _5555_ (.A(net1882),
    .B(_1174_),
    .Y(_1392_));
 sg13g2_nor4_1 _5556_ (.A(_0959_),
    .B(_0982_),
    .C(_1013_),
    .D(_1017_),
    .Y(_1393_));
 sg13g2_nor2_1 _5557_ (.A(_0989_),
    .B(_1011_),
    .Y(_1394_));
 sg13g2_nand2_1 _5558_ (.Y(_1395_),
    .A(_0919_),
    .B(_1394_));
 sg13g2_a21o_1 _5559_ (.A2(_1001_),
    .A1(\z80.tv80s.i_tv80_core.NMICycle ),
    .B1(_0971_),
    .X(_1396_));
 sg13g2_nor4_1 _5560_ (.A(_0923_),
    .B(_1301_),
    .C(_1395_),
    .D(_1396_),
    .Y(_1397_));
 sg13g2_nand3_1 _5561_ (.B(_1393_),
    .C(_1397_),
    .A(_1389_),
    .Y(_1398_));
 sg13g2_o21ai_1 _5562_ (.B1(_1366_),
    .Y(_1399_),
    .A1(_1391_),
    .A2(_1398_));
 sg13g2_nor2_1 _5563_ (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .B(_1034_),
    .Y(_1400_));
 sg13g2_a21oi_1 _5564_ (.A1(\z80.tv80s.i_tv80_core.F[0] ),
    .A2(net1878),
    .Y(_1401_),
    .B1(_1400_));
 sg13g2_nor2_1 _5565_ (.A(_0662_),
    .B(_1038_),
    .Y(_1402_));
 sg13g2_a21oi_1 _5566_ (.A1(_0662_),
    .A2(_1050_),
    .Y(_1403_),
    .B1(_1402_));
 sg13g2_a21oi_1 _5567_ (.A1(_1401_),
    .A2(_1403_),
    .Y(_1404_),
    .B1(_1381_));
 sg13g2_nand2_1 _5568_ (.Y(_1405_),
    .A(_0860_),
    .B(_1189_));
 sg13g2_a221oi_1 _5569_ (.B2(_1405_),
    .C1(_1404_),
    .B1(_1365_),
    .A1(net631),
    .Y(_1406_),
    .A2(net1980));
 sg13g2_nand3_1 _5570_ (.B(net1996),
    .C(_1180_),
    .A(net2167),
    .Y(_1407_));
 sg13g2_nor2_1 _5571_ (.A(net1864),
    .B(_1258_),
    .Y(_1408_));
 sg13g2_and2_1 _5572_ (.A(net2111),
    .B(_1018_),
    .X(_1409_));
 sg13g2_o21ai_1 _5573_ (.B1(_1366_),
    .Y(_1410_),
    .A1(_1408_),
    .A2(_1409_));
 sg13g2_nand4_1 _5574_ (.B(_1406_),
    .C(_1407_),
    .A(_1399_),
    .Y(_0015_),
    .D(_1410_));
 sg13g2_nor3_1 _5575_ (.A(_0835_),
    .B(_0836_),
    .C(_0842_),
    .Y(_1411_));
 sg13g2_a21o_1 _5576_ (.A2(_0835_),
    .A1(net526),
    .B1(_1411_),
    .X(_0000_));
 sg13g2_nor4_1 _5577_ (.A(net2063),
    .B(net1949),
    .C(net1885),
    .D(_1041_),
    .Y(_1412_));
 sg13g2_nor3_1 _5578_ (.A(net2081),
    .B(_0851_),
    .C(net1934),
    .Y(_1413_));
 sg13g2_o21ai_1 _5579_ (.B1(_1365_),
    .Y(_1414_),
    .A1(_1412_),
    .A2(_1413_));
 sg13g2_nand2_1 _5580_ (.Y(_1415_),
    .A(_1365_),
    .B(_1372_));
 sg13g2_nand3_1 _5581_ (.B(_1365_),
    .C(_1372_),
    .A(net2021),
    .Y(_1416_));
 sg13g2_nand3_1 _5582_ (.B(_1414_),
    .C(_1416_),
    .A(net484),
    .Y(_1417_));
 sg13g2_o21ai_1 _5583_ (.B1(_1417_),
    .Y(_0004_),
    .A1(_1034_),
    .A2(_1415_));
 sg13g2_o21ai_1 _5584_ (.B1(net490),
    .Y(_1418_),
    .A1(net1877),
    .A2(_1415_));
 sg13g2_nand2_1 _5585_ (.Y(_0003_),
    .A(_1414_),
    .B(_1418_));
 sg13g2_nor2b_1 _5586_ (.A(_0834_),
    .B_N(net258),
    .Y(_0002_));
 sg13g2_nor4_1 _5587_ (.A(_0669_),
    .B(_0825_),
    .C(_0837_),
    .D(_0841_),
    .Y(_1419_));
 sg13g2_nand3_1 _5588_ (.B(_0833_),
    .C(_1366_),
    .A(_0818_),
    .Y(_1420_));
 sg13g2_a21oi_1 _5589_ (.A1(net2166),
    .A2(_0835_),
    .Y(_1421_),
    .B1(_1419_));
 sg13g2_nand2_1 _5590_ (.Y(_0001_),
    .A(_1420_),
    .B(net621));
 sg13g2_nor2_2 _5591_ (.A(net2014),
    .B(net1946),
    .Y(_1422_));
 sg13g2_nand2_2 _5592_ (.Y(_1423_),
    .A(net2109),
    .B(_0861_));
 sg13g2_nand2_1 _5593_ (.Y(_1424_),
    .A(_1192_),
    .B(net1922));
 sg13g2_nor2_2 _5594_ (.A(_1083_),
    .B(_1351_),
    .Y(_1425_));
 sg13g2_nor2_1 _5595_ (.A(net2080),
    .B(_1200_),
    .Y(_1426_));
 sg13g2_o21ai_1 _5596_ (.B1(_1424_),
    .Y(_1427_),
    .A1(_0872_),
    .A2(_0885_));
 sg13g2_a221oi_1 _5597_ (.B2(_1426_),
    .C1(_1427_),
    .B1(_1425_),
    .A1(_1108_),
    .Y(_1428_),
    .A2(_1422_));
 sg13g2_a21o_1 _5598_ (.A2(_1369_),
    .A1(_0677_),
    .B1(net1843),
    .X(_1429_));
 sg13g2_nor2_2 _5599_ (.A(net2082),
    .B(_0927_),
    .Y(_1430_));
 sg13g2_o21ai_1 _5600_ (.B1(_1004_),
    .Y(_1431_),
    .A1(net2080),
    .A2(_0927_));
 sg13g2_o21ai_1 _5601_ (.B1(_1425_),
    .Y(_1432_),
    .A1(net1884),
    .A2(_1431_));
 sg13g2_nand2b_1 _5602_ (.Y(_1433_),
    .B(_1312_),
    .A_N(_0917_));
 sg13g2_o21ai_1 _5603_ (.B1(_1433_),
    .Y(_1434_),
    .A1(_0872_),
    .A2(_0916_));
 sg13g2_a221oi_1 _5604_ (.B2(net1889),
    .C1(_1434_),
    .B1(_1174_),
    .A1(_0984_),
    .Y(_1435_),
    .A2(_1094_));
 sg13g2_o21ai_1 _5605_ (.B1(_1408_),
    .Y(_1436_),
    .A1(net1883),
    .A2(_1422_));
 sg13g2_a21oi_1 _5606_ (.A1(_0021_),
    .A2(net1883),
    .Y(_1437_),
    .B1(_1436_));
 sg13g2_nor3_1 _5607_ (.A(net2088),
    .B(net2111),
    .C(_0896_),
    .Y(_1438_));
 sg13g2_a21o_1 _5608_ (.A2(_1028_),
    .A1(_0021_),
    .B1(net1946),
    .X(_1439_));
 sg13g2_nor2_1 _5609_ (.A(_1165_),
    .B(_1439_),
    .Y(_1440_));
 sg13g2_nor3_1 _5610_ (.A(_1002_),
    .B(_1064_),
    .C(_1095_),
    .Y(_1441_));
 sg13g2_nor4_1 _5611_ (.A(_1437_),
    .B(_1438_),
    .C(_1440_),
    .D(_1441_),
    .Y(_1442_));
 sg13g2_nand4_1 _5612_ (.B(_1432_),
    .C(_1435_),
    .A(net1843),
    .Y(_1443_),
    .D(_1442_));
 sg13g2_nand3_1 _5613_ (.B(_1429_),
    .C(_1443_),
    .A(net2169),
    .Y(_1444_));
 sg13g2_nand4_1 _5614_ (.B(_0852_),
    .C(net1889),
    .A(net2167),
    .Y(_1445_),
    .D(_1180_));
 sg13g2_and2_1 _5615_ (.A(net1892),
    .B(_1445_),
    .X(_1446_));
 sg13g2_a22oi_1 _5616_ (.Y(doe),
    .B1(_1444_),
    .B2(_1446_),
    .A2(_1428_),
    .A1(net1954));
 sg13g2_nand2_1 _5617_ (.Y(_1447_),
    .A(\addr_bus[8] ),
    .B(net2188));
 sg13g2_o21ai_1 _5618_ (.B1(_1447_),
    .Y(_1448_),
    .A1(_0752_),
    .A2(net2188));
 sg13g2_mux2_2 _5619_ (.A0(_1448_),
    .A1(\z80.m1_n ),
    .S(net2185),
    .X(uo_out[0]));
 sg13g2_nand2b_1 _5620_ (.Y(_1449_),
    .B(\addr_bus[1] ),
    .A_N(net2188));
 sg13g2_a21oi_1 _5621_ (.A1(net2188),
    .A2(\addr_bus[9] ),
    .Y(_1450_),
    .B1(net2185));
 sg13g2_a22oi_1 _5622_ (.Y(uo_out[1]),
    .B1(_1449_),
    .B2(_1450_),
    .A2(_0753_),
    .A1(net2185));
 sg13g2_nand2b_1 _5623_ (.Y(_1451_),
    .B(\addr_bus[2] ),
    .A_N(net2186));
 sg13g2_a21oi_1 _5624_ (.A1(net2186),
    .A2(\addr_bus[10] ),
    .Y(_1452_),
    .B1(net2184));
 sg13g2_a22oi_1 _5625_ (.Y(uo_out[2]),
    .B1(_1451_),
    .B2(_1452_),
    .A2(_0754_),
    .A1(net2185));
 sg13g2_nand2b_1 _5626_ (.Y(_1453_),
    .B(\addr_bus[3] ),
    .A_N(net2186));
 sg13g2_a21oi_1 _5627_ (.A1(net2187),
    .A2(\addr_bus[11] ),
    .Y(_1454_),
    .B1(net2185));
 sg13g2_a22oi_1 _5628_ (.Y(uo_out[3]),
    .B1(_1453_),
    .B2(_1454_),
    .A2(_0755_),
    .A1(net2184));
 sg13g2_nand2b_1 _5629_ (.Y(_1455_),
    .B(\addr_bus[4] ),
    .A_N(net2186));
 sg13g2_a21oi_1 _5630_ (.A1(net2187),
    .A2(\addr_bus[12] ),
    .Y(_1456_),
    .B1(net2185));
 sg13g2_a22oi_1 _5631_ (.Y(uo_out[4]),
    .B1(_1455_),
    .B2(_1456_),
    .A2(_0756_),
    .A1(net2184));
 sg13g2_nand2b_1 _5632_ (.Y(_1457_),
    .B(\addr_bus[5] ),
    .A_N(net2186));
 sg13g2_a21oi_1 _5633_ (.A1(net2187),
    .A2(\addr_bus[13] ),
    .Y(_1458_),
    .B1(net2184));
 sg13g2_a22oi_1 _5634_ (.Y(uo_out[5]),
    .B1(_1457_),
    .B2(_1458_),
    .A2(_0757_),
    .A1(net2184));
 sg13g2_nand2_1 _5635_ (.Y(_1459_),
    .A(net2187),
    .B(\addr_bus[14] ));
 sg13g2_o21ai_1 _5636_ (.B1(_1459_),
    .Y(_1460_),
    .A1(net2186),
    .A2(_0758_));
 sg13g2_mux2_2 _5637_ (.A0(_1460_),
    .A1(_0167_),
    .S(net2184),
    .X(uo_out[6]));
 sg13g2_nand2b_1 _5638_ (.Y(_1461_),
    .B(\addr_bus[7] ),
    .A_N(net2186));
 sg13g2_a21oi_1 _5639_ (.A1(net2186),
    .A2(\addr_bus[15] ),
    .Y(_1462_),
    .B1(net2184));
 sg13g2_a22oi_1 _5640_ (.Y(uo_out[7]),
    .B1(_1461_),
    .B2(_1462_),
    .A2(_0759_),
    .A1(net2184));
 sg13g2_and3_2 _5641_ (.X(_1463_),
    .A(net2142),
    .B(_1037_),
    .C(_1116_));
 sg13g2_nand2_1 _5642_ (.Y(_1464_),
    .A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .B(_1463_));
 sg13g2_nand2_2 _5643_ (.Y(_1465_),
    .A(net1984),
    .B(net1862));
 sg13g2_inv_1 _5644_ (.Y(_1466_),
    .A(_1465_));
 sg13g2_nand4_1 _5645_ (.B(net1907),
    .C(_0820_),
    .A(net563),
    .Y(_1467_),
    .D(net1993));
 sg13g2_nand2_1 _5646_ (.Y(_1468_),
    .A(_1465_),
    .B(_1467_));
 sg13g2_nor2_1 _5647_ (.A(net563),
    .B(_0834_),
    .Y(_1469_));
 sg13g2_a22oi_1 _5648_ (.Y(_0297_),
    .B1(_1469_),
    .B2(_1465_),
    .A2(_1468_),
    .A1(_1464_));
 sg13g2_nor2_1 _5649_ (.A(net502),
    .B(_1468_),
    .Y(_1470_));
 sg13g2_nand2_1 _5650_ (.Y(_1471_),
    .A(\z80.tv80s.i_tv80_core.ACC[1] ),
    .B(_1463_));
 sg13g2_nand2_1 _5651_ (.Y(_1472_),
    .A(\z80.tv80s.i_tv80_core.R[0] ),
    .B(\z80.tv80s.i_tv80_core.R[1] ));
 sg13g2_o21ai_1 _5652_ (.B1(_1465_),
    .Y(_1473_),
    .A1(_0835_),
    .A2(_1472_));
 sg13g2_inv_1 _5653_ (.Y(_1474_),
    .A(_1473_));
 sg13g2_a21oi_1 _5654_ (.A1(_1471_),
    .A2(_1473_),
    .Y(_0298_),
    .B1(net503));
 sg13g2_o21ai_1 _5655_ (.B1(_1473_),
    .Y(_1475_),
    .A1(net540),
    .A2(net1862));
 sg13g2_a21oi_1 _5656_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(net1862),
    .Y(_1476_),
    .B1(_1475_));
 sg13g2_a21oi_1 _5657_ (.A1(_0772_),
    .A2(_1474_),
    .Y(_0299_),
    .B1(_1476_));
 sg13g2_a21oi_1 _5658_ (.A1(\z80.tv80s.i_tv80_core.R[2] ),
    .A2(net537),
    .Y(_1477_),
    .B1(net1862));
 sg13g2_nor2_1 _5659_ (.A(_1474_),
    .B(_1477_),
    .Y(_1478_));
 sg13g2_nand2_1 _5660_ (.Y(_1479_),
    .A(net2146),
    .B(net1862));
 sg13g2_a22oi_1 _5661_ (.Y(_0300_),
    .B1(_1478_),
    .B2(_1479_),
    .A2(_1475_),
    .A1(_0774_));
 sg13g2_nor2_1 _5662_ (.A(net520),
    .B(_1478_),
    .Y(_1480_));
 sg13g2_and3_1 _5663_ (.X(_1481_),
    .A(\z80.tv80s.i_tv80_core.R[2] ),
    .B(\z80.tv80s.i_tv80_core.R[3] ),
    .C(\z80.tv80s.i_tv80_core.R[4] ));
 sg13g2_o21ai_1 _5664_ (.B1(_1473_),
    .Y(_1482_),
    .A1(_1466_),
    .A2(_1481_));
 sg13g2_a21oi_1 _5665_ (.A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(net1862),
    .Y(_1483_),
    .B1(_1482_));
 sg13g2_nor2_1 _5666_ (.A(net521),
    .B(_1483_),
    .Y(_0301_));
 sg13g2_nand2_1 _5667_ (.Y(_1484_),
    .A(net2145),
    .B(net1862));
 sg13g2_a21oi_1 _5668_ (.A1(_0775_),
    .A2(_1465_),
    .Y(_1485_),
    .B1(_1482_));
 sg13g2_a22oi_1 _5669_ (.Y(_0302_),
    .B1(_1484_),
    .B2(_1485_),
    .A2(_1482_),
    .A1(_0775_));
 sg13g2_nor2_1 _5670_ (.A(net523),
    .B(_1485_),
    .Y(_1486_));
 sg13g2_nand2b_1 _5671_ (.Y(_1487_),
    .B(_1463_),
    .A_N(\z80.tv80s.i_tv80_core.ACC[6] ));
 sg13g2_nor3_1 _5672_ (.A(_0775_),
    .B(net1997),
    .C(_1472_),
    .Y(_1488_));
 sg13g2_nand4_1 _5673_ (.B(net1905),
    .C(_1481_),
    .A(net523),
    .Y(_1489_),
    .D(_1488_));
 sg13g2_o21ai_1 _5674_ (.B1(_1487_),
    .Y(_1490_),
    .A1(net1862),
    .A2(_1489_));
 sg13g2_a21oi_1 _5675_ (.A1(net1984),
    .A2(_1490_),
    .Y(_0303_),
    .B1(net524));
 sg13g2_o21ai_1 _5676_ (.B1(_1245_),
    .Y(_1491_),
    .A1(net2101),
    .A2(net1883));
 sg13g2_nor3_1 _5677_ (.A(_0863_),
    .B(_1164_),
    .C(_1491_),
    .Y(_1492_));
 sg13g2_nand2_2 _5678_ (.Y(_1493_),
    .A(net2101),
    .B(_1008_));
 sg13g2_a21oi_1 _5679_ (.A1(net2101),
    .A2(_1008_),
    .Y(_1494_),
    .B1(_1001_));
 sg13g2_and4_2 _5680_ (.A(_1254_),
    .B(_1392_),
    .C(_1492_),
    .D(_1494_),
    .X(_1495_));
 sg13g2_o21ai_1 _5681_ (.B1(net1950),
    .Y(_1496_),
    .A1(net2067),
    .A2(_0831_));
 sg13g2_o21ai_1 _5682_ (.B1(_0931_),
    .Y(_1497_),
    .A1(net2023),
    .A2(_0896_));
 sg13g2_nor2_1 _5683_ (.A(_1496_),
    .B(_1497_),
    .Y(_1498_));
 sg13g2_nand2b_1 _5684_ (.Y(_1499_),
    .B(_1498_),
    .A_N(_1265_));
 sg13g2_nand2_2 _5685_ (.Y(_1500_),
    .A(net2067),
    .B(_0828_));
 sg13g2_o21ai_1 _5686_ (.B1(_1500_),
    .Y(_1501_),
    .A1(net1935),
    .A2(_0983_));
 sg13g2_or2_1 _5687_ (.X(_1502_),
    .B(_1501_),
    .A(_1499_));
 sg13g2_a22oi_1 _5688_ (.Y(_1503_),
    .B1(_0926_),
    .B2(net2086),
    .A2(net1888),
    .A1(_0894_));
 sg13g2_or2_1 _5689_ (.X(_1504_),
    .B(_1301_),
    .A(_0932_));
 sg13g2_nor3_1 _5690_ (.A(_0966_),
    .B(_1430_),
    .C(_1504_),
    .Y(_1505_));
 sg13g2_and2_1 _5691_ (.A(_1503_),
    .B(_1505_),
    .X(_1506_));
 sg13g2_inv_1 _5692_ (.Y(_1507_),
    .A(_1506_));
 sg13g2_o21ai_1 _5693_ (.B1(_1263_),
    .Y(_1508_),
    .A1(net1933),
    .A2(_0983_));
 sg13g2_nand3_1 _5694_ (.B(_0899_),
    .C(net1888),
    .A(net2022),
    .Y(_1509_));
 sg13g2_o21ai_1 _5695_ (.B1(net1888),
    .Y(_1510_),
    .A1(_0906_),
    .A2(_0925_));
 sg13g2_nand3_1 _5696_ (.B(net1928),
    .C(_1151_),
    .A(_0900_),
    .Y(_1511_));
 sg13g2_nand2_1 _5697_ (.Y(_1512_),
    .A(_1510_),
    .B(_1511_));
 sg13g2_nor3_1 _5698_ (.A(_1507_),
    .B(_1508_),
    .C(_1512_),
    .Y(_1513_));
 sg13g2_nor2b_1 _5699_ (.A(_1502_),
    .B_N(_1513_),
    .Y(_1514_));
 sg13g2_nand3_1 _5700_ (.B(_1495_),
    .C(_1514_),
    .A(net2171),
    .Y(_1515_));
 sg13g2_nor3_2 _5701_ (.A(_0950_),
    .B(_1240_),
    .C(_1515_),
    .Y(_1516_));
 sg13g2_and2_1 _5702_ (.A(_0976_),
    .B(_1516_),
    .X(_1517_));
 sg13g2_nand2_2 _5703_ (.Y(_1518_),
    .A(_0976_),
    .B(_1516_));
 sg13g2_nand2_1 _5704_ (.Y(_1519_),
    .A(_1495_),
    .B(_1506_));
 sg13g2_inv_1 _5705_ (.Y(_1520_),
    .A(_1519_));
 sg13g2_or2_1 _5706_ (.X(_1521_),
    .B(_1512_),
    .A(_1499_));
 sg13g2_a21oi_1 _5707_ (.A1(net2087),
    .A2(_0950_),
    .Y(_1522_),
    .B1(net1881));
 sg13g2_a221oi_1 _5708_ (.B2(net2087),
    .C1(net1881),
    .B1(_0950_),
    .A1(_0906_),
    .Y(_1523_),
    .A2(_0942_));
 sg13g2_o21ai_1 _5709_ (.B1(_1522_),
    .Y(_1524_),
    .A1(_0907_),
    .A2(_0943_));
 sg13g2_nor2_1 _5710_ (.A(net2082),
    .B(_0951_),
    .Y(_1525_));
 sg13g2_nor4_2 _5711_ (.A(net2005),
    .B(net1937),
    .C(net1933),
    .Y(_1526_),
    .D(net1929));
 sg13g2_nor3_2 _5712_ (.A(net2082),
    .B(net1944),
    .C(_0949_),
    .Y(_1527_));
 sg13g2_nor4_1 _5713_ (.A(_0941_),
    .B(_0944_),
    .C(_1526_),
    .D(_1527_),
    .Y(_1528_));
 sg13g2_nand2_2 _5714_ (.Y(_1529_),
    .A(_1523_),
    .B(_1528_));
 sg13g2_nor3_2 _5715_ (.A(_0818_),
    .B(_1021_),
    .C(_1255_),
    .Y(_1530_));
 sg13g2_and2_1 _5716_ (.A(_1260_),
    .B(_1530_),
    .X(_1531_));
 sg13g2_nand2_2 _5717_ (.Y(_1532_),
    .A(_1260_),
    .B(_1530_));
 sg13g2_nor2_2 _5718_ (.A(net2017),
    .B(_1532_),
    .Y(_1533_));
 sg13g2_nor3_1 _5719_ (.A(_0945_),
    .B(_0982_),
    .C(_1005_),
    .Y(_1534_));
 sg13g2_nand3_1 _5720_ (.B(_1533_),
    .C(_1534_),
    .A(_1500_),
    .Y(_1535_));
 sg13g2_or4_2 _5721_ (.A(_1519_),
    .B(_1521_),
    .C(_1529_),
    .D(_1535_),
    .X(_1536_));
 sg13g2_nand2_1 _5722_ (.Y(_1537_),
    .A(_1518_),
    .B(net1835));
 sg13g2_or2_1 _5723_ (.X(_1538_),
    .B(_1537_),
    .A(net2106));
 sg13g2_nor3_1 _5724_ (.A(net1978),
    .B(_1321_),
    .C(_1538_),
    .Y(_1539_));
 sg13g2_a21oi_1 _5725_ (.A1(_0760_),
    .A2(net1977),
    .Y(_0304_),
    .B1(_1539_));
 sg13g2_a21oi_1 _5726_ (.A1(_1140_),
    .A2(_1537_),
    .Y(_1540_),
    .B1(net2106));
 sg13g2_a221oi_1 _5727_ (.B2(net532),
    .C1(net1978),
    .B1(_1540_),
    .A1(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .Y(_1541_),
    .A2(_1538_));
 sg13g2_a21oi_1 _5728_ (.A1(net2006),
    .A2(net1977),
    .Y(_0305_),
    .B1(_1541_));
 sg13g2_nand2_1 _5729_ (.Y(_1542_),
    .A(net193),
    .B(net1977));
 sg13g2_a21oi_1 _5730_ (.A1(net2097),
    .A2(net2166),
    .Y(_1543_),
    .B1(net1952));
 sg13g2_nand2_1 _5731_ (.Y(_1544_),
    .A(_1175_),
    .B(_1245_));
 sg13g2_nand3_1 _5732_ (.B(_0930_),
    .C(net1875),
    .A(net2118),
    .Y(_1545_));
 sg13g2_a22oi_1 _5733_ (.Y(_1546_),
    .B1(_1544_),
    .B2(net2118),
    .A2(_1264_),
    .A1(net2127));
 sg13g2_nand2_1 _5734_ (.Y(_1547_),
    .A(_1545_),
    .B(_1546_));
 sg13g2_nor2_1 _5735_ (.A(net2114),
    .B(net1885),
    .Y(_1548_));
 sg13g2_nand2_1 _5736_ (.Y(_1549_),
    .A(net1886),
    .B(_1313_));
 sg13g2_nand2_1 _5737_ (.Y(_1550_),
    .A(_0863_),
    .B(_1549_));
 sg13g2_a21oi_1 _5738_ (.A1(_0024_),
    .A2(net1885),
    .Y(_1551_),
    .B1(_1550_));
 sg13g2_nand2_2 _5739_ (.Y(_1552_),
    .A(net1876),
    .B(_1313_));
 sg13g2_nand2_1 _5740_ (.Y(_1553_),
    .A(_1008_),
    .B(_1552_));
 sg13g2_nand2_2 _5741_ (.Y(_1554_),
    .A(net2131),
    .B(_1011_));
 sg13g2_nand2_1 _5742_ (.Y(_1555_),
    .A(_1553_),
    .B(_1554_));
 sg13g2_nand2_1 _5743_ (.Y(_1556_),
    .A(_0886_),
    .B(_0915_));
 sg13g2_nor2_1 _5744_ (.A(net2118),
    .B(_0684_),
    .Y(_1557_));
 sg13g2_nand2b_1 _5745_ (.Y(_1558_),
    .B(_0021_),
    .A_N(net2120));
 sg13g2_nor2_2 _5746_ (.A(net1932),
    .B(_1557_),
    .Y(_1559_));
 sg13g2_nor2_1 _5747_ (.A(net2022),
    .B(_1292_),
    .Y(_1560_));
 sg13g2_a22oi_1 _5748_ (.Y(_1561_),
    .B1(_1560_),
    .B2(_0981_),
    .A2(_1559_),
    .A1(net1882));
 sg13g2_nand2_1 _5749_ (.Y(_1562_),
    .A(_1556_),
    .B(_1561_));
 sg13g2_nor4_2 _5750_ (.A(_1547_),
    .B(_1551_),
    .C(_1555_),
    .Y(_1563_),
    .D(_1562_));
 sg13g2_nand2_1 _5751_ (.Y(_1564_),
    .A(net1843),
    .B(_1563_));
 sg13g2_nand3_1 _5752_ (.B(net2126),
    .C(_1369_),
    .A(net2097),
    .Y(_1565_));
 sg13g2_o21ai_1 _5753_ (.B1(_1565_),
    .Y(_1566_),
    .A1(_0024_),
    .A2(_1238_));
 sg13g2_o21ai_1 _5754_ (.B1(_1564_),
    .Y(_1567_),
    .A1(net1843),
    .A2(_1566_));
 sg13g2_o21ai_1 _5755_ (.B1(_1543_),
    .Y(_1568_),
    .A1(net2015),
    .A2(_1567_));
 sg13g2_o21ai_1 _5756_ (.B1(net1954),
    .Y(_1569_),
    .A1(_0885_),
    .A2(_0887_));
 sg13g2_a21oi_1 _5757_ (.A1(_0879_),
    .A2(net1922),
    .Y(_1570_),
    .B1(_1569_));
 sg13g2_nand2_1 _5758_ (.Y(_1571_),
    .A(net1954),
    .B(_1229_));
 sg13g2_nor2b_1 _5759_ (.A(_1569_),
    .B_N(_1229_),
    .Y(_1572_));
 sg13g2_nand2_1 _5760_ (.Y(_1573_),
    .A(_1229_),
    .B(_1570_));
 sg13g2_o21ai_1 _5761_ (.B1(_1426_),
    .Y(_1574_),
    .A1(net2109),
    .A2(_0680_));
 sg13g2_nand2b_1 _5762_ (.Y(_1575_),
    .B(net2075),
    .A_N(net2121));
 sg13g2_nor3_1 _5763_ (.A(net2068),
    .B(_1574_),
    .C(_1575_),
    .Y(_1576_));
 sg13g2_nand2_1 _5764_ (.Y(_1577_),
    .A(net2102),
    .B(net2123));
 sg13g2_and2_1 _5765_ (.A(net2124),
    .B(_1192_),
    .X(_1578_));
 sg13g2_a22oi_1 _5766_ (.Y(_1579_),
    .B1(_1578_),
    .B2(net2075),
    .A2(_1559_),
    .A1(_0859_));
 sg13g2_o21ai_1 _5767_ (.B1(_1579_),
    .Y(_1580_),
    .A1(_0861_),
    .A2(_1106_));
 sg13g2_nor3_1 _5768_ (.A(_1573_),
    .B(_1576_),
    .C(_1580_),
    .Y(_1581_));
 sg13g2_nor2_1 _5769_ (.A(net2105),
    .B(_1581_),
    .Y(_1582_));
 sg13g2_a22oi_1 _5770_ (.Y(_1583_),
    .B1(_1568_),
    .B2(_1582_),
    .A2(net2097),
    .A1(net2105));
 sg13g2_inv_2 _5771_ (.Y(_1584_),
    .A(_1583_));
 sg13g2_a21oi_1 _5772_ (.A1(net2093),
    .A2(net2166),
    .Y(_1585_),
    .B1(_0845_));
 sg13g2_a22oi_1 _5773_ (.Y(_1586_),
    .B1(_1289_),
    .B2(_1390_),
    .A2(_0982_),
    .A1(net1946));
 sg13g2_a21oi_1 _5774_ (.A1(_0027_),
    .A2(net1885),
    .Y(_1587_),
    .B1(_1550_));
 sg13g2_a21o_1 _5775_ (.A2(_1431_),
    .A1(_0881_),
    .B1(_1587_),
    .X(_1588_));
 sg13g2_nor2_1 _5776_ (.A(net2022),
    .B(net2131),
    .Y(_1589_));
 sg13g2_nor2_1 _5777_ (.A(net1956),
    .B(_1557_),
    .Y(_1590_));
 sg13g2_nand2_1 _5778_ (.Y(_1591_),
    .A(net1882),
    .B(_1590_));
 sg13g2_nand2_2 _5779_ (.Y(_1592_),
    .A(_0681_),
    .B(_0028_));
 sg13g2_nand3_1 _5780_ (.B(_1001_),
    .C(_1592_),
    .A(net1946),
    .Y(_1593_));
 sg13g2_a21oi_1 _5781_ (.A1(net2112),
    .A2(_0871_),
    .Y(_1594_),
    .B1(_1298_));
 sg13g2_nor2_1 _5782_ (.A(_1292_),
    .B(_1589_),
    .Y(_1595_));
 sg13g2_nand4_1 _5783_ (.B(net2002),
    .C(_0980_),
    .A(net2066),
    .Y(_1596_),
    .D(_1595_));
 sg13g2_nand4_1 _5784_ (.B(_1591_),
    .C(_1593_),
    .A(_1556_),
    .Y(_1597_),
    .D(_1596_));
 sg13g2_nor4_1 _5785_ (.A(_1547_),
    .B(_1588_),
    .C(_1594_),
    .D(_1597_),
    .Y(_1598_));
 sg13g2_nand3_1 _5786_ (.B(_1586_),
    .C(_1598_),
    .A(net1844),
    .Y(_1599_));
 sg13g2_nand3_1 _5787_ (.B(net2126),
    .C(_1369_),
    .A(net2093),
    .Y(_1600_));
 sg13g2_o21ai_1 _5788_ (.B1(_1600_),
    .Y(_1601_),
    .A1(_0027_),
    .A2(_1238_));
 sg13g2_o21ai_1 _5789_ (.B1(_1599_),
    .Y(_1602_),
    .A1(net1843),
    .A2(_1601_));
 sg13g2_o21ai_1 _5790_ (.B1(_1585_),
    .Y(_1603_),
    .A1(net2015),
    .A2(_1602_));
 sg13g2_nand3_1 _5791_ (.B(_0865_),
    .C(net1922),
    .A(_0671_),
    .Y(_1604_));
 sg13g2_nor3_1 _5792_ (.A(net2114),
    .B(net1956),
    .C(_1574_),
    .Y(_1605_));
 sg13g2_a221oi_1 _5793_ (.B2(_0859_),
    .C1(_1605_),
    .B1(_1590_),
    .A1(net2068),
    .Y(_1606_),
    .A2(_1578_));
 sg13g2_nand3_1 _5794_ (.B(_1604_),
    .C(_1606_),
    .A(_1572_),
    .Y(_1607_));
 sg13g2_nand3_1 _5795_ (.B(_1603_),
    .C(_1607_),
    .A(net2025),
    .Y(_1608_));
 sg13g2_o21ai_1 _5796_ (.B1(_1608_),
    .Y(_1609_),
    .A1(net2025),
    .A2(_0027_));
 sg13g2_nand2_1 _5797_ (.Y(_1610_),
    .A(_1141_),
    .B(_1609_));
 sg13g2_nor2_1 _5798_ (.A(_1584_),
    .B(_1610_),
    .Y(_1611_));
 sg13g2_nor3_1 _5799_ (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .B(_1584_),
    .C(_1610_),
    .Y(_1612_));
 sg13g2_o21ai_1 _5800_ (.B1(net1988),
    .Y(_1613_),
    .A1(\z80.tv80s.i_tv80_core.Alternate ),
    .A2(_1611_));
 sg13g2_o21ai_1 _5801_ (.B1(_1542_),
    .Y(_0306_),
    .A1(_1612_),
    .A2(_1613_));
 sg13g2_nand2_1 _5802_ (.Y(_1614_),
    .A(net187),
    .B(net1976));
 sg13g2_and2_1 _5803_ (.A(net2119),
    .B(_1373_),
    .X(_1615_));
 sg13g2_o21ai_1 _5804_ (.B1(net2075),
    .Y(_1616_),
    .A1(_1268_),
    .A2(_1615_));
 sg13g2_nor3_1 _5805_ (.A(_1136_),
    .B(_1369_),
    .C(_1548_),
    .Y(_1617_));
 sg13g2_nor2_1 _5806_ (.A(net1843),
    .B(_1617_),
    .Y(_1618_));
 sg13g2_nor2_1 _5807_ (.A(net2112),
    .B(_1245_),
    .Y(_1619_));
 sg13g2_o21ai_1 _5808_ (.B1(_1550_),
    .Y(_1620_),
    .A1(net2112),
    .A2(_1245_));
 sg13g2_or2_1 _5809_ (.X(_1621_),
    .B(_1620_),
    .A(_1257_));
 sg13g2_a22oi_1 _5810_ (.Y(_1622_),
    .B1(_0933_),
    .B2(_1589_),
    .A2(net1888),
    .A1(_0906_));
 sg13g2_nor2_1 _5811_ (.A(_1557_),
    .B(_1622_),
    .Y(_1623_));
 sg13g2_a21oi_1 _5812_ (.A1(_0026_),
    .A2(net1864),
    .Y(_1624_),
    .B1(_1553_));
 sg13g2_nor3_1 _5813_ (.A(_1621_),
    .B(_1623_),
    .C(_1624_),
    .Y(_1625_));
 sg13g2_o21ai_1 _5814_ (.B1(_1625_),
    .Y(_1626_),
    .A1(_1616_),
    .A2(_1618_));
 sg13g2_nand2_1 _5815_ (.Y(_1627_),
    .A(net2169),
    .B(_1626_));
 sg13g2_nor3_2 _5816_ (.A(net2124),
    .B(net2113),
    .C(_1230_),
    .Y(_1628_));
 sg13g2_nand3_1 _5817_ (.B(net1864),
    .C(_1628_),
    .A(net2072),
    .Y(_1629_));
 sg13g2_nor2_1 _5818_ (.A(net2023),
    .B(_1200_),
    .Y(_1630_));
 sg13g2_nand2b_1 _5819_ (.Y(_1631_),
    .B(_0025_),
    .A_N(net2107));
 sg13g2_and3_1 _5820_ (.X(_1632_),
    .A(net1942),
    .B(_1630_),
    .C(_1631_));
 sg13g2_nand3_1 _5821_ (.B(_1630_),
    .C(_1631_),
    .A(net1942),
    .Y(_1633_));
 sg13g2_a21oi_1 _5822_ (.A1(_0904_),
    .A2(_1632_),
    .Y(_1634_),
    .B1(_1573_));
 sg13g2_a22oi_1 _5823_ (.Y(_1635_),
    .B1(_1629_),
    .B2(_1634_),
    .A2(_1627_),
    .A1(_1543_));
 sg13g2_nand2_1 _5824_ (.Y(_1636_),
    .A(net2063),
    .B(_1034_));
 sg13g2_and2_1 _5825_ (.A(net2063),
    .B(_1034_),
    .X(_1637_));
 sg13g2_o21ai_1 _5826_ (.B1(_1268_),
    .Y(_1638_),
    .A1(_1548_),
    .A2(_1636_));
 sg13g2_nor2b_1 _5827_ (.A(net2125),
    .B_N(net2063),
    .Y(_1639_));
 sg13g2_nand2_1 _5828_ (.Y(_1640_),
    .A(net2068),
    .B(net2018));
 sg13g2_a21oi_1 _5829_ (.A1(net2116),
    .A2(_1639_),
    .Y(_1641_),
    .B1(_1034_));
 sg13g2_nor3_1 _5830_ (.A(net2061),
    .B(net1883),
    .C(_1641_),
    .Y(_1642_));
 sg13g2_nor3_1 _5831_ (.A(_1594_),
    .B(_1620_),
    .C(_1642_),
    .Y(_1643_));
 sg13g2_nor3_1 _5832_ (.A(_0924_),
    .B(_1038_),
    .C(_1351_),
    .Y(_1644_));
 sg13g2_a22oi_1 _5833_ (.Y(_1645_),
    .B1(_1644_),
    .B2(net1943),
    .A2(_1615_),
    .A1(net2068));
 sg13g2_nor2_1 _5834_ (.A(net1943),
    .B(_1014_),
    .Y(_1646_));
 sg13g2_nand2_2 _5835_ (.Y(_1647_),
    .A(net2019),
    .B(_0933_));
 sg13g2_nor2b_1 _5836_ (.A(net2120),
    .B_N(net2066),
    .Y(_1648_));
 sg13g2_nor2_1 _5837_ (.A(_0838_),
    .B(_1648_),
    .Y(_1649_));
 sg13g2_o21ai_1 _5838_ (.B1(_1509_),
    .Y(_1650_),
    .A1(_1647_),
    .A2(_1649_));
 sg13g2_a221oi_1 _5839_ (.B2(_1650_),
    .C1(_1257_),
    .B1(_1558_),
    .A1(_0870_),
    .Y(_1651_),
    .A2(net1882));
 sg13g2_nand4_1 _5840_ (.B(_1643_),
    .C(_1645_),
    .A(net1844),
    .Y(_1652_),
    .D(_1651_));
 sg13g2_nand3_1 _5841_ (.B(_1638_),
    .C(_1652_),
    .A(net2169),
    .Y(_1653_));
 sg13g2_nor2_2 _5842_ (.A(_0860_),
    .B(net1942),
    .Y(_1654_));
 sg13g2_nand2_1 _5843_ (.Y(_1655_),
    .A(_0859_),
    .B(_0870_));
 sg13g2_a221oi_1 _5844_ (.B2(_1628_),
    .C1(_1654_),
    .B1(_1637_),
    .A1(_0838_),
    .Y(_1656_),
    .A2(_1632_));
 sg13g2_a22oi_1 _5845_ (.Y(_1657_),
    .B1(_1656_),
    .B2(_1570_),
    .A2(_1653_),
    .A1(_1585_));
 sg13g2_nand2_2 _5846_ (.Y(_1658_),
    .A(_1141_),
    .B(_1657_));
 sg13g2_nor2_1 _5847_ (.A(_1635_),
    .B(_1658_),
    .Y(_1659_));
 sg13g2_nor3_1 _5848_ (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .B(_1635_),
    .C(_1658_),
    .Y(_1660_));
 sg13g2_o21ai_1 _5849_ (.B1(net1991),
    .Y(_1661_),
    .A1(\z80.tv80s.i_tv80_core.Alternate ),
    .A2(_1659_));
 sg13g2_o21ai_1 _5850_ (.B1(_1614_),
    .Y(_0307_),
    .A1(_1660_),
    .A2(_1661_));
 sg13g2_nand4_1 _5851_ (.B(_0983_),
    .C(_1498_),
    .A(_0909_),
    .Y(_1662_),
    .D(_1500_));
 sg13g2_o21ai_1 _5852_ (.B1(_1511_),
    .Y(_1663_),
    .A1(net2082),
    .A2(_1233_));
 sg13g2_nor4_1 _5853_ (.A(_0972_),
    .B(net1884),
    .C(_1662_),
    .D(_1663_),
    .Y(_1664_));
 sg13g2_nand2_1 _5854_ (.Y(_1665_),
    .A(_1241_),
    .B(_1664_));
 sg13g2_nand2_2 _5855_ (.Y(_1666_),
    .A(_1503_),
    .B(_1510_));
 sg13g2_nor4_2 _5856_ (.A(_1430_),
    .B(_1504_),
    .C(_1665_),
    .Y(_1667_),
    .D(_1666_));
 sg13g2_nand2_2 _5857_ (.Y(_1668_),
    .A(_0965_),
    .B(_1234_));
 sg13g2_a21oi_2 _5858_ (.B1(_1001_),
    .Y(_1669_),
    .A2(net1886),
    .A1(net2002));
 sg13g2_nand4_1 _5859_ (.B(_1392_),
    .C(_1552_),
    .A(net2170),
    .Y(_1670_),
    .D(_1669_));
 sg13g2_nor3_1 _5860_ (.A(_1163_),
    .B(_1668_),
    .C(_1670_),
    .Y(_1671_));
 sg13g2_nand3_1 _5861_ (.B(_1667_),
    .C(_1671_),
    .A(_1254_),
    .Y(_1672_));
 sg13g2_nand2_2 _5862_ (.Y(_1673_),
    .A(net1952),
    .B(net1922));
 sg13g2_nor2_1 _5863_ (.A(_1110_),
    .B(_1673_),
    .Y(_1674_));
 sg13g2_nor2_1 _5864_ (.A(net1980),
    .B(_1674_),
    .Y(_1675_));
 sg13g2_a22oi_1 _5865_ (.Y(_0308_),
    .B1(_1672_),
    .B2(_1675_),
    .A2(net1980),
    .A1(_0800_));
 sg13g2_a22oi_1 _5866_ (.Y(_1676_),
    .B1(_1289_),
    .B2(_1390_),
    .A2(_0984_),
    .A1(net1946));
 sg13g2_nor2_1 _5867_ (.A(net2127),
    .B(_0998_),
    .Y(_1677_));
 sg13g2_a21oi_1 _5868_ (.A1(_0934_),
    .A2(_0998_),
    .Y(_1678_),
    .B1(_1095_));
 sg13g2_a221oi_1 _5869_ (.B2(_1390_),
    .C1(_1678_),
    .B1(_1289_),
    .A1(net1946),
    .Y(_1679_),
    .A2(_0984_));
 sg13g2_o21ai_1 _5870_ (.B1(_1593_),
    .Y(_1680_),
    .A1(_1004_),
    .A2(_1296_));
 sg13g2_a221oi_1 _5871_ (.B2(_1000_),
    .C1(_1680_),
    .B1(_1024_),
    .A1(net2075),
    .Y(_1681_),
    .A2(net1881));
 sg13g2_a221oi_1 _5872_ (.B2(_1681_),
    .C1(net2016),
    .B1(_1679_),
    .A1(_1026_),
    .Y(_1682_),
    .A2(_1439_));
 sg13g2_nor2_1 _5873_ (.A(_1095_),
    .B(_1189_),
    .Y(_1683_));
 sg13g2_nand2_1 _5874_ (.Y(_1684_),
    .A(net1952),
    .B(_1683_));
 sg13g2_nor2_2 _5875_ (.A(net1891),
    .B(_1423_),
    .Y(_1685_));
 sg13g2_nand2_2 _5876_ (.Y(_1686_),
    .A(_1104_),
    .B(_1685_));
 sg13g2_nand2_2 _5877_ (.Y(_1687_),
    .A(_1684_),
    .B(_1686_));
 sg13g2_and2_1 _5878_ (.A(_0879_),
    .B(_1685_),
    .X(_1688_));
 sg13g2_nor2_2 _5879_ (.A(_1682_),
    .B(_1687_),
    .Y(_1689_));
 sg13g2_a21o_1 _5880_ (.A2(net1881),
    .A1(net2080),
    .B1(_1680_),
    .X(_1690_));
 sg13g2_a21oi_1 _5881_ (.A1(_1000_),
    .A2(_1024_),
    .Y(_1691_),
    .B1(_1690_));
 sg13g2_a221oi_1 _5882_ (.B2(_1000_),
    .C1(_1690_),
    .B1(_1024_),
    .A1(net2023),
    .Y(_1692_),
    .A2(net1881));
 sg13g2_a221oi_1 _5883_ (.B2(_1692_),
    .C1(net2016),
    .B1(_1679_),
    .A1(_1026_),
    .Y(_1693_),
    .A2(_1439_));
 sg13g2_nor2_1 _5884_ (.A(net1952),
    .B(_1693_),
    .Y(_1694_));
 sg13g2_nor3_2 _5885_ (.A(_0858_),
    .B(net1890),
    .C(_1423_),
    .Y(_1695_));
 sg13g2_nor3_1 _5886_ (.A(net1891),
    .B(_1683_),
    .C(_1695_),
    .Y(_1696_));
 sg13g2_nand2b_1 _5887_ (.Y(_1697_),
    .B(_1104_),
    .A_N(_1066_));
 sg13g2_a22oi_1 _5888_ (.Y(_1698_),
    .B1(net1922),
    .B2(_0868_),
    .A2(_1109_),
    .A1(net1946));
 sg13g2_nand3_1 _5889_ (.B(_1697_),
    .C(_1698_),
    .A(_1696_),
    .Y(_1699_));
 sg13g2_nor2b_2 _5890_ (.A(_1694_),
    .B_N(_1699_),
    .Y(_1700_));
 sg13g2_o21ai_1 _5891_ (.B1(_1699_),
    .Y(_1701_),
    .A1(net1952),
    .A2(_1693_));
 sg13g2_nand2_1 _5892_ (.Y(_1702_),
    .A(net2020),
    .B(_0031_));
 sg13g2_a21oi_2 _5893_ (.B1(_0688_),
    .Y(_1703_),
    .A2(net2142),
    .A1(net2123));
 sg13g2_or2_1 _5894_ (.X(_1704_),
    .B(_1703_),
    .A(_1140_));
 sg13g2_a21oi_2 _5895_ (.B1(_1704_),
    .Y(_1705_),
    .A2(_1701_),
    .A1(_0031_));
 sg13g2_a21o_2 _5896_ (.A2(_1701_),
    .A1(_0031_),
    .B1(_1704_),
    .X(_1706_));
 sg13g2_and2_1 _5897_ (.A(_1689_),
    .B(_1705_),
    .X(_1707_));
 sg13g2_nand2_2 _5898_ (.Y(_1708_),
    .A(_1689_),
    .B(_1705_));
 sg13g2_a21oi_1 _5899_ (.A1(_0942_),
    .A2(_0948_),
    .Y(_1709_),
    .B1(net1884));
 sg13g2_o21ai_1 _5900_ (.B1(_1006_),
    .Y(_1710_),
    .A1(_0943_),
    .A2(_0949_));
 sg13g2_nor4_2 _5901_ (.A(_0945_),
    .B(_0972_),
    .C(_1529_),
    .Y(_1711_),
    .D(_1710_));
 sg13g2_and3_1 _5902_ (.X(_1712_),
    .A(_1146_),
    .B(_1169_),
    .C(_1711_));
 sg13g2_nor3_1 _5903_ (.A(net1951),
    .B(_0930_),
    .C(_1172_),
    .Y(_1713_));
 sg13g2_and2_1 _5904_ (.A(_0922_),
    .B(_1713_),
    .X(_1714_));
 sg13g2_nand2_1 _5905_ (.Y(_1715_),
    .A(_1712_),
    .B(_1714_));
 sg13g2_and4_2 _5906_ (.A(_1495_),
    .B(_1533_),
    .C(_1712_),
    .D(_1714_),
    .X(_1716_));
 sg13g2_nor2_2 _5907_ (.A(_0966_),
    .B(_1301_),
    .Y(_1717_));
 sg13g2_nand4_1 _5908_ (.B(_0928_),
    .C(_1716_),
    .A(net2144),
    .Y(_1718_),
    .D(_1717_));
 sg13g2_and4_2 _5909_ (.A(\z80.tv80s.i_tv80_core.ts[4] ),
    .B(_0928_),
    .C(_1716_),
    .D(_1717_),
    .X(_1719_));
 sg13g2_nand4_1 _5910_ (.B(_0928_),
    .C(_1716_),
    .A(\z80.tv80s.i_tv80_core.ts[4] ),
    .Y(_1720_),
    .D(_1717_));
 sg13g2_o21ai_1 _5911_ (.B1(net1829),
    .Y(_1721_),
    .A1(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .A2(_1719_));
 sg13g2_a221oi_1 _5912_ (.B2(_1000_),
    .C1(_1680_),
    .B1(_1024_),
    .A1(net2068),
    .Y(_1722_),
    .A2(net1881));
 sg13g2_a221oi_1 _5913_ (.B2(_1722_),
    .C1(net2016),
    .B1(_1679_),
    .A1(_1026_),
    .Y(_1723_),
    .A2(_1439_));
 sg13g2_nor3_2 _5914_ (.A(net1890),
    .B(net1945),
    .C(_1095_),
    .Y(_1724_));
 sg13g2_a21oi_1 _5915_ (.A1(_0879_),
    .A2(net1922),
    .Y(_1725_),
    .B1(_1724_));
 sg13g2_nand2_1 _5916_ (.Y(_1726_),
    .A(_1696_),
    .B(_1725_));
 sg13g2_o21ai_1 _5917_ (.B1(_1726_),
    .Y(_1727_),
    .A1(net1952),
    .A2(_1723_));
 sg13g2_nor3_2 _5918_ (.A(_1682_),
    .B(_1687_),
    .C(_1703_),
    .Y(_1728_));
 sg13g2_or3_2 _5919_ (.A(_1682_),
    .B(_1687_),
    .C(_1703_),
    .X(_1729_));
 sg13g2_nand2b_1 _5920_ (.Y(_1730_),
    .B(_1728_),
    .A_N(net1824));
 sg13g2_and3_1 _5921_ (.X(_1731_),
    .A(_1706_),
    .B(_1721_),
    .C(_1730_));
 sg13g2_nand3_1 _5922_ (.B(_1721_),
    .C(_1730_),
    .A(_1706_),
    .Y(_1732_));
 sg13g2_nor2_2 _5923_ (.A(_1707_),
    .B(_1731_),
    .Y(_1733_));
 sg13g2_nand2_1 _5924_ (.Y(_1734_),
    .A(_1708_),
    .B(_1732_));
 sg13g2_nand2_2 _5925_ (.Y(_1735_),
    .A(_1705_),
    .B(net1824));
 sg13g2_nand2_1 _5926_ (.Y(_1736_),
    .A(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .B(net1826));
 sg13g2_nand4_1 _5927_ (.B(net1829),
    .C(_1730_),
    .A(_1706_),
    .Y(_1737_),
    .D(_1736_));
 sg13g2_and2_1 _5928_ (.A(net1829),
    .B(net1826),
    .X(_1738_));
 sg13g2_nand2_1 _5929_ (.Y(_1739_),
    .A(net1829),
    .B(net1825));
 sg13g2_o21ai_1 _5930_ (.B1(_0695_),
    .Y(_1740_),
    .A1(net1824),
    .A2(_1729_));
 sg13g2_nand3b_1 _5931_ (.B(_1728_),
    .C(_0696_),
    .Y(_1741_),
    .A_N(net1824));
 sg13g2_or3_1 _5932_ (.A(_0696_),
    .B(net1824),
    .C(_1729_),
    .X(_1742_));
 sg13g2_o21ai_1 _5933_ (.B1(_0040_),
    .Y(_1743_),
    .A1(net1824),
    .A2(_1729_));
 sg13g2_nand4_1 _5934_ (.B(_1738_),
    .C(_1740_),
    .A(_1706_),
    .Y(_1744_),
    .D(_1741_));
 sg13g2_o21ai_1 _5935_ (.B1(_0020_),
    .Y(_1745_),
    .A1(_1705_),
    .A2(_1739_));
 sg13g2_nand4_1 _5936_ (.B(_1738_),
    .C(_1742_),
    .A(_1706_),
    .Y(_1746_),
    .D(_1743_));
 sg13g2_a21o_1 _5937_ (.A2(_1738_),
    .A1(_1706_),
    .B1(_0020_),
    .X(_1747_));
 sg13g2_nand4_1 _5938_ (.B(_1737_),
    .C(_1744_),
    .A(_1735_),
    .Y(_1748_),
    .D(_1745_));
 sg13g2_nor2_2 _5939_ (.A(net1765),
    .B(_1748_),
    .Y(_1749_));
 sg13g2_or2_1 _5940_ (.X(_1750_),
    .B(_1727_),
    .A(_1689_));
 sg13g2_nand2_2 _5941_ (.Y(_1751_),
    .A(net2123),
    .B(_0023_));
 sg13g2_nand2_1 _5942_ (.Y(_1752_),
    .A(net2020),
    .B(net1997));
 sg13g2_nand4_1 _5943_ (.B(_1750_),
    .C(_1751_),
    .A(_1700_),
    .Y(_1753_),
    .D(_1752_));
 sg13g2_and2_1 _5944_ (.A(_1738_),
    .B(_1753_),
    .X(_1754_));
 sg13g2_nor2_1 _5945_ (.A(_0790_),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .Y(_1755_));
 sg13g2_nand2_1 _5946_ (.Y(_1756_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .B(_1755_));
 sg13g2_nor2_1 _5947_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .B(_1756_),
    .Y(_1757_));
 sg13g2_nor2_1 _5948_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .Y(_1758_));
 sg13g2_o21ai_1 _5949_ (.B1(_0790_),
    .Y(_1759_),
    .A1(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .A2(_1758_));
 sg13g2_a21oi_1 _5950_ (.A1(_0228_),
    .A2(_1758_),
    .Y(_1760_),
    .B1(_1759_));
 sg13g2_a21oi_1 _5951_ (.A1(_0791_),
    .A2(_1760_),
    .Y(_1761_),
    .B1(_1757_));
 sg13g2_and2_1 _5952_ (.A(net2041),
    .B(net2038),
    .X(_1762_));
 sg13g2_nand2_2 _5953_ (.Y(_1763_),
    .A(net2040),
    .B(net2038));
 sg13g2_nand3_1 _5954_ (.B(net2036),
    .C(_1762_),
    .A(_0778_),
    .Y(_1764_));
 sg13g2_nor2_1 _5955_ (.A(_0683_),
    .B(net2033),
    .Y(_1765_));
 sg13g2_a22oi_1 _5956_ (.Y(_1766_),
    .B1(_1765_),
    .B2(_0227_),
    .A2(_1764_),
    .A1(net2033));
 sg13g2_nor2_2 _5957_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .B(_1766_),
    .Y(_1767_));
 sg13g2_nand2b_2 _5958_ (.Y(_1768_),
    .B(_1767_),
    .A_N(_1761_));
 sg13g2_a21oi_2 _5959_ (.B1(net1961),
    .Y(_1769_),
    .A2(_1768_),
    .A1(_1754_));
 sg13g2_and2_2 _5960_ (.A(net1748),
    .B(_1769_),
    .X(_1770_));
 sg13g2_and3_2 _5961_ (.X(_1771_),
    .A(_1700_),
    .B(_1702_),
    .C(_1751_));
 sg13g2_nand3_1 _5962_ (.B(_1702_),
    .C(_1751_),
    .A(_1700_),
    .Y(_1772_));
 sg13g2_nor4_1 _5963_ (.A(_1172_),
    .B(_1265_),
    .C(_1497_),
    .D(_1512_),
    .Y(_1773_));
 sg13g2_nand4_1 _5964_ (.B(_1533_),
    .C(_1712_),
    .A(_1520_),
    .Y(_1774_),
    .D(_1773_));
 sg13g2_nor2_2 _5965_ (.A(_1238_),
    .B(_1774_),
    .Y(_1775_));
 sg13g2_nor2_1 _5966_ (.A(_0778_),
    .B(net2036),
    .Y(_1776_));
 sg13g2_nand2_2 _5967_ (.Y(_1777_),
    .A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0779_));
 sg13g2_nand3_1 _5968_ (.B(net2036),
    .C(_1763_),
    .A(net2034),
    .Y(_1778_));
 sg13g2_o21ai_1 _5969_ (.B1(net2035),
    .Y(_1779_),
    .A1(_0779_),
    .A2(_1763_));
 sg13g2_nand2_2 _5970_ (.Y(_1780_),
    .A(_1777_),
    .B(_1778_));
 sg13g2_xnor2_1 _5971_ (.Y(_1781_),
    .A(net2039),
    .B(\z80.tv80s.i_tv80_core.BusB[0] ));
 sg13g2_nor2_1 _5972_ (.A(_0212_),
    .B(_1781_),
    .Y(_1782_));
 sg13g2_xor2_1 _5973_ (.B(_1781_),
    .A(_0212_),
    .X(_1783_));
 sg13g2_nand3b_1 _5974_ (.B(net2040),
    .C(net2151),
    .Y(_1784_),
    .A_N(net2036));
 sg13g2_xnor2_1 _5975_ (.Y(_1785_),
    .A(_0789_),
    .B(_1784_));
 sg13g2_and2_1 _5976_ (.A(_1783_),
    .B(_1785_),
    .X(_1786_));
 sg13g2_nand2_1 _5977_ (.Y(_1787_),
    .A(net2040),
    .B(_0789_));
 sg13g2_a22oi_1 _5978_ (.Y(_1788_),
    .B1(_1763_),
    .B2(_0779_),
    .A2(_0789_),
    .A1(net2040));
 sg13g2_o21ai_1 _5979_ (.B1(_1787_),
    .Y(_1789_),
    .A1(net2036),
    .A2(_1762_));
 sg13g2_nor2_1 _5980_ (.A(_1783_),
    .B(_1785_),
    .Y(_1790_));
 sg13g2_nor3_1 _5981_ (.A(_1786_),
    .B(net1873),
    .C(_1790_),
    .Y(_1791_));
 sg13g2_and2_1 _5982_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_1792_));
 sg13g2_nand2_2 _5983_ (.Y(_1793_),
    .A(net2039),
    .B(net1873));
 sg13g2_nand2_2 _5984_ (.Y(_1794_),
    .A(net2040),
    .B(_0780_));
 sg13g2_nor2_2 _5985_ (.A(_0226_),
    .B(_1794_),
    .Y(_1795_));
 sg13g2_o21ai_1 _5986_ (.B1(_1793_),
    .Y(_1796_),
    .A1(_0226_),
    .A2(_1794_));
 sg13g2_nor2_2 _5987_ (.A(net2040),
    .B(net2038),
    .Y(_1797_));
 sg13g2_or2_2 _5988_ (.X(_1798_),
    .B(net2038),
    .A(net2040));
 sg13g2_nor2_2 _5989_ (.A(_0226_),
    .B(_1798_),
    .Y(_1799_));
 sg13g2_nand2b_1 _5990_ (.Y(_1800_),
    .B(_1797_),
    .A_N(_0226_));
 sg13g2_nand2_2 _5991_ (.Y(_1801_),
    .A(_1793_),
    .B(_1800_));
 sg13g2_xor2_1 _5992_ (.B(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(_1802_));
 sg13g2_a221oi_1 _5993_ (.B2(_1796_),
    .C1(_1791_),
    .B1(_1802_),
    .A1(_1792_),
    .Y(_1803_),
    .A2(_1801_));
 sg13g2_nand2_2 _5994_ (.Y(_1804_),
    .A(_1776_),
    .B(_1797_));
 sg13g2_nor2_1 _5995_ (.A(net2062),
    .B(_1051_),
    .Y(_1805_));
 sg13g2_o21ai_1 _5996_ (.B1(net1864),
    .Y(_1806_),
    .A1(net2024),
    .A2(_0209_));
 sg13g2_a221oi_1 _5997_ (.B2(_0781_),
    .C1(_1806_),
    .B1(_1805_),
    .A1(net2151),
    .Y(_1807_),
    .A2(net1880));
 sg13g2_nor2_2 _5998_ (.A(_1778_),
    .B(_1797_),
    .Y(_1808_));
 sg13g2_nand2b_2 _5999_ (.Y(_1809_),
    .B(_1798_),
    .A_N(_1778_));
 sg13g2_mux2_2 _6000_ (.A0(_0217_),
    .A1(_0221_),
    .S(net2042),
    .X(_1810_));
 sg13g2_nor2_1 _6001_ (.A(_1809_),
    .B(_1810_),
    .Y(_1811_));
 sg13g2_nor2_2 _6002_ (.A(_1777_),
    .B(_1794_),
    .Y(_1812_));
 sg13g2_or2_2 _6003_ (.X(_1813_),
    .B(_1794_),
    .A(_1777_));
 sg13g2_nor3_1 _6004_ (.A(net2062),
    .B(_0217_),
    .C(_1051_),
    .Y(_1814_));
 sg13g2_and2_1 _6005_ (.A(_1812_),
    .B(_1814_),
    .X(_1815_));
 sg13g2_nor3_2 _6006_ (.A(_0778_),
    .B(_0779_),
    .C(_1798_),
    .Y(_1816_));
 sg13g2_nand3_1 _6007_ (.B(net2036),
    .C(_1797_),
    .A(net2034),
    .Y(_1817_));
 sg13g2_o21ai_1 _6008_ (.B1(_1780_),
    .Y(_1818_),
    .A1(_0212_),
    .A2(_1817_));
 sg13g2_o21ai_1 _6009_ (.B1(_0217_),
    .Y(_1819_),
    .A1(net2062),
    .A2(_1051_));
 sg13g2_nor2_1 _6010_ (.A(net2040),
    .B(_0780_),
    .Y(_1820_));
 sg13g2_and2_2 _6011_ (.A(_1776_),
    .B(_1820_),
    .X(_1821_));
 sg13g2_inv_2 _6012_ (.Y(_1822_),
    .A(_1821_));
 sg13g2_nor2_2 _6013_ (.A(_1763_),
    .B(_1777_),
    .Y(_1823_));
 sg13g2_o21ai_1 _6014_ (.B1(_1823_),
    .Y(_1824_),
    .A1(net2062),
    .A2(_1051_));
 sg13g2_inv_1 _6015_ (.Y(_1825_),
    .A(_1824_));
 sg13g2_o21ai_1 _6016_ (.B1(_1819_),
    .Y(_1826_),
    .A1(_1821_),
    .A2(_1825_));
 sg13g2_o21ai_1 _6017_ (.B1(_1826_),
    .Y(_1827_),
    .A1(net1863),
    .A2(_1807_));
 sg13g2_nor4_1 _6018_ (.A(_1811_),
    .B(_1815_),
    .C(_1818_),
    .D(_1827_),
    .Y(_1828_));
 sg13g2_a21oi_1 _6019_ (.A1(net1874),
    .A2(_1803_),
    .Y(_1829_),
    .B1(_1828_));
 sg13g2_mux2_1 _6020_ (.A0(net2051),
    .A1(_1829_),
    .S(net2033),
    .X(_1830_));
 sg13g2_mux2_2 _6021_ (.A0(_1830_),
    .A1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .S(net1787),
    .X(_1831_));
 sg13g2_a21oi_1 _6022_ (.A1(net1789),
    .A2(_1831_),
    .Y(_1832_),
    .B1(_1719_));
 sg13g2_nand2_1 _6023_ (.Y(_1833_),
    .A(_0021_),
    .B(_1029_));
 sg13g2_nor2_1 _6024_ (.A(net2128),
    .B(_1833_),
    .Y(_1834_));
 sg13g2_inv_1 _6025_ (.Y(_1835_),
    .A(_1834_));
 sg13g2_a221oi_1 _6026_ (.B2(_1026_),
    .C1(net2015),
    .B1(_1835_),
    .A1(_1676_),
    .Y(_1836_),
    .A2(_1691_));
 sg13g2_nand2b_1 _6027_ (.Y(_1837_),
    .B(net2088),
    .A_N(net2120));
 sg13g2_nor2_1 _6028_ (.A(net2088),
    .B(net2120),
    .Y(_1838_));
 sg13g2_a21oi_2 _6029_ (.B1(_1838_),
    .Y(_1839_),
    .A2(_0034_),
    .A1(net2121));
 sg13g2_nor2_2 _6030_ (.A(net2081),
    .B(net2125),
    .Y(_1840_));
 sg13g2_or3_1 _6031_ (.A(_0861_),
    .B(_1110_),
    .C(_1840_),
    .X(_1841_));
 sg13g2_nor2_1 _6032_ (.A(net1942),
    .B(_1105_),
    .Y(_1842_));
 sg13g2_o21ai_1 _6033_ (.B1(_1839_),
    .Y(_1843_),
    .A1(_1724_),
    .A2(_1842_));
 sg13g2_a22oi_1 _6034_ (.Y(_1844_),
    .B1(_1695_),
    .B2(net2081),
    .A2(_1104_),
    .A1(net2124));
 sg13g2_and2_1 _6035_ (.A(_1843_),
    .B(_1844_),
    .X(_1845_));
 sg13g2_a21oi_2 _6036_ (.B1(net1892),
    .Y(_1846_),
    .A2(_1845_),
    .A1(_1841_));
 sg13g2_or2_2 _6037_ (.X(_1847_),
    .B(_1846_),
    .A(_1836_));
 sg13g2_inv_1 _6038_ (.Y(_1848_),
    .A(net1823));
 sg13g2_nor2_1 _6039_ (.A(net1764),
    .B(_1748_),
    .Y(_1849_));
 sg13g2_a22oi_1 _6040_ (.Y(_1850_),
    .B1(_1744_),
    .B2(_1745_),
    .A2(_1737_),
    .A1(_1735_));
 sg13g2_and2_1 _6041_ (.A(net1765),
    .B(_1850_),
    .X(_1851_));
 sg13g2_nand3_1 _6042_ (.B(net1765),
    .C(_1850_),
    .A(_0078_),
    .Y(_1852_));
 sg13g2_and4_2 _6043_ (.A(_1735_),
    .B(_1737_),
    .C(_1746_),
    .D(_1747_),
    .X(_1853_));
 sg13g2_nand4_1 _6044_ (.B(_1737_),
    .C(_1746_),
    .A(_1735_),
    .Y(_1854_),
    .D(_1747_));
 sg13g2_nor2_2 _6045_ (.A(net1764),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_nand3_1 _6046_ (.B(net1765),
    .C(_1853_),
    .A(_0080_),
    .Y(_1856_));
 sg13g2_a22oi_1 _6047_ (.Y(_1857_),
    .B1(_1746_),
    .B2(_1747_),
    .A2(_1737_),
    .A1(_1735_));
 sg13g2_and2_1 _6048_ (.A(_1733_),
    .B(_1857_),
    .X(_1858_));
 sg13g2_nand3_1 _6049_ (.B(net1765),
    .C(_1857_),
    .A(_0082_),
    .Y(_1859_));
 sg13g2_nor2_1 _6050_ (.A(_1733_),
    .B(_1854_),
    .Y(_1860_));
 sg13g2_and2_2 _6051_ (.A(_1734_),
    .B(_1850_),
    .X(_1861_));
 sg13g2_and2_1 _6052_ (.A(net1764),
    .B(_1857_),
    .X(_1862_));
 sg13g2_nand3_1 _6053_ (.B(net1764),
    .C(_1857_),
    .A(_0081_),
    .Y(_1863_));
 sg13g2_a22oi_1 _6054_ (.Y(_1864_),
    .B1(net1737),
    .B2(_0077_),
    .A2(net1739),
    .A1(_0079_));
 sg13g2_a22oi_1 _6055_ (.Y(_1865_),
    .B1(net1747),
    .B2(_0084_),
    .A2(net1749),
    .A1(_0083_));
 sg13g2_and4_1 _6056_ (.A(_1852_),
    .B(_1856_),
    .C(_1859_),
    .D(_1863_),
    .X(_1866_));
 sg13g2_nand3_1 _6057_ (.B(_1865_),
    .C(_1866_),
    .A(_1864_),
    .Y(_1867_));
 sg13g2_xnor2_1 _6058_ (.Y(_1868_),
    .A(net1822),
    .B(_1867_));
 sg13g2_o21ai_1 _6059_ (.B1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .Y(_1869_),
    .A1(_1707_),
    .A2(_1731_));
 sg13g2_nand3_1 _6060_ (.B(_1708_),
    .C(_1732_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .Y(_1870_));
 sg13g2_a21o_1 _6061_ (.A2(_1870_),
    .A1(_1869_),
    .B1(_1748_),
    .X(_1871_));
 sg13g2_a21oi_1 _6062_ (.A1(_1708_),
    .A2(_1732_),
    .Y(_1872_),
    .B1(_0700_));
 sg13g2_and3_1 _6063_ (.X(_1873_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .B(_1708_),
    .C(_1732_));
 sg13g2_o21ai_1 _6064_ (.B1(_1857_),
    .Y(_1874_),
    .A1(_1872_),
    .A2(_1873_));
 sg13g2_o21ai_1 _6065_ (.B1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .Y(_1875_),
    .A1(_1707_),
    .A2(_1731_));
 sg13g2_nand3_1 _6066_ (.B(_1708_),
    .C(_1732_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .Y(_1876_));
 sg13g2_a21o_1 _6067_ (.A2(_1876_),
    .A1(_1875_),
    .B1(_1854_),
    .X(_1877_));
 sg13g2_a21oi_1 _6068_ (.A1(_1708_),
    .A2(_1732_),
    .Y(_1878_),
    .B1(_0699_));
 sg13g2_and3_1 _6069_ (.X(_1879_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .B(_1708_),
    .C(_1732_));
 sg13g2_o21ai_1 _6070_ (.B1(_1850_),
    .Y(_1880_),
    .A1(_1878_),
    .A2(_1879_));
 sg13g2_nand4_1 _6071_ (.B(_1874_),
    .C(_1877_),
    .A(_1871_),
    .Y(_1881_),
    .D(_1880_));
 sg13g2_nand2_1 _6072_ (.Y(_1882_),
    .A(net1823),
    .B(_1881_));
 sg13g2_a22oi_1 _6073_ (.Y(_1883_),
    .B1(net1737),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .A2(net1743),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ));
 sg13g2_a22oi_1 _6074_ (.Y(_1884_),
    .B1(net1741),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A2(net1749),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ));
 sg13g2_a22oi_1 _6075_ (.Y(_1885_),
    .B1(net1739),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .A2(net1745),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ));
 sg13g2_a22oi_1 _6076_ (.Y(_1886_),
    .B1(net1735),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .A2(net1747),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ));
 sg13g2_and4_2 _6077_ (.A(_1883_),
    .B(_1884_),
    .C(_1885_),
    .D(_1886_),
    .X(_1887_));
 sg13g2_nand4_1 _6078_ (.B(_1884_),
    .C(_1885_),
    .A(_1883_),
    .Y(_1888_),
    .D(_1886_));
 sg13g2_xnor2_1 _6079_ (.Y(_1889_),
    .A(net1822),
    .B(_1881_));
 sg13g2_nand2b_1 _6080_ (.Y(_1890_),
    .B(_1888_),
    .A_N(_1889_));
 sg13g2_o21ai_1 _6081_ (.B1(_1882_),
    .Y(_1891_),
    .A1(_1887_),
    .A2(_1889_));
 sg13g2_a22oi_1 _6082_ (.Y(_1892_),
    .B1(net1747),
    .B2(_0068_),
    .A2(net1749),
    .A1(_0067_));
 sg13g2_nand2_1 _6083_ (.Y(_1893_),
    .A(_0065_),
    .B(net1735));
 sg13g2_and3_1 _6084_ (.X(_1894_),
    .A(_0066_),
    .B(_1733_),
    .C(_1857_));
 sg13g2_a22oi_1 _6085_ (.Y(_1895_),
    .B1(net1737),
    .B2(_0061_),
    .A2(net1743),
    .A1(_0064_));
 sg13g2_a221oi_1 _6086_ (.B2(_0063_),
    .C1(_1894_),
    .B1(net1739),
    .A1(_0062_),
    .Y(_1896_),
    .A2(net1745));
 sg13g2_nand4_1 _6087_ (.B(_1893_),
    .C(_1895_),
    .A(_1892_),
    .Y(_1897_),
    .D(_1896_));
 sg13g2_nor2_1 _6088_ (.A(net1817),
    .B(_1897_),
    .Y(_1898_));
 sg13g2_xnor2_1 _6089_ (.Y(_1899_),
    .A(net1822),
    .B(_1897_));
 sg13g2_xnor2_1 _6090_ (.Y(_1900_),
    .A(net1817),
    .B(_1897_));
 sg13g2_and2_1 _6091_ (.A(_1891_),
    .B(_1899_),
    .X(_1901_));
 sg13g2_nand3_1 _6092_ (.B(_1891_),
    .C(_1899_),
    .A(_1868_),
    .Y(_1902_));
 sg13g2_a21o_1 _6093_ (.A2(_1897_),
    .A1(_1867_),
    .B1(net1817),
    .X(_1903_));
 sg13g2_and2_1 _6094_ (.A(_1902_),
    .B(_1903_),
    .X(_1904_));
 sg13g2_a22oi_1 _6095_ (.Y(_1905_),
    .B1(net1735),
    .B2(_0145_),
    .A2(net1745),
    .A1(_0142_));
 sg13g2_nand2_1 _6096_ (.Y(_1906_),
    .A(_0144_),
    .B(net1743));
 sg13g2_nor3_1 _6097_ (.A(_0729_),
    .B(net1765),
    .C(_1854_),
    .Y(_1907_));
 sg13g2_a22oi_1 _6098_ (.Y(_1908_),
    .B1(net1737),
    .B2(_0141_),
    .A2(net1741),
    .A1(_0146_));
 sg13g2_a221oi_1 _6099_ (.B2(_0148_),
    .C1(_1907_),
    .B1(net1747),
    .A1(_0147_),
    .Y(_1909_),
    .A2(net1749));
 sg13g2_nand4_1 _6100_ (.B(_1906_),
    .C(_1908_),
    .A(_1905_),
    .Y(_1910_),
    .D(_1909_));
 sg13g2_xnor2_1 _6101_ (.Y(_1911_),
    .A(net1822),
    .B(_1910_));
 sg13g2_nand3_1 _6102_ (.B(net1764),
    .C(_1853_),
    .A(_0127_),
    .Y(_1912_));
 sg13g2_nand3_1 _6103_ (.B(net1765),
    .C(_1857_),
    .A(_0130_),
    .Y(_1913_));
 sg13g2_nand3_1 _6104_ (.B(net1764),
    .C(_1857_),
    .A(_0129_),
    .Y(_1914_));
 sg13g2_a22oi_1 _6105_ (.Y(_1915_),
    .B1(net1747),
    .B2(_0132_),
    .A2(net1749),
    .A1(_0131_));
 sg13g2_nand3_1 _6106_ (.B(net1765),
    .C(_1850_),
    .A(_0126_),
    .Y(_1916_));
 sg13g2_and4_1 _6107_ (.A(_1912_),
    .B(_1913_),
    .C(_1914_),
    .D(_1916_),
    .X(_1917_));
 sg13g2_a22oi_1 _6108_ (.Y(_1918_),
    .B1(net1737),
    .B2(_0125_),
    .A2(net1743),
    .A1(_0128_));
 sg13g2_nand3_1 _6109_ (.B(_1917_),
    .C(_1918_),
    .A(_1915_),
    .Y(_1919_));
 sg13g2_nand2b_1 _6110_ (.Y(_1920_),
    .B(net1822),
    .A_N(_1919_));
 sg13g2_xnor2_1 _6111_ (.Y(_1921_),
    .A(net1822),
    .B(_1919_));
 sg13g2_inv_1 _6112_ (.Y(_1922_),
    .A(_1921_));
 sg13g2_a22oi_1 _6113_ (.Y(_1923_),
    .B1(net1735),
    .B2(_0113_),
    .A2(net1737),
    .A1(_0109_));
 sg13g2_nand2_1 _6114_ (.Y(_1924_),
    .A(_0111_),
    .B(net1739));
 sg13g2_nor3_1 _6115_ (.A(_0716_),
    .B(net1764),
    .C(_1748_),
    .Y(_1925_));
 sg13g2_a22oi_1 _6116_ (.Y(_1926_),
    .B1(net1741),
    .B2(_0114_),
    .A2(net1743),
    .A1(_0112_));
 sg13g2_a221oi_1 _6117_ (.B2(_0110_),
    .C1(_1925_),
    .B1(net1745),
    .A1(_0115_),
    .Y(_1927_),
    .A2(net1749));
 sg13g2_nand4_1 _6118_ (.B(_1924_),
    .C(_1926_),
    .A(_1923_),
    .Y(_1928_),
    .D(_1927_));
 sg13g2_xnor2_1 _6119_ (.Y(_1929_),
    .A(net1822),
    .B(_1928_));
 sg13g2_a22oi_1 _6120_ (.Y(_1930_),
    .B1(net1739),
    .B2(_0095_),
    .A2(net1743),
    .A1(_0096_));
 sg13g2_nand2_1 _6121_ (.Y(_1931_),
    .A(_0097_),
    .B(net1735));
 sg13g2_nor3_1 _6122_ (.A(_0713_),
    .B(net1764),
    .C(_1748_),
    .Y(_1932_));
 sg13g2_a22oi_1 _6123_ (.Y(_1933_),
    .B1(net1741),
    .B2(_0098_),
    .A2(net1745),
    .A1(_0094_));
 sg13g2_a221oi_1 _6124_ (.B2(_0093_),
    .C1(_1932_),
    .B1(net1737),
    .A1(_0099_),
    .Y(_1934_),
    .A2(net1749));
 sg13g2_nand4_1 _6125_ (.B(_1931_),
    .C(_1933_),
    .A(_1930_),
    .Y(_1935_),
    .D(_1934_));
 sg13g2_nor2_1 _6126_ (.A(net1817),
    .B(_1935_),
    .Y(_1936_));
 sg13g2_xnor2_1 _6127_ (.Y(_1937_),
    .A(net1822),
    .B(_1935_));
 sg13g2_nand4_1 _6128_ (.B(_1921_),
    .C(_1929_),
    .A(_1911_),
    .Y(_1938_),
    .D(_1937_));
 sg13g2_a21oi_1 _6129_ (.A1(_1902_),
    .A2(_1903_),
    .Y(_1939_),
    .B1(_1938_));
 sg13g2_a21oi_1 _6130_ (.A1(_1928_),
    .A2(_1935_),
    .Y(_1940_),
    .B1(net1817));
 sg13g2_nand3_1 _6131_ (.B(_1921_),
    .C(_1940_),
    .A(_1911_),
    .Y(_1941_));
 sg13g2_a21oi_1 _6132_ (.A1(_1910_),
    .A2(_1919_),
    .Y(_1942_),
    .B1(net1817));
 sg13g2_nand2b_1 _6133_ (.Y(_1943_),
    .B(_1941_),
    .A_N(_1942_));
 sg13g2_nor2_1 _6134_ (.A(_1939_),
    .B(_1943_),
    .Y(_1944_));
 sg13g2_a22oi_1 _6135_ (.Y(_1945_),
    .B1(net1740),
    .B2(_0042_),
    .A2(net1747),
    .A1(_0044_));
 sg13g2_a22oi_1 _6136_ (.Y(_1946_),
    .B1(net1734),
    .B2(_0041_),
    .A2(net1736),
    .A1(_0035_));
 sg13g2_a22oi_1 _6137_ (.Y(_1947_),
    .B1(net1738),
    .B2(_0037_),
    .A2(net1748),
    .A1(_0043_));
 sg13g2_a22oi_1 _6138_ (.Y(_1948_),
    .B1(net1742),
    .B2(_0038_),
    .A2(net1744),
    .A1(_0036_));
 sg13g2_and2_1 _6139_ (.A(_1945_),
    .B(_1948_),
    .X(_1949_));
 sg13g2_nand3_1 _6140_ (.B(_1947_),
    .C(_1949_),
    .A(_1946_),
    .Y(_1950_));
 sg13g2_xnor2_1 _6141_ (.Y(_1951_),
    .A(net1817),
    .B(_1950_));
 sg13g2_inv_1 _6142_ (.Y(_1952_),
    .A(_1951_));
 sg13g2_o21ai_1 _6143_ (.B1(_1952_),
    .Y(_1953_),
    .A1(_1939_),
    .A2(_1943_));
 sg13g2_xnor2_1 _6144_ (.Y(_1954_),
    .A(_1944_),
    .B(_1951_));
 sg13g2_o21ai_1 _6145_ (.B1(_1832_),
    .Y(_1955_),
    .A1(_1772_),
    .A2(_1954_));
 sg13g2_and2_1 _6146_ (.A(net2009),
    .B(net1831),
    .X(_1956_));
 sg13g2_nand2_1 _6147_ (.Y(_1957_),
    .A(net2010),
    .B(net1831));
 sg13g2_nor2_1 _6148_ (.A(_0035_),
    .B(net1809),
    .Y(_1958_));
 sg13g2_nand2b_1 _6149_ (.Y(_1959_),
    .B(net1832),
    .A_N(_0150_));
 sg13g2_o21ai_1 _6150_ (.B1(_1959_),
    .Y(_1960_),
    .A1(_0020_),
    .A2(net1831));
 sg13g2_mux2_1 _6151_ (.A0(_0020_),
    .A1(_0150_),
    .S(net1831),
    .X(_1961_));
 sg13g2_and2_1 _6152_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(net1833),
    .X(_1962_));
 sg13g2_nand2_2 _6153_ (.Y(_1963_),
    .A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(net1833));
 sg13g2_mux4_1 _6154_ (.S0(net1814),
    .A0(_0042_),
    .A1(_0041_),
    .A2(_0044_),
    .A3(_0043_),
    .S1(net1800),
    .X(_1964_));
 sg13g2_o21ai_1 _6155_ (.B1(_1963_),
    .Y(_1965_),
    .A1(_0036_),
    .A2(net1813));
 sg13g2_mux2_1 _6156_ (.A0(_0038_),
    .A1(_0037_),
    .S(net1813),
    .X(_1966_));
 sg13g2_a21oi_1 _6157_ (.A1(net1800),
    .A2(_1966_),
    .Y(_1967_),
    .B1(_1960_));
 sg13g2_o21ai_1 _6158_ (.B1(_1967_),
    .Y(_1968_),
    .A1(_1958_),
    .A2(_1965_));
 sg13g2_o21ai_1 _6159_ (.B1(_1968_),
    .Y(_1969_),
    .A1(net1805),
    .A2(_1964_));
 sg13g2_o21ai_1 _6160_ (.B1(_1955_),
    .Y(_1970_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[8] ),
    .A2(net1827));
 sg13g2_nor2_1 _6161_ (.A(net1833),
    .B(_1969_),
    .Y(_1971_));
 sg13g2_a21oi_2 _6162_ (.B1(_1971_),
    .Y(_1972_),
    .A2(_1970_),
    .A1(net1833));
 sg13g2_mux2_1 _6163_ (.A0(net353),
    .A1(_1972_),
    .S(_1770_),
    .X(_0309_));
 sg13g2_nand2_1 _6164_ (.Y(_1973_),
    .A(\z80.tv80s.i_tv80_core.BusB[1] ),
    .B(net1787));
 sg13g2_nor2_1 _6165_ (.A(_1782_),
    .B(_1786_),
    .Y(_1974_));
 sg13g2_xor2_1 _6166_ (.B(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A(net2037),
    .X(_1975_));
 sg13g2_xnor2_1 _6167_ (.Y(_1976_),
    .A(_0209_),
    .B(_1975_));
 sg13g2_o21ai_1 _6168_ (.B1(_1976_),
    .Y(_1977_),
    .A1(_1782_),
    .A2(_1786_));
 sg13g2_xnor2_1 _6169_ (.Y(_1978_),
    .A(_1974_),
    .B(_1976_));
 sg13g2_nor2_1 _6170_ (.A(net2027),
    .B(\z80.tv80s.i_tv80_core.BusB[1] ),
    .Y(_1979_));
 sg13g2_nand2_1 _6171_ (.Y(_1980_),
    .A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(\z80.tv80s.i_tv80_core.BusB[1] ));
 sg13g2_a22oi_1 _6172_ (.Y(_1981_),
    .B1(_1795_),
    .B2(_1980_),
    .A2(net1873),
    .A1(net2039));
 sg13g2_or2_1 _6173_ (.X(_1982_),
    .B(_1980_),
    .A(_1800_));
 sg13g2_o21ai_1 _6174_ (.B1(_1982_),
    .Y(_1983_),
    .A1(_1979_),
    .A2(_1981_));
 sg13g2_a21oi_2 _6175_ (.B1(_1983_),
    .Y(_1984_),
    .A2(_1978_),
    .A1(_1789_));
 sg13g2_nand2_1 _6176_ (.Y(_1985_),
    .A(net1874),
    .B(_1984_));
 sg13g2_nor2_1 _6177_ (.A(net2027),
    .B(\z80.tv80s.i_tv80_core.BusA[2] ),
    .Y(_1986_));
 sg13g2_o21ai_1 _6178_ (.B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .Y(_1987_),
    .A1(net2027),
    .A2(net2028));
 sg13g2_nand2b_2 _6179_ (.Y(_1988_),
    .B(_1987_),
    .A_N(\z80.tv80s.i_tv80_core.F[4] ));
 sg13g2_xor2_1 _6180_ (.B(_1988_),
    .A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(_1989_));
 sg13g2_nand2_1 _6181_ (.Y(_1990_),
    .A(net2060),
    .B(_1037_));
 sg13g2_nand2_1 _6182_ (.Y(_1991_),
    .A(_1823_),
    .B(_1990_));
 sg13g2_a22oi_1 _6183_ (.Y(_1992_),
    .B1(_1991_),
    .B2(_1822_),
    .A2(_1990_),
    .A1(_0218_));
 sg13g2_nor2_1 _6184_ (.A(_0218_),
    .B(_1990_),
    .Y(_1993_));
 sg13g2_mux2_2 _6185_ (.A0(_0218_),
    .A1(_0222_),
    .S(net2042),
    .X(_1994_));
 sg13g2_mux2_1 _6186_ (.A0(_0212_),
    .A1(_0211_),
    .S(net2076),
    .X(_1995_));
 sg13g2_or2_1 _6187_ (.X(_1996_),
    .B(_1995_),
    .A(net1863));
 sg13g2_o21ai_1 _6188_ (.B1(_1996_),
    .Y(_1997_),
    .A1(_1809_),
    .A2(_1994_));
 sg13g2_a21oi_1 _6189_ (.A1(_1812_),
    .A2(_1993_),
    .Y(_1998_),
    .B1(net1874));
 sg13g2_a21oi_1 _6190_ (.A1(_1816_),
    .A2(_1989_),
    .Y(_1999_),
    .B1(_1997_));
 sg13g2_nand2_1 _6191_ (.Y(_2000_),
    .A(_1998_),
    .B(_1999_));
 sg13g2_o21ai_1 _6192_ (.B1(_1985_),
    .Y(_2001_),
    .A1(_1992_),
    .A2(_2000_));
 sg13g2_inv_1 _6193_ (.Y(_2002_),
    .A(_2001_));
 sg13g2_nand2_1 _6194_ (.Y(_2003_),
    .A(net2032),
    .B(_2001_));
 sg13g2_o21ai_1 _6195_ (.B1(_2003_),
    .Y(_2004_),
    .A1(net2032),
    .A2(net2050));
 sg13g2_o21ai_1 _6196_ (.B1(_1973_),
    .Y(_2005_),
    .A1(net1787),
    .A2(_2004_));
 sg13g2_a21oi_2 _6197_ (.B1(_1719_),
    .Y(_2006_),
    .A2(_2005_),
    .A1(net1789));
 sg13g2_a22oi_1 _6198_ (.Y(_2007_),
    .B1(net1738),
    .B2(_0047_),
    .A2(net1748),
    .A1(_0051_));
 sg13g2_a22oi_1 _6199_ (.Y(_2008_),
    .B1(net1734),
    .B2(_0049_),
    .A2(net1746),
    .A1(_0052_));
 sg13g2_and2_1 _6200_ (.A(_2007_),
    .B(_2008_),
    .X(_2009_));
 sg13g2_a22oi_1 _6201_ (.Y(_2010_),
    .B1(net1740),
    .B2(_0050_),
    .A2(net1744),
    .A1(_0046_));
 sg13g2_a22oi_1 _6202_ (.Y(_2011_),
    .B1(_1861_),
    .B2(_0045_),
    .A2(_1855_),
    .A1(_0048_));
 sg13g2_nand3_1 _6203_ (.B(_2010_),
    .C(_2011_),
    .A(_2009_),
    .Y(_2012_));
 sg13g2_xnor2_1 _6204_ (.Y(_2013_),
    .A(net1816),
    .B(_2012_));
 sg13g2_o21ai_1 _6205_ (.B1(_1953_),
    .Y(_2014_),
    .A1(net1816),
    .A2(_1950_));
 sg13g2_xnor2_1 _6206_ (.Y(_2015_),
    .A(_2013_),
    .B(_2014_));
 sg13g2_nand2_1 _6207_ (.Y(_2016_),
    .A(net1791),
    .B(_2015_));
 sg13g2_a22oi_1 _6208_ (.Y(_2017_),
    .B1(_2006_),
    .B2(_2016_),
    .A2(_1719_),
    .A1(_0803_));
 sg13g2_mux4_1 _6209_ (.S0(net1810),
    .A0(_0049_),
    .A1(_0050_),
    .A2(_0045_),
    .A3(_0046_),
    .S1(net1805),
    .X(_2018_));
 sg13g2_nor2_1 _6210_ (.A(net1799),
    .B(_2018_),
    .Y(_2019_));
 sg13g2_mux2_2 _6211_ (.A0(_2019_),
    .A1(_2017_),
    .S(net1834),
    .X(_2020_));
 sg13g2_mux2_1 _6212_ (.A0(net271),
    .A1(_2020_),
    .S(_1770_),
    .X(_0310_));
 sg13g2_nand3_1 _6213_ (.B(\z80.tv80s.i_tv80_core.BusB[2] ),
    .C(_1799_),
    .A(net2028),
    .Y(_2021_));
 sg13g2_nor3_1 _6214_ (.A(_0780_),
    .B(net2028),
    .C(\z80.tv80s.i_tv80_core.BusB[2] ),
    .Y(_2022_));
 sg13g2_nand2_1 _6215_ (.Y(_2023_),
    .A(net2027),
    .B(_1975_));
 sg13g2_xnor2_1 _6216_ (.Y(_2024_),
    .A(net2037),
    .B(\z80.tv80s.i_tv80_core.BusB[2] ));
 sg13g2_xnor2_1 _6217_ (.Y(_2025_),
    .A(net2028),
    .B(_2024_));
 sg13g2_inv_1 _6218_ (.Y(_2026_),
    .A(_2025_));
 sg13g2_a21oi_1 _6219_ (.A1(_1977_),
    .A2(_2023_),
    .Y(_2027_),
    .B1(_2026_));
 sg13g2_nand3_1 _6220_ (.B(_2023_),
    .C(_2026_),
    .A(_1977_),
    .Y(_2028_));
 sg13g2_nor2b_1 _6221_ (.A(_2027_),
    .B_N(_2028_),
    .Y(_2029_));
 sg13g2_a22oi_1 _6222_ (.Y(_2030_),
    .B1(_1795_),
    .B2(_2025_),
    .A2(net1873),
    .A1(net2037));
 sg13g2_a22oi_1 _6223_ (.Y(_2031_),
    .B1(_2030_),
    .B2(_2021_),
    .A2(_2022_),
    .A1(net1873));
 sg13g2_a21oi_2 _6224_ (.B1(_2031_),
    .Y(_2032_),
    .A2(_2029_),
    .A1(_1789_));
 sg13g2_nand2_2 _6225_ (.Y(_2033_),
    .A(net2027),
    .B(net2028));
 sg13g2_nor2b_1 _6226_ (.A(_1986_),
    .B_N(_2033_),
    .Y(_2034_));
 sg13g2_xnor2_1 _6227_ (.Y(_2035_),
    .A(net2149),
    .B(_2034_));
 sg13g2_nor2_1 _6228_ (.A(_0211_),
    .B(_1988_),
    .Y(_2036_));
 sg13g2_a21oi_2 _6229_ (.B1(_2036_),
    .Y(_2037_),
    .A2(_2035_),
    .A1(_1988_));
 sg13g2_nand2_1 _6230_ (.Y(_2038_),
    .A(_1035_),
    .B(_1823_));
 sg13g2_a22oi_1 _6231_ (.Y(_2039_),
    .B1(_1822_),
    .B2(_2038_),
    .A2(_1035_),
    .A1(_0219_));
 sg13g2_mux2_1 _6232_ (.A0(_0219_),
    .A1(_0223_),
    .S(net2041),
    .X(_2040_));
 sg13g2_nor2_1 _6233_ (.A(_1809_),
    .B(_2040_),
    .Y(_2041_));
 sg13g2_nor3_1 _6234_ (.A(_0219_),
    .B(_1035_),
    .C(_1813_),
    .Y(_2042_));
 sg13g2_mux2_1 _6235_ (.A0(_0209_),
    .A1(_0213_),
    .S(net2076),
    .X(_2043_));
 sg13g2_o21ai_1 _6236_ (.B1(_1780_),
    .Y(_2044_),
    .A1(net1863),
    .A2(_2043_));
 sg13g2_nor4_1 _6237_ (.A(_2039_),
    .B(_2041_),
    .C(_2042_),
    .D(_2044_),
    .Y(_2045_));
 sg13g2_o21ai_1 _6238_ (.B1(_2045_),
    .Y(_2046_),
    .A1(_1817_),
    .A2(_2037_));
 sg13g2_a21oi_1 _6239_ (.A1(_1779_),
    .A2(_2032_),
    .Y(_2047_),
    .B1(_0690_));
 sg13g2_nand2_1 _6240_ (.Y(_2048_),
    .A(_2046_),
    .B(_2047_));
 sg13g2_a21oi_1 _6241_ (.A1(_0690_),
    .A2(net2049),
    .Y(_2049_),
    .B1(net1787));
 sg13g2_a22oi_1 _6242_ (.Y(_2050_),
    .B1(_2048_),
    .B2(_2049_),
    .A2(net1788),
    .A1(_0784_));
 sg13g2_a21o_1 _6243_ (.A2(_2050_),
    .A1(net1789),
    .B1(_1719_),
    .X(_2051_));
 sg13g2_a22oi_1 _6244_ (.Y(_2052_),
    .B1(net1738),
    .B2(_0055_),
    .A2(net1744),
    .A1(_0054_));
 sg13g2_a22oi_1 _6245_ (.Y(_2053_),
    .B1(net1736),
    .B2(_0053_),
    .A2(net1740),
    .A1(_0058_));
 sg13g2_a22oi_1 _6246_ (.Y(_2054_),
    .B1(net1742),
    .B2(_0056_),
    .A2(net1746),
    .A1(_0060_));
 sg13g2_a22oi_1 _6247_ (.Y(_2055_),
    .B1(net1734),
    .B2(_0057_),
    .A2(net1748),
    .A1(_0059_));
 sg13g2_nand4_1 _6248_ (.B(_2053_),
    .C(_2054_),
    .A(_2052_),
    .Y(_2056_),
    .D(_2055_));
 sg13g2_nand2b_1 _6249_ (.Y(_2057_),
    .B(net1823),
    .A_N(_2056_));
 sg13g2_inv_1 _6250_ (.Y(_2058_),
    .A(_2057_));
 sg13g2_nand2_1 _6251_ (.Y(_2059_),
    .A(net1815),
    .B(_2056_));
 sg13g2_nand2_1 _6252_ (.Y(_2060_),
    .A(_2057_),
    .B(_2059_));
 sg13g2_a21o_1 _6253_ (.A2(_2012_),
    .A1(_1950_),
    .B1(net1815),
    .X(_2061_));
 sg13g2_a22oi_1 _6254_ (.Y(_2062_),
    .B1(_2061_),
    .B2(_1953_),
    .A2(_2012_),
    .A1(net1815));
 sg13g2_xnor2_1 _6255_ (.Y(_2063_),
    .A(_2060_),
    .B(_2062_));
 sg13g2_a21oi_2 _6256_ (.B1(_2051_),
    .Y(_2064_),
    .A2(_2063_),
    .A1(net1791));
 sg13g2_o21ai_1 _6257_ (.B1(net1833),
    .Y(_2065_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[10] ),
    .A2(net1827));
 sg13g2_mux4_1 _6258_ (.S0(net1810),
    .A0(_0057_),
    .A1(_0058_),
    .A2(_0053_),
    .A3(_0054_),
    .S1(net1805),
    .X(_2066_));
 sg13g2_nor2_1 _6259_ (.A(net1799),
    .B(_2066_),
    .Y(_2067_));
 sg13g2_or2_1 _6260_ (.X(_2068_),
    .B(_2066_),
    .A(net1832));
 sg13g2_o21ai_1 _6261_ (.B1(_2068_),
    .Y(_2069_),
    .A1(_2064_),
    .A2(_2065_));
 sg13g2_mux2_1 _6262_ (.A0(net322),
    .A1(_2069_),
    .S(_1770_),
    .X(_0311_));
 sg13g2_xor2_1 _6263_ (.B(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A(net2037),
    .X(_2070_));
 sg13g2_inv_1 _6264_ (.Y(_2071_),
    .A(_2070_));
 sg13g2_xnor2_1 _6265_ (.Y(_2072_),
    .A(_0783_),
    .B(_2070_));
 sg13g2_nor2_1 _6266_ (.A(_0211_),
    .B(_2024_),
    .Y(_2073_));
 sg13g2_o21ai_1 _6267_ (.B1(_2072_),
    .Y(_2074_),
    .A1(_2027_),
    .A2(_2073_));
 sg13g2_nor3_1 _6268_ (.A(_2027_),
    .B(_2072_),
    .C(_2073_),
    .Y(_2075_));
 sg13g2_nor2_1 _6269_ (.A(net1873),
    .B(_2075_),
    .Y(_2076_));
 sg13g2_and2_1 _6270_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(_2077_));
 sg13g2_nor3_1 _6271_ (.A(_0780_),
    .B(\z80.tv80s.i_tv80_core.BusA[3] ),
    .C(\z80.tv80s.i_tv80_core.BusB[3] ),
    .Y(_2078_));
 sg13g2_a22oi_1 _6272_ (.Y(_2079_),
    .B1(_2077_),
    .B2(_1799_),
    .A2(_2072_),
    .A1(_1795_));
 sg13g2_a21oi_1 _6273_ (.A1(_1793_),
    .A2(_2079_),
    .Y(_2080_),
    .B1(_2078_));
 sg13g2_a21oi_2 _6274_ (.B1(_2080_),
    .Y(_2081_),
    .A2(_2076_),
    .A1(_2074_));
 sg13g2_nor2_1 _6275_ (.A(_1780_),
    .B(_2081_),
    .Y(_2082_));
 sg13g2_nor2_1 _6276_ (.A(net2148),
    .B(_1986_),
    .Y(_2083_));
 sg13g2_a21oi_1 _6277_ (.A1(net2148),
    .A2(_2033_),
    .Y(_2084_),
    .B1(_2083_));
 sg13g2_xnor2_1 _6278_ (.Y(_2085_),
    .A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B(_2084_));
 sg13g2_nor2_1 _6279_ (.A(_0213_),
    .B(_1988_),
    .Y(_2086_));
 sg13g2_a21oi_2 _6280_ (.B1(_2086_),
    .Y(_2087_),
    .A2(_2085_),
    .A1(_1988_));
 sg13g2_mux2_1 _6281_ (.A0(_0211_),
    .A1(_0214_),
    .S(net2076),
    .X(_2088_));
 sg13g2_nor2_1 _6282_ (.A(net1863),
    .B(_2088_),
    .Y(_2089_));
 sg13g2_mux2_1 _6283_ (.A0(_0220_),
    .A1(_0224_),
    .S(net2041),
    .X(_2090_));
 sg13g2_inv_1 _6284_ (.Y(_2091_),
    .A(_2090_));
 sg13g2_a21oi_1 _6285_ (.A1(_1808_),
    .A2(_2091_),
    .Y(_2092_),
    .B1(_2089_));
 sg13g2_o21ai_1 _6286_ (.B1(_2092_),
    .Y(_2093_),
    .A1(_1817_),
    .A2(_2087_));
 sg13g2_nor2_1 _6287_ (.A(_0220_),
    .B(_1042_),
    .Y(_2094_));
 sg13g2_a221oi_1 _6288_ (.B2(_1812_),
    .C1(_1821_),
    .B1(_2094_),
    .A1(_1042_),
    .Y(_2095_),
    .A2(_1823_));
 sg13g2_a21oi_1 _6289_ (.A1(_0220_),
    .A2(_1042_),
    .Y(_2096_),
    .B1(_2095_));
 sg13g2_nor3_2 _6290_ (.A(_2082_),
    .B(_2093_),
    .C(_2096_),
    .Y(_2097_));
 sg13g2_nand2_1 _6291_ (.Y(_2098_),
    .A(net2032),
    .B(_2097_));
 sg13g2_a21oi_1 _6292_ (.A1(_0690_),
    .A2(_0705_),
    .Y(_2099_),
    .B1(net1787));
 sg13g2_a22oi_1 _6293_ (.Y(_2100_),
    .B1(_2098_),
    .B2(_2099_),
    .A2(net1787),
    .A1(\z80.tv80s.i_tv80_core.BusB[3] ));
 sg13g2_inv_1 _6294_ (.Y(_2101_),
    .A(_2100_));
 sg13g2_o21ai_1 _6295_ (.B1(net1825),
    .Y(_2102_),
    .A1(net1790),
    .A2(_2100_));
 sg13g2_a22oi_1 _6296_ (.Y(_2103_),
    .B1(net1742),
    .B2(_0072_),
    .A2(net1744),
    .A1(_0070_));
 sg13g2_a22oi_1 _6297_ (.Y(_2104_),
    .B1(net1746),
    .B2(_0076_),
    .A2(net1748),
    .A1(_0075_));
 sg13g2_a22oi_1 _6298_ (.Y(_2105_),
    .B1(net1736),
    .B2(_0069_),
    .A2(net1740),
    .A1(_0074_));
 sg13g2_a22oi_1 _6299_ (.Y(_2106_),
    .B1(net1734),
    .B2(_0073_),
    .A2(net1738),
    .A1(_0071_));
 sg13g2_nand4_1 _6300_ (.B(_2104_),
    .C(_2105_),
    .A(_2103_),
    .Y(_2107_),
    .D(_2106_));
 sg13g2_xnor2_1 _6301_ (.Y(_2108_),
    .A(net1816),
    .B(_2107_));
 sg13g2_a21oi_1 _6302_ (.A1(_2059_),
    .A2(_2062_),
    .Y(_2109_),
    .B1(_2058_));
 sg13g2_xor2_1 _6303_ (.B(_2109_),
    .A(_2108_),
    .X(_2110_));
 sg13g2_a21oi_1 _6304_ (.A1(net1791),
    .A2(_2110_),
    .Y(_2111_),
    .B1(_2102_));
 sg13g2_o21ai_1 _6305_ (.B1(net1832),
    .Y(_2112_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[11] ),
    .A2(net1827));
 sg13g2_or2_1 _6306_ (.X(_2113_),
    .B(_2112_),
    .A(_2111_));
 sg13g2_mux4_1 _6307_ (.S0(net1813),
    .A0(_0074_),
    .A1(_0073_),
    .A2(_0076_),
    .A3(_0075_),
    .S1(net1799),
    .X(_2114_));
 sg13g2_nor2_1 _6308_ (.A(net1805),
    .B(_2114_),
    .Y(_2115_));
 sg13g2_a21oi_1 _6309_ (.A1(_0706_),
    .A2(net1809),
    .Y(_2116_),
    .B1(net1800));
 sg13g2_o21ai_1 _6310_ (.B1(_2116_),
    .Y(_2117_),
    .A1(_0069_),
    .A2(net1809));
 sg13g2_mux2_1 _6311_ (.A0(_0072_),
    .A1(_0071_),
    .S(net1813),
    .X(_2118_));
 sg13g2_a21oi_1 _6312_ (.A1(net1799),
    .A2(_2118_),
    .Y(_2119_),
    .B1(net1786));
 sg13g2_a21oi_2 _6313_ (.B1(_2115_),
    .Y(_2120_),
    .A2(_2119_),
    .A1(_2117_));
 sg13g2_o21ai_1 _6314_ (.B1(_2113_),
    .Y(_2121_),
    .A1(net1833),
    .A2(_2120_));
 sg13g2_mux2_1 _6315_ (.A0(net274),
    .A1(_2121_),
    .S(_1770_),
    .X(_0312_));
 sg13g2_o21ai_1 _6316_ (.B1(_2074_),
    .Y(_2122_),
    .A1(_0213_),
    .A2(_2071_));
 sg13g2_xor2_1 _6317_ (.B(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A(net2039),
    .X(_2123_));
 sg13g2_nand2b_1 _6318_ (.Y(_2124_),
    .B(_2123_),
    .A_N(_0214_));
 sg13g2_xnor2_1 _6319_ (.Y(_2125_),
    .A(_0214_),
    .B(_2123_));
 sg13g2_nand2_1 _6320_ (.Y(_2126_),
    .A(_2122_),
    .B(_2125_));
 sg13g2_o21ai_1 _6321_ (.B1(_1789_),
    .Y(_2127_),
    .A1(_2122_),
    .A2(_2125_));
 sg13g2_nor2b_1 _6322_ (.A(_2127_),
    .B_N(_2126_),
    .Y(_2128_));
 sg13g2_and2_1 _6323_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(\z80.tv80s.i_tv80_core.BusB[4] ),
    .X(_2129_));
 sg13g2_xor2_1 _6324_ (.B(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .X(_2130_));
 sg13g2_a221oi_1 _6325_ (.B2(_1796_),
    .C1(_2128_),
    .B1(_2130_),
    .A1(_1801_),
    .Y(_2131_),
    .A2(_2129_));
 sg13g2_nand2_1 _6326_ (.Y(_2132_),
    .A(_1779_),
    .B(_2131_));
 sg13g2_nand4_1 _6327_ (.B(_0213_),
    .C(_1988_),
    .A(net2148),
    .Y(_2133_),
    .D(_2033_));
 sg13g2_o21ai_1 _6328_ (.B1(_2133_),
    .Y(_2134_),
    .A1(net2148),
    .A2(_1987_));
 sg13g2_xor2_1 _6329_ (.B(_2134_),
    .A(_0214_),
    .X(_2135_));
 sg13g2_nand2_1 _6330_ (.Y(_2136_),
    .A(_1054_),
    .B(_1823_));
 sg13g2_a22oi_1 _6331_ (.Y(_2137_),
    .B1(_1822_),
    .B2(_2136_),
    .A2(_1054_),
    .A1(_0221_));
 sg13g2_nand2_1 _6332_ (.Y(_2138_),
    .A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_1808_));
 sg13g2_or2_1 _6333_ (.X(_2139_),
    .B(_1054_),
    .A(_0221_));
 sg13g2_nor2_1 _6334_ (.A(_1813_),
    .B(_2139_),
    .Y(_2140_));
 sg13g2_mux2_1 _6335_ (.A0(_0213_),
    .A1(_0215_),
    .S(net2076),
    .X(_2141_));
 sg13g2_o21ai_1 _6336_ (.B1(_2138_),
    .Y(_2142_),
    .A1(net1863),
    .A2(_2141_));
 sg13g2_nor4_1 _6337_ (.A(net1874),
    .B(_2137_),
    .C(_2140_),
    .D(_2142_),
    .Y(_2143_));
 sg13g2_o21ai_1 _6338_ (.B1(_2143_),
    .Y(_2144_),
    .A1(_1817_),
    .A2(_2135_));
 sg13g2_nand3_1 _6339_ (.B(_2132_),
    .C(_2144_),
    .A(net2032),
    .Y(_2145_));
 sg13g2_a21oi_1 _6340_ (.A1(_0690_),
    .A2(\z80.tv80s.di_reg[4] ),
    .Y(_2146_),
    .B1(net1788));
 sg13g2_a22oi_1 _6341_ (.Y(_2147_),
    .B1(_2145_),
    .B2(_2146_),
    .A2(net1788),
    .A1(_0785_));
 sg13g2_a21o_1 _6342_ (.A2(_2147_),
    .A1(net1789),
    .B1(_1719_),
    .X(_2148_));
 sg13g2_nor4_1 _6343_ (.A(_1951_),
    .B(_2013_),
    .C(_2060_),
    .D(_2108_),
    .Y(_2149_));
 sg13g2_o21ai_1 _6344_ (.B1(_2149_),
    .Y(_2150_),
    .A1(_1939_),
    .A2(_1943_));
 sg13g2_or3_1 _6345_ (.A(_2060_),
    .B(_2061_),
    .C(_2108_),
    .X(_2151_));
 sg13g2_a21oi_1 _6346_ (.A1(_2056_),
    .A2(_2107_),
    .Y(_2152_),
    .B1(net1815));
 sg13g2_nor2b_1 _6347_ (.A(_2152_),
    .B_N(_2151_),
    .Y(_2153_));
 sg13g2_a22oi_1 _6348_ (.Y(_2154_),
    .B1(net1740),
    .B2(_0090_),
    .A2(net1746),
    .A1(_0092_));
 sg13g2_a22oi_1 _6349_ (.Y(_2155_),
    .B1(net1734),
    .B2(_0089_),
    .A2(net1744),
    .A1(_0086_));
 sg13g2_a22oi_1 _6350_ (.Y(_2156_),
    .B1(net1738),
    .B2(_0087_),
    .A2(net1748),
    .A1(_0091_));
 sg13g2_a22oi_1 _6351_ (.Y(_2157_),
    .B1(net1736),
    .B2(_0085_),
    .A2(net1742),
    .A1(_0088_));
 sg13g2_and2_1 _6352_ (.A(_2154_),
    .B(_2157_),
    .X(_2158_));
 sg13g2_nand3_1 _6353_ (.B(_2156_),
    .C(_2158_),
    .A(_2155_),
    .Y(_2159_));
 sg13g2_inv_1 _6354_ (.Y(_2160_),
    .A(_2159_));
 sg13g2_xnor2_1 _6355_ (.Y(_2161_),
    .A(net1816),
    .B(_2159_));
 sg13g2_a21oi_1 _6356_ (.A1(_2150_),
    .A2(_2153_),
    .Y(_2162_),
    .B1(_2161_));
 sg13g2_nand3_1 _6357_ (.B(_2153_),
    .C(_2161_),
    .A(_2150_),
    .Y(_2163_));
 sg13g2_nor2b_1 _6358_ (.A(_2162_),
    .B_N(_2163_),
    .Y(_2164_));
 sg13g2_a21oi_2 _6359_ (.B1(_2148_),
    .Y(_2165_),
    .A2(_2164_),
    .A1(net1791));
 sg13g2_o21ai_1 _6360_ (.B1(net1831),
    .Y(_2166_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[12] ),
    .A2(net1827));
 sg13g2_a21oi_1 _6361_ (.A1(_0711_),
    .A2(net1809),
    .Y(_2167_),
    .B1(net1804));
 sg13g2_o21ai_1 _6362_ (.B1(_2167_),
    .Y(_2168_),
    .A1(_0091_),
    .A2(net2163));
 sg13g2_nor2_1 _6363_ (.A(_0087_),
    .B(net2163),
    .Y(_2169_));
 sg13g2_o21ai_1 _6364_ (.B1(net1804),
    .Y(_2170_),
    .A1(_0088_),
    .A2(net1813));
 sg13g2_o21ai_1 _6365_ (.B1(_2168_),
    .Y(_2171_),
    .A1(_2169_),
    .A2(_2170_));
 sg13g2_mux4_1 _6366_ (.S0(net1810),
    .A0(_0089_),
    .A1(_0090_),
    .A2(_0085_),
    .A3(_0086_),
    .S1(net1804),
    .X(_2172_));
 sg13g2_mux2_1 _6367_ (.A0(_2171_),
    .A1(_2172_),
    .S(_1963_),
    .X(_2173_));
 sg13g2_or2_1 _6368_ (.X(_2174_),
    .B(_2172_),
    .A(net1831));
 sg13g2_o21ai_1 _6369_ (.B1(_2174_),
    .Y(_2175_),
    .A1(_2165_),
    .A2(_2166_));
 sg13g2_mux2_1 _6370_ (.A0(net279),
    .A1(_2175_),
    .S(_1770_),
    .X(_0313_));
 sg13g2_xor2_1 _6371_ (.B(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A(net2037),
    .X(_2176_));
 sg13g2_nor2b_1 _6372_ (.A(_0215_),
    .B_N(_2176_),
    .Y(_2177_));
 sg13g2_xor2_1 _6373_ (.B(_2176_),
    .A(_0215_),
    .X(_2178_));
 sg13g2_nand3_1 _6374_ (.B(_2126_),
    .C(_2178_),
    .A(_2124_),
    .Y(_2179_));
 sg13g2_a21oi_1 _6375_ (.A1(_2124_),
    .A2(_2126_),
    .Y(_2180_),
    .B1(_2178_));
 sg13g2_nor2_1 _6376_ (.A(net1873),
    .B(_2180_),
    .Y(_2181_));
 sg13g2_and3_1 _6377_ (.X(_2182_),
    .A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(\z80.tv80s.i_tv80_core.BusB[5] ),
    .C(_1801_));
 sg13g2_xor2_1 _6378_ (.B(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A(net2029),
    .X(_2183_));
 sg13g2_a221oi_1 _6379_ (.B2(_1796_),
    .C1(_2182_),
    .B1(_2183_),
    .A1(_2179_),
    .Y(_2184_),
    .A2(_2181_));
 sg13g2_inv_1 _6380_ (.Y(_2185_),
    .A(_2184_));
 sg13g2_nand2_1 _6381_ (.Y(_2186_),
    .A(_1779_),
    .B(_2184_));
 sg13g2_nand3b_1 _6382_ (.B(\z80.tv80s.i_tv80_core.BusA[4] ),
    .C(\z80.tv80s.i_tv80_core.BusA[3] ),
    .Y(_2187_),
    .A_N(_1986_));
 sg13g2_nor2_1 _6383_ (.A(net2029),
    .B(net2030),
    .Y(_2188_));
 sg13g2_nand2_1 _6384_ (.Y(_2189_),
    .A(_2187_),
    .B(_2188_));
 sg13g2_a21oi_2 _6385_ (.B1(net2151),
    .Y(_2190_),
    .A2(_2189_),
    .A1(\z80.tv80s.i_tv80_core.BusA[7] ));
 sg13g2_nand2_1 _6386_ (.Y(_2191_),
    .A(\z80.tv80s.i_tv80_core.F[4] ),
    .B(_2033_));
 sg13g2_nor3_1 _6387_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B(\z80.tv80s.i_tv80_core.BusA[4] ),
    .C(_2191_),
    .Y(_2192_));
 sg13g2_xnor2_1 _6388_ (.Y(_2193_),
    .A(_0215_),
    .B(_2192_));
 sg13g2_nor2b_1 _6389_ (.A(_2190_),
    .B_N(_2193_),
    .Y(_2194_));
 sg13g2_xor2_1 _6390_ (.B(_2193_),
    .A(_2190_),
    .X(_2195_));
 sg13g2_nor2_1 _6391_ (.A(_0215_),
    .B(_2187_),
    .Y(_2196_));
 sg13g2_xor2_1 _6392_ (.B(_2187_),
    .A(_0215_),
    .X(_2197_));
 sg13g2_nand2_1 _6393_ (.Y(_2198_),
    .A(net2029),
    .B(net2030));
 sg13g2_nor2_1 _6394_ (.A(_2187_),
    .B(_2198_),
    .Y(_2199_));
 sg13g2_nand2_1 _6395_ (.Y(_2200_),
    .A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .B(_2199_));
 sg13g2_xnor2_1 _6396_ (.Y(_2201_),
    .A(_0216_),
    .B(_2196_));
 sg13g2_nor2_1 _6397_ (.A(_2197_),
    .B(_2201_),
    .Y(_2202_));
 sg13g2_xnor2_1 _6398_ (.Y(_2203_),
    .A(_0781_),
    .B(_2199_));
 sg13g2_or2_1 _6399_ (.X(_2204_),
    .B(_2203_),
    .A(_2202_));
 sg13g2_and3_1 _6400_ (.X(_2205_),
    .A(_0665_),
    .B(_2200_),
    .C(_2204_));
 sg13g2_nor2_1 _6401_ (.A(_2197_),
    .B(_2205_),
    .Y(_2206_));
 sg13g2_a21oi_1 _6402_ (.A1(_2197_),
    .A2(_2205_),
    .Y(_2207_),
    .B1(net2149));
 sg13g2_nor2b_1 _6403_ (.A(_2206_),
    .B_N(_2207_),
    .Y(_2208_));
 sg13g2_a21oi_2 _6404_ (.B1(_2208_),
    .Y(_2209_),
    .A2(_2195_),
    .A1(net2148));
 sg13g2_a22oi_1 _6405_ (.Y(_2210_),
    .B1(_1816_),
    .B2(_2209_),
    .A2(_1808_),
    .A1(net2029));
 sg13g2_nand2_1 _6406_ (.Y(_2211_),
    .A(_1044_),
    .B(_1823_));
 sg13g2_a22oi_1 _6407_ (.Y(_2212_),
    .B1(_1822_),
    .B2(_2211_),
    .A2(_1044_),
    .A1(_0222_));
 sg13g2_nor3_1 _6408_ (.A(_0222_),
    .B(_1044_),
    .C(_1813_),
    .Y(_2213_));
 sg13g2_mux2_1 _6409_ (.A0(_0214_),
    .A1(_0216_),
    .S(net2076),
    .X(_2214_));
 sg13g2_nor2_1 _6410_ (.A(_1804_),
    .B(_2214_),
    .Y(_2215_));
 sg13g2_nor4_1 _6411_ (.A(net1874),
    .B(_2212_),
    .C(_2213_),
    .D(_2215_),
    .Y(_2216_));
 sg13g2_a21oi_1 _6412_ (.A1(_2210_),
    .A2(_2216_),
    .Y(_2217_),
    .B1(_0690_));
 sg13g2_a22oi_1 _6413_ (.Y(_2218_),
    .B1(_2186_),
    .B2(_2217_),
    .A2(net2046),
    .A1(_0690_));
 sg13g2_mux2_2 _6414_ (.A0(_2218_),
    .A1(_0786_),
    .S(net1788),
    .X(_2219_));
 sg13g2_inv_1 _6415_ (.Y(_2220_),
    .A(_2219_));
 sg13g2_o21ai_1 _6416_ (.B1(net1826),
    .Y(_2221_),
    .A1(net1790),
    .A2(_2219_));
 sg13g2_a22oi_1 _6417_ (.Y(_2222_),
    .B1(net1738),
    .B2(_0103_),
    .A2(net1748),
    .A1(_0107_));
 sg13g2_a22oi_1 _6418_ (.Y(_2223_),
    .B1(net1740),
    .B2(_0106_),
    .A2(net1744),
    .A1(_0102_));
 sg13g2_a22oi_1 _6419_ (.Y(_2224_),
    .B1(net1736),
    .B2(_0101_),
    .A2(net1742),
    .A1(_0104_));
 sg13g2_a22oi_1 _6420_ (.Y(_2225_),
    .B1(net1734),
    .B2(_0105_),
    .A2(net1746),
    .A1(_0108_));
 sg13g2_and2_1 _6421_ (.A(_2222_),
    .B(_2225_),
    .X(_2226_));
 sg13g2_nand3_1 _6422_ (.B(_2224_),
    .C(_2226_),
    .A(_2223_),
    .Y(_2227_));
 sg13g2_nor2_1 _6423_ (.A(net1815),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_xnor2_1 _6424_ (.Y(_2229_),
    .A(net1815),
    .B(_2227_));
 sg13g2_inv_1 _6425_ (.Y(_2230_),
    .A(_2229_));
 sg13g2_a21o_1 _6426_ (.A2(_2160_),
    .A1(net1823),
    .B1(_2162_),
    .X(_2231_));
 sg13g2_xnor2_1 _6427_ (.Y(_2232_),
    .A(_2229_),
    .B(_2231_));
 sg13g2_a21oi_1 _6428_ (.A1(net1791),
    .A2(_2232_),
    .Y(_2233_),
    .B1(_2221_));
 sg13g2_o21ai_1 _6429_ (.B1(net1832),
    .Y(_2234_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[13] ),
    .A2(net1827));
 sg13g2_mux4_1 _6430_ (.S0(net1810),
    .A0(_0105_),
    .A1(_0106_),
    .A2(_0101_),
    .A3(_0102_),
    .S1(net1804),
    .X(_2235_));
 sg13g2_nor2_1 _6431_ (.A(net1799),
    .B(_2235_),
    .Y(_2236_));
 sg13g2_or2_1 _6432_ (.X(_2237_),
    .B(_2235_),
    .A(net1832));
 sg13g2_o21ai_1 _6433_ (.B1(_2237_),
    .Y(_2238_),
    .A1(_2233_),
    .A2(_2234_));
 sg13g2_mux2_1 _6434_ (.A0(net280),
    .A1(_2238_),
    .S(_1770_),
    .X(_0314_));
 sg13g2_mux4_1 _6435_ (.S0(net1809),
    .A0(_0121_),
    .A1(_0122_),
    .A2(_0117_),
    .A3(_0118_),
    .S1(net1805),
    .X(_2239_));
 sg13g2_nor2_1 _6436_ (.A(net1800),
    .B(_2239_),
    .Y(_2240_));
 sg13g2_or2_1 _6437_ (.X(_2241_),
    .B(_2239_),
    .A(net1833));
 sg13g2_nand2_1 _6438_ (.Y(_2242_),
    .A(_0787_),
    .B(net1788));
 sg13g2_xor2_1 _6439_ (.B(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A(net2037),
    .X(_2243_));
 sg13g2_xnor2_1 _6440_ (.Y(_2244_),
    .A(_0216_),
    .B(_2243_));
 sg13g2_nor3_1 _6441_ (.A(_2177_),
    .B(_2180_),
    .C(_2244_),
    .Y(_2245_));
 sg13g2_o21ai_1 _6442_ (.B1(_2244_),
    .Y(_2246_),
    .A1(_2177_),
    .A2(_2180_));
 sg13g2_nor2_1 _6443_ (.A(net1873),
    .B(_2245_),
    .Y(_2247_));
 sg13g2_and3_1 _6444_ (.X(_2248_),
    .A(net2030),
    .B(\z80.tv80s.i_tv80_core.BusB[6] ),
    .C(_1801_));
 sg13g2_xor2_1 _6445_ (.B(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A(net2030),
    .X(_2249_));
 sg13g2_a221oi_1 _6446_ (.B2(_1796_),
    .C1(_2248_),
    .B1(_2249_),
    .A1(_2246_),
    .Y(_2250_),
    .A2(_2247_));
 sg13g2_nand2_1 _6447_ (.Y(_2251_),
    .A(net1874),
    .B(_2250_));
 sg13g2_nand2b_1 _6448_ (.Y(_2252_),
    .B(_2192_),
    .A_N(net2029));
 sg13g2_xor2_1 _6449_ (.B(_2252_),
    .A(_0216_),
    .X(_2253_));
 sg13g2_or2_1 _6450_ (.X(_2254_),
    .B(_2253_),
    .A(_2194_));
 sg13g2_a21oi_1 _6451_ (.A1(_2194_),
    .A2(_2253_),
    .Y(_2255_),
    .B1(_0664_));
 sg13g2_xor2_1 _6452_ (.B(_2206_),
    .A(_2201_),
    .X(_2256_));
 sg13g2_a22oi_1 _6453_ (.Y(_2257_),
    .B1(_2256_),
    .B2(_0664_),
    .A2(_2255_),
    .A1(_2254_));
 sg13g2_nand2b_1 _6454_ (.Y(_2258_),
    .B(_1816_),
    .A_N(_2257_));
 sg13g2_a21oi_1 _6455_ (.A1(net1864),
    .A2(_1823_),
    .Y(_2259_),
    .B1(_1821_));
 sg13g2_a21o_1 _6456_ (.A2(net1864),
    .A1(_0223_),
    .B1(_2259_),
    .X(_2260_));
 sg13g2_nor2_1 _6457_ (.A(_0223_),
    .B(net1864),
    .Y(_2261_));
 sg13g2_nor2_1 _6458_ (.A(net2076),
    .B(_0215_),
    .Y(_2262_));
 sg13g2_a21oi_2 _6459_ (.B1(_2262_),
    .Y(_2263_),
    .A2(_0781_),
    .A1(net2076));
 sg13g2_inv_1 _6460_ (.Y(_2264_),
    .A(_2263_));
 sg13g2_o21ai_1 _6461_ (.B1(_1780_),
    .Y(_2265_),
    .A1(net1863),
    .A2(_2263_));
 sg13g2_a221oi_1 _6462_ (.B2(_2261_),
    .C1(_2265_),
    .B1(_1812_),
    .A1(net2031),
    .Y(_2266_),
    .A2(_1808_));
 sg13g2_nand3_1 _6463_ (.B(_2260_),
    .C(_2266_),
    .A(_2258_),
    .Y(_2267_));
 sg13g2_nand3_1 _6464_ (.B(_2251_),
    .C(_2267_),
    .A(net2032),
    .Y(_2268_));
 sg13g2_o21ai_1 _6465_ (.B1(_2268_),
    .Y(_2269_),
    .A1(net2032),
    .A2(_0719_));
 sg13g2_o21ai_1 _6466_ (.B1(_2242_),
    .Y(_2270_),
    .A1(net1788),
    .A2(_2269_));
 sg13g2_inv_1 _6467_ (.Y(_2271_),
    .A(_2270_));
 sg13g2_o21ai_1 _6468_ (.B1(net1825),
    .Y(_2272_),
    .A1(net1790),
    .A2(_2270_));
 sg13g2_a22oi_1 _6469_ (.Y(_2273_),
    .B1(net1735),
    .B2(_0121_),
    .A2(net1741),
    .A1(_0122_));
 sg13g2_a22oi_1 _6470_ (.Y(_2274_),
    .B1(net1736),
    .B2(_0117_),
    .A2(net1739),
    .A1(_0119_));
 sg13g2_and2_1 _6471_ (.A(_2273_),
    .B(_2274_),
    .X(_2275_));
 sg13g2_a22oi_1 _6472_ (.Y(_2276_),
    .B1(net1746),
    .B2(_0124_),
    .A2(_1749_),
    .A1(_0123_));
 sg13g2_a22oi_1 _6473_ (.Y(_2277_),
    .B1(net1742),
    .B2(_0120_),
    .A2(net1745),
    .A1(_0118_));
 sg13g2_nand3_1 _6474_ (.B(_2276_),
    .C(_2277_),
    .A(_2275_),
    .Y(_2278_));
 sg13g2_nand2b_1 _6475_ (.Y(_2279_),
    .B(net1823),
    .A_N(_2278_));
 sg13g2_and2_1 _6476_ (.A(net1815),
    .B(_2278_),
    .X(_2280_));
 sg13g2_xnor2_1 _6477_ (.Y(_2281_),
    .A(net1823),
    .B(_2278_));
 sg13g2_a221oi_1 _6478_ (.B2(_2230_),
    .C1(_2228_),
    .B1(_2162_),
    .A1(net1823),
    .Y(_2282_),
    .A2(_2160_));
 sg13g2_xnor2_1 _6479_ (.Y(_2283_),
    .A(_2281_),
    .B(_2282_));
 sg13g2_a21oi_2 _6480_ (.B1(_2272_),
    .Y(_2284_),
    .A2(_2283_),
    .A1(net1790));
 sg13g2_o21ai_1 _6481_ (.B1(net1833),
    .Y(_2285_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[14] ),
    .A2(net1827));
 sg13g2_o21ai_1 _6482_ (.B1(_2241_),
    .Y(_2286_),
    .A1(_2284_),
    .A2(_2285_));
 sg13g2_mux2_1 _6483_ (.A0(net312),
    .A1(_2286_),
    .S(_1770_),
    .X(_0315_));
 sg13g2_nand2_1 _6484_ (.Y(_2287_),
    .A(net2030),
    .B(_2243_));
 sg13g2_nand2_2 _6485_ (.Y(_2288_),
    .A(_2246_),
    .B(_2287_));
 sg13g2_xnor2_1 _6486_ (.Y(_2289_),
    .A(_0781_),
    .B(_2288_));
 sg13g2_xnor2_1 _6487_ (.Y(_2290_),
    .A(net2037),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ));
 sg13g2_nand2_1 _6488_ (.Y(_2291_),
    .A(_2289_),
    .B(_2290_));
 sg13g2_nor2_1 _6489_ (.A(_2289_),
    .B(_2290_),
    .Y(_2292_));
 sg13g2_nor2_1 _6490_ (.A(_1788_),
    .B(_2292_),
    .Y(_2293_));
 sg13g2_nand2_1 _6491_ (.Y(_2294_),
    .A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ));
 sg13g2_nor2_1 _6492_ (.A(_1799_),
    .B(_2294_),
    .Y(_2295_));
 sg13g2_o21ai_1 _6493_ (.B1(_1796_),
    .Y(_2296_),
    .A1(\z80.tv80s.i_tv80_core.BusA[7] ),
    .A2(\z80.tv80s.i_tv80_core.BusB[7] ));
 sg13g2_a22oi_1 _6494_ (.Y(_2297_),
    .B1(_2296_),
    .B2(_2294_),
    .A2(_2295_),
    .A1(_1793_));
 sg13g2_a21oi_2 _6495_ (.B1(_2297_),
    .Y(_2298_),
    .A2(_2293_),
    .A1(_2291_));
 sg13g2_o21ai_1 _6496_ (.B1(_2203_),
    .Y(_2299_),
    .A1(_2202_),
    .A2(_2205_));
 sg13g2_nand3_1 _6497_ (.B(_2204_),
    .C(_2299_),
    .A(_0664_),
    .Y(_2300_));
 sg13g2_nor2_1 _6498_ (.A(net2030),
    .B(_2252_),
    .Y(_2301_));
 sg13g2_xnor2_1 _6499_ (.Y(_2302_),
    .A(_0781_),
    .B(_2301_));
 sg13g2_a21o_1 _6500_ (.A2(_2253_),
    .A1(_2193_),
    .B1(_2190_),
    .X(_2303_));
 sg13g2_a21oi_1 _6501_ (.A1(_2302_),
    .A2(_2303_),
    .Y(_2304_),
    .B1(_0664_));
 sg13g2_o21ai_1 _6502_ (.B1(_2304_),
    .Y(_2305_),
    .A1(_2302_),
    .A2(_2303_));
 sg13g2_nand2_1 _6503_ (.Y(_2306_),
    .A(_2300_),
    .B(_2305_));
 sg13g2_a21oi_1 _6504_ (.A1(_2300_),
    .A2(_2305_),
    .Y(_2307_),
    .B1(_1817_));
 sg13g2_a22oi_1 _6505_ (.Y(_2308_),
    .B1(_1052_),
    .B2(net2062),
    .A2(net1878),
    .A1(_0678_));
 sg13g2_nor2_1 _6506_ (.A(_0224_),
    .B(_2308_),
    .Y(_2309_));
 sg13g2_a221oi_1 _6507_ (.B2(_2309_),
    .C1(_2307_),
    .B1(_1812_),
    .A1(\z80.tv80s.i_tv80_core.BusA[7] ),
    .Y(_2310_),
    .A2(_1808_));
 sg13g2_nand2_1 _6508_ (.Y(_2311_),
    .A(_1823_),
    .B(_2308_));
 sg13g2_a22oi_1 _6509_ (.Y(_2312_),
    .B1(_2311_),
    .B2(_1822_),
    .A2(_2308_),
    .A1(_0224_));
 sg13g2_nor2b_1 _6510_ (.A(net2079),
    .B_N(net2031),
    .Y(_2313_));
 sg13g2_nand3_1 _6511_ (.B(\z80.tv80s.i_tv80_core.BusA[0] ),
    .C(_0815_),
    .A(net2077),
    .Y(_2314_));
 sg13g2_o21ai_1 _6512_ (.B1(_2314_),
    .Y(_2315_),
    .A1(_0210_),
    .A2(_1044_));
 sg13g2_nor3_1 _6513_ (.A(_1043_),
    .B(_2313_),
    .C(_2315_),
    .Y(_2316_));
 sg13g2_a21oi_2 _6514_ (.B1(_2316_),
    .Y(_2317_),
    .A2(net1936),
    .A1(net2077));
 sg13g2_nor2b_1 _6515_ (.A(net1863),
    .B_N(_2317_),
    .Y(_2318_));
 sg13g2_nor3_1 _6516_ (.A(net1874),
    .B(_2312_),
    .C(_2318_),
    .Y(_2319_));
 sg13g2_a22oi_1 _6517_ (.Y(_2320_),
    .B1(_2310_),
    .B2(_2319_),
    .A2(_2298_),
    .A1(net1874));
 sg13g2_nand2_1 _6518_ (.Y(_2321_),
    .A(net2032),
    .B(_2320_));
 sg13g2_a21oi_1 _6519_ (.A1(_0690_),
    .A2(net2043),
    .Y(_2322_),
    .B1(net1787));
 sg13g2_a22oi_1 _6520_ (.Y(_2323_),
    .B1(_2321_),
    .B2(_2322_),
    .A2(net1787),
    .A1(_0788_));
 sg13g2_a21o_1 _6521_ (.A2(_2323_),
    .A1(net1789),
    .B1(_1719_),
    .X(_2324_));
 sg13g2_o21ai_1 _6522_ (.B1(_2279_),
    .Y(_2325_),
    .A1(_2280_),
    .A2(_2282_));
 sg13g2_a22oi_1 _6523_ (.Y(_2326_),
    .B1(net1734),
    .B2(_0137_),
    .A2(net1748),
    .A1(_0139_));
 sg13g2_a22oi_1 _6524_ (.Y(_2327_),
    .B1(net1738),
    .B2(_0135_),
    .A2(net1740),
    .A1(_0138_));
 sg13g2_and2_1 _6525_ (.A(_2326_),
    .B(_2327_),
    .X(_2328_));
 sg13g2_a22oi_1 _6526_ (.Y(_2329_),
    .B1(net1744),
    .B2(_0134_),
    .A2(net1746),
    .A1(_0140_));
 sg13g2_a22oi_1 _6527_ (.Y(_2330_),
    .B1(net1736),
    .B2(_0133_),
    .A2(net1742),
    .A1(_0136_));
 sg13g2_nand3_1 _6528_ (.B(_2329_),
    .C(_2330_),
    .A(_2328_),
    .Y(_2331_));
 sg13g2_xnor2_1 _6529_ (.Y(_2332_),
    .A(net1815),
    .B(_2331_));
 sg13g2_xnor2_1 _6530_ (.Y(_2333_),
    .A(_2325_),
    .B(_2332_));
 sg13g2_a21oi_1 _6531_ (.A1(net1790),
    .A2(_2333_),
    .Y(_2334_),
    .B1(_2324_));
 sg13g2_o21ai_1 _6532_ (.B1(net1831),
    .Y(_2335_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[15] ),
    .A2(net1827));
 sg13g2_mux4_1 _6533_ (.S0(net1810),
    .A0(_0137_),
    .A1(_0138_),
    .A2(_0133_),
    .A3(_0134_),
    .S1(net1804),
    .X(_2336_));
 sg13g2_or2_1 _6534_ (.X(_2337_),
    .B(_2336_),
    .A(net1831));
 sg13g2_o21ai_1 _6535_ (.B1(_2337_),
    .Y(_2338_),
    .A1(_2334_),
    .A2(_2335_));
 sg13g2_mux2_1 _6536_ (.A0(net268),
    .A1(_2338_),
    .S(_1770_),
    .X(_0316_));
 sg13g2_nand2_2 _6537_ (.Y(_2339_),
    .A(_1769_),
    .B(net1740));
 sg13g2_mux2_1 _6538_ (.A0(_1972_),
    .A1(net442),
    .S(_2339_),
    .X(_0317_));
 sg13g2_mux2_1 _6539_ (.A0(_2020_),
    .A1(net411),
    .S(_2339_),
    .X(_0318_));
 sg13g2_mux2_1 _6540_ (.A0(_2069_),
    .A1(net439),
    .S(_2339_),
    .X(_0319_));
 sg13g2_mux2_1 _6541_ (.A0(_2121_),
    .A1(net365),
    .S(_2339_),
    .X(_0320_));
 sg13g2_mux2_1 _6542_ (.A0(_2175_),
    .A1(net424),
    .S(_2339_),
    .X(_0321_));
 sg13g2_mux2_1 _6543_ (.A0(_2238_),
    .A1(net361),
    .S(_2339_),
    .X(_0322_));
 sg13g2_mux2_1 _6544_ (.A0(_2286_),
    .A1(net379),
    .S(_2339_),
    .X(_0323_));
 sg13g2_mux2_1 _6545_ (.A0(_2338_),
    .A1(net400),
    .S(_2339_),
    .X(_0324_));
 sg13g2_nand2_2 _6546_ (.Y(_2340_),
    .A(_1769_),
    .B(net1734));
 sg13g2_mux2_1 _6547_ (.A0(_1972_),
    .A1(net402),
    .S(_2340_),
    .X(_0325_));
 sg13g2_mux2_1 _6548_ (.A0(_2020_),
    .A1(net431),
    .S(_2340_),
    .X(_0326_));
 sg13g2_mux2_1 _6549_ (.A0(_2069_),
    .A1(net403),
    .S(_2340_),
    .X(_0327_));
 sg13g2_mux2_1 _6550_ (.A0(_2121_),
    .A1(net374),
    .S(_2340_),
    .X(_0328_));
 sg13g2_mux2_1 _6551_ (.A0(_2175_),
    .A1(net416),
    .S(_2340_),
    .X(_0329_));
 sg13g2_mux2_1 _6552_ (.A0(_2238_),
    .A1(net393),
    .S(_2340_),
    .X(_0330_));
 sg13g2_mux2_1 _6553_ (.A0(_2286_),
    .A1(net429),
    .S(_2340_),
    .X(_0331_));
 sg13g2_mux2_1 _6554_ (.A0(_2338_),
    .A1(net435),
    .S(_2340_),
    .X(_0332_));
 sg13g2_and2_2 _6555_ (.A(_1769_),
    .B(net1742),
    .X(_2341_));
 sg13g2_mux2_1 _6556_ (.A0(net332),
    .A1(_1972_),
    .S(_2341_),
    .X(_0333_));
 sg13g2_mux2_1 _6557_ (.A0(net331),
    .A1(_2020_),
    .S(_2341_),
    .X(_0334_));
 sg13g2_mux2_1 _6558_ (.A0(net245),
    .A1(_2069_),
    .S(_2341_),
    .X(_0335_));
 sg13g2_mux2_1 _6559_ (.A0(net246),
    .A1(_2121_),
    .S(_2341_),
    .X(_0336_));
 sg13g2_mux2_1 _6560_ (.A0(net275),
    .A1(_2175_),
    .S(_2341_),
    .X(_0337_));
 sg13g2_mux2_1 _6561_ (.A0(net293),
    .A1(_2238_),
    .S(_2341_),
    .X(_0338_));
 sg13g2_mux2_1 _6562_ (.A0(net291),
    .A1(_2286_),
    .S(_2341_),
    .X(_0339_));
 sg13g2_mux2_1 _6563_ (.A0(net286),
    .A1(_2338_),
    .S(_2341_),
    .X(_0340_));
 sg13g2_nand2_2 _6564_ (.Y(_2342_),
    .A(_0032_),
    .B(_1133_));
 sg13g2_nand2_1 _6565_ (.Y(_2343_),
    .A(doe),
    .B(_2342_));
 sg13g2_nand2_1 _6566_ (.Y(_2344_),
    .A(net2020),
    .B(net2227));
 sg13g2_nand2_1 _6567_ (.Y(_2345_),
    .A(net228),
    .B(net2181));
 sg13g2_o21ai_1 _6568_ (.B1(_2345_),
    .Y(_0341_),
    .A1(_2343_),
    .A2(_2344_));
 sg13g2_nand2_1 _6569_ (.Y(_2346_),
    .A(net2123),
    .B(net2227));
 sg13g2_nor2_1 _6570_ (.A(_0028_),
    .B(_2346_),
    .Y(_2347_));
 sg13g2_a22oi_1 _6571_ (.Y(_2348_),
    .B1(_2342_),
    .B2(_2347_),
    .A2(net2181),
    .A1(net459));
 sg13g2_and2_1 _6572_ (.A(_1492_),
    .B(_1513_),
    .X(_2349_));
 sg13g2_nand4_1 _6573_ (.B(_0991_),
    .C(_0996_),
    .A(_0969_),
    .Y(_2350_),
    .D(_1252_));
 sg13g2_or2_1 _6574_ (.X(_2351_),
    .B(_2350_),
    .A(_1019_));
 sg13g2_nor2_1 _6575_ (.A(_0959_),
    .B(_1019_),
    .Y(_2352_));
 sg13g2_nor2_1 _6576_ (.A(_0959_),
    .B(_2351_),
    .Y(_2353_));
 sg13g2_nand2_1 _6577_ (.Y(_2354_),
    .A(_1012_),
    .B(_1494_));
 sg13g2_nor3_1 _6578_ (.A(_1242_),
    .B(_1502_),
    .C(_2354_),
    .Y(_2355_));
 sg13g2_nand3_1 _6579_ (.B(_2353_),
    .C(_2355_),
    .A(_2349_),
    .Y(_2356_));
 sg13g2_o21ai_1 _6580_ (.B1(_1097_),
    .Y(_2357_),
    .A1(_1012_),
    .A2(_1423_));
 sg13g2_nor2_2 _6581_ (.A(net2017),
    .B(_0887_),
    .Y(_2358_));
 sg13g2_mux2_2 _6582_ (.A0(_0870_),
    .A1(_2357_),
    .S(_2356_),
    .X(_2359_));
 sg13g2_nor2_2 _6583_ (.A(net2129),
    .B(_0872_),
    .Y(_2360_));
 sg13g2_nand2_1 _6584_ (.Y(_2361_),
    .A(net2080),
    .B(_0884_));
 sg13g2_o21ai_1 _6585_ (.B1(_1655_),
    .Y(_2362_),
    .A1(net2113),
    .A2(_2361_));
 sg13g2_a221oi_1 _6586_ (.B2(_1108_),
    .C1(_2362_),
    .B1(_2360_),
    .A1(_1281_),
    .Y(_2363_),
    .A2(_1295_));
 sg13g2_nand3_1 _6587_ (.B(_0033_),
    .C(_1138_),
    .A(net2103),
    .Y(_2364_));
 sg13g2_o21ai_1 _6588_ (.B1(_2342_),
    .Y(_2365_),
    .A1(net1893),
    .A2(_2363_));
 sg13g2_a21oi_1 _6589_ (.A1(net2169),
    .A2(_2359_),
    .Y(_2366_),
    .B1(_2365_));
 sg13g2_nand2_1 _6590_ (.Y(_2367_),
    .A(_2364_),
    .B(_2366_));
 sg13g2_nand2_1 _6591_ (.Y(_2368_),
    .A(_2343_),
    .B(_2367_));
 sg13g2_nand4_1 _6592_ (.B(_1062_),
    .C(_1246_),
    .A(_0998_),
    .Y(_2369_),
    .D(_1252_));
 sg13g2_nand4_1 _6593_ (.B(net1883),
    .C(_1245_),
    .A(_1002_),
    .Y(_2370_),
    .D(_2358_));
 sg13g2_nor2_1 _6594_ (.A(_1316_),
    .B(_1673_),
    .Y(_2371_));
 sg13g2_nor4_2 _6595_ (.A(_1163_),
    .B(_1668_),
    .C(_2369_),
    .Y(_2372_),
    .D(_2370_));
 sg13g2_a221oi_1 _6596_ (.B2(_1667_),
    .C1(_2371_),
    .B1(_2372_),
    .A1(_0868_),
    .Y(_2373_),
    .A2(_1685_));
 sg13g2_nor2_1 _6597_ (.A(_2344_),
    .B(_2373_),
    .Y(_2374_));
 sg13g2_and2_1 _6598_ (.A(_2368_),
    .B(_2374_),
    .X(_2375_));
 sg13g2_nand2b_1 _6599_ (.Y(_0342_),
    .B(_2348_),
    .A_N(_2375_));
 sg13g2_or3_1 _6600_ (.A(doe),
    .B(_2344_),
    .C(_2367_),
    .X(_2376_));
 sg13g2_nand2_1 _6601_ (.Y(_2377_),
    .A(net460),
    .B(net2181));
 sg13g2_nand4_1 _6602_ (.B(net2227),
    .C(_0028_),
    .A(net2123),
    .Y(_2378_),
    .D(_2342_));
 sg13g2_nand3_1 _6603_ (.B(_2377_),
    .C(_2378_),
    .A(_2376_),
    .Y(_0343_));
 sg13g2_a21oi_1 _6604_ (.A1(_2368_),
    .A2(_2373_),
    .Y(_2379_),
    .B1(net2132));
 sg13g2_a21oi_1 _6605_ (.A1(_0028_),
    .A2(_2342_),
    .Y(_2380_),
    .B1(_1751_));
 sg13g2_nor3_1 _6606_ (.A(net2181),
    .B(_2379_),
    .C(_2380_),
    .Y(_2381_));
 sg13g2_a21o_1 _6607_ (.A2(net2181),
    .A1(net326),
    .B1(_2381_),
    .X(_0344_));
 sg13g2_nor2b_2 _6608_ (.A(_1766_),
    .B_N(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .Y(_2382_));
 sg13g2_nand2b_2 _6609_ (.Y(_2383_),
    .B(_2382_),
    .A_N(_1761_));
 sg13g2_a21oi_2 _6610_ (.B1(net1961),
    .Y(_2384_),
    .A2(_2383_),
    .A1(_1754_));
 sg13g2_and2_2 _6611_ (.A(net1749),
    .B(_2384_),
    .X(_2385_));
 sg13g2_o21ai_1 _6612_ (.B1(_1832_),
    .Y(_2386_),
    .A1(_1772_),
    .A2(_1888_));
 sg13g2_mux4_1 _6613_ (.S0(net1811),
    .A0(_0155_),
    .A1(_0156_),
    .A2(_0151_),
    .A3(_0152_),
    .S1(net1803),
    .X(_2387_));
 sg13g2_o21ai_1 _6614_ (.B1(net1830),
    .Y(_2388_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[0] ),
    .A2(net1826));
 sg13g2_nand2b_1 _6615_ (.Y(_2389_),
    .B(_2386_),
    .A_N(_2388_));
 sg13g2_o21ai_1 _6616_ (.B1(_2389_),
    .Y(_2390_),
    .A1(net1830),
    .A2(_2387_));
 sg13g2_mux2_1 _6617_ (.A0(net329),
    .A1(_2390_),
    .S(_2385_),
    .X(_0345_));
 sg13g2_nand2_1 _6618_ (.Y(_2391_),
    .A(_1887_),
    .B(_1889_));
 sg13g2_nand3_1 _6619_ (.B(_1890_),
    .C(_2391_),
    .A(net1790),
    .Y(_2392_));
 sg13g2_nand2_1 _6620_ (.Y(_2393_),
    .A(_2006_),
    .B(_2392_));
 sg13g2_o21ai_1 _6621_ (.B1(_2393_),
    .Y(_2394_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[1] ),
    .A2(net1825));
 sg13g2_mux2_1 _6622_ (.A0(_0160_),
    .A1(_0159_),
    .S(net1812),
    .X(_2395_));
 sg13g2_nand2_1 _6623_ (.Y(_2396_),
    .A(_0163_),
    .B(net1812));
 sg13g2_a21oi_1 _6624_ (.A1(_0164_),
    .A2(net1807),
    .Y(_2397_),
    .B1(net1802));
 sg13g2_a21oi_1 _6625_ (.A1(_2396_),
    .A2(_2397_),
    .Y(_2398_),
    .B1(net1797));
 sg13g2_o21ai_1 _6626_ (.B1(_2398_),
    .Y(_2399_),
    .A1(net1785),
    .A2(_2395_));
 sg13g2_nor2_1 _6627_ (.A(net1829),
    .B(_2399_),
    .Y(_2400_));
 sg13g2_a21oi_2 _6628_ (.B1(_2400_),
    .Y(_2401_),
    .A2(_2394_),
    .A1(net1829));
 sg13g2_mux2_1 _6629_ (.A0(net359),
    .A1(_2401_),
    .S(_2385_),
    .X(_0346_));
 sg13g2_nor2_1 _6630_ (.A(_1891_),
    .B(_1899_),
    .Y(_2402_));
 sg13g2_nor3_1 _6631_ (.A(net1789),
    .B(_1901_),
    .C(_2402_),
    .Y(_2403_));
 sg13g2_nand2b_1 _6632_ (.Y(_2404_),
    .B(_1719_),
    .A_N(\z80.tv80s.i_tv80_core.RegBusA_r[2] ));
 sg13g2_mux4_1 _6633_ (.S0(net1808),
    .A0(_0065_),
    .A1(_0066_),
    .A2(_0061_),
    .A3(_0062_),
    .S1(net1803),
    .X(_2405_));
 sg13g2_nor2_1 _6634_ (.A(net1798),
    .B(_2405_),
    .Y(_2406_));
 sg13g2_nor2_1 _6635_ (.A(_0064_),
    .B(_1956_),
    .Y(_2407_));
 sg13g2_o21ai_1 _6636_ (.B1(net1803),
    .Y(_2408_),
    .A1(_0063_),
    .A2(net2164));
 sg13g2_a22oi_1 _6637_ (.Y(_2409_),
    .B1(net1808),
    .B2(_0703_),
    .A2(net2009),
    .A1(_0704_));
 sg13g2_o21ai_1 _6638_ (.B1(net1798),
    .Y(_2410_),
    .A1(_2407_),
    .A2(_2408_));
 sg13g2_a21oi_1 _6639_ (.A1(net1786),
    .A2(_2409_),
    .Y(_2411_),
    .B1(_2410_));
 sg13g2_o21ai_1 _6640_ (.B1(_2404_),
    .Y(_2412_),
    .A1(_2051_),
    .A2(_2403_));
 sg13g2_nor2_1 _6641_ (.A(net1830),
    .B(_2406_),
    .Y(_2413_));
 sg13g2_a21oi_2 _6642_ (.B1(_2413_),
    .Y(_2414_),
    .A2(_2412_),
    .A1(net1830));
 sg13g2_mux2_1 _6643_ (.A0(net237),
    .A1(_2414_),
    .S(_2385_),
    .X(_0347_));
 sg13g2_nor2_1 _6644_ (.A(_1898_),
    .B(_1901_),
    .Y(_2415_));
 sg13g2_xnor2_1 _6645_ (.Y(_2416_),
    .A(_1868_),
    .B(_2415_));
 sg13g2_a21oi_1 _6646_ (.A1(net1790),
    .A2(_2416_),
    .Y(_2417_),
    .B1(_2102_));
 sg13g2_o21ai_1 _6647_ (.B1(net1828),
    .Y(_2418_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[3] ),
    .A2(net1825));
 sg13g2_mux4_1 _6648_ (.S0(net1808),
    .A0(_0081_),
    .A1(_0082_),
    .A2(_0077_),
    .A3(_0078_),
    .S1(net1803),
    .X(_2419_));
 sg13g2_or2_1 _6649_ (.X(_2420_),
    .B(_2419_),
    .A(net1828));
 sg13g2_nor2_1 _6650_ (.A(_0080_),
    .B(net1812),
    .Y(_2421_));
 sg13g2_o21ai_1 _6651_ (.B1(_2420_),
    .Y(_2422_),
    .A1(_2417_),
    .A2(_2418_));
 sg13g2_mux2_1 _6652_ (.A0(net254),
    .A1(_2422_),
    .S(_2385_),
    .X(_0348_));
 sg13g2_mux4_1 _6653_ (.S0(net1807),
    .A0(_0097_),
    .A1(_0098_),
    .A2(_0093_),
    .A3(_0094_),
    .S1(net1802),
    .X(_2423_));
 sg13g2_or2_1 _6654_ (.X(_2424_),
    .B(_2423_),
    .A(net1828));
 sg13g2_nor2b_1 _6655_ (.A(_1904_),
    .B_N(_1937_),
    .Y(_2425_));
 sg13g2_xor2_1 _6656_ (.B(_1937_),
    .A(_1904_),
    .X(_2426_));
 sg13g2_nor2_1 _6657_ (.A(net1789),
    .B(_2426_),
    .Y(_2427_));
 sg13g2_nor2_1 _6658_ (.A(_2148_),
    .B(_2427_),
    .Y(_2428_));
 sg13g2_o21ai_1 _6659_ (.B1(net1828),
    .Y(_2429_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[4] ),
    .A2(net1825));
 sg13g2_o21ai_1 _6660_ (.B1(_2424_),
    .Y(_2430_),
    .A1(_2428_),
    .A2(_2429_));
 sg13g2_mux2_1 _6661_ (.A0(net313),
    .A1(_2430_),
    .S(_2385_),
    .X(_0349_));
 sg13g2_nor2_1 _6662_ (.A(_1936_),
    .B(_2425_),
    .Y(_2431_));
 sg13g2_xor2_1 _6663_ (.B(_2431_),
    .A(_1929_),
    .X(_2432_));
 sg13g2_nor2_1 _6664_ (.A(net1789),
    .B(_2432_),
    .Y(_2433_));
 sg13g2_nor2_1 _6665_ (.A(_2221_),
    .B(_2433_),
    .Y(_2434_));
 sg13g2_a22oi_1 _6666_ (.Y(_2435_),
    .B1(net1807),
    .B2(_0716_),
    .A2(net2009),
    .A1(_0717_));
 sg13g2_nor2_1 _6667_ (.A(_0112_),
    .B(net1812),
    .Y(_2436_));
 sg13g2_o21ai_1 _6668_ (.B1(net1802),
    .Y(_2437_),
    .A1(_0111_),
    .A2(net2164));
 sg13g2_a21oi_1 _6669_ (.A1(net1785),
    .A2(_2435_),
    .Y(_2438_),
    .B1(_1963_));
 sg13g2_o21ai_1 _6670_ (.B1(_2438_),
    .Y(_2439_),
    .A1(_2436_),
    .A2(_2437_));
 sg13g2_mux4_1 _6671_ (.S0(net1807),
    .A0(_0113_),
    .A1(_0114_),
    .A2(_0109_),
    .A3(_0110_),
    .S1(net1802),
    .X(_2440_));
 sg13g2_o21ai_1 _6672_ (.B1(_2439_),
    .Y(_2441_),
    .A1(net1797),
    .A2(_2440_));
 sg13g2_o21ai_1 _6673_ (.B1(net1828),
    .Y(_2442_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[5] ),
    .A2(net1825));
 sg13g2_or2_1 _6674_ (.X(_2443_),
    .B(_2440_),
    .A(net1828));
 sg13g2_o21ai_1 _6675_ (.B1(_2443_),
    .Y(_2444_),
    .A1(_2434_),
    .A2(_2442_));
 sg13g2_mux2_1 _6676_ (.A0(net299),
    .A1(_2444_),
    .S(_2385_),
    .X(_0350_));
 sg13g2_mux4_1 _6677_ (.S0(net1808),
    .A0(_0129_),
    .A1(_0130_),
    .A2(_0125_),
    .A3(_0126_),
    .S1(net1803),
    .X(_2445_));
 sg13g2_or2_1 _6678_ (.X(_2446_),
    .B(_2445_),
    .A(net1829));
 sg13g2_a21oi_1 _6679_ (.A1(_1929_),
    .A2(_2425_),
    .Y(_2447_),
    .B1(_1940_));
 sg13g2_xnor2_1 _6680_ (.Y(_2448_),
    .A(_1921_),
    .B(_2447_));
 sg13g2_a21oi_1 _6681_ (.A1(net1790),
    .A2(_2448_),
    .Y(_2449_),
    .B1(_2272_));
 sg13g2_o21ai_1 _6682_ (.B1(net1828),
    .Y(_2450_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[6] ),
    .A2(net1825));
 sg13g2_o21ai_1 _6683_ (.B1(_2446_),
    .Y(_2451_),
    .A1(_2449_),
    .A2(_2450_));
 sg13g2_mux2_1 _6684_ (.A0(net308),
    .A1(_2451_),
    .S(_2385_),
    .X(_0351_));
 sg13g2_o21ai_1 _6685_ (.B1(_1920_),
    .Y(_2452_),
    .A1(_1922_),
    .A2(_2447_));
 sg13g2_xor2_1 _6686_ (.B(_2452_),
    .A(_1911_),
    .X(_2453_));
 sg13g2_a21oi_1 _6687_ (.A1(net1791),
    .A2(_2453_),
    .Y(_2454_),
    .B1(_2324_));
 sg13g2_mux4_1 _6688_ (.S0(net1811),
    .A0(_0145_),
    .A1(_0146_),
    .A2(_0141_),
    .A3(_0142_),
    .S1(net1806),
    .X(_2455_));
 sg13g2_or2_1 _6689_ (.X(_2456_),
    .B(_2455_),
    .A(net1830));
 sg13g2_o21ai_1 _6690_ (.B1(net1828),
    .Y(_2457_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[7] ),
    .A2(net1826));
 sg13g2_o21ai_1 _6691_ (.B1(_2456_),
    .Y(_2458_),
    .A1(_2454_),
    .A2(_2457_));
 sg13g2_mux2_1 _6692_ (.A0(net297),
    .A1(_2458_),
    .S(_2385_),
    .X(_0352_));
 sg13g2_and2_2 _6693_ (.A(_1769_),
    .B(net1746),
    .X(_2459_));
 sg13g2_mux2_1 _6694_ (.A0(net321),
    .A1(_1972_),
    .S(_2459_),
    .X(_0353_));
 sg13g2_mux2_1 _6695_ (.A0(net256),
    .A1(_2020_),
    .S(_2459_),
    .X(_0354_));
 sg13g2_mux2_1 _6696_ (.A0(net320),
    .A1(_2069_),
    .S(_2459_),
    .X(_0355_));
 sg13g2_mux2_1 _6697_ (.A0(net287),
    .A1(_2121_),
    .S(_2459_),
    .X(_0356_));
 sg13g2_mux2_1 _6698_ (.A0(net272),
    .A1(_2175_),
    .S(_2459_),
    .X(_0357_));
 sg13g2_mux2_1 _6699_ (.A0(net257),
    .A1(_2238_),
    .S(_2459_),
    .X(_0358_));
 sg13g2_mux2_1 _6700_ (.A0(net288),
    .A1(_2286_),
    .S(_2459_),
    .X(_0359_));
 sg13g2_mux2_1 _6701_ (.A0(net270),
    .A1(_2338_),
    .S(_2459_),
    .X(_0360_));
 sg13g2_nand2_2 _6702_ (.Y(_2460_),
    .A(net1741),
    .B(_2384_));
 sg13g2_mux2_1 _6703_ (.A0(_2390_),
    .A1(net447),
    .S(_2460_),
    .X(_0361_));
 sg13g2_mux2_1 _6704_ (.A0(_2401_),
    .A1(net483),
    .S(_2460_),
    .X(_0362_));
 sg13g2_mux2_1 _6705_ (.A0(_2414_),
    .A1(net426),
    .S(_2460_),
    .X(_0363_));
 sg13g2_mux2_1 _6706_ (.A0(_2422_),
    .A1(net392),
    .S(_2460_),
    .X(_0364_));
 sg13g2_mux2_1 _6707_ (.A0(_2430_),
    .A1(net385),
    .S(_2460_),
    .X(_0365_));
 sg13g2_mux2_1 _6708_ (.A0(_2444_),
    .A1(net398),
    .S(_2460_),
    .X(_0366_));
 sg13g2_mux2_1 _6709_ (.A0(_2451_),
    .A1(net409),
    .S(_2460_),
    .X(_0367_));
 sg13g2_mux2_1 _6710_ (.A0(_2458_),
    .A1(net420),
    .S(_2460_),
    .X(_0368_));
 sg13g2_nand2_2 _6711_ (.Y(_2461_),
    .A(_1769_),
    .B(net1744));
 sg13g2_mux2_1 _6712_ (.A0(_1972_),
    .A1(net441),
    .S(_2461_),
    .X(_0369_));
 sg13g2_mux2_1 _6713_ (.A0(_2020_),
    .A1(net438),
    .S(_2461_),
    .X(_0370_));
 sg13g2_mux2_1 _6714_ (.A0(_2069_),
    .A1(net373),
    .S(_2461_),
    .X(_0371_));
 sg13g2_mux2_1 _6715_ (.A0(_2121_),
    .A1(net406),
    .S(_2461_),
    .X(_0372_));
 sg13g2_mux2_1 _6716_ (.A0(_2175_),
    .A1(net378),
    .S(_2461_),
    .X(_0373_));
 sg13g2_mux2_1 _6717_ (.A0(_2238_),
    .A1(net414),
    .S(_2461_),
    .X(_0374_));
 sg13g2_mux2_1 _6718_ (.A0(_2286_),
    .A1(net405),
    .S(_2461_),
    .X(_0375_));
 sg13g2_mux2_1 _6719_ (.A0(_2338_),
    .A1(net410),
    .S(_2461_),
    .X(_0376_));
 sg13g2_nand2_1 _6720_ (.Y(_2462_),
    .A(net1737),
    .B(_2384_));
 sg13g2_mux2_1 _6721_ (.A0(_2390_),
    .A1(net454),
    .S(_2462_),
    .X(_0377_));
 sg13g2_nor2_1 _6722_ (.A(_2401_),
    .B(net1729),
    .Y(_2463_));
 sg13g2_a21oi_1 _6723_ (.A1(_0699_),
    .A2(net1729),
    .Y(_0378_),
    .B1(_2463_));
 sg13g2_mux2_1 _6724_ (.A0(_2414_),
    .A1(net401),
    .S(net1729),
    .X(_0379_));
 sg13g2_mux2_1 _6725_ (.A0(_2422_),
    .A1(net423),
    .S(net1729),
    .X(_0380_));
 sg13g2_mux2_1 _6726_ (.A0(_2430_),
    .A1(net380),
    .S(net1729),
    .X(_0381_));
 sg13g2_mux2_1 _6727_ (.A0(_2444_),
    .A1(net436),
    .S(net1729),
    .X(_0382_));
 sg13g2_mux2_1 _6728_ (.A0(_2451_),
    .A1(net391),
    .S(net1729),
    .X(_0383_));
 sg13g2_mux2_1 _6729_ (.A0(_2458_),
    .A1(net417),
    .S(net1729),
    .X(_0384_));
 sg13g2_nand2_2 _6730_ (.Y(_2464_),
    .A(net1745),
    .B(_2384_));
 sg13g2_mux2_1 _6731_ (.A0(_2390_),
    .A1(net452),
    .S(_2464_),
    .X(_0385_));
 sg13g2_mux2_1 _6732_ (.A0(_2401_),
    .A1(net455),
    .S(_2464_),
    .X(_0386_));
 sg13g2_mux2_1 _6733_ (.A0(_2414_),
    .A1(net418),
    .S(_2464_),
    .X(_0387_));
 sg13g2_mux2_1 _6734_ (.A0(_2422_),
    .A1(net407),
    .S(_2464_),
    .X(_0388_));
 sg13g2_mux2_1 _6735_ (.A0(_2430_),
    .A1(net376),
    .S(_2464_),
    .X(_0389_));
 sg13g2_mux2_1 _6736_ (.A0(_2444_),
    .A1(net384),
    .S(_2464_),
    .X(_0390_));
 sg13g2_mux2_1 _6737_ (.A0(_2451_),
    .A1(net427),
    .S(_2464_),
    .X(_0391_));
 sg13g2_mux2_1 _6738_ (.A0(_2458_),
    .A1(net415),
    .S(_2464_),
    .X(_0392_));
 sg13g2_and2_2 _6739_ (.A(_1769_),
    .B(net1738),
    .X(_2465_));
 sg13g2_mux2_1 _6740_ (.A0(net307),
    .A1(_1972_),
    .S(_2465_),
    .X(_0393_));
 sg13g2_mux2_1 _6741_ (.A0(net289),
    .A1(_2020_),
    .S(_2465_),
    .X(_0394_));
 sg13g2_mux2_1 _6742_ (.A0(net234),
    .A1(_2069_),
    .S(_2465_),
    .X(_0395_));
 sg13g2_mux2_1 _6743_ (.A0(net273),
    .A1(_2121_),
    .S(_2465_),
    .X(_0396_));
 sg13g2_mux2_1 _6744_ (.A0(net281),
    .A1(_2175_),
    .S(_2465_),
    .X(_0397_));
 sg13g2_mux2_1 _6745_ (.A0(net292),
    .A1(_2238_),
    .S(_2465_),
    .X(_0398_));
 sg13g2_mux2_1 _6746_ (.A0(net296),
    .A1(_2286_),
    .S(_2465_),
    .X(_0399_));
 sg13g2_mux2_1 _6747_ (.A0(net255),
    .A1(_2338_),
    .S(_2465_),
    .X(_0400_));
 sg13g2_and2_2 _6748_ (.A(net1743),
    .B(_2384_),
    .X(_2466_));
 sg13g2_mux2_1 _6749_ (.A0(net350),
    .A1(_2390_),
    .S(_2466_),
    .X(_0401_));
 sg13g2_mux2_1 _6750_ (.A0(net395),
    .A1(_2401_),
    .S(_2466_),
    .X(_0402_));
 sg13g2_mux2_1 _6751_ (.A0(net238),
    .A1(_2414_),
    .S(_2466_),
    .X(_0403_));
 sg13g2_mux2_1 _6752_ (.A0(net261),
    .A1(_2422_),
    .S(_2466_),
    .X(_0404_));
 sg13g2_mux2_1 _6753_ (.A0(net298),
    .A1(_2430_),
    .S(_2466_),
    .X(_0405_));
 sg13g2_mux2_1 _6754_ (.A0(net259),
    .A1(_2444_),
    .S(_2466_),
    .X(_0406_));
 sg13g2_mux2_1 _6755_ (.A0(net302),
    .A1(_2451_),
    .S(_2466_),
    .X(_0407_));
 sg13g2_mux2_1 _6756_ (.A0(net300),
    .A1(_2458_),
    .S(_2466_),
    .X(_0408_));
 sg13g2_nand2_1 _6757_ (.Y(_2467_),
    .A(net1735),
    .B(_2384_));
 sg13g2_mux2_1 _6758_ (.A0(_2390_),
    .A1(net456),
    .S(_2467_),
    .X(_0409_));
 sg13g2_nor2_1 _6759_ (.A(_2401_),
    .B(net1728),
    .Y(_2468_));
 sg13g2_a21oi_1 _6760_ (.A1(_0700_),
    .A2(net1728),
    .Y(_0410_),
    .B1(_2468_));
 sg13g2_mux2_1 _6761_ (.A0(_2414_),
    .A1(net371),
    .S(net1728),
    .X(_0411_));
 sg13g2_mux2_1 _6762_ (.A0(_2422_),
    .A1(net389),
    .S(net1728),
    .X(_0412_));
 sg13g2_mux2_1 _6763_ (.A0(_2430_),
    .A1(net390),
    .S(net1728),
    .X(_0413_));
 sg13g2_mux2_1 _6764_ (.A0(_2444_),
    .A1(net386),
    .S(net1728),
    .X(_0414_));
 sg13g2_mux2_1 _6765_ (.A0(_2451_),
    .A1(net428),
    .S(net1728),
    .X(_0415_));
 sg13g2_mux2_1 _6766_ (.A0(_2458_),
    .A1(net432),
    .S(net1728),
    .X(_0416_));
 sg13g2_and2_2 _6767_ (.A(net1747),
    .B(_2384_),
    .X(_2469_));
 sg13g2_mux2_1 _6768_ (.A0(net352),
    .A1(_2390_),
    .S(_2469_),
    .X(_0417_));
 sg13g2_mux2_1 _6769_ (.A0(net364),
    .A1(_2401_),
    .S(_2469_),
    .X(_0418_));
 sg13g2_mux2_1 _6770_ (.A0(net294),
    .A1(_2414_),
    .S(_2469_),
    .X(_0419_));
 sg13g2_mux2_1 _6771_ (.A0(net301),
    .A1(_2422_),
    .S(_2469_),
    .X(_0420_));
 sg13g2_mux2_1 _6772_ (.A0(net285),
    .A1(_2430_),
    .S(_2469_),
    .X(_0421_));
 sg13g2_mux2_1 _6773_ (.A0(net290),
    .A1(_2444_),
    .S(_2469_),
    .X(_0422_));
 sg13g2_mux2_1 _6774_ (.A0(net262),
    .A1(_2451_),
    .S(_2469_),
    .X(_0423_));
 sg13g2_mux2_1 _6775_ (.A0(net295),
    .A1(_2458_),
    .S(_2469_),
    .X(_0424_));
 sg13g2_nand2_2 _6776_ (.Y(_2470_),
    .A(_1769_),
    .B(net1736));
 sg13g2_mux2_1 _6777_ (.A0(_1972_),
    .A1(net433),
    .S(_2470_),
    .X(_0425_));
 sg13g2_mux2_1 _6778_ (.A0(_2020_),
    .A1(net412),
    .S(_2470_),
    .X(_0426_));
 sg13g2_mux2_1 _6779_ (.A0(_2069_),
    .A1(net437),
    .S(_2470_),
    .X(_0427_));
 sg13g2_mux2_1 _6780_ (.A0(_2121_),
    .A1(net425),
    .S(_2470_),
    .X(_0428_));
 sg13g2_mux2_1 _6781_ (.A0(_2175_),
    .A1(net419),
    .S(_2470_),
    .X(_0429_));
 sg13g2_mux2_1 _6782_ (.A0(_2238_),
    .A1(net360),
    .S(_2470_),
    .X(_0430_));
 sg13g2_mux2_1 _6783_ (.A0(_2286_),
    .A1(net388),
    .S(_2470_),
    .X(_0431_));
 sg13g2_mux2_1 _6784_ (.A0(_2338_),
    .A1(net413),
    .S(_2470_),
    .X(_0432_));
 sg13g2_and2_2 _6785_ (.A(net1739),
    .B(_2384_),
    .X(_2471_));
 sg13g2_mux2_1 _6786_ (.A0(net372),
    .A1(_2390_),
    .S(_2471_),
    .X(_0433_));
 sg13g2_mux2_1 _6787_ (.A0(net440),
    .A1(_2401_),
    .S(_2471_),
    .X(_0434_));
 sg13g2_mux2_1 _6788_ (.A0(net247),
    .A1(_2414_),
    .S(_2471_),
    .X(_0435_));
 sg13g2_mux2_1 _6789_ (.A0(net284),
    .A1(_2422_),
    .S(_2471_),
    .X(_0436_));
 sg13g2_mux2_1 _6790_ (.A0(net263),
    .A1(_2430_),
    .S(_2471_),
    .X(_0437_));
 sg13g2_mux2_1 _6791_ (.A0(net239),
    .A1(_2444_),
    .S(_2471_),
    .X(_0438_));
 sg13g2_mux2_1 _6792_ (.A0(net305),
    .A1(_2451_),
    .S(_2471_),
    .X(_0439_));
 sg13g2_mux2_1 _6793_ (.A0(net269),
    .A1(_2458_),
    .S(_2471_),
    .X(_0440_));
 sg13g2_nand2_1 _6794_ (.Y(_2472_),
    .A(net2183),
    .B(net485));
 sg13g2_o21ai_1 _6795_ (.B1(net2123),
    .Y(_2473_),
    .A1(\z80.tv80s.i_tv80_core.IntCycle ),
    .A2(\z80.tv80s.i_tv80_core.NMICycle ));
 sg13g2_o21ai_1 _6796_ (.B1(_2473_),
    .Y(_2474_),
    .A1(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .A2(_2373_));
 sg13g2_nand2_1 _6797_ (.Y(_2475_),
    .A(net2227),
    .B(_2474_));
 sg13g2_o21ai_1 _6798_ (.B1(_2472_),
    .Y(_0441_),
    .A1(net1689),
    .A2(_2475_));
 sg13g2_nand2_1 _6799_ (.Y(_2476_),
    .A(\z80.tv80s.i_tv80_core.BusReq_s ),
    .B(net1689));
 sg13g2_o21ai_1 _6800_ (.B1(net491),
    .Y(_2477_),
    .A1(net2182),
    .A2(\z80.tv80s.i_tv80_core.BusReq_s ));
 sg13g2_o21ai_1 _6801_ (.B1(net492),
    .Y(_0442_),
    .A1(_1346_),
    .A2(_2476_));
 sg13g2_a21oi_2 _6802_ (.B1(_1303_),
    .Y(_2478_),
    .A2(net1886),
    .A1(net2055));
 sg13g2_nor2_2 _6803_ (.A(_0961_),
    .B(_1164_),
    .Y(_2479_));
 sg13g2_nand3_1 _6804_ (.B(_2478_),
    .C(_2479_),
    .A(_1176_),
    .Y(_2480_));
 sg13g2_or2_1 _6805_ (.X(_2481_),
    .B(_1504_),
    .A(_0964_));
 sg13g2_nor3_2 _6806_ (.A(_0923_),
    .B(_0926_),
    .C(_2481_),
    .Y(_2482_));
 sg13g2_nand2b_2 _6807_ (.Y(_2483_),
    .B(_2482_),
    .A_N(_2480_));
 sg13g2_inv_1 _6808_ (.Y(_2484_),
    .A(_2483_));
 sg13g2_nand2_1 _6809_ (.Y(_2485_),
    .A(_1014_),
    .B(_1149_));
 sg13g2_nand4_1 _6810_ (.B(_1014_),
    .C(_1149_),
    .A(net1947),
    .Y(_2486_),
    .D(_1533_));
 sg13g2_nor4_2 _6811_ (.A(_1715_),
    .B(_2351_),
    .C(_2483_),
    .Y(_2487_),
    .D(_2486_));
 sg13g2_and3_1 _6812_ (.X(_2488_),
    .A(_0677_),
    .B(\z80.tv80s.i_tv80_core.IncDecZ ),
    .C(_2487_));
 sg13g2_nand2b_1 _6813_ (.Y(_2489_),
    .B(net2125),
    .A_N(\z80.tv80s.i_tv80_core.mcycles[1] ));
 sg13g2_nor4_1 _6814_ (.A(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .B(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .C(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .D(_2489_),
    .Y(_2490_));
 sg13g2_a22oi_1 _6815_ (.Y(_2491_),
    .B1(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .B2(net2116),
    .A2(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ));
 sg13g2_a221oi_1 _6816_ (.B2(net2110),
    .C1(_2490_),
    .B1(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .A1(net2107),
    .Y(_2492_),
    .A2(\z80.tv80s.i_tv80_core.mcycles[1] ));
 sg13g2_nand2_1 _6817_ (.Y(_2493_),
    .A(_2491_),
    .B(_2492_));
 sg13g2_nor3_2 _6818_ (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .B(_2488_),
    .C(_2493_),
    .Y(_2494_));
 sg13g2_nor2_1 _6819_ (.A(net2103),
    .B(_2494_),
    .Y(_2495_));
 sg13g2_nor3_1 _6820_ (.A(net625),
    .B(_1131_),
    .C(_1338_),
    .Y(_2496_));
 sg13g2_and2_1 _6821_ (.A(_2495_),
    .B(_2496_),
    .X(_2497_));
 sg13g2_nand2_2 _6822_ (.Y(_2498_),
    .A(_1134_),
    .B(_2497_));
 sg13g2_and2_1 _6823_ (.A(net580),
    .B(_0843_),
    .X(_2499_));
 sg13g2_nor2_1 _6824_ (.A(_2498_),
    .B(_2499_),
    .Y(_2500_));
 sg13g2_a21oi_1 _6825_ (.A1(_0681_),
    .A2(_2498_),
    .Y(_0443_),
    .B1(_2500_));
 sg13g2_nor3_1 _6826_ (.A(net2183),
    .B(net471),
    .C(net1689),
    .Y(_2501_));
 sg13g2_a21o_1 _6827_ (.A2(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .A1(net2183),
    .B1(_2501_),
    .X(_0444_));
 sg13g2_nor2_1 _6828_ (.A(net2228),
    .B(net558),
    .Y(_2502_));
 sg13g2_a21oi_1 _6829_ (.A1(net2228),
    .A2(net4),
    .Y(_0445_),
    .B1(_2502_));
 sg13g2_nor2_1 _6830_ (.A(net2181),
    .B(net3),
    .Y(_2503_));
 sg13g2_a21oi_1 _6831_ (.A1(net225),
    .A2(_2503_),
    .Y(_2504_),
    .B1(\z80.tv80s.i_tv80_core.NMI_s ));
 sg13g2_a21oi_1 _6832_ (.A1(net2228),
    .A2(_0692_),
    .Y(_0446_),
    .B1(net226));
 sg13g2_nor2_1 _6833_ (.A(net2228),
    .B(net430),
    .Y(_2505_));
 sg13g2_a21oi_1 _6834_ (.A1(net2228),
    .A2(net2),
    .Y(_0447_),
    .B1(_2505_));
 sg13g2_a21oi_1 _6835_ (.A1(net2181),
    .A2(_0691_),
    .Y(_0448_),
    .B1(_2503_));
 sg13g2_a21oi_1 _6836_ (.A1(_0023_),
    .A2(net1997),
    .Y(_2506_),
    .B1(_2346_));
 sg13g2_a21o_1 _6837_ (.A2(net2181),
    .A1(net351),
    .B1(_2506_),
    .X(_0449_));
 sg13g2_nor2_1 _6838_ (.A(net1961),
    .B(_1635_),
    .Y(_2507_));
 sg13g2_a22oi_1 _6839_ (.Y(_0450_),
    .B1(_1658_),
    .B2(_2507_),
    .A2(net1961),
    .A1(_0694_));
 sg13g2_mux2_1 _6840_ (.A0(net404),
    .A1(_1657_),
    .S(net1984),
    .X(_0451_));
 sg13g2_nand3_1 _6841_ (.B(_1583_),
    .C(_1610_),
    .A(net1986),
    .Y(_2508_));
 sg13g2_o21ai_1 _6842_ (.B1(_2508_),
    .Y(_2509_),
    .A1(net2163),
    .A2(net1986));
 sg13g2_inv_1 _6843_ (.Y(_0452_),
    .A(_2509_));
 sg13g2_mux2_1 _6844_ (.A0(net515),
    .A1(_1609_),
    .S(net1990),
    .X(_0453_));
 sg13g2_nand3_1 _6845_ (.B(_1518_),
    .C(net1835),
    .A(_1333_),
    .Y(_2510_));
 sg13g2_nand3_1 _6846_ (.B(_1540_),
    .C(_2510_),
    .A(net1990),
    .Y(_2511_));
 sg13g2_o21ai_1 _6847_ (.B1(_2511_),
    .Y(_2512_),
    .A1(net2161),
    .A2(net1988));
 sg13g2_inv_1 _6848_ (.Y(_0454_),
    .A(_2512_));
 sg13g2_nor2_1 _6849_ (.A(net325),
    .B(net1986),
    .Y(_2513_));
 sg13g2_a21oi_1 _6850_ (.A1(net1986),
    .A2(_1887_),
    .Y(_0455_),
    .B1(_2513_));
 sg13g2_mux2_1 _6851_ (.A0(net434),
    .A1(_1881_),
    .S(net1985),
    .X(_0456_));
 sg13g2_nor2_1 _6852_ (.A(net330),
    .B(net1986),
    .Y(_2514_));
 sg13g2_a21oi_1 _6853_ (.A1(net1986),
    .A2(_1897_),
    .Y(_0457_),
    .B1(_2514_));
 sg13g2_nor2_1 _6854_ (.A(net366),
    .B(net1983),
    .Y(_2515_));
 sg13g2_a21oi_1 _6855_ (.A1(net1983),
    .A2(_1867_),
    .Y(_0458_),
    .B1(_2515_));
 sg13g2_nor2_1 _6856_ (.A(net362),
    .B(net1983),
    .Y(_2516_));
 sg13g2_a21oi_1 _6857_ (.A1(net1983),
    .A2(_1935_),
    .Y(_0459_),
    .B1(_2516_));
 sg13g2_nor2_1 _6858_ (.A(net354),
    .B(net1983),
    .Y(_2517_));
 sg13g2_a21oi_1 _6859_ (.A1(net1983),
    .A2(_1928_),
    .Y(_0460_),
    .B1(_2517_));
 sg13g2_nor2_1 _6860_ (.A(net421),
    .B(net1985),
    .Y(_2518_));
 sg13g2_a21oi_1 _6861_ (.A1(net1983),
    .A2(_1919_),
    .Y(_0461_),
    .B1(_2518_));
 sg13g2_nor2_1 _6862_ (.A(net444),
    .B(net1987),
    .Y(_2519_));
 sg13g2_a21oi_1 _6863_ (.A1(net1983),
    .A2(_1910_),
    .Y(_0462_),
    .B1(_2519_));
 sg13g2_nor2_1 _6864_ (.A(net357),
    .B(net1989),
    .Y(_2520_));
 sg13g2_a21oi_1 _6865_ (.A1(net1988),
    .A2(_1950_),
    .Y(_0463_),
    .B1(_2520_));
 sg13g2_nor2_1 _6866_ (.A(net369),
    .B(net1987),
    .Y(_2521_));
 sg13g2_a21oi_1 _6867_ (.A1(net1986),
    .A2(_2012_),
    .Y(_0464_),
    .B1(_2521_));
 sg13g2_nor2_1 _6868_ (.A(net396),
    .B(net1989),
    .Y(_2522_));
 sg13g2_a21oi_1 _6869_ (.A1(net1989),
    .A2(_2056_),
    .Y(_0465_),
    .B1(_2522_));
 sg13g2_nor2_1 _6870_ (.A(net399),
    .B(net1989),
    .Y(_2523_));
 sg13g2_a21oi_1 _6871_ (.A1(net1988),
    .A2(_2107_),
    .Y(_0466_),
    .B1(_2523_));
 sg13g2_nor2_1 _6872_ (.A(net347),
    .B(net1988),
    .Y(_2524_));
 sg13g2_a21oi_1 _6873_ (.A1(net1988),
    .A2(_2159_),
    .Y(_0467_),
    .B1(_2524_));
 sg13g2_nor2_1 _6874_ (.A(net318),
    .B(net1987),
    .Y(_2525_));
 sg13g2_a21oi_1 _6875_ (.A1(net1986),
    .A2(_2227_),
    .Y(_0468_),
    .B1(_2525_));
 sg13g2_nor2_1 _6876_ (.A(net328),
    .B(net1988),
    .Y(_2526_));
 sg13g2_a21oi_1 _6877_ (.A1(net1988),
    .A2(_2278_),
    .Y(_0469_),
    .B1(_2526_));
 sg13g2_nor2_1 _6878_ (.A(net303),
    .B(net1987),
    .Y(_2527_));
 sg13g2_a21oi_1 _6879_ (.A1(net1987),
    .A2(_2331_),
    .Y(_0470_),
    .B1(_2527_));
 sg13g2_nand2_1 _6880_ (.Y(_2528_),
    .A(net2033),
    .B(_2487_));
 sg13g2_and3_1 _6881_ (.X(_2529_),
    .A(_1700_),
    .B(net1824),
    .C(_1728_));
 sg13g2_nand3_1 _6882_ (.B(net1824),
    .C(_1728_),
    .A(_1700_),
    .Y(_2530_));
 sg13g2_a21oi_1 _6883_ (.A1(_2528_),
    .A2(_2530_),
    .Y(_2531_),
    .B1(net1970));
 sg13g2_nand2b_1 _6884_ (.Y(_2532_),
    .B(net494),
    .A_N(_2531_));
 sg13g2_and3_2 _6885_ (.X(_2533_),
    .A(net2034),
    .B(net2038),
    .C(_1778_));
 sg13g2_nand3_1 _6886_ (.B(net2038),
    .C(_1778_),
    .A(net2035),
    .Y(_2534_));
 sg13g2_nand2_1 _6887_ (.Y(_2535_),
    .A(_2032_),
    .B(_2081_));
 sg13g2_nand2_1 _6888_ (.Y(_2536_),
    .A(_0662_),
    .B(\z80.tv80s.i_tv80_core.Z16_r ));
 sg13g2_nand3_1 _6889_ (.B(_1984_),
    .C(_2536_),
    .A(_1803_),
    .Y(_2537_));
 sg13g2_nand4_1 _6890_ (.B(_2184_),
    .C(_2250_),
    .A(_2131_),
    .Y(_2538_),
    .D(_2298_));
 sg13g2_nor3_1 _6891_ (.A(_2535_),
    .B(_2537_),
    .C(_2538_),
    .Y(_2539_));
 sg13g2_a21oi_1 _6892_ (.A1(_0662_),
    .A2(\z80.tv80s.i_tv80_core.Arith16_r ),
    .Y(_2540_),
    .B1(net2035));
 sg13g2_o21ai_1 _6893_ (.B1(_2540_),
    .Y(_2541_),
    .A1(\z80.tv80s.i_tv80_core.Arith16_r ),
    .A2(_2539_));
 sg13g2_nand2_1 _6894_ (.Y(_2542_),
    .A(_1807_),
    .B(_1995_));
 sg13g2_o21ai_1 _6895_ (.B1(_1812_),
    .Y(_2543_),
    .A1(_0219_),
    .A2(_1035_));
 sg13g2_o21ai_1 _6896_ (.B1(_2139_),
    .Y(_2544_),
    .A1(_0222_),
    .A2(_1044_));
 sg13g2_or4_1 _6897_ (.A(_1814_),
    .B(_1993_),
    .C(_2094_),
    .D(_2261_),
    .X(_2545_));
 sg13g2_nor4_1 _6898_ (.A(_2309_),
    .B(_2543_),
    .C(_2544_),
    .D(_2545_),
    .Y(_2546_));
 sg13g2_nor2_1 _6899_ (.A(_2533_),
    .B(_2546_),
    .Y(_2547_));
 sg13g2_nor4_1 _6900_ (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .B(\z80.tv80s.i_tv80_core.BusA[4] ),
    .C(net2029),
    .D(net2031),
    .Y(_2548_));
 sg13g2_and4_1 _6901_ (.A(_1810_),
    .B(_1994_),
    .C(_2040_),
    .D(_2090_),
    .X(_2549_));
 sg13g2_nand3_1 _6902_ (.B(_2548_),
    .C(_2549_),
    .A(_1808_),
    .Y(_2550_));
 sg13g2_nand4_1 _6903_ (.B(_2088_),
    .C(_2141_),
    .A(_2043_),
    .Y(_2551_),
    .D(_2214_));
 sg13g2_nor4_1 _6904_ (.A(_2264_),
    .B(_2317_),
    .C(_2542_),
    .D(_2551_),
    .Y(_2552_));
 sg13g2_a21oi_1 _6905_ (.A1(_0662_),
    .A2(net2172),
    .Y(_2553_),
    .B1(_1804_));
 sg13g2_o21ai_1 _6906_ (.B1(_2553_),
    .Y(_2554_),
    .A1(net2172),
    .A2(_2552_));
 sg13g2_nand3_1 _6907_ (.B(_2550_),
    .C(_2554_),
    .A(_2547_),
    .Y(_2555_));
 sg13g2_and3_1 _6908_ (.X(_2556_),
    .A(_2257_),
    .B(_2300_),
    .C(_2305_));
 sg13g2_nand3_1 _6909_ (.B(_2037_),
    .C(_2087_),
    .A(_0212_),
    .Y(_2557_));
 sg13g2_nand2b_1 _6910_ (.Y(_2558_),
    .B(_2135_),
    .A_N(_2209_));
 sg13g2_nor4_1 _6911_ (.A(_1817_),
    .B(_1989_),
    .C(_2557_),
    .D(_2558_),
    .Y(_2559_));
 sg13g2_a21oi_1 _6912_ (.A1(_2556_),
    .A2(_2559_),
    .Y(_2560_),
    .B1(_2555_));
 sg13g2_a22oi_1 _6913_ (.Y(_2561_),
    .B1(_2541_),
    .B2(_2560_),
    .A2(_2533_),
    .A1(_0662_));
 sg13g2_o21ai_1 _6914_ (.B1(_2531_),
    .Y(_2562_),
    .A1(_2529_),
    .A2(_2561_));
 sg13g2_nor4_1 _6915_ (.A(_1890_),
    .B(_1900_),
    .C(_2416_),
    .D(_2530_),
    .Y(_2563_));
 sg13g2_nand4_1 _6916_ (.B(_2426_),
    .C(_2432_),
    .A(_1954_),
    .Y(_2564_),
    .D(_2563_));
 sg13g2_or4_1 _6917_ (.A(_2015_),
    .B(_2164_),
    .C(_2448_),
    .D(_2564_),
    .X(_2565_));
 sg13g2_or4_1 _6918_ (.A(_2063_),
    .B(_2232_),
    .C(_2453_),
    .D(_2565_),
    .X(_2566_));
 sg13g2_nor4_2 _6919_ (.A(_2110_),
    .B(_2283_),
    .C(_2333_),
    .Y(_2567_),
    .D(_2566_));
 sg13g2_o21ai_1 _6920_ (.B1(_2532_),
    .Y(_0471_),
    .A1(_2562_),
    .A2(_2567_));
 sg13g2_or2_2 _6921_ (.X(_2568_),
    .B(_1774_),
    .A(_1137_));
 sg13g2_nor2_1 _6922_ (.A(_1345_),
    .B(_2568_),
    .Y(_2569_));
 sg13g2_nand2b_1 _6923_ (.Y(_2570_),
    .B(_1064_),
    .A_N(net467));
 sg13g2_a21oi_1 _6924_ (.A1(net1689),
    .A2(_2569_),
    .Y(_2571_),
    .B1(net2183));
 sg13g2_a22oi_1 _6925_ (.Y(_0472_),
    .B1(_2570_),
    .B2(_2571_),
    .A2(_0693_),
    .A1(net2183));
 sg13g2_nand2_2 _6926_ (.Y(_2572_),
    .A(_1188_),
    .B(_1685_));
 sg13g2_nor3_1 _6927_ (.A(_0971_),
    .B(_1019_),
    .C(_2485_),
    .Y(_2573_));
 sg13g2_nand4_1 _6928_ (.B(_1175_),
    .C(_1493_),
    .A(_1004_),
    .Y(_2574_),
    .D(_2573_));
 sg13g2_nor4_1 _6929_ (.A(_1242_),
    .B(_1251_),
    .C(_1502_),
    .D(_2574_),
    .Y(_2575_));
 sg13g2_nand2_1 _6930_ (.Y(_2576_),
    .A(_2349_),
    .B(_2575_));
 sg13g2_nor2_2 _6931_ (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(_0028_),
    .Y(_2577_));
 sg13g2_a21oi_1 _6932_ (.A1(_1834_),
    .A2(_2577_),
    .Y(_2578_),
    .B1(_2576_));
 sg13g2_nand3b_1 _6933_ (.B(_0684_),
    .C(_1057_),
    .Y(_2579_),
    .A_N(net2118));
 sg13g2_inv_1 _6934_ (.Y(_2580_),
    .A(_2579_));
 sg13g2_a22oi_1 _6935_ (.Y(_2581_),
    .B1(_0970_),
    .B2(_2580_),
    .A2(_0968_),
    .A1(_0684_));
 sg13g2_nand2_1 _6936_ (.Y(_2582_),
    .A(_2576_),
    .B(_2581_));
 sg13g2_a22oi_1 _6937_ (.Y(_2583_),
    .B1(_2582_),
    .B2(net2170),
    .A2(_2358_),
    .A1(_1677_));
 sg13g2_o21ai_1 _6938_ (.B1(_2572_),
    .Y(_2584_),
    .A1(_2578_),
    .A2(_2583_));
 sg13g2_and2_1 _6939_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(net1725),
    .X(_2585_));
 sg13g2_a21oi_1 _6940_ (.A1(_0737_),
    .A2(net2155),
    .Y(_2586_),
    .B1(net2177));
 sg13g2_o21ai_1 _6941_ (.B1(_2586_),
    .Y(_2587_),
    .A1(_0155_),
    .A2(net2155));
 sg13g2_o21ai_1 _6942_ (.B1(net2177),
    .Y(_2588_),
    .A1(_0157_),
    .A2(net2155));
 sg13g2_a21oi_1 _6943_ (.A1(_0738_),
    .A2(net2156),
    .Y(_2589_),
    .B1(_2588_));
 sg13g2_nor2_1 _6944_ (.A(net2007),
    .B(_2589_),
    .Y(_2590_));
 sg13g2_mux4_1 _6945_ (.S0(net2180),
    .A0(_0151_),
    .A1(_0153_),
    .A2(_0152_),
    .A3(_0154_),
    .S1(net2155),
    .X(_2591_));
 sg13g2_nor2_1 _6946_ (.A(net2174),
    .B(_2591_),
    .Y(_2592_));
 sg13g2_a21oi_2 _6947_ (.B1(_2592_),
    .Y(_2593_),
    .A2(_2590_),
    .A1(_2587_));
 sg13g2_or2_1 _6948_ (.X(_2594_),
    .B(_2593_),
    .A(net1840));
 sg13g2_nand4_1 _6949_ (.B(_1263_),
    .C(_1422_),
    .A(net2170),
    .Y(_2595_),
    .D(_1500_));
 sg13g2_or4_1 _6950_ (.A(_1242_),
    .B(_1519_),
    .C(_1521_),
    .D(_2595_),
    .X(_2596_));
 sg13g2_nand2_1 _6951_ (.Y(_2597_),
    .A(net2170),
    .B(_1162_));
 sg13g2_nand3_1 _6952_ (.B(_1169_),
    .C(_1241_),
    .A(_1147_),
    .Y(_2598_));
 sg13g2_nor3_1 _6953_ (.A(_0971_),
    .B(_1253_),
    .C(_2485_),
    .Y(_2599_));
 sg13g2_nand3_1 _6954_ (.B(_2484_),
    .C(_2599_),
    .A(_1714_),
    .Y(_2600_));
 sg13g2_or4_2 _6955_ (.A(_1833_),
    .B(_2597_),
    .C(_2598_),
    .D(_2600_),
    .X(_2601_));
 sg13g2_nand2_1 _6956_ (.Y(_2602_),
    .A(_2596_),
    .B(_2601_));
 sg13g2_and2_1 _6957_ (.A(net2136),
    .B(net1783),
    .X(_2603_));
 sg13g2_nand2_2 _6958_ (.Y(_2604_),
    .A(\z80.tv80s.i_tv80_core.IntCycle ),
    .B(\z80.tv80s.i_tv80_core.IStatus[1] ));
 sg13g2_nor2_2 _6959_ (.A(net2014),
    .B(_2604_),
    .Y(_2605_));
 sg13g2_nand3_1 _6960_ (.B(\z80.tv80s.i_tv80_core.IntCycle ),
    .C(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .A(net2110),
    .Y(_2606_));
 sg13g2_and2_1 _6961_ (.A(_1321_),
    .B(_1333_),
    .X(_2607_));
 sg13g2_inv_2 _6962_ (.Y(_2608_),
    .A(net1712));
 sg13g2_nor2_1 _6963_ (.A(_0194_),
    .B(_2608_),
    .Y(_2609_));
 sg13g2_nor2_1 _6964_ (.A(_1288_),
    .B(_1321_),
    .Y(_2610_));
 sg13g2_nor3_1 _6965_ (.A(_1288_),
    .B(_1321_),
    .C(_2593_),
    .Y(_2611_));
 sg13g2_nand2b_1 _6966_ (.Y(_2612_),
    .B(_1287_),
    .A_N(_1321_));
 sg13g2_nor2_2 _6967_ (.A(_1332_),
    .B(_2612_),
    .Y(_2613_));
 sg13g2_nor2b_1 _6968_ (.A(_2612_),
    .B_N(_1332_),
    .Y(_2614_));
 sg13g2_and3_1 _6969_ (.X(_2615_),
    .A(_1288_),
    .B(_1321_),
    .C(_1334_));
 sg13g2_nand2_1 _6970_ (.Y(_2616_),
    .A(_1177_),
    .B(_1510_));
 sg13g2_nor4_1 _6971_ (.A(_0923_),
    .B(_1301_),
    .C(_1665_),
    .D(_2616_),
    .Y(_2617_));
 sg13g2_and4_1 _6972_ (.A(net2170),
    .B(_1162_),
    .C(_1495_),
    .D(_2617_),
    .X(_2618_));
 sg13g2_o21ai_1 _6973_ (.B1(_0873_),
    .Y(_2619_),
    .A1(_1277_),
    .A2(_2618_));
 sg13g2_xnor2_1 _6974_ (.Y(_2620_),
    .A(net2136),
    .B(net1763));
 sg13g2_and2_1 _6975_ (.A(net1700),
    .B(_2620_),
    .X(_2621_));
 sg13g2_nand2b_1 _6976_ (.Y(_2622_),
    .B(net2053),
    .A_N(_0193_));
 sg13g2_a21oi_1 _6977_ (.A1(net2012),
    .A2(_0770_),
    .Y(_2623_),
    .B1(net1926));
 sg13g2_a221oi_1 _6978_ (.B2(_2623_),
    .C1(net1702),
    .B1(_2622_),
    .A1(net1926),
    .Y(_2624_),
    .A2(_2593_));
 sg13g2_a221oi_1 _6979_ (.B2(\z80.tv80s.i_tv80_core.SP[0] ),
    .C1(_2621_),
    .B1(net1705),
    .A1(\z80.tv80s.di_reg[0] ),
    .Y(_2625_),
    .A2(net1707));
 sg13g2_nor4_1 _6980_ (.A(net1872),
    .B(_2609_),
    .C(_2611_),
    .D(_2624_),
    .Y(_2626_));
 sg13g2_a21oi_2 _6981_ (.B1(_0681_),
    .Y(_2627_),
    .A2(_2492_),
    .A1(_2491_));
 sg13g2_or2_1 _6982_ (.X(_2628_),
    .B(_2627_),
    .A(net1783));
 sg13g2_a221oi_1 _6983_ (.B2(_2626_),
    .C1(net1758),
    .B1(_2625_),
    .A1(_0193_),
    .Y(_2629_),
    .A2(net1872));
 sg13g2_o21ai_1 _6984_ (.B1(net1841),
    .Y(_2630_),
    .A1(_2603_),
    .A2(_2629_));
 sg13g2_a21oi_1 _6985_ (.A1(_2594_),
    .A2(_2630_),
    .Y(_2631_),
    .B1(net1724));
 sg13g2_o21ai_1 _6986_ (.B1(net1903),
    .Y(_2632_),
    .A1(_2585_),
    .A2(_2631_));
 sg13g2_nand2_2 _6987_ (.Y(_2633_),
    .A(net1993),
    .B(net1688));
 sg13g2_nand2b_1 _6988_ (.Y(_2634_),
    .B(net1694),
    .A_N(_0825_));
 sg13g2_and2_1 _6989_ (.A(_0835_),
    .B(net1686),
    .X(_2635_));
 sg13g2_nand2_1 _6990_ (.Y(_2636_),
    .A(_0835_),
    .B(net1686));
 sg13g2_a21oi_1 _6991_ (.A1(\z80.tv80s.i_tv80_core.R[0] ),
    .A2(net1907),
    .Y(_2637_),
    .B1(net1685));
 sg13g2_a22oi_1 _6992_ (.Y(_0473_),
    .B1(_2637_),
    .B2(_2632_),
    .A2(net1685),
    .A1(_0752_));
 sg13g2_nand2_1 _6993_ (.Y(_2638_),
    .A(net244),
    .B(net1685));
 sg13g2_a21oi_1 _6994_ (.A1(net2135),
    .A2(net1872),
    .Y(_2639_),
    .B1(_2627_));
 sg13g2_nand2_2 _6995_ (.Y(_2640_),
    .A(net2135),
    .B(net2136));
 sg13g2_or2_1 _6996_ (.X(_2641_),
    .B(net2136),
    .A(net2135));
 sg13g2_a21oi_1 _6997_ (.A1(_2640_),
    .A2(_2641_),
    .Y(_2642_),
    .B1(net1762));
 sg13g2_a21oi_1 _6998_ (.A1(_0195_),
    .A2(net1762),
    .Y(_2643_),
    .B1(_2642_));
 sg13g2_mux2_1 _6999_ (.A0(_0163_),
    .A1(_0164_),
    .S(net2154),
    .X(_2644_));
 sg13g2_nand2_1 _7000_ (.Y(_2645_),
    .A(net2008),
    .B(_2644_));
 sg13g2_mux2_1 _7001_ (.A0(_0165_),
    .A1(_0166_),
    .S(net2154),
    .X(_2646_));
 sg13g2_a21oi_1 _7002_ (.A1(net2176),
    .A2(_2646_),
    .Y(_2647_),
    .B1(net2007));
 sg13g2_mux4_1 _7003_ (.S0(net2176),
    .A0(_0159_),
    .A1(_0161_),
    .A2(_0160_),
    .A3(_0162_),
    .S1(net2154),
    .X(_2648_));
 sg13g2_nor2_1 _7004_ (.A(net2174),
    .B(_2648_),
    .Y(_2649_));
 sg13g2_a21oi_2 _7005_ (.B1(_2649_),
    .Y(_2650_),
    .A2(_2647_),
    .A1(_2645_));
 sg13g2_inv_1 _7006_ (.Y(_2651_),
    .A(_2650_));
 sg13g2_a221oi_1 _7007_ (.B2(net1709),
    .C1(net1712),
    .B1(_2651_),
    .A1(_2615_),
    .Y(_2652_),
    .A2(_2643_));
 sg13g2_nand2b_1 _7008_ (.Y(_2653_),
    .B(net2053),
    .A_N(_0195_));
 sg13g2_a21oi_1 _7009_ (.A1(net2011),
    .A2(_0771_),
    .Y(_2654_),
    .B1(net1926));
 sg13g2_a221oi_1 _7010_ (.B2(_2654_),
    .C1(net1702),
    .B1(_2653_),
    .A1(net1927),
    .Y(_2655_),
    .A2(_2650_));
 sg13g2_a221oi_1 _7011_ (.B2(\z80.tv80s.i_tv80_core.SP[1] ),
    .C1(_2655_),
    .B1(net1705),
    .A1(\z80.tv80s.di_reg[1] ),
    .Y(_2656_),
    .A2(net1707));
 sg13g2_a22oi_1 _7012_ (.Y(_2657_),
    .B1(_2652_),
    .B2(_2656_),
    .A2(net1712),
    .A1(_0741_));
 sg13g2_nand2_1 _7013_ (.Y(_2658_),
    .A(net1920),
    .B(_2657_));
 sg13g2_a21oi_1 _7014_ (.A1(_2639_),
    .A2(_2658_),
    .Y(_2659_),
    .B1(net1783));
 sg13g2_a21oi_1 _7015_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .A2(net1782),
    .Y(_2660_),
    .B1(_2659_));
 sg13g2_mux2_1 _7016_ (.A0(_2650_),
    .A1(_2660_),
    .S(net1841),
    .X(_2661_));
 sg13g2_a21oi_1 _7017_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .A2(net1724),
    .Y(_2662_),
    .B1(net1913));
 sg13g2_o21ai_1 _7018_ (.B1(_2662_),
    .Y(_2663_),
    .A1(net1724),
    .A2(_2661_));
 sg13g2_o21ai_1 _7019_ (.B1(_2663_),
    .Y(_2664_),
    .A1(\z80.tv80s.i_tv80_core.R[1] ),
    .A2(net1899));
 sg13g2_o21ai_1 _7020_ (.B1(_2638_),
    .Y(_0474_),
    .A1(net1684),
    .A2(_2664_));
 sg13g2_a21oi_1 _7021_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .A2(net1867),
    .Y(_2665_),
    .B1(_2627_));
 sg13g2_nand2b_1 _7022_ (.Y(_2666_),
    .B(net2156),
    .A_N(_0066_));
 sg13g2_o21ai_1 _7023_ (.B1(_2666_),
    .Y(_2667_),
    .A1(_0065_),
    .A2(net2155));
 sg13g2_nor2_1 _7024_ (.A(_0067_),
    .B(net2155),
    .Y(_2668_));
 sg13g2_a21oi_1 _7025_ (.A1(_0703_),
    .A2(net2155),
    .Y(_2669_),
    .B1(_2668_));
 sg13g2_a21oi_1 _7026_ (.A1(net2177),
    .A2(_2669_),
    .Y(_2670_),
    .B1(net2007));
 sg13g2_o21ai_1 _7027_ (.B1(_2670_),
    .Y(_2671_),
    .A1(net2177),
    .A2(_2667_));
 sg13g2_mux4_1 _7028_ (.S0(net2177),
    .A0(_0061_),
    .A1(_0063_),
    .A2(_0062_),
    .A3(_0064_),
    .S1(net2155),
    .X(_2672_));
 sg13g2_o21ai_1 _7029_ (.B1(_2671_),
    .Y(_2673_),
    .A1(net2174),
    .A2(_2672_));
 sg13g2_nand2_1 _7030_ (.Y(_2674_),
    .A(net2054),
    .B(_0197_));
 sg13g2_a21oi_2 _7031_ (.B1(net1926),
    .Y(_2675_),
    .A2(_0198_),
    .A1(net2012));
 sg13g2_a22oi_1 _7032_ (.Y(_2676_),
    .B1(_2674_),
    .B2(_2675_),
    .A2(_2673_),
    .A1(net1923));
 sg13g2_nor2_1 _7033_ (.A(net1701),
    .B(_2676_),
    .Y(_2677_));
 sg13g2_nor2_1 _7034_ (.A(net1762),
    .B(_2640_),
    .Y(_2678_));
 sg13g2_nor3_1 _7035_ (.A(_0197_),
    .B(net1762),
    .C(_2640_),
    .Y(_2679_));
 sg13g2_xnor2_1 _7036_ (.Y(_2680_),
    .A(_0197_),
    .B(_2678_));
 sg13g2_a22oi_1 _7037_ (.Y(_2681_),
    .B1(_2673_),
    .B2(net1708),
    .A2(net1706),
    .A1(\z80.tv80s.di_reg[2] ));
 sg13g2_a221oi_1 _7038_ (.B2(_2680_),
    .C1(_2677_),
    .B1(net1699),
    .A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .Y(_2682_),
    .A2(net1704));
 sg13g2_nand3_1 _7039_ (.B(_2681_),
    .C(_2682_),
    .A(_2608_),
    .Y(_2683_));
 sg13g2_o21ai_1 _7040_ (.B1(_2683_),
    .Y(_2684_),
    .A1(\z80.tv80s.i_tv80_core.PC[2] ),
    .A2(_2608_));
 sg13g2_o21ai_1 _7041_ (.B1(_2665_),
    .Y(_2685_),
    .A1(net1868),
    .A2(_2684_));
 sg13g2_mux2_1 _7042_ (.A0(_2685_),
    .A1(net2134),
    .S(net1781),
    .X(_2686_));
 sg13g2_nor2b_1 _7043_ (.A(net1839),
    .B_N(_2673_),
    .Y(_2687_));
 sg13g2_a21oi_1 _7044_ (.A1(net1839),
    .A2(_2686_),
    .Y(_2688_),
    .B1(_2687_));
 sg13g2_a21oi_1 _7045_ (.A1(net2134),
    .A2(net1720),
    .Y(_2689_),
    .B1(net1909));
 sg13g2_o21ai_1 _7046_ (.B1(_2689_),
    .Y(_2690_),
    .A1(net1720),
    .A2(_2688_));
 sg13g2_o21ai_1 _7047_ (.B1(_2690_),
    .Y(_2691_),
    .A1(\z80.tv80s.i_tv80_core.R[2] ),
    .A2(net1896));
 sg13g2_nor2_1 _7048_ (.A(net375),
    .B(net1681),
    .Y(_2692_));
 sg13g2_a21oi_1 _7049_ (.A1(net1681),
    .A2(_2691_),
    .Y(_0475_),
    .B1(_2692_));
 sg13g2_a21oi_1 _7050_ (.A1(_0708_),
    .A2(net2153),
    .Y(_2693_),
    .B1(net2175));
 sg13g2_o21ai_1 _7051_ (.B1(_2693_),
    .Y(_2694_),
    .A1(_0081_),
    .A2(net2153));
 sg13g2_o21ai_1 _7052_ (.B1(net2175),
    .Y(_2695_),
    .A1(_0083_),
    .A2(net2153));
 sg13g2_a21oi_1 _7053_ (.A1(_0709_),
    .A2(net2153),
    .Y(_2696_),
    .B1(_2695_));
 sg13g2_nor2_1 _7054_ (.A(net2007),
    .B(_2696_),
    .Y(_2697_));
 sg13g2_mux4_1 _7055_ (.S0(net2175),
    .A0(_0077_),
    .A1(_0079_),
    .A2(_0078_),
    .A3(_0080_),
    .S1(net2153),
    .X(_2698_));
 sg13g2_nor2_1 _7056_ (.A(net2174),
    .B(_2698_),
    .Y(_2699_));
 sg13g2_a21oi_2 _7057_ (.B1(_2699_),
    .Y(_2700_),
    .A2(_2697_),
    .A1(_2694_));
 sg13g2_inv_1 _7058_ (.Y(_2701_),
    .A(_2700_));
 sg13g2_nor2_1 _7059_ (.A(net1838),
    .B(_2700_),
    .Y(_2702_));
 sg13g2_nand2_1 _7060_ (.Y(_2703_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .B(net1781));
 sg13g2_nand2b_1 _7061_ (.Y(_2704_),
    .B(net2052),
    .A_N(_0199_));
 sg13g2_a21oi_1 _7062_ (.A1(net2013),
    .A2(_0773_),
    .Y(_2705_),
    .B1(net1923));
 sg13g2_a221oi_1 _7063_ (.B2(_2705_),
    .C1(net1702),
    .B1(_2704_),
    .A1(net1923),
    .Y(_2706_),
    .A2(_2700_));
 sg13g2_xnor2_1 _7064_ (.Y(_2707_),
    .A(_0199_),
    .B(_2679_));
 sg13g2_a221oi_1 _7065_ (.B2(net1708),
    .C1(net1713),
    .B1(_2701_),
    .A1(\z80.tv80s.di_reg[3] ),
    .Y(_2708_),
    .A2(net1707));
 sg13g2_a221oi_1 _7066_ (.B2(_2707_),
    .C1(_2706_),
    .B1(net1699),
    .A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .Y(_2709_),
    .A2(net1705));
 sg13g2_a22oi_1 _7067_ (.Y(_2710_),
    .B1(_2708_),
    .B2(_2709_),
    .A2(net1713),
    .A1(_0200_));
 sg13g2_a21oi_1 _7068_ (.A1(_0199_),
    .A2(net1867),
    .Y(_2711_),
    .B1(net1756));
 sg13g2_o21ai_1 _7069_ (.B1(_2711_),
    .Y(_2712_),
    .A1(net1867),
    .A2(_2710_));
 sg13g2_nand2_1 _7070_ (.Y(_2713_),
    .A(_2703_),
    .B(_2712_));
 sg13g2_a21oi_1 _7071_ (.A1(net1838),
    .A2(_2713_),
    .Y(_2714_),
    .B1(_2702_));
 sg13g2_a21oi_1 _7072_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net1719),
    .Y(_2715_),
    .B1(net1909));
 sg13g2_o21ai_1 _7073_ (.B1(_2715_),
    .Y(_2716_),
    .A1(net1719),
    .A2(_2714_));
 sg13g2_o21ai_1 _7074_ (.B1(_2716_),
    .Y(_2717_),
    .A1(\z80.tv80s.i_tv80_core.R[3] ),
    .A2(net1895));
 sg13g2_nor2_1 _7075_ (.A(net377),
    .B(net1681),
    .Y(_2718_));
 sg13g2_a21oi_1 _7076_ (.A1(net1681),
    .A2(_2717_),
    .Y(_0476_),
    .B1(_2718_));
 sg13g2_and2_1 _7077_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .B(net1781),
    .X(_2719_));
 sg13g2_nand2b_1 _7078_ (.Y(_2720_),
    .B(net2152),
    .A_N(_0098_));
 sg13g2_o21ai_1 _7079_ (.B1(_2720_),
    .Y(_2721_),
    .A1(_0097_),
    .A2(net2152));
 sg13g2_o21ai_1 _7080_ (.B1(net2175),
    .Y(_2722_),
    .A1(_0099_),
    .A2(net2152));
 sg13g2_a21oi_1 _7081_ (.A1(_0713_),
    .A2(net2152),
    .Y(_2723_),
    .B1(_2722_));
 sg13g2_nor2_1 _7082_ (.A(net2007),
    .B(_2723_),
    .Y(_2724_));
 sg13g2_o21ai_1 _7083_ (.B1(_2724_),
    .Y(_2725_),
    .A1(net2175),
    .A2(_2721_));
 sg13g2_mux4_1 _7084_ (.S0(net2175),
    .A0(_0093_),
    .A1(_0095_),
    .A2(_0094_),
    .A3(_0096_),
    .S1(net2152),
    .X(_2726_));
 sg13g2_o21ai_1 _7085_ (.B1(_2725_),
    .Y(_2727_),
    .A1(net2174),
    .A2(_2726_));
 sg13g2_o21ai_1 _7086_ (.B1(net1921),
    .Y(_2728_),
    .A1(_0202_),
    .A2(_2608_));
 sg13g2_nand3_1 _7087_ (.B(net2134),
    .C(_2678_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .Y(_2729_));
 sg13g2_nor2_1 _7088_ (.A(_0201_),
    .B(_2729_),
    .Y(_2730_));
 sg13g2_xor2_1 _7089_ (.B(_2729_),
    .A(_0201_),
    .X(_2731_));
 sg13g2_nand2_1 _7090_ (.Y(_2732_),
    .A(net2054),
    .B(_0201_));
 sg13g2_a21oi_1 _7091_ (.A1(net2013),
    .A2(_0202_),
    .Y(_2733_),
    .B1(net1923));
 sg13g2_a22oi_1 _7092_ (.Y(_2734_),
    .B1(_2732_),
    .B2(_2733_),
    .A2(_2727_),
    .A1(net1923));
 sg13g2_nor2_1 _7093_ (.A(net1701),
    .B(_2734_),
    .Y(_2735_));
 sg13g2_a221oi_1 _7094_ (.B2(_2731_),
    .C1(_2735_),
    .B1(net1699),
    .A1(net2047),
    .Y(_2736_),
    .A2(net1707));
 sg13g2_a221oi_1 _7095_ (.B2(net1708),
    .C1(_2728_),
    .B1(_2727_),
    .A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .Y(_2737_),
    .A2(net1704));
 sg13g2_a221oi_1 _7096_ (.B2(_2737_),
    .C1(net1759),
    .B1(_2736_),
    .A1(_0201_),
    .Y(_2738_),
    .A2(net1867));
 sg13g2_o21ai_1 _7097_ (.B1(net1838),
    .Y(_2739_),
    .A1(_2719_),
    .A2(_2738_));
 sg13g2_nand2b_1 _7098_ (.Y(_2740_),
    .B(_2727_),
    .A_N(net1838));
 sg13g2_a21oi_1 _7099_ (.A1(_2739_),
    .A2(_2740_),
    .Y(_2741_),
    .B1(net1727));
 sg13g2_a21oi_2 _7100_ (.B1(_2741_),
    .Y(_2742_),
    .A2(net1720),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sg13g2_o21ai_1 _7101_ (.B1(net1683),
    .Y(_2743_),
    .A1(\z80.tv80s.i_tv80_core.R[4] ),
    .A2(net1895));
 sg13g2_a21oi_2 _7102_ (.B1(_2743_),
    .Y(_2744_),
    .A2(_2742_),
    .A1(net1895));
 sg13g2_a21o_1 _7103_ (.A2(net1685),
    .A1(net453),
    .B1(_2744_),
    .X(_0477_));
 sg13g2_a21oi_1 _7104_ (.A1(_0715_),
    .A2(net2153),
    .Y(_2745_),
    .B1(net2176));
 sg13g2_o21ai_1 _7105_ (.B1(_2745_),
    .Y(_2746_),
    .A1(_0113_),
    .A2(net2152));
 sg13g2_o21ai_1 _7106_ (.B1(net2175),
    .Y(_2747_),
    .A1(_0115_),
    .A2(net2152));
 sg13g2_a21oi_1 _7107_ (.A1(_0716_),
    .A2(net2152),
    .Y(_2748_),
    .B1(_2747_));
 sg13g2_nor2_1 _7108_ (.A(net2007),
    .B(_2748_),
    .Y(_2749_));
 sg13g2_mux4_1 _7109_ (.S0(net2175),
    .A0(_0109_),
    .A1(_0111_),
    .A2(_0110_),
    .A3(_0112_),
    .S1(net2153),
    .X(_2750_));
 sg13g2_nor2_1 _7110_ (.A(net2174),
    .B(_2750_),
    .Y(_2751_));
 sg13g2_a21oi_2 _7111_ (.B1(_2751_),
    .Y(_2752_),
    .A2(_2749_),
    .A1(_2746_));
 sg13g2_inv_1 _7112_ (.Y(_2753_),
    .A(_2752_));
 sg13g2_nor2_1 _7113_ (.A(net1839),
    .B(_2752_),
    .Y(_2754_));
 sg13g2_a21oi_1 _7114_ (.A1(net2133),
    .A2(net1868),
    .Y(_2755_),
    .B1(_2627_));
 sg13g2_a22oi_1 _7115_ (.Y(_2756_),
    .B1(_2753_),
    .B2(net1709),
    .A2(net1704),
    .A1(\z80.tv80s.i_tv80_core.SP[5] ));
 sg13g2_nand2_1 _7116_ (.Y(_2757_),
    .A(net2013),
    .B(\z80.tv80s.i_tv80_core.PC[5] ));
 sg13g2_a21oi_1 _7117_ (.A1(net2054),
    .A2(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .Y(_2758_),
    .B1(net1923));
 sg13g2_a221oi_1 _7118_ (.B2(_2758_),
    .C1(net1701),
    .B1(_2757_),
    .A1(net1923),
    .Y(_2759_),
    .A2(_2752_));
 sg13g2_xnor2_1 _7119_ (.Y(_2760_),
    .A(_0203_),
    .B(_2730_));
 sg13g2_a221oi_1 _7120_ (.B2(_2760_),
    .C1(_2759_),
    .B1(net1699),
    .A1(\z80.tv80s.di_reg[5] ),
    .Y(_2761_),
    .A2(net1706));
 sg13g2_nand3_1 _7121_ (.B(_2756_),
    .C(_2761_),
    .A(_2608_),
    .Y(_2762_));
 sg13g2_o21ai_1 _7122_ (.B1(_2762_),
    .Y(_2763_),
    .A1(\z80.tv80s.i_tv80_core.PC[5] ),
    .A2(_2608_));
 sg13g2_o21ai_1 _7123_ (.B1(_2755_),
    .Y(_2764_),
    .A1(net1867),
    .A2(_2763_));
 sg13g2_mux2_1 _7124_ (.A0(_2764_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net1781),
    .X(_2765_));
 sg13g2_a21oi_1 _7125_ (.A1(net1839),
    .A2(_2765_),
    .Y(_2766_),
    .B1(_2754_));
 sg13g2_nand2_1 _7126_ (.Y(_2767_),
    .A(net2133),
    .B(net1726));
 sg13g2_a21oi_1 _7127_ (.A1(net2133),
    .A2(net1726),
    .Y(_2768_),
    .B1(net1912));
 sg13g2_o21ai_1 _7128_ (.B1(_2768_),
    .Y(_2769_),
    .A1(net1726),
    .A2(_2766_));
 sg13g2_o21ai_1 _7129_ (.B1(_2769_),
    .Y(_2770_),
    .A1(\z80.tv80s.i_tv80_core.R[5] ),
    .A2(net1895));
 sg13g2_nor2_1 _7130_ (.A(net383),
    .B(net1681),
    .Y(_2771_));
 sg13g2_a21oi_1 _7131_ (.A1(net1681),
    .A2(_2770_),
    .Y(_0478_),
    .B1(_2771_));
 sg13g2_and2_1 _7132_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .B(net1724),
    .X(_2772_));
 sg13g2_a21oi_1 _7133_ (.A1(_0721_),
    .A2(net2154),
    .Y(_2773_),
    .B1(net2176));
 sg13g2_o21ai_1 _7134_ (.B1(_2773_),
    .Y(_2774_),
    .A1(_0129_),
    .A2(net2154));
 sg13g2_o21ai_1 _7135_ (.B1(net2176),
    .Y(_2775_),
    .A1(_0131_),
    .A2(net2162));
 sg13g2_a21oi_1 _7136_ (.A1(_0722_),
    .A2(net2154),
    .Y(_2776_),
    .B1(_2775_));
 sg13g2_nor2_1 _7137_ (.A(net2007),
    .B(_2776_),
    .Y(_2777_));
 sg13g2_mux4_1 _7138_ (.S0(net2176),
    .A0(_0125_),
    .A1(_0127_),
    .A2(_0126_),
    .A3(_0128_),
    .S1(net2154),
    .X(_2778_));
 sg13g2_nor2_1 _7139_ (.A(net2174),
    .B(_2778_),
    .Y(_2779_));
 sg13g2_a21oi_2 _7140_ (.B1(_2779_),
    .Y(_2780_),
    .A2(_2777_),
    .A1(_2774_));
 sg13g2_inv_2 _7141_ (.Y(_2781_),
    .A(_2780_));
 sg13g2_nand2b_1 _7142_ (.Y(_2782_),
    .B(_2781_),
    .A_N(net1838));
 sg13g2_and2_1 _7143_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .B(net1781),
    .X(_2783_));
 sg13g2_a21oi_1 _7144_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A2(net1872),
    .Y(_2784_),
    .B1(_2627_));
 sg13g2_nand4_1 _7145_ (.B(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .C(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A(net2133),
    .Y(_2785_),
    .D(net2134));
 sg13g2_nor3_1 _7146_ (.A(net1762),
    .B(_2640_),
    .C(_2785_),
    .Y(_2786_));
 sg13g2_nand2b_1 _7147_ (.Y(_2787_),
    .B(net2054),
    .A_N(_0204_));
 sg13g2_a21oi_1 _7148_ (.A1(net2012),
    .A2(_0776_),
    .Y(_2788_),
    .B1(net1926));
 sg13g2_a221oi_1 _7149_ (.B2(_2788_),
    .C1(net1701),
    .B1(_2787_),
    .A1(net1923),
    .Y(_2789_),
    .A2(_2780_));
 sg13g2_a221oi_1 _7150_ (.B2(net1708),
    .C1(net1710),
    .B1(_2781_),
    .A1(\z80.tv80s.i_tv80_core.SP[6] ),
    .Y(_2790_),
    .A2(net1705));
 sg13g2_nor2b_1 _7151_ (.A(_0204_),
    .B_N(_2786_),
    .Y(_2791_));
 sg13g2_xnor2_1 _7152_ (.Y(_2792_),
    .A(_0204_),
    .B(_2786_));
 sg13g2_a221oi_1 _7153_ (.B2(_2792_),
    .C1(_2789_),
    .B1(net1699),
    .A1(net2045),
    .Y(_2793_),
    .A2(net1706));
 sg13g2_a22oi_1 _7154_ (.Y(_2794_),
    .B1(_2790_),
    .B2(_2793_),
    .A2(net1712),
    .A1(_0749_));
 sg13g2_nand2_1 _7155_ (.Y(_2795_),
    .A(net1921),
    .B(_2794_));
 sg13g2_a21oi_1 _7156_ (.A1(_2784_),
    .A2(_2795_),
    .Y(_2796_),
    .B1(net1782));
 sg13g2_o21ai_1 _7157_ (.B1(net1841),
    .Y(_2797_),
    .A1(_2783_),
    .A2(_2796_));
 sg13g2_a21oi_1 _7158_ (.A1(_2782_),
    .A2(_2797_),
    .Y(_2798_),
    .B1(net1724));
 sg13g2_o21ai_1 _7159_ (.B1(net1903),
    .Y(_2799_),
    .A1(_2772_),
    .A2(_2798_));
 sg13g2_a21oi_1 _7160_ (.A1(\z80.tv80s.i_tv80_core.R[6] ),
    .A2(net1907),
    .Y(_2800_),
    .B1(net1685));
 sg13g2_a22oi_1 _7161_ (.Y(_0479_),
    .B1(_2799_),
    .B2(_2800_),
    .A2(net1685),
    .A1(_0758_));
 sg13g2_nand2_1 _7162_ (.Y(_2801_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .B(net1782));
 sg13g2_a21oi_1 _7163_ (.A1(_0730_),
    .A2(net2156),
    .Y(_2802_),
    .B1(net2177));
 sg13g2_o21ai_1 _7164_ (.B1(_2802_),
    .Y(_2803_),
    .A1(_0145_),
    .A2(net2156));
 sg13g2_o21ai_1 _7165_ (.B1(net2177),
    .Y(_2804_),
    .A1(_0147_),
    .A2(net2156));
 sg13g2_a21oi_1 _7166_ (.A1(_0731_),
    .A2(net2156),
    .Y(_2805_),
    .B1(_2804_));
 sg13g2_nor2_1 _7167_ (.A(net2007),
    .B(_2805_),
    .Y(_2806_));
 sg13g2_mux4_1 _7168_ (.S0(net2177),
    .A0(_0141_),
    .A1(_0143_),
    .A2(_0142_),
    .A3(_0144_),
    .S1(net2156),
    .X(_2807_));
 sg13g2_nor2_1 _7169_ (.A(net2174),
    .B(_2807_),
    .Y(_2808_));
 sg13g2_a21oi_2 _7170_ (.B1(_2808_),
    .Y(_2809_),
    .A2(_2806_),
    .A1(_2803_));
 sg13g2_inv_1 _7171_ (.Y(_2810_),
    .A(_2809_));
 sg13g2_a221oi_1 _7172_ (.B2(_2810_),
    .C1(_2605_),
    .B1(net1709),
    .A1(_0777_),
    .Y(_2811_),
    .A2(net1712));
 sg13g2_nand2b_1 _7173_ (.Y(_2812_),
    .B(net2053),
    .A_N(_0206_));
 sg13g2_a21oi_1 _7174_ (.A1(net2013),
    .A2(_0777_),
    .Y(_2813_),
    .B1(net1927));
 sg13g2_a22oi_1 _7175_ (.Y(_2814_),
    .B1(_2812_),
    .B2(_2813_),
    .A2(_2809_),
    .A1(net1924));
 sg13g2_xnor2_1 _7176_ (.Y(_2815_),
    .A(_0206_),
    .B(_2791_));
 sg13g2_a22oi_1 _7177_ (.Y(_2816_),
    .B1(_2815_),
    .B2(net1699),
    .A2(_2814_),
    .A1(_1336_));
 sg13g2_a22oi_1 _7178_ (.Y(_2817_),
    .B1(net1704),
    .B2(\z80.tv80s.i_tv80_core.SP[7] ),
    .A2(net1706),
    .A1(net2044));
 sg13g2_nand3_1 _7179_ (.B(_2816_),
    .C(_2817_),
    .A(_2811_),
    .Y(_2818_));
 sg13g2_a21oi_1 _7180_ (.A1(_0206_),
    .A2(net1872),
    .Y(_2819_),
    .B1(net1758));
 sg13g2_a22oi_1 _7181_ (.Y(_2820_),
    .B1(_2818_),
    .B2(_2819_),
    .A2(net1782),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sg13g2_inv_1 _7182_ (.Y(_2821_),
    .A(_2820_));
 sg13g2_nor2_1 _7183_ (.A(net1840),
    .B(_2809_),
    .Y(_2822_));
 sg13g2_a21oi_1 _7184_ (.A1(net1840),
    .A2(_2821_),
    .Y(_2823_),
    .B1(_2822_));
 sg13g2_nand2_1 _7185_ (.Y(_2824_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .B(net1725));
 sg13g2_o21ai_1 _7186_ (.B1(_2824_),
    .Y(_2825_),
    .A1(net1724),
    .A2(_2823_));
 sg13g2_nor2_1 _7187_ (.A(net1908),
    .B(_2825_),
    .Y(_2826_));
 sg13g2_o21ai_1 _7188_ (.B1(net1683),
    .Y(_2827_),
    .A1(\z80.tv80s.i_tv80_core.R[7] ),
    .A2(net1899));
 sg13g2_nand2_1 _7189_ (.Y(_2828_),
    .A(net457),
    .B(net1685));
 sg13g2_o21ai_1 _7190_ (.B1(_2828_),
    .Y(_0480_),
    .A1(_2826_),
    .A2(_2827_));
 sg13g2_nand2_1 _7191_ (.Y(_2829_),
    .A(net479),
    .B(net1685));
 sg13g2_mux2_1 _7192_ (.A0(_0041_),
    .A1(_0042_),
    .S(net2160),
    .X(_2830_));
 sg13g2_nand2b_1 _7193_ (.Y(_2831_),
    .B(net2160),
    .A_N(_0044_));
 sg13g2_o21ai_1 _7194_ (.B1(_2831_),
    .Y(_2832_),
    .A1(_0043_),
    .A2(net2160));
 sg13g2_a21oi_1 _7195_ (.A1(net2008),
    .A2(_2830_),
    .Y(_2833_),
    .B1(net2006));
 sg13g2_o21ai_1 _7196_ (.B1(_2833_),
    .Y(_2834_),
    .A1(net2008),
    .A2(_2832_));
 sg13g2_mux4_1 _7197_ (.S0(net2178),
    .A0(_0035_),
    .A1(_0037_),
    .A2(_0036_),
    .A3(_0038_),
    .S1(net2160),
    .X(_2835_));
 sg13g2_o21ai_1 _7198_ (.B1(_2834_),
    .Y(_2836_),
    .A1(net2173),
    .A2(_2835_));
 sg13g2_nand2b_1 _7199_ (.Y(_2837_),
    .B(_2836_),
    .A_N(net1840));
 sg13g2_and2_1 _7200_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .B(net1782),
    .X(_2838_));
 sg13g2_nand2_1 _7201_ (.Y(_2839_),
    .A(\z80.tv80s.i_tv80_core.I[0] ),
    .B(net1870));
 sg13g2_nand2_1 _7202_ (.Y(_2840_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sg13g2_nor3_2 _7203_ (.A(_2640_),
    .B(_2785_),
    .C(_2840_),
    .Y(_2841_));
 sg13g2_nor2b_1 _7204_ (.A(_0170_),
    .B_N(_2841_),
    .Y(_2842_));
 sg13g2_xnor2_1 _7205_ (.Y(_2843_),
    .A(_0170_),
    .B(_2841_));
 sg13g2_nor2_1 _7206_ (.A(net1762),
    .B(_2843_),
    .Y(_2844_));
 sg13g2_a21oi_1 _7207_ (.A1(_0169_),
    .A2(net1762),
    .Y(_2845_),
    .B1(_2844_));
 sg13g2_nand2_1 _7208_ (.Y(_2846_),
    .A(net2012),
    .B(_0171_));
 sg13g2_a21oi_1 _7209_ (.A1(net2053),
    .A2(_0170_),
    .Y(_2847_),
    .B1(net1927));
 sg13g2_a22oi_1 _7210_ (.Y(_2848_),
    .B1(_2846_),
    .B2(_2847_),
    .A2(_2836_),
    .A1(net1926));
 sg13g2_nor2_1 _7211_ (.A(_1335_),
    .B(_2848_),
    .Y(_2849_));
 sg13g2_a221oi_1 _7212_ (.B2(net1709),
    .C1(net1711),
    .B1(_2836_),
    .A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .Y(_2850_),
    .A2(_2614_));
 sg13g2_a221oi_1 _7213_ (.B2(_2845_),
    .C1(_2849_),
    .B1(net1699),
    .A1(\z80.tv80s.i_tv80_core.ACC[0] ),
    .Y(_2851_),
    .A2(net1707));
 sg13g2_a221oi_1 _7214_ (.B2(_2851_),
    .C1(net1870),
    .B1(_2850_),
    .A1(_0734_),
    .Y(_2852_),
    .A2(net1711));
 sg13g2_a21oi_1 _7215_ (.A1(\z80.tv80s.i_tv80_core.I[0] ),
    .A2(net1872),
    .Y(_2853_),
    .B1(_2852_));
 sg13g2_nor2_1 _7216_ (.A(net1758),
    .B(_2853_),
    .Y(_2854_));
 sg13g2_o21ai_1 _7217_ (.B1(net1840),
    .Y(_2855_),
    .A1(_2838_),
    .A2(_2854_));
 sg13g2_a21oi_1 _7218_ (.A1(_2837_),
    .A2(_2855_),
    .Y(_2856_),
    .B1(net1723));
 sg13g2_and2_1 _7219_ (.A(\z80.tv80s.di_reg[0] ),
    .B(net1723),
    .X(_2857_));
 sg13g2_nor3_2 _7220_ (.A(net1911),
    .B(_2856_),
    .C(_2857_),
    .Y(_2858_));
 sg13g2_o21ai_1 _7221_ (.B1(net1683),
    .Y(_2859_),
    .A1(\z80.tv80s.i_tv80_core.I[0] ),
    .A2(net1899));
 sg13g2_o21ai_1 _7222_ (.B1(_2829_),
    .Y(_0481_),
    .A1(_2858_),
    .A2(_2859_));
 sg13g2_nand2_1 _7223_ (.Y(_2860_),
    .A(net241),
    .B(net1684));
 sg13g2_mux2_1 _7224_ (.A0(_0049_),
    .A1(_0050_),
    .S(net2159),
    .X(_2861_));
 sg13g2_o21ai_1 _7225_ (.B1(net2180),
    .Y(_2862_),
    .A1(_0051_),
    .A2(net2159));
 sg13g2_a21oi_1 _7226_ (.A1(_0698_),
    .A2(net2159),
    .Y(_2863_),
    .B1(_2862_));
 sg13g2_a21oi_1 _7227_ (.A1(net2008),
    .A2(_2861_),
    .Y(_2864_),
    .B1(net2006));
 sg13g2_nand2b_1 _7228_ (.Y(_2865_),
    .B(_2864_),
    .A_N(_2863_));
 sg13g2_mux4_1 _7229_ (.S0(net2180),
    .A0(_0045_),
    .A1(_0047_),
    .A2(_0046_),
    .A3(_0048_),
    .S1(net2158),
    .X(_2866_));
 sg13g2_o21ai_1 _7230_ (.B1(_2865_),
    .Y(_2867_),
    .A1(net2173),
    .A2(_2866_));
 sg13g2_nor2b_1 _7231_ (.A(net1836),
    .B_N(_2867_),
    .Y(_2868_));
 sg13g2_nand2_1 _7232_ (.Y(_2869_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .B(net1784));
 sg13g2_xnor2_1 _7233_ (.Y(_2870_),
    .A(_0173_),
    .B(_2842_));
 sg13g2_nor2_1 _7234_ (.A(net1763),
    .B(_2870_),
    .Y(_2871_));
 sg13g2_a21oi_1 _7235_ (.A1(_0172_),
    .A2(net1762),
    .Y(_2872_),
    .B1(_2871_));
 sg13g2_nand2_1 _7236_ (.Y(_2873_),
    .A(net1699),
    .B(_2872_));
 sg13g2_nand2_1 _7237_ (.Y(_2874_),
    .A(net2053),
    .B(_0173_));
 sg13g2_a21oi_1 _7238_ (.A1(net2011),
    .A2(_0174_),
    .Y(_2875_),
    .B1(net1925));
 sg13g2_a22oi_1 _7239_ (.Y(_2876_),
    .B1(_2874_),
    .B2(_2875_),
    .A2(_2867_),
    .A1(net1925));
 sg13g2_nor2_1 _7240_ (.A(net1702),
    .B(_2876_),
    .Y(_2877_));
 sg13g2_a22oi_1 _7241_ (.Y(_2878_),
    .B1(net1704),
    .B2(\z80.tv80s.i_tv80_core.SP[9] ),
    .A2(net1706),
    .A1(\z80.tv80s.i_tv80_core.ACC[1] ));
 sg13g2_a21oi_1 _7242_ (.A1(net1709),
    .A2(_2867_),
    .Y(_2879_),
    .B1(_2877_));
 sg13g2_nand4_1 _7243_ (.B(_2873_),
    .C(_2878_),
    .A(_2608_),
    .Y(_2880_),
    .D(_2879_));
 sg13g2_a21oi_1 _7244_ (.A1(_0740_),
    .A2(net1711),
    .Y(_2881_),
    .B1(net1870));
 sg13g2_a22oi_1 _7245_ (.Y(_2882_),
    .B1(_2880_),
    .B2(_2881_),
    .A2(net1869),
    .A1(\z80.tv80s.i_tv80_core.I[1] ));
 sg13g2_o21ai_1 _7246_ (.B1(_2869_),
    .Y(_2883_),
    .A1(net1757),
    .A2(_2882_));
 sg13g2_a21oi_2 _7247_ (.B1(_2868_),
    .Y(_2884_),
    .A2(_2883_),
    .A1(net1836));
 sg13g2_nand2_1 _7248_ (.Y(_2885_),
    .A(\z80.tv80s.di_reg[1] ),
    .B(net1722));
 sg13g2_a21oi_1 _7249_ (.A1(net2050),
    .A2(net1718),
    .Y(_2886_),
    .B1(net1906));
 sg13g2_o21ai_1 _7250_ (.B1(_2886_),
    .Y(_2887_),
    .A1(net1718),
    .A2(_2884_));
 sg13g2_o21ai_1 _7251_ (.B1(_2887_),
    .Y(_2888_),
    .A1(\z80.tv80s.i_tv80_core.I[1] ),
    .A2(net1897));
 sg13g2_o21ai_1 _7252_ (.B1(_2860_),
    .Y(_0482_),
    .A1(net1684),
    .A2(_2888_));
 sg13g2_and2_1 _7253_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .B(net1784),
    .X(_2889_));
 sg13g2_nand2_1 _7254_ (.Y(_2890_),
    .A(\z80.tv80s.i_tv80_core.I[2] ),
    .B(net1871));
 sg13g2_and3_1 _7255_ (.X(_2891_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .C(_2841_));
 sg13g2_nor2b_1 _7256_ (.A(_0176_),
    .B_N(_2891_),
    .Y(_2892_));
 sg13g2_xnor2_1 _7257_ (.Y(_2893_),
    .A(_0176_),
    .B(_2891_));
 sg13g2_nor2_1 _7258_ (.A(net1761),
    .B(_2893_),
    .Y(_2894_));
 sg13g2_a21oi_1 _7259_ (.A1(_0175_),
    .A2(net1761),
    .Y(_2895_),
    .B1(_2894_));
 sg13g2_mux2_1 _7260_ (.A0(_0057_),
    .A1(_0058_),
    .S(net2160),
    .X(_2896_));
 sg13g2_nand2_1 _7261_ (.Y(_2897_),
    .A(net2008),
    .B(_2896_));
 sg13g2_mux2_1 _7262_ (.A0(_0059_),
    .A1(_0060_),
    .S(net2160),
    .X(_2898_));
 sg13g2_a21oi_1 _7263_ (.A1(net2178),
    .A2(_2898_),
    .Y(_2899_),
    .B1(net2006));
 sg13g2_mux4_1 _7264_ (.S0(net2180),
    .A0(_0053_),
    .A1(_0055_),
    .A2(_0054_),
    .A3(_0056_),
    .S1(net2160),
    .X(_2900_));
 sg13g2_nor2_1 _7265_ (.A(net2173),
    .B(_2900_),
    .Y(_2901_));
 sg13g2_a21oi_2 _7266_ (.B1(_2901_),
    .Y(_2902_),
    .A2(_2899_),
    .A1(_2897_));
 sg13g2_inv_1 _7267_ (.Y(_2903_),
    .A(_2902_));
 sg13g2_nand2b_1 _7268_ (.Y(_2904_),
    .B(net2053),
    .A_N(_0176_));
 sg13g2_a21oi_1 _7269_ (.A1(net2011),
    .A2(_0765_),
    .Y(_2905_),
    .B1(net1925));
 sg13g2_a221oi_1 _7270_ (.B2(_2905_),
    .C1(net1702),
    .B1(_2904_),
    .A1(net1926),
    .Y(_2906_),
    .A2(_2902_));
 sg13g2_a221oi_1 _7271_ (.B2(net1709),
    .C1(net1711),
    .B1(_2903_),
    .A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .Y(_2907_),
    .A2(net1707));
 sg13g2_a221oi_1 _7272_ (.B2(_2895_),
    .C1(_2906_),
    .B1(net1700),
    .A1(\z80.tv80s.i_tv80_core.SP[10] ),
    .Y(_2908_),
    .A2(net1705));
 sg13g2_a22oi_1 _7273_ (.Y(_2909_),
    .B1(_2907_),
    .B2(_2908_),
    .A2(net1711),
    .A1(_0744_));
 sg13g2_nand2_1 _7274_ (.Y(_2910_),
    .A(net1920),
    .B(_2909_));
 sg13g2_a21oi_1 _7275_ (.A1(_2890_),
    .A2(_2910_),
    .Y(_2911_),
    .B1(net1757));
 sg13g2_o21ai_1 _7276_ (.B1(net1836),
    .Y(_2912_),
    .A1(_2889_),
    .A2(_2911_));
 sg13g2_nand2b_1 _7277_ (.Y(_2913_),
    .B(_2903_),
    .A_N(net1836));
 sg13g2_a21oi_2 _7278_ (.B1(net1722),
    .Y(_2914_),
    .A2(_2913_),
    .A1(_2912_));
 sg13g2_a21oi_1 _7279_ (.A1(net2049),
    .A2(net1719),
    .Y(_2915_),
    .B1(_2914_));
 sg13g2_o21ai_1 _7280_ (.B1(net1683),
    .Y(_2916_),
    .A1(\z80.tv80s.i_tv80_core.I[2] ),
    .A2(net1897));
 sg13g2_a21oi_2 _7281_ (.B1(_2916_),
    .Y(_2917_),
    .A2(_2915_),
    .A1(net1897));
 sg13g2_a21o_1 _7282_ (.A2(net1684),
    .A1(net451),
    .B1(_2917_),
    .X(_0483_));
 sg13g2_a21oi_1 _7283_ (.A1(_0707_),
    .A2(net2158),
    .Y(_2918_),
    .B1(net2178));
 sg13g2_o21ai_1 _7284_ (.B1(_2918_),
    .Y(_2919_),
    .A1(_0073_),
    .A2(net2158));
 sg13g2_mux2_1 _7285_ (.A0(_0075_),
    .A1(_0076_),
    .S(net2158),
    .X(_2920_));
 sg13g2_a21oi_1 _7286_ (.A1(net2178),
    .A2(_2920_),
    .Y(_2921_),
    .B1(net2006));
 sg13g2_mux4_1 _7287_ (.S0(net2178),
    .A0(_0069_),
    .A1(_0071_),
    .A2(_0070_),
    .A3(_0072_),
    .S1(net2158),
    .X(_2922_));
 sg13g2_nor2_1 _7288_ (.A(net2173),
    .B(_2922_),
    .Y(_2923_));
 sg13g2_a21oi_2 _7289_ (.B1(_2923_),
    .Y(_2924_),
    .A2(_2921_),
    .A1(_2919_));
 sg13g2_inv_1 _7290_ (.Y(_2925_),
    .A(_2924_));
 sg13g2_nor2_1 _7291_ (.A(net1835),
    .B(_2924_),
    .Y(_2926_));
 sg13g2_nand2_1 _7292_ (.Y(_2927_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .B(net1784));
 sg13g2_xnor2_1 _7293_ (.Y(_2928_),
    .A(_0179_),
    .B(_2892_));
 sg13g2_nor2_1 _7294_ (.A(net1761),
    .B(_2928_),
    .Y(_2929_));
 sg13g2_a21oi_1 _7295_ (.A1(_0178_),
    .A2(net1760),
    .Y(_2930_),
    .B1(_2929_));
 sg13g2_nand2b_1 _7296_ (.Y(_2931_),
    .B(net2052),
    .A_N(_0179_));
 sg13g2_a21oi_1 _7297_ (.A1(net2011),
    .A2(_0766_),
    .Y(_2932_),
    .B1(net1925));
 sg13g2_a221oi_1 _7298_ (.B2(_2932_),
    .C1(net1702),
    .B1(_2931_),
    .A1(net1925),
    .Y(_2933_),
    .A2(_2924_));
 sg13g2_a221oi_1 _7299_ (.B2(net1708),
    .C1(net1710),
    .B1(_2925_),
    .A1(\z80.tv80s.i_tv80_core.SP[11] ),
    .Y(_2934_),
    .A2(net1704));
 sg13g2_a221oi_1 _7300_ (.B2(_2930_),
    .C1(_2933_),
    .B1(net1700),
    .A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .Y(_2935_),
    .A2(_2613_));
 sg13g2_a221oi_1 _7301_ (.B2(_2935_),
    .C1(net1869),
    .B1(_2934_),
    .A1(_0745_),
    .Y(_2936_),
    .A2(net1711));
 sg13g2_a21oi_1 _7302_ (.A1(\z80.tv80s.i_tv80_core.I[3] ),
    .A2(net1869),
    .Y(_2937_),
    .B1(_2936_));
 sg13g2_o21ai_1 _7303_ (.B1(_2927_),
    .Y(_2938_),
    .A1(net1757),
    .A2(_2937_));
 sg13g2_a21oi_2 _7304_ (.B1(_2926_),
    .Y(_2939_),
    .A2(_2938_),
    .A1(net1836));
 sg13g2_nand2_1 _7305_ (.Y(_2940_),
    .A(\z80.tv80s.di_reg[3] ),
    .B(net1722));
 sg13g2_a21oi_1 _7306_ (.A1(net2048),
    .A2(net1718),
    .Y(_2941_),
    .B1(net1906));
 sg13g2_o21ai_1 _7307_ (.B1(_2941_),
    .Y(_2942_),
    .A1(net1718),
    .A2(_2939_));
 sg13g2_o21ai_1 _7308_ (.B1(_2942_),
    .Y(_2943_),
    .A1(\z80.tv80s.i_tv80_core.I[3] ),
    .A2(net1897));
 sg13g2_nor2_1 _7309_ (.A(net368),
    .B(net1682),
    .Y(_2944_));
 sg13g2_a21oi_1 _7310_ (.A1(net1681),
    .A2(_2943_),
    .Y(_0484_),
    .B1(_2944_));
 sg13g2_nand2_1 _7311_ (.Y(_2945_),
    .A(net314),
    .B(net1684));
 sg13g2_nand2_1 _7312_ (.Y(_2946_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .B(net1784));
 sg13g2_nand3_1 _7313_ (.B(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .C(_2891_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .Y(_2947_));
 sg13g2_inv_1 _7314_ (.Y(_2948_),
    .A(_2947_));
 sg13g2_nor2_1 _7315_ (.A(_0182_),
    .B(_2947_),
    .Y(_2949_));
 sg13g2_xor2_1 _7316_ (.B(_2947_),
    .A(_0182_),
    .X(_2950_));
 sg13g2_nor2_1 _7317_ (.A(net1760),
    .B(_2950_),
    .Y(_2951_));
 sg13g2_a21oi_1 _7318_ (.A1(_0181_),
    .A2(net1760),
    .Y(_2952_),
    .B1(_2951_));
 sg13g2_mux2_1 _7319_ (.A0(_0089_),
    .A1(_0090_),
    .S(net2157),
    .X(_2953_));
 sg13g2_nand2_1 _7320_ (.Y(_2954_),
    .A(net2008),
    .B(_2953_));
 sg13g2_mux2_1 _7321_ (.A0(_0091_),
    .A1(_0092_),
    .S(net2157),
    .X(_2955_));
 sg13g2_a21oi_1 _7322_ (.A1(net2178),
    .A2(_2955_),
    .Y(_2956_),
    .B1(_0761_));
 sg13g2_mux4_1 _7323_ (.S0(net2179),
    .A0(_0085_),
    .A1(_0087_),
    .A2(_0086_),
    .A3(_0088_),
    .S1(net2157),
    .X(_2957_));
 sg13g2_nor2_1 _7324_ (.A(net2173),
    .B(_2957_),
    .Y(_2958_));
 sg13g2_a21oi_2 _7325_ (.B1(_2958_),
    .Y(_2959_),
    .A2(_2956_),
    .A1(_2954_));
 sg13g2_inv_1 _7326_ (.Y(_2960_),
    .A(_2959_));
 sg13g2_nand2_1 _7327_ (.Y(_2961_),
    .A(net2011),
    .B(_0183_));
 sg13g2_a21oi_1 _7328_ (.A1(net2052),
    .A2(_0182_),
    .Y(_2962_),
    .B1(net1924));
 sg13g2_a22oi_1 _7329_ (.Y(_2963_),
    .B1(_2961_),
    .B2(_2962_),
    .A2(_2960_),
    .A1(net1924));
 sg13g2_nor2_1 _7330_ (.A(net1701),
    .B(_2963_),
    .Y(_2964_));
 sg13g2_a221oi_1 _7331_ (.B2(net1708),
    .C1(net1710),
    .B1(_2960_),
    .A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .Y(_2965_),
    .A2(net1706));
 sg13g2_a221oi_1 _7332_ (.B2(_2952_),
    .C1(_2964_),
    .B1(net1700),
    .A1(\z80.tv80s.i_tv80_core.SP[12] ),
    .Y(_2966_),
    .A2(net1705));
 sg13g2_a221oi_1 _7333_ (.B2(_2966_),
    .C1(net1866),
    .B1(_2965_),
    .A1(_0746_),
    .Y(_2967_),
    .A2(net1710));
 sg13g2_a21oi_1 _7334_ (.A1(\z80.tv80s.i_tv80_core.I[4] ),
    .A2(net1866),
    .Y(_2968_),
    .B1(_2967_));
 sg13g2_o21ai_1 _7335_ (.B1(_2946_),
    .Y(_2969_),
    .A1(net1756),
    .A2(_2968_));
 sg13g2_nor2_1 _7336_ (.A(net1837),
    .B(_2959_),
    .Y(_2970_));
 sg13g2_a21oi_2 _7337_ (.B1(_2970_),
    .Y(_2971_),
    .A2(_2969_),
    .A1(net1837));
 sg13g2_nand2_1 _7338_ (.Y(_2972_),
    .A(net2047),
    .B(net1721));
 sg13g2_a21oi_1 _7339_ (.A1(net2047),
    .A2(net1717),
    .Y(_2973_),
    .B1(net1906));
 sg13g2_o21ai_1 _7340_ (.B1(_2973_),
    .Y(_2974_),
    .A1(net1717),
    .A2(_2971_));
 sg13g2_o21ai_1 _7341_ (.B1(_2974_),
    .Y(_2975_),
    .A1(\z80.tv80s.i_tv80_core.I[4] ),
    .A2(net1896));
 sg13g2_o21ai_1 _7342_ (.B1(_2945_),
    .Y(_0485_),
    .A1(net1684),
    .A2(_2975_));
 sg13g2_nand2_1 _7343_ (.Y(_2976_),
    .A(net306),
    .B(net1684));
 sg13g2_mux2_1 _7344_ (.A0(_0105_),
    .A1(_0106_),
    .S(net2161),
    .X(_2977_));
 sg13g2_nand2_1 _7345_ (.Y(_2978_),
    .A(net2008),
    .B(_2977_));
 sg13g2_mux2_1 _7346_ (.A0(_0107_),
    .A1(_0108_),
    .S(net2161),
    .X(_2979_));
 sg13g2_a21oi_1 _7347_ (.A1(net2179),
    .A2(_2979_),
    .Y(_2980_),
    .B1(net2006));
 sg13g2_mux4_1 _7348_ (.S0(net2179),
    .A0(_0101_),
    .A1(_0103_),
    .A2(_0102_),
    .A3(_0104_),
    .S1(net2157),
    .X(_2981_));
 sg13g2_nor2_1 _7349_ (.A(net2173),
    .B(_2981_),
    .Y(_2982_));
 sg13g2_a21oi_2 _7350_ (.B1(_2982_),
    .Y(_2983_),
    .A2(_2980_),
    .A1(_2978_));
 sg13g2_inv_1 _7351_ (.Y(_2984_),
    .A(_2983_));
 sg13g2_nor2_1 _7352_ (.A(net1835),
    .B(_2983_),
    .Y(_2985_));
 sg13g2_nand2_1 _7353_ (.Y(_2986_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .B(net1784));
 sg13g2_xnor2_1 _7354_ (.Y(_2987_),
    .A(_0185_),
    .B(_2949_));
 sg13g2_nor2_1 _7355_ (.A(net1760),
    .B(_2987_),
    .Y(_2988_));
 sg13g2_a21oi_1 _7356_ (.A1(_0184_),
    .A2(net1761),
    .Y(_2989_),
    .B1(_2988_));
 sg13g2_nand2b_1 _7357_ (.Y(_2990_),
    .B(net2052),
    .A_N(_0185_));
 sg13g2_a21oi_1 _7358_ (.A1(net2011),
    .A2(_0767_),
    .Y(_2991_),
    .B1(net1925));
 sg13g2_a221oi_1 _7359_ (.B2(_2991_),
    .C1(net1702),
    .B1(_2990_),
    .A1(net1925),
    .Y(_2992_),
    .A2(_2983_));
 sg13g2_a221oi_1 _7360_ (.B2(net1709),
    .C1(net1711),
    .B1(_2984_),
    .A1(\z80.tv80s.i_tv80_core.SP[13] ),
    .Y(_2993_),
    .A2(net1705));
 sg13g2_a221oi_1 _7361_ (.B2(_2989_),
    .C1(_2992_),
    .B1(net1700),
    .A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .Y(_2994_),
    .A2(net1707));
 sg13g2_a221oi_1 _7362_ (.B2(_2994_),
    .C1(net1871),
    .B1(_2993_),
    .A1(_0747_),
    .Y(_2995_),
    .A2(net1711));
 sg13g2_a21oi_1 _7363_ (.A1(\z80.tv80s.i_tv80_core.I[5] ),
    .A2(net1869),
    .Y(_2996_),
    .B1(_2995_));
 sg13g2_o21ai_1 _7364_ (.B1(_2986_),
    .Y(_2997_),
    .A1(net1757),
    .A2(_2996_));
 sg13g2_a21oi_2 _7365_ (.B1(_2985_),
    .Y(_2998_),
    .A2(_2997_),
    .A1(net1835));
 sg13g2_nand2_1 _7366_ (.Y(_2999_),
    .A(net2046),
    .B(net1722));
 sg13g2_a21oi_1 _7367_ (.A1(net2046),
    .A2(net1717),
    .Y(_3000_),
    .B1(net1906));
 sg13g2_o21ai_1 _7368_ (.B1(_3000_),
    .Y(_3001_),
    .A1(net1717),
    .A2(_2998_));
 sg13g2_o21ai_1 _7369_ (.B1(_3001_),
    .Y(_3002_),
    .A1(\z80.tv80s.i_tv80_core.I[5] ),
    .A2(net1897));
 sg13g2_o21ai_1 _7370_ (.B1(_2976_),
    .Y(_0486_),
    .A1(net1684),
    .A2(_3002_));
 sg13g2_nand2_1 _7371_ (.Y(_3003_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .B(net1784));
 sg13g2_nand3_1 _7372_ (.B(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .C(_2948_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .Y(_3004_));
 sg13g2_nor2_1 _7373_ (.A(_0188_),
    .B(_3004_),
    .Y(_3005_));
 sg13g2_xor2_1 _7374_ (.B(_3004_),
    .A(_0188_),
    .X(_3006_));
 sg13g2_nor2_1 _7375_ (.A(net1760),
    .B(_3006_),
    .Y(_3007_));
 sg13g2_a21oi_1 _7376_ (.A1(_0187_),
    .A2(net1760),
    .Y(_3008_),
    .B1(_3007_));
 sg13g2_mux2_1 _7377_ (.A0(_0121_),
    .A1(_0122_),
    .S(net2159),
    .X(_3009_));
 sg13g2_nand2_1 _7378_ (.Y(_3010_),
    .A(net2008),
    .B(_3009_));
 sg13g2_o21ai_1 _7379_ (.B1(net2178),
    .Y(_3011_),
    .A1(_0123_),
    .A2(net2158));
 sg13g2_a21oi_1 _7380_ (.A1(_0720_),
    .A2(net2158),
    .Y(_3012_),
    .B1(_3011_));
 sg13g2_nor2_1 _7381_ (.A(net2006),
    .B(_3012_),
    .Y(_3013_));
 sg13g2_mux4_1 _7382_ (.S0(net2178),
    .A0(_0117_),
    .A1(_0119_),
    .A2(_0118_),
    .A3(_0120_),
    .S1(net2158),
    .X(_3014_));
 sg13g2_nor2_1 _7383_ (.A(net2173),
    .B(_3014_),
    .Y(_3015_));
 sg13g2_a21oi_2 _7384_ (.B1(_3015_),
    .Y(_3016_),
    .A2(_3013_),
    .A1(_3010_));
 sg13g2_inv_1 _7385_ (.Y(_3017_),
    .A(_3016_));
 sg13g2_nand2_1 _7386_ (.Y(_3018_),
    .A(net2011),
    .B(_0189_));
 sg13g2_a21oi_1 _7387_ (.A1(net2052),
    .A2(_0188_),
    .Y(_3019_),
    .B1(net1924));
 sg13g2_a22oi_1 _7388_ (.Y(_3020_),
    .B1(_3018_),
    .B2(_3019_),
    .A2(_3017_),
    .A1(net1924));
 sg13g2_nor2_1 _7389_ (.A(net1701),
    .B(_3020_),
    .Y(_3021_));
 sg13g2_a221oi_1 _7390_ (.B2(net1708),
    .C1(net1710),
    .B1(_3017_),
    .A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .Y(_3022_),
    .A2(net1706));
 sg13g2_a221oi_1 _7391_ (.B2(_3008_),
    .C1(_3021_),
    .B1(net1700),
    .A1(\z80.tv80s.i_tv80_core.SP[14] ),
    .Y(_3023_),
    .A2(net1704));
 sg13g2_a221oi_1 _7392_ (.B2(_3023_),
    .C1(net1865),
    .B1(_3022_),
    .A1(_0748_),
    .Y(_3024_),
    .A2(net1710));
 sg13g2_a21oi_1 _7393_ (.A1(\z80.tv80s.i_tv80_core.I[6] ),
    .A2(net1865),
    .Y(_3025_),
    .B1(_3024_));
 sg13g2_o21ai_1 _7394_ (.B1(_3003_),
    .Y(_3026_),
    .A1(net1756),
    .A2(_3025_));
 sg13g2_nor2_1 _7395_ (.A(net1837),
    .B(_3016_),
    .Y(_3027_));
 sg13g2_a21oi_2 _7396_ (.B1(_3027_),
    .Y(_3028_),
    .A2(_3026_),
    .A1(net1837));
 sg13g2_nand2_1 _7397_ (.Y(_3029_),
    .A(net2045),
    .B(net1721));
 sg13g2_a21oi_1 _7398_ (.A1(net2045),
    .A2(net1717),
    .Y(_3030_),
    .B1(net1906));
 sg13g2_o21ai_1 _7399_ (.B1(_3030_),
    .Y(_3031_),
    .A1(net1717),
    .A2(_3028_));
 sg13g2_o21ai_1 _7400_ (.B1(_3031_),
    .Y(_3032_),
    .A1(\z80.tv80s.i_tv80_core.I[6] ),
    .A2(net1896));
 sg13g2_nor2_1 _7401_ (.A(net394),
    .B(net1682),
    .Y(_3033_));
 sg13g2_a21oi_1 _7402_ (.A1(net1681),
    .A2(_3032_),
    .Y(_0487_),
    .B1(_3033_));
 sg13g2_a21oi_1 _7403_ (.A1(_0726_),
    .A2(net2157),
    .Y(_3034_),
    .B1(net2179));
 sg13g2_o21ai_1 _7404_ (.B1(_3034_),
    .Y(_3035_),
    .A1(_0137_),
    .A2(net2157));
 sg13g2_mux2_1 _7405_ (.A0(_0139_),
    .A1(_0140_),
    .S(net2157),
    .X(_3036_));
 sg13g2_a21oi_1 _7406_ (.A1(net2179),
    .A2(_3036_),
    .Y(_3037_),
    .B1(net2006));
 sg13g2_mux4_1 _7407_ (.S0(net2179),
    .A0(_0133_),
    .A1(_0135_),
    .A2(_0134_),
    .A3(_0136_),
    .S1(net2157),
    .X(_3038_));
 sg13g2_nor2_1 _7408_ (.A(net2173),
    .B(_3038_),
    .Y(_3039_));
 sg13g2_a21oi_2 _7409_ (.B1(_3039_),
    .Y(_3040_),
    .A2(_3037_),
    .A1(_3035_));
 sg13g2_inv_1 _7410_ (.Y(_3041_),
    .A(_3040_));
 sg13g2_nor2_1 _7411_ (.A(net1837),
    .B(_3040_),
    .Y(_3042_));
 sg13g2_nand2_1 _7412_ (.Y(_3043_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .B(net1784));
 sg13g2_xnor2_1 _7413_ (.Y(_3044_),
    .A(_0191_),
    .B(_3005_));
 sg13g2_nor2_1 _7414_ (.A(net1760),
    .B(_3044_),
    .Y(_3045_));
 sg13g2_a21oi_1 _7415_ (.A1(_0190_),
    .A2(net1760),
    .Y(_3046_),
    .B1(_3045_));
 sg13g2_nand2b_1 _7416_ (.Y(_3047_),
    .B(net2052),
    .A_N(_0191_));
 sg13g2_a21oi_1 _7417_ (.A1(net2011),
    .A2(_0769_),
    .Y(_3048_),
    .B1(net1925));
 sg13g2_a221oi_1 _7418_ (.B2(_3048_),
    .C1(net1701),
    .B1(_3047_),
    .A1(net1924),
    .Y(_3049_),
    .A2(_3040_));
 sg13g2_a221oi_1 _7419_ (.B2(net1708),
    .C1(net1710),
    .B1(_3041_),
    .A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .Y(_3050_),
    .A2(net1706));
 sg13g2_a221oi_1 _7420_ (.B2(_3046_),
    .C1(_3049_),
    .B1(net1700),
    .A1(\z80.tv80s.i_tv80_core.SP[15] ),
    .Y(_3051_),
    .A2(net1704));
 sg13g2_a221oi_1 _7421_ (.B2(_3051_),
    .C1(net1865),
    .B1(_3050_),
    .A1(_0750_),
    .Y(_3052_),
    .A2(net1710));
 sg13g2_a21oi_1 _7422_ (.A1(\z80.tv80s.i_tv80_core.I[7] ),
    .A2(net1865),
    .Y(_3053_),
    .B1(_3052_));
 sg13g2_o21ai_1 _7423_ (.B1(_3043_),
    .Y(_3054_),
    .A1(net1756),
    .A2(_3053_));
 sg13g2_a21oi_2 _7424_ (.B1(_3042_),
    .Y(_3055_),
    .A2(_3054_),
    .A1(net1837));
 sg13g2_nand2_1 _7425_ (.Y(_3056_),
    .A(net2044),
    .B(net1721));
 sg13g2_a21oi_1 _7426_ (.A1(net2043),
    .A2(net1717),
    .Y(_3057_),
    .B1(net1906));
 sg13g2_o21ai_1 _7427_ (.B1(_3057_),
    .Y(_3058_),
    .A1(net1717),
    .A2(_3055_));
 sg13g2_o21ai_1 _7428_ (.B1(_3058_),
    .Y(_3059_),
    .A1(\z80.tv80s.i_tv80_core.I[7] ),
    .A2(net1896));
 sg13g2_nor2_1 _7429_ (.A(net356),
    .B(net1682),
    .Y(_3060_));
 sg13g2_a21oi_1 _7430_ (.A1(net1682),
    .A2(_3059_),
    .Y(_0488_),
    .B1(_3060_));
 sg13g2_nand2_2 _7431_ (.Y(_3061_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .B(_2382_));
 sg13g2_nand3_1 _7432_ (.B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .C(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .A(_0790_),
    .Y(_3062_));
 sg13g2_nor2_2 _7433_ (.A(_3061_),
    .B(_3062_),
    .Y(_3063_));
 sg13g2_or2_2 _7434_ (.X(_3064_),
    .B(_3062_),
    .A(_3061_));
 sg13g2_a21oi_1 _7435_ (.A1(_0781_),
    .A2(_2288_),
    .Y(_3065_),
    .B1(_2292_));
 sg13g2_nor2_2 _7436_ (.A(_0226_),
    .B(_1763_),
    .Y(_3066_));
 sg13g2_a22oi_1 _7437_ (.Y(_3067_),
    .B1(_1820_),
    .B2(_0226_),
    .A2(_1762_),
    .A1(_0779_));
 sg13g2_nor2b_1 _7438_ (.A(_3066_),
    .B_N(_3067_),
    .Y(_3068_));
 sg13g2_nor2_1 _7439_ (.A(net2036),
    .B(net2038),
    .Y(_3069_));
 sg13g2_nand2_1 _7440_ (.Y(_3070_),
    .A(_0779_),
    .B(_0780_));
 sg13g2_mux2_1 _7441_ (.A0(_3070_),
    .A1(_3068_),
    .S(_3065_),
    .X(_3071_));
 sg13g2_xor2_1 _7442_ (.B(_2204_),
    .A(_2200_),
    .X(_3072_));
 sg13g2_o21ai_1 _7443_ (.B1(_2255_),
    .Y(_3073_),
    .A1(_2190_),
    .A2(_2302_));
 sg13g2_o21ai_1 _7444_ (.B1(_3073_),
    .Y(_3074_),
    .A1(net2148),
    .A2(_3072_));
 sg13g2_a21oi_1 _7445_ (.A1(_0665_),
    .A2(_3074_),
    .Y(_3075_),
    .B1(_1817_));
 sg13g2_nand2_1 _7446_ (.Y(_3076_),
    .A(net2076),
    .B(_0212_));
 sg13g2_a21oi_1 _7447_ (.A1(net2024),
    .A2(_0210_),
    .Y(_3077_),
    .B1(_1777_));
 sg13g2_a221oi_1 _7448_ (.B2(_3077_),
    .C1(_3075_),
    .B1(_3076_),
    .A1(net2034),
    .Y(_3078_),
    .A2(_1798_));
 sg13g2_o21ai_1 _7449_ (.B1(_3078_),
    .Y(_3079_),
    .A1(net2034),
    .A2(_3071_));
 sg13g2_nand3_1 _7450_ (.B(net2034),
    .C(_1798_),
    .A(_0665_),
    .Y(_3080_));
 sg13g2_o21ai_1 _7451_ (.B1(_1813_),
    .Y(_3081_),
    .A1(_0208_),
    .A2(_2487_));
 sg13g2_and4_1 _7452_ (.A(_0800_),
    .B(_3079_),
    .C(_3080_),
    .D(net1796),
    .X(_3082_));
 sg13g2_nand2_2 _7453_ (.Y(_3083_),
    .A(_1516_),
    .B(_1530_));
 sg13g2_nor3_2 _7454_ (.A(_1261_),
    .B(_1526_),
    .C(_3083_),
    .Y(_3084_));
 sg13g2_a21o_1 _7455_ (.A2(_3084_),
    .A1(net1689),
    .B1(_0665_),
    .X(_3085_));
 sg13g2_o21ai_1 _7456_ (.B1(net2151),
    .Y(_3086_),
    .A1(_1259_),
    .A2(_3083_));
 sg13g2_nor2_2 _7457_ (.A(_1261_),
    .B(_3083_),
    .Y(_3087_));
 sg13g2_nand2_1 _7458_ (.Y(_3088_),
    .A(net1688),
    .B(_3087_));
 sg13g2_nand3_1 _7459_ (.B(_3086_),
    .C(_3087_),
    .A(net1688),
    .Y(_3089_));
 sg13g2_nor4_2 _7460_ (.A(_0923_),
    .B(_0926_),
    .C(_0961_),
    .Y(_3090_),
    .D(_1504_));
 sg13g2_nand2_2 _7461_ (.Y(_3091_),
    .A(_1716_),
    .B(_3090_));
 sg13g2_a21oi_1 _7462_ (.A1(_1716_),
    .A2(_3090_),
    .Y(_3092_),
    .B1(_0808_));
 sg13g2_and2_1 _7463_ (.A(_3089_),
    .B(net1821),
    .X(_3093_));
 sg13g2_nor2_2 _7464_ (.A(net1908),
    .B(_3091_),
    .Y(_3094_));
 sg13g2_nand3_1 _7465_ (.B(_1716_),
    .C(_3090_),
    .A(net1895),
    .Y(_3095_));
 sg13g2_nand2_1 _7466_ (.Y(_3096_),
    .A(_0665_),
    .B(net1908));
 sg13g2_o21ai_1 _7467_ (.B1(_3096_),
    .Y(_3097_),
    .A1(\z80.tv80s.i_tv80_core.Fp[0] ),
    .A2(net1819));
 sg13g2_a221oi_1 _7468_ (.B2(_3093_),
    .C1(_3097_),
    .B1(_3085_),
    .A1(_0800_),
    .Y(_3098_),
    .A2(net1796));
 sg13g2_o21ai_1 _7469_ (.B1(_3064_),
    .Y(_3099_),
    .A1(_3082_),
    .A2(_3098_));
 sg13g2_a21oi_1 _7470_ (.A1(_1831_),
    .A2(_3063_),
    .Y(_3100_),
    .B1(net1965));
 sg13g2_a22oi_1 _7471_ (.Y(_3101_),
    .B1(_3099_),
    .B2(_3100_),
    .A2(net1966),
    .A1(net251));
 sg13g2_inv_1 _7472_ (.Y(_0489_),
    .A(_3101_));
 sg13g2_nand4_1 _7473_ (.B(net2035),
    .C(_1809_),
    .A(net2149),
    .Y(_3102_),
    .D(_3070_));
 sg13g2_o21ai_1 _7474_ (.B1(_3102_),
    .Y(_3103_),
    .A1(net2034),
    .A2(_3068_));
 sg13g2_or2_2 _7475_ (.X(_3104_),
    .B(_3083_),
    .A(_0947_));
 sg13g2_nor2_1 _7476_ (.A(net1687),
    .B(_3104_),
    .Y(_3105_));
 sg13g2_o21ai_1 _7477_ (.B1(_3088_),
    .Y(_3106_),
    .A1(net2150),
    .A2(net1680));
 sg13g2_nor2_1 _7478_ (.A(net2150),
    .B(net1895),
    .Y(_3107_));
 sg13g2_and3_1 _7479_ (.X(_3108_),
    .A(net2070),
    .B(net2142),
    .C(_1116_));
 sg13g2_nor3_1 _7480_ (.A(net1795),
    .B(_3107_),
    .C(net1860),
    .Y(_3109_));
 sg13g2_o21ai_1 _7481_ (.B1(_3109_),
    .Y(_3110_),
    .A1(\z80.tv80s.i_tv80_core.Fp[1] ),
    .A2(net1819));
 sg13g2_a21oi_1 _7482_ (.A1(net1821),
    .A2(_3106_),
    .Y(_3111_),
    .B1(_3110_));
 sg13g2_a21o_1 _7483_ (.A2(_3103_),
    .A1(net1795),
    .B1(_3111_),
    .X(_3112_));
 sg13g2_nor2_2 _7484_ (.A(_0032_),
    .B(_1686_),
    .Y(_3113_));
 sg13g2_nor3_2 _7485_ (.A(_1131_),
    .B(_1230_),
    .C(_1673_),
    .Y(_3114_));
 sg13g2_nor3_1 _7486_ (.A(_3063_),
    .B(_3113_),
    .C(_3114_),
    .Y(_3115_));
 sg13g2_a221oi_1 _7487_ (.B2(_3115_),
    .C1(net1966),
    .B1(_3112_),
    .A1(_2005_),
    .Y(_3116_),
    .A2(_3063_));
 sg13g2_a21o_1 _7488_ (.A2(net1965),
    .A1(net324),
    .B1(_3116_),
    .X(_0490_));
 sg13g2_xor2_1 _7489_ (.B(_3065_),
    .A(_2288_),
    .X(_3117_));
 sg13g2_nand2_1 _7490_ (.Y(_3118_),
    .A(_1789_),
    .B(_3117_));
 sg13g2_xor2_1 _7491_ (.B(_2298_),
    .A(_2250_),
    .X(_3119_));
 sg13g2_xor2_1 _7492_ (.B(_2184_),
    .A(_2131_),
    .X(_3120_));
 sg13g2_xor2_1 _7493_ (.B(_2081_),
    .A(_2032_),
    .X(_3121_));
 sg13g2_xor2_1 _7494_ (.B(_1984_),
    .A(_1803_),
    .X(_3122_));
 sg13g2_xnor2_1 _7495_ (.Y(_3123_),
    .A(_3121_),
    .B(_3122_));
 sg13g2_xnor2_1 _7496_ (.Y(_3124_),
    .A(_3120_),
    .B(_3123_));
 sg13g2_a21oi_1 _7497_ (.A1(_3119_),
    .A2(_3124_),
    .Y(_3125_),
    .B1(_1789_));
 sg13g2_o21ai_1 _7498_ (.B1(_3125_),
    .Y(_3126_),
    .A1(_3119_),
    .A2(_3124_));
 sg13g2_a21oi_1 _7499_ (.A1(_3118_),
    .A2(_3126_),
    .Y(_3127_),
    .B1(\z80.tv80s.i_tv80_core.Arith16_r ));
 sg13g2_nor2b_1 _7500_ (.A(net2147),
    .B_N(\z80.tv80s.i_tv80_core.Arith16_r ),
    .Y(_3128_));
 sg13g2_nor3_1 _7501_ (.A(net2034),
    .B(_3127_),
    .C(_3128_),
    .Y(_3129_));
 sg13g2_xor2_1 _7502_ (.B(_2306_),
    .A(_2257_),
    .X(_3130_));
 sg13g2_xnor2_1 _7503_ (.Y(_3131_),
    .A(_2135_),
    .B(_2209_));
 sg13g2_xor2_1 _7504_ (.B(_2087_),
    .A(_2037_),
    .X(_3132_));
 sg13g2_xnor2_1 _7505_ (.Y(_3133_),
    .A(_0782_),
    .B(_1989_));
 sg13g2_xnor2_1 _7506_ (.Y(_3134_),
    .A(_3132_),
    .B(_3133_));
 sg13g2_xnor2_1 _7507_ (.Y(_3135_),
    .A(_3074_),
    .B(_3134_));
 sg13g2_xnor2_1 _7508_ (.Y(_3136_),
    .A(_3131_),
    .B(_3135_));
 sg13g2_o21ai_1 _7509_ (.B1(_1816_),
    .Y(_3137_),
    .A1(_3130_),
    .A2(_3136_));
 sg13g2_a21oi_1 _7510_ (.A1(_3130_),
    .A2(_3136_),
    .Y(_3138_),
    .B1(_3137_));
 sg13g2_xor2_1 _7511_ (.B(_2088_),
    .A(_2043_),
    .X(_3139_));
 sg13g2_xor2_1 _7512_ (.B(_1995_),
    .A(_1807_),
    .X(_3140_));
 sg13g2_xnor2_1 _7513_ (.Y(_3141_),
    .A(_3139_),
    .B(_3140_));
 sg13g2_xnor2_1 _7514_ (.Y(_3142_),
    .A(_2263_),
    .B(_2317_));
 sg13g2_xor2_1 _7515_ (.B(_2214_),
    .A(_2141_),
    .X(_3143_));
 sg13g2_xnor2_1 _7516_ (.Y(_3144_),
    .A(_3142_),
    .B(_3143_));
 sg13g2_a21oi_1 _7517_ (.A1(_3141_),
    .A2(_3144_),
    .Y(_3145_),
    .B1(net2172));
 sg13g2_o21ai_1 _7518_ (.B1(_3145_),
    .Y(_3146_),
    .A1(_3141_),
    .A2(_3144_));
 sg13g2_o21ai_1 _7519_ (.B1(_3146_),
    .Y(_3147_),
    .A1(net2147),
    .A2(_0676_));
 sg13g2_xor2_1 _7520_ (.B(net2030),
    .A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .X(_3148_));
 sg13g2_xor2_1 _7521_ (.B(net2029),
    .A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .X(_3149_));
 sg13g2_xnor2_1 _7522_ (.Y(_3150_),
    .A(_3148_),
    .B(_3149_));
 sg13g2_xnor2_1 _7523_ (.Y(_3151_),
    .A(_2040_),
    .B(_2090_));
 sg13g2_xor2_1 _7524_ (.B(_1994_),
    .A(_1810_),
    .X(_3152_));
 sg13g2_xnor2_1 _7525_ (.Y(_3153_),
    .A(_3151_),
    .B(_3152_));
 sg13g2_o21ai_1 _7526_ (.B1(_1808_),
    .Y(_3154_),
    .A1(_3150_),
    .A2(_3153_));
 sg13g2_a21oi_1 _7527_ (.A1(_3150_),
    .A2(_3153_),
    .Y(_3155_),
    .B1(_3154_));
 sg13g2_o21ai_1 _7528_ (.B1(_2547_),
    .Y(_3156_),
    .A1(net1863),
    .A2(_3147_));
 sg13g2_nor4_2 _7529_ (.A(_3129_),
    .B(_3138_),
    .C(_3155_),
    .Y(_3157_),
    .D(_3156_));
 sg13g2_o21ai_1 _7530_ (.B1(net1796),
    .Y(_3158_),
    .A1(net2147),
    .A2(_2534_));
 sg13g2_nand2_1 _7531_ (.Y(_3159_),
    .A(\z80.tv80s.i_tv80_core.Fp[2] ),
    .B(_3094_));
 sg13g2_a21oi_1 _7532_ (.A1(net2147),
    .A2(net1819),
    .Y(_3160_),
    .B1(net1860));
 sg13g2_a221oi_1 _7533_ (.B2(_3160_),
    .C1(net1796),
    .B1(_3159_),
    .A1(_0799_),
    .Y(_3161_),
    .A2(net1860));
 sg13g2_nor2_1 _7534_ (.A(_3114_),
    .B(_3161_),
    .Y(_3162_));
 sg13g2_o21ai_1 _7535_ (.B1(_3162_),
    .Y(_3163_),
    .A1(_3157_),
    .A2(_3158_));
 sg13g2_xor2_1 _7536_ (.B(net2043),
    .A(net2045),
    .X(_3164_));
 sg13g2_xor2_1 _7537_ (.B(net2046),
    .A(\z80.tv80s.di_reg[4] ),
    .X(_3165_));
 sg13g2_xnor2_1 _7538_ (.Y(_3166_),
    .A(_3164_),
    .B(_3165_));
 sg13g2_xnor2_1 _7539_ (.Y(_3167_),
    .A(net2051),
    .B(net2050));
 sg13g2_xor2_1 _7540_ (.B(net2048),
    .A(net2049),
    .X(_3168_));
 sg13g2_xnor2_1 _7541_ (.Y(_3169_),
    .A(_3167_),
    .B(_3168_));
 sg13g2_xnor2_1 _7542_ (.Y(_3170_),
    .A(_3166_),
    .B(_3169_));
 sg13g2_a21oi_1 _7543_ (.A1(_3114_),
    .A2(_3170_),
    .Y(_3171_),
    .B1(_1688_));
 sg13g2_a22oi_1 _7544_ (.Y(_3172_),
    .B1(_3163_),
    .B2(_3171_),
    .A2(_1688_),
    .A1(\z80.tv80s.i_tv80_core.IncDecZ ));
 sg13g2_a21oi_1 _7545_ (.A1(_2050_),
    .A2(_3063_),
    .Y(_3173_),
    .B1(net1970));
 sg13g2_o21ai_1 _7546_ (.B1(_3173_),
    .Y(_3174_),
    .A1(_3063_),
    .A2(_3172_));
 sg13g2_o21ai_1 _7547_ (.B1(_3174_),
    .Y(_0491_),
    .A1(_0667_),
    .A2(net1994));
 sg13g2_nand2_1 _7548_ (.Y(_3175_),
    .A(net206),
    .B(net1960));
 sg13g2_nand2_1 _7549_ (.Y(_3176_),
    .A(net2146),
    .B(_3087_));
 sg13g2_nor2_1 _7550_ (.A(net2146),
    .B(_3104_),
    .Y(_3177_));
 sg13g2_a21oi_1 _7551_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_3104_),
    .Y(_3178_),
    .B1(_3177_));
 sg13g2_o21ai_1 _7552_ (.B1(_3176_),
    .Y(_3179_),
    .A1(_3087_),
    .A2(_3178_));
 sg13g2_o21ai_1 _7553_ (.B1(net1821),
    .Y(_3180_),
    .A1(_0663_),
    .A2(net1688));
 sg13g2_a21oi_1 _7554_ (.A1(net1688),
    .A2(_3179_),
    .Y(_3181_),
    .B1(_3180_));
 sg13g2_nor2_1 _7555_ (.A(\z80.tv80s.i_tv80_core.Fp[3] ),
    .B(net1819),
    .Y(_3182_));
 sg13g2_nor2_1 _7556_ (.A(\z80.tv80s.i_tv80_core.F[3] ),
    .B(net1895),
    .Y(_3183_));
 sg13g2_or4_1 _7557_ (.A(net1795),
    .B(_3181_),
    .C(_3182_),
    .D(_3183_),
    .X(_3184_));
 sg13g2_mux2_1 _7558_ (.A0(_2081_),
    .A1(_0220_),
    .S(_3066_),
    .X(_3185_));
 sg13g2_nor3_1 _7559_ (.A(_0220_),
    .B(net1887),
    .C(_1813_),
    .Y(_3186_));
 sg13g2_nor3_1 _7560_ (.A(_2093_),
    .B(_2533_),
    .C(_3186_),
    .Y(_3187_));
 sg13g2_o21ai_1 _7561_ (.B1(_3187_),
    .Y(_3188_),
    .A1(net2035),
    .A2(_3185_));
 sg13g2_nand2_1 _7562_ (.Y(_3189_),
    .A(net1796),
    .B(_3188_));
 sg13g2_a21oi_1 _7563_ (.A1(_0663_),
    .A2(_2533_),
    .Y(_3190_),
    .B1(_3189_));
 sg13g2_nor2_1 _7564_ (.A(_3113_),
    .B(_3190_),
    .Y(_3191_));
 sg13g2_a221oi_1 _7565_ (.B2(_3191_),
    .C1(_3063_),
    .B1(_3184_),
    .A1(_2097_),
    .Y(_3192_),
    .A2(_3113_));
 sg13g2_o21ai_1 _7566_ (.B1(net1993),
    .Y(_3193_),
    .A1(_2100_),
    .A2(_3064_));
 sg13g2_o21ai_1 _7567_ (.B1(_3175_),
    .Y(_0492_),
    .A1(_3192_),
    .A2(_3193_));
 sg13g2_a21oi_1 _7568_ (.A1(_2122_),
    .A2(_3069_),
    .Y(_3194_),
    .B1(_1799_));
 sg13g2_o21ai_1 _7569_ (.B1(_3194_),
    .Y(_3195_),
    .A1(_2122_),
    .A2(_3068_));
 sg13g2_nand4_1 _7570_ (.B(net2148),
    .C(_0783_),
    .A(\z80.tv80s.i_tv80_core.F[4] ),
    .Y(_3196_),
    .D(_2033_));
 sg13g2_o21ai_1 _7571_ (.B1(_3196_),
    .Y(_3197_),
    .A1(net2149),
    .A2(_1987_));
 sg13g2_nand2_1 _7572_ (.Y(_3198_),
    .A(_1813_),
    .B(_2534_));
 sg13g2_a221oi_1 _7573_ (.B2(_1816_),
    .C1(_3198_),
    .B1(_3197_),
    .A1(_0778_),
    .Y(_3199_),
    .A2(_3195_));
 sg13g2_o21ai_1 _7574_ (.B1(net1796),
    .Y(_3200_),
    .A1(\z80.tv80s.i_tv80_core.F[4] ),
    .A2(_2534_));
 sg13g2_a21oi_1 _7575_ (.A1(net1688),
    .A2(_3084_),
    .Y(_3201_),
    .B1(\z80.tv80s.i_tv80_core.F[4] ));
 sg13g2_o21ai_1 _7576_ (.B1(_3201_),
    .Y(_3202_),
    .A1(net1687),
    .A2(_3104_));
 sg13g2_nand3_1 _7577_ (.B(_3091_),
    .C(_3202_),
    .A(_3089_),
    .Y(_3203_));
 sg13g2_o21ai_1 _7578_ (.B1(_3203_),
    .Y(_3204_),
    .A1(_0801_),
    .A2(_3091_));
 sg13g2_nor2_1 _7579_ (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .B(net1895),
    .Y(_3205_));
 sg13g2_nor3_1 _7580_ (.A(net1795),
    .B(net1860),
    .C(_3205_),
    .Y(_3206_));
 sg13g2_o21ai_1 _7581_ (.B1(_3206_),
    .Y(_3207_),
    .A1(net1908),
    .A2(_3204_));
 sg13g2_o21ai_1 _7582_ (.B1(_3207_),
    .Y(_3208_),
    .A1(_3199_),
    .A2(_3200_));
 sg13g2_a221oi_1 _7583_ (.B2(_3208_),
    .C1(net1966),
    .B1(_3115_),
    .A1(_2147_),
    .Y(_3209_),
    .A2(_3063_));
 sg13g2_a21o_1 _7584_ (.A2(net1965),
    .A1(net317),
    .B1(_3209_),
    .X(_0493_));
 sg13g2_nand2_1 _7585_ (.Y(_3210_),
    .A(net209),
    .B(net1965));
 sg13g2_nor2_1 _7586_ (.A(net2145),
    .B(_3104_),
    .Y(_3211_));
 sg13g2_a21oi_1 _7587_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_3104_),
    .Y(_3212_),
    .B1(_3211_));
 sg13g2_nor2_1 _7588_ (.A(_3087_),
    .B(_3212_),
    .Y(_3213_));
 sg13g2_a21oi_1 _7589_ (.A1(net2145),
    .A2(_3087_),
    .Y(_3214_),
    .B1(_3213_));
 sg13g2_o21ai_1 _7590_ (.B1(net1820),
    .Y(_3215_),
    .A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(net1688));
 sg13g2_a21o_1 _7591_ (.A2(_3214_),
    .A1(net1688),
    .B1(_3215_),
    .X(_3216_));
 sg13g2_a221oi_1 _7592_ (.B2(\z80.tv80s.i_tv80_core.Fp[5] ),
    .C1(net1795),
    .B1(_3094_),
    .A1(\z80.tv80s.i_tv80_core.F[5] ),
    .Y(_3217_),
    .A2(net1908));
 sg13g2_a21oi_1 _7593_ (.A1(_0222_),
    .A2(_3066_),
    .Y(_3218_),
    .B1(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sg13g2_o21ai_1 _7594_ (.B1(_3218_),
    .Y(_3219_),
    .A1(_2185_),
    .A2(_3066_));
 sg13g2_nor3_1 _7595_ (.A(_0222_),
    .B(net1887),
    .C(_1813_),
    .Y(_3220_));
 sg13g2_nor3_1 _7596_ (.A(_2215_),
    .B(_2533_),
    .C(_3220_),
    .Y(_3221_));
 sg13g2_nand3_1 _7597_ (.B(_3219_),
    .C(_3221_),
    .A(_2210_),
    .Y(_3222_));
 sg13g2_o21ai_1 _7598_ (.B1(_3222_),
    .Y(_3223_),
    .A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_2534_));
 sg13g2_a221oi_1 _7599_ (.B2(net1795),
    .C1(_3113_),
    .B1(_3223_),
    .A1(_3216_),
    .Y(_3224_),
    .A2(_3217_));
 sg13g2_a21oi_1 _7600_ (.A1(_2002_),
    .A2(_3113_),
    .Y(_3225_),
    .B1(_3224_));
 sg13g2_nor2_1 _7601_ (.A(_3063_),
    .B(_3225_),
    .Y(_3226_));
 sg13g2_o21ai_1 _7602_ (.B1(net1993),
    .Y(_3227_),
    .A1(_2219_),
    .A2(_3064_));
 sg13g2_o21ai_1 _7603_ (.B1(_3210_),
    .Y(_0494_),
    .A1(_3226_),
    .A2(_3227_));
 sg13g2_or2_1 _7604_ (.X(_3228_),
    .B(net1819),
    .A(\z80.tv80s.i_tv80_core.Fp[6] ));
 sg13g2_o21ai_1 _7605_ (.B1(_3228_),
    .Y(_3229_),
    .A1(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(_3094_));
 sg13g2_nand2b_1 _7606_ (.Y(_3230_),
    .B(_3229_),
    .A_N(net1861));
 sg13g2_nor4_1 _7607_ (.A(\z80.tv80s.i_tv80_core.I[4] ),
    .B(\z80.tv80s.i_tv80_core.I[5] ),
    .C(\z80.tv80s.i_tv80_core.I[6] ),
    .D(\z80.tv80s.i_tv80_core.I[7] ),
    .Y(_3231_));
 sg13g2_nor4_1 _7608_ (.A(\z80.tv80s.i_tv80_core.I[0] ),
    .B(\z80.tv80s.i_tv80_core.I[1] ),
    .C(\z80.tv80s.i_tv80_core.I[2] ),
    .D(\z80.tv80s.i_tv80_core.I[3] ),
    .Y(_3232_));
 sg13g2_nand2_1 _7609_ (.Y(_3233_),
    .A(_3231_),
    .B(_3232_));
 sg13g2_a21oi_1 _7610_ (.A1(net1861),
    .A2(_3233_),
    .Y(_3234_),
    .B1(net1796));
 sg13g2_a221oi_1 _7611_ (.B2(_3234_),
    .C1(_3114_),
    .B1(_3230_),
    .A1(_2561_),
    .Y(_3235_),
    .A2(net1795));
 sg13g2_nor4_1 _7612_ (.A(\z80.tv80s.di_reg[4] ),
    .B(net2046),
    .C(net2045),
    .D(net2043),
    .Y(_3236_));
 sg13g2_nor4_1 _7613_ (.A(net2051),
    .B(net2050),
    .C(net2049),
    .D(net2048),
    .Y(_3237_));
 sg13g2_nand2_1 _7614_ (.Y(_3238_),
    .A(_3236_),
    .B(_3237_));
 sg13g2_a21oi_1 _7615_ (.A1(_3114_),
    .A2(_3238_),
    .Y(_3239_),
    .B1(_3235_));
 sg13g2_o21ai_1 _7616_ (.B1(net1993),
    .Y(_3240_),
    .A1(_2270_),
    .A2(_3064_));
 sg13g2_a21oi_1 _7617_ (.A1(_3064_),
    .A2(_3239_),
    .Y(_3241_),
    .B1(_3240_));
 sg13g2_a21o_1 _7618_ (.A2(net1970),
    .A1(net335),
    .B1(_3241_),
    .X(_0495_));
 sg13g2_nand2b_1 _7619_ (.Y(_3242_),
    .B(_2298_),
    .A_N(\z80.tv80s.i_tv80_core.Arith16_r ));
 sg13g2_a21oi_1 _7620_ (.A1(_0661_),
    .A2(\z80.tv80s.i_tv80_core.Arith16_r ),
    .Y(_3243_),
    .B1(net2035));
 sg13g2_nand2_1 _7621_ (.Y(_3244_),
    .A(\z80.tv80s.i_tv80_core.F[7] ),
    .B(_2533_));
 sg13g2_a21oi_1 _7622_ (.A1(_0661_),
    .A2(net2172),
    .Y(_3245_),
    .B1(_1804_));
 sg13g2_o21ai_1 _7623_ (.B1(_3245_),
    .Y(_3246_),
    .A1(net2172),
    .A2(_2317_));
 sg13g2_nand4_1 _7624_ (.B(_3081_),
    .C(_3244_),
    .A(_2310_),
    .Y(_3247_),
    .D(_3246_));
 sg13g2_a21oi_1 _7625_ (.A1(_3242_),
    .A2(_3243_),
    .Y(_3248_),
    .B1(_3247_));
 sg13g2_nand2_1 _7626_ (.Y(_3249_),
    .A(_0661_),
    .B(net1818));
 sg13g2_a21oi_1 _7627_ (.A1(_0802_),
    .A2(_3094_),
    .Y(_3250_),
    .B1(net1860));
 sg13g2_a221oi_1 _7628_ (.B2(_3250_),
    .C1(net1795),
    .B1(_3249_),
    .A1(\z80.tv80s.i_tv80_core.I[7] ),
    .Y(_3251_),
    .A2(net1860));
 sg13g2_nor3_1 _7629_ (.A(_3114_),
    .B(_3248_),
    .C(_3251_),
    .Y(_3252_));
 sg13g2_a21oi_1 _7630_ (.A1(net2043),
    .A2(_3114_),
    .Y(_3253_),
    .B1(_3252_));
 sg13g2_o21ai_1 _7631_ (.B1(net1993),
    .Y(_3254_),
    .A1(_2323_),
    .A2(_3064_));
 sg13g2_a21oi_1 _7632_ (.A1(_3064_),
    .A2(_3253_),
    .Y(_3255_),
    .B1(_3254_));
 sg13g2_a21oi_1 _7633_ (.A1(_0666_),
    .A2(net1965),
    .Y(_0496_),
    .B1(_3255_));
 sg13g2_nor2_1 _7634_ (.A(_0023_),
    .B(net1971),
    .Y(_3256_));
 sg13g2_nand3_1 _7635_ (.B(_1116_),
    .C(_3256_),
    .A(_1050_),
    .Y(_3257_));
 sg13g2_mux2_1 _7636_ (.A0(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A1(net614),
    .S(_3257_),
    .X(_0497_));
 sg13g2_mux2_1 _7637_ (.A0(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A1(net610),
    .S(_3257_),
    .X(_0498_));
 sg13g2_mux2_1 _7638_ (.A0(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A1(net604),
    .S(_3257_),
    .X(_0499_));
 sg13g2_mux2_1 _7639_ (.A0(net2146),
    .A1(net618),
    .S(_3257_),
    .X(_0500_));
 sg13g2_mux2_1 _7640_ (.A0(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A1(net615),
    .S(_3257_),
    .X(_0501_));
 sg13g2_mux2_1 _7641_ (.A0(net2145),
    .A1(net613),
    .S(_3257_),
    .X(_0502_));
 sg13g2_mux2_1 _7642_ (.A0(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A1(net608),
    .S(_3257_),
    .X(_0503_));
 sg13g2_mux2_1 _7643_ (.A0(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A1(net633),
    .S(_3257_),
    .X(_0504_));
 sg13g2_nor4_2 _7644_ (.A(_1240_),
    .B(_1515_),
    .C(_1525_),
    .Y(_3258_),
    .D(_1532_));
 sg13g2_nand3_1 _7645_ (.B(net430),
    .C(_0843_),
    .A(net478),
    .Y(_3259_));
 sg13g2_nor2_1 _7646_ (.A(_3258_),
    .B(_3259_),
    .Y(_3260_));
 sg13g2_nor3_1 _7647_ (.A(_2499_),
    .B(_3258_),
    .C(_3259_),
    .Y(_3261_));
 sg13g2_nor2b_1 _7648_ (.A(_1345_),
    .B_N(_2497_),
    .Y(_3262_));
 sg13g2_nand2_1 _7649_ (.Y(_3263_),
    .A(net2144),
    .B(_1522_));
 sg13g2_or4_2 _7650_ (.A(_0946_),
    .B(_1526_),
    .C(_1532_),
    .D(_3263_),
    .X(_3264_));
 sg13g2_o21ai_1 _7651_ (.B1(net2229),
    .Y(_3265_),
    .A1(_1515_),
    .A2(_3264_));
 sg13g2_nand2_1 _7652_ (.Y(_3266_),
    .A(\z80.tv80s.i_tv80_core.ts[2] ),
    .B(_3258_));
 sg13g2_a221oi_1 _7653_ (.B2(net473),
    .C1(_3265_),
    .B1(_3266_),
    .A1(_3261_),
    .Y(_3267_),
    .A2(_3262_));
 sg13g2_a21o_1 _7654_ (.A2(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .A1(net2182),
    .B1(_3267_),
    .X(_0505_));
 sg13g2_nand3_1 _7655_ (.B(_1116_),
    .C(_3256_),
    .A(_1037_),
    .Y(_3268_));
 sg13g2_mux2_1 _7656_ (.A0(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A1(net511),
    .S(_3268_),
    .X(_0506_));
 sg13g2_mux2_1 _7657_ (.A0(_3261_),
    .A1(net596),
    .S(_2498_),
    .X(_0507_));
 sg13g2_and4_2 _7658_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .C(_1755_),
    .D(_1767_),
    .X(_3269_));
 sg13g2_nand4_1 _7659_ (.B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .C(_1755_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .Y(_3270_),
    .D(_1767_));
 sg13g2_nor2_1 _7660_ (.A(net2080),
    .B(_0885_),
    .Y(_3271_));
 sg13g2_nand3_1 _7661_ (.B(_0873_),
    .C(_3271_),
    .A(net1954),
    .Y(_3272_));
 sg13g2_nor3_2 _7662_ (.A(net1892),
    .B(_0872_),
    .C(_2361_),
    .Y(_3273_));
 sg13g2_nor2_1 _7663_ (.A(\z80.tv80s.i_tv80_core.BusB[0] ),
    .B(_3273_),
    .Y(_3274_));
 sg13g2_a21oi_1 _7664_ (.A1(_0782_),
    .A2(_3273_),
    .Y(_3275_),
    .B1(_3274_));
 sg13g2_nor2_2 _7665_ (.A(_0683_),
    .B(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .Y(_3276_));
 sg13g2_nand2b_2 _7666_ (.Y(_3277_),
    .B(\z80.tv80s.i_tv80_core.ts[1] ),
    .A_N(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ));
 sg13g2_a21oi_1 _7667_ (.A1(net1857),
    .A2(_3275_),
    .Y(_3278_),
    .B1(_3277_));
 sg13g2_o21ai_1 _7668_ (.B1(_3278_),
    .Y(_3279_),
    .A1(_0785_),
    .A2(_3272_));
 sg13g2_o21ai_1 _7669_ (.B1(_3279_),
    .Y(_3280_),
    .A1(uio_out[0]),
    .A2(_3276_));
 sg13g2_a21oi_1 _7670_ (.A1(_3270_),
    .A2(_3280_),
    .Y(_3281_),
    .B1(net1968));
 sg13g2_o21ai_1 _7671_ (.B1(_3281_),
    .Y(_3282_),
    .A1(_1831_),
    .A2(net1853));
 sg13g2_o21ai_1 _7672_ (.B1(_3282_),
    .Y(_0508_),
    .A1(_0795_),
    .A2(net1996));
 sg13g2_mux2_1 _7673_ (.A0(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A1(net2027),
    .S(net1852),
    .X(_3283_));
 sg13g2_a21oi_1 _7674_ (.A1(net1856),
    .A2(_3283_),
    .Y(_3284_),
    .B1(_3277_));
 sg13g2_o21ai_1 _7675_ (.B1(_3284_),
    .Y(_3285_),
    .A1(_0786_),
    .A2(net1857));
 sg13g2_o21ai_1 _7676_ (.B1(_3285_),
    .Y(_3286_),
    .A1(uio_out[1]),
    .A2(_3276_));
 sg13g2_a21oi_1 _7677_ (.A1(net1853),
    .A2(_3286_),
    .Y(_3287_),
    .B1(net1968));
 sg13g2_o21ai_1 _7678_ (.B1(_3287_),
    .Y(_3288_),
    .A1(_2005_),
    .A2(net1853));
 sg13g2_o21ai_1 _7679_ (.B1(_3288_),
    .Y(_0509_),
    .A1(_0796_),
    .A2(net1994));
 sg13g2_mux2_1 _7680_ (.A0(\z80.tv80s.i_tv80_core.BusB[2] ),
    .A1(net2028),
    .S(net1852),
    .X(_3289_));
 sg13g2_a21oi_1 _7681_ (.A1(net1857),
    .A2(_3289_),
    .Y(_3290_),
    .B1(_3277_));
 sg13g2_o21ai_1 _7682_ (.B1(_3290_),
    .Y(_3291_),
    .A1(_0787_),
    .A2(net1857));
 sg13g2_o21ai_1 _7683_ (.B1(_3291_),
    .Y(_3292_),
    .A1(uio_out[2]),
    .A2(_3276_));
 sg13g2_a21oi_1 _7684_ (.A1(_3270_),
    .A2(_3292_),
    .Y(_3293_),
    .B1(net1968));
 sg13g2_o21ai_1 _7685_ (.B1(_3293_),
    .Y(_3294_),
    .A1(_2050_),
    .A2(net1853));
 sg13g2_o21ai_1 _7686_ (.B1(_3294_),
    .Y(_0510_),
    .A1(_0797_),
    .A2(net1994));
 sg13g2_nand2_1 _7687_ (.Y(_3295_),
    .A(_0783_),
    .B(net1852));
 sg13g2_o21ai_1 _7688_ (.B1(_3295_),
    .Y(_3296_),
    .A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A2(net1852));
 sg13g2_o21ai_1 _7689_ (.B1(_3276_),
    .Y(_3297_),
    .A1(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A2(net1856));
 sg13g2_a21o_1 _7690_ (.A2(_3296_),
    .A1(net1856),
    .B1(_3297_),
    .X(_3298_));
 sg13g2_a21oi_1 _7691_ (.A1(net496),
    .A2(_3277_),
    .Y(_3299_),
    .B1(_3269_));
 sg13g2_a221oi_1 _7692_ (.B2(_3299_),
    .C1(net1967),
    .B1(_3298_),
    .A1(_2100_),
    .Y(_3300_),
    .A2(_3269_));
 sg13g2_a21o_1 _7693_ (.A2(net1967),
    .A1(net496),
    .B1(_3300_),
    .X(_0511_));
 sg13g2_mux2_1 _7694_ (.A0(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .S(net1852),
    .X(_3301_));
 sg13g2_a21oi_1 _7695_ (.A1(net1857),
    .A2(_3301_),
    .Y(_3302_),
    .B1(_3277_));
 sg13g2_o21ai_1 _7696_ (.B1(_3302_),
    .Y(_3303_),
    .A1(_0782_),
    .A2(net1856));
 sg13g2_o21ai_1 _7697_ (.B1(_3303_),
    .Y(_3304_),
    .A1(net465),
    .A2(_3276_));
 sg13g2_a21oi_1 _7698_ (.A1(net1853),
    .A2(_3304_),
    .Y(_3305_),
    .B1(net1967));
 sg13g2_o21ai_1 _7699_ (.B1(_3305_),
    .Y(_3306_),
    .A1(_2147_),
    .A2(net1853));
 sg13g2_o21ai_1 _7700_ (.B1(_3306_),
    .Y(_0512_),
    .A1(_0792_),
    .A2(net1994));
 sg13g2_nand2b_1 _7701_ (.Y(_3307_),
    .B(net1852),
    .A_N(\z80.tv80s.i_tv80_core.BusB[1] ));
 sg13g2_o21ai_1 _7702_ (.B1(_3307_),
    .Y(_3308_),
    .A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A2(net1852));
 sg13g2_o21ai_1 _7703_ (.B1(_3276_),
    .Y(_3309_),
    .A1(net2027),
    .A2(net1856));
 sg13g2_a21o_1 _7704_ (.A2(_3308_),
    .A1(net1856),
    .B1(_3309_),
    .X(_3310_));
 sg13g2_a21oi_1 _7705_ (.A1(net497),
    .A2(_3277_),
    .Y(_3311_),
    .B1(_3269_));
 sg13g2_a221oi_1 _7706_ (.B2(_3311_),
    .C1(net1967),
    .B1(_3310_),
    .A1(_2219_),
    .Y(_3312_),
    .A2(_3269_));
 sg13g2_a21o_1 _7707_ (.A2(net1967),
    .A1(net497),
    .B1(_3312_),
    .X(_0513_));
 sg13g2_mux2_1 _7708_ (.A0(_0787_),
    .A1(_0784_),
    .S(_3273_),
    .X(_3313_));
 sg13g2_o21ai_1 _7709_ (.B1(_3276_),
    .Y(_3314_),
    .A1(net2028),
    .A2(net1857));
 sg13g2_a21o_1 _7710_ (.A2(_3313_),
    .A1(net1857),
    .B1(_3314_),
    .X(_3315_));
 sg13g2_a21oi_1 _7711_ (.A1(net487),
    .A2(_3277_),
    .Y(_3316_),
    .B1(_3269_));
 sg13g2_a221oi_1 _7712_ (.B2(_3316_),
    .C1(net1968),
    .B1(_3315_),
    .A1(_2270_),
    .Y(_3317_),
    .A2(_3269_));
 sg13g2_a21o_1 _7713_ (.A2(net1967),
    .A1(net487),
    .B1(_3317_),
    .X(_0514_));
 sg13g2_mux2_1 _7714_ (.A0(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .S(net1852),
    .X(_3318_));
 sg13g2_a21oi_1 _7715_ (.A1(net1856),
    .A2(_3318_),
    .Y(_3319_),
    .B1(_3277_));
 sg13g2_o21ai_1 _7716_ (.B1(_3319_),
    .Y(_3320_),
    .A1(_0783_),
    .A2(net1856));
 sg13g2_o21ai_1 _7717_ (.B1(_3320_),
    .Y(_3321_),
    .A1(net475),
    .A2(_3276_));
 sg13g2_a21oi_1 _7718_ (.A1(net1853),
    .A2(_3321_),
    .Y(_3322_),
    .B1(net1968));
 sg13g2_o21ai_1 _7719_ (.B1(_3322_),
    .Y(_3323_),
    .A1(_2323_),
    .A2(net1853));
 sg13g2_o21ai_1 _7720_ (.B1(_3323_),
    .Y(_0515_),
    .A1(_0793_),
    .A2(net1994));
 sg13g2_xnor2_1 _7721_ (.Y(_3324_),
    .A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .B(_3105_));
 sg13g2_nand2b_1 _7722_ (.Y(_3325_),
    .B(net1905),
    .A_N(\z80.tv80s.i_tv80_core.ACC[0] ));
 sg13g2_o21ai_1 _7723_ (.B1(_3325_),
    .Y(_3326_),
    .A1(\z80.tv80s.i_tv80_core.Ap[0] ),
    .A2(net1818));
 sg13g2_a21oi_1 _7724_ (.A1(net1820),
    .A2(_3324_),
    .Y(_3327_),
    .B1(_3326_));
 sg13g2_nor4_2 _7725_ (.A(_0790_),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .C(_0228_),
    .Y(_3328_),
    .D(_3061_));
 sg13g2_a22oi_1 _7726_ (.Y(_3329_),
    .B1(net1877),
    .B2(\z80.tv80s.i_tv80_core.R[0] ),
    .A2(net1879),
    .A1(\z80.tv80s.i_tv80_core.I[0] ));
 sg13g2_a21oi_1 _7727_ (.A1(net1859),
    .A2(_3329_),
    .Y(_3330_),
    .B1(net1848));
 sg13g2_o21ai_1 _7728_ (.B1(_3330_),
    .Y(_3331_),
    .A1(net1859),
    .A2(_3327_));
 sg13g2_a21oi_1 _7729_ (.A1(_1831_),
    .A2(_3328_),
    .Y(_3332_),
    .B1(net1973));
 sg13g2_a22oi_1 _7730_ (.Y(_3333_),
    .B1(_3331_),
    .B2(_3332_),
    .A2(net1960),
    .A1(net339));
 sg13g2_inv_1 _7731_ (.Y(_0516_),
    .A(net340));
 sg13g2_xnor2_1 _7732_ (.Y(_3334_),
    .A(\z80.tv80s.i_tv80_core.ACC[1] ),
    .B(net1680));
 sg13g2_nand2b_1 _7733_ (.Y(_3335_),
    .B(net1908),
    .A_N(\z80.tv80s.i_tv80_core.ACC[1] ));
 sg13g2_o21ai_1 _7734_ (.B1(_3335_),
    .Y(_3336_),
    .A1(\z80.tv80s.i_tv80_core.Ap[1] ),
    .A2(net1818));
 sg13g2_a21oi_1 _7735_ (.A1(net1820),
    .A2(_3334_),
    .Y(_3337_),
    .B1(_3336_));
 sg13g2_a22oi_1 _7736_ (.Y(_3338_),
    .B1(net1877),
    .B2(\z80.tv80s.i_tv80_core.R[1] ),
    .A2(net1879),
    .A1(\z80.tv80s.i_tv80_core.I[1] ));
 sg13g2_a21oi_1 _7737_ (.A1(net1858),
    .A2(_3338_),
    .Y(_3339_),
    .B1(net1848));
 sg13g2_o21ai_1 _7738_ (.B1(_3339_),
    .Y(_3340_),
    .A1(net1858),
    .A2(_3337_));
 sg13g2_a21oi_1 _7739_ (.A1(_2005_),
    .A2(net1848),
    .Y(_3341_),
    .B1(net1960));
 sg13g2_a22oi_1 _7740_ (.Y(_3342_),
    .B1(_3340_),
    .B2(_3341_),
    .A2(net1960),
    .A1(net315));
 sg13g2_inv_1 _7741_ (.Y(_0517_),
    .A(net316));
 sg13g2_xnor2_1 _7742_ (.Y(_3343_),
    .A(\z80.tv80s.i_tv80_core.ACC[2] ),
    .B(net1680));
 sg13g2_nand2b_1 _7743_ (.Y(_3344_),
    .B(net1905),
    .A_N(\z80.tv80s.i_tv80_core.ACC[2] ));
 sg13g2_o21ai_1 _7744_ (.B1(_3344_),
    .Y(_3345_),
    .A1(\z80.tv80s.i_tv80_core.Ap[2] ),
    .A2(net1818));
 sg13g2_a21oi_1 _7745_ (.A1(net1820),
    .A2(_3343_),
    .Y(_3346_),
    .B1(_3345_));
 sg13g2_a22oi_1 _7746_ (.Y(_3347_),
    .B1(net1877),
    .B2(\z80.tv80s.i_tv80_core.R[2] ),
    .A2(net1879),
    .A1(\z80.tv80s.i_tv80_core.I[2] ));
 sg13g2_a21oi_1 _7747_ (.A1(net1858),
    .A2(_3347_),
    .Y(_3348_),
    .B1(net1847));
 sg13g2_o21ai_1 _7748_ (.B1(_3348_),
    .Y(_3349_),
    .A1(net1858),
    .A2(_3346_));
 sg13g2_a21oi_1 _7749_ (.A1(_2050_),
    .A2(net1847),
    .Y(_3350_),
    .B1(net1959));
 sg13g2_a22oi_1 _7750_ (.Y(_3351_),
    .B1(_3349_),
    .B2(_3350_),
    .A2(net1959),
    .A1(net336));
 sg13g2_inv_1 _7751_ (.Y(_0518_),
    .A(net337));
 sg13g2_xnor2_1 _7752_ (.Y(_3352_),
    .A(net2146),
    .B(net1680));
 sg13g2_nand2b_1 _7753_ (.Y(_3353_),
    .B(net1905),
    .A_N(net2146));
 sg13g2_o21ai_1 _7754_ (.B1(_3353_),
    .Y(_3354_),
    .A1(\z80.tv80s.i_tv80_core.Ap[3] ),
    .A2(net1818));
 sg13g2_a21oi_1 _7755_ (.A1(net1820),
    .A2(_3352_),
    .Y(_3355_),
    .B1(_3354_));
 sg13g2_a22oi_1 _7756_ (.Y(_3356_),
    .B1(net1877),
    .B2(\z80.tv80s.i_tv80_core.R[3] ),
    .A2(net1879),
    .A1(\z80.tv80s.i_tv80_core.I[3] ));
 sg13g2_a21oi_1 _7757_ (.A1(net1859),
    .A2(_3356_),
    .Y(_3357_),
    .B1(net1848));
 sg13g2_o21ai_1 _7758_ (.B1(_3357_),
    .Y(_3358_),
    .A1(net1858),
    .A2(_3355_));
 sg13g2_a21oi_1 _7759_ (.A1(_2101_),
    .A2(net1847),
    .Y(_3359_),
    .B1(net1959));
 sg13g2_a22oi_1 _7760_ (.Y(_3360_),
    .B1(_3358_),
    .B2(_3359_),
    .A2(net1959),
    .A1(net232));
 sg13g2_inv_1 _7761_ (.Y(_0519_),
    .A(net233));
 sg13g2_xnor2_1 _7762_ (.Y(_3361_),
    .A(\z80.tv80s.i_tv80_core.ACC[4] ),
    .B(net1680));
 sg13g2_nand2b_1 _7763_ (.Y(_3362_),
    .B(net1905),
    .A_N(\z80.tv80s.i_tv80_core.ACC[4] ));
 sg13g2_o21ai_1 _7764_ (.B1(_3362_),
    .Y(_3363_),
    .A1(\z80.tv80s.i_tv80_core.Ap[4] ),
    .A2(net1818));
 sg13g2_a21oi_1 _7765_ (.A1(net1820),
    .A2(_3361_),
    .Y(_3364_),
    .B1(_3363_));
 sg13g2_a22oi_1 _7766_ (.Y(_3365_),
    .B1(net1877),
    .B2(\z80.tv80s.i_tv80_core.R[4] ),
    .A2(net1879),
    .A1(\z80.tv80s.i_tv80_core.I[4] ));
 sg13g2_a21oi_1 _7767_ (.A1(net1858),
    .A2(_3365_),
    .Y(_3366_),
    .B1(net1847));
 sg13g2_o21ai_1 _7768_ (.B1(_3366_),
    .Y(_3367_),
    .A1(net1858),
    .A2(_3364_));
 sg13g2_a21oi_1 _7769_ (.A1(_2147_),
    .A2(net1847),
    .Y(_3368_),
    .B1(net1960));
 sg13g2_a22oi_1 _7770_ (.Y(_3369_),
    .B1(_3367_),
    .B2(_3368_),
    .A2(net1959),
    .A1(net381));
 sg13g2_inv_1 _7771_ (.Y(_0520_),
    .A(net382));
 sg13g2_xnor2_1 _7772_ (.Y(_3370_),
    .A(net2145),
    .B(net1680));
 sg13g2_nand2b_1 _7773_ (.Y(_3371_),
    .B(net1905),
    .A_N(net2145));
 sg13g2_o21ai_1 _7774_ (.B1(_3371_),
    .Y(_3372_),
    .A1(\z80.tv80s.i_tv80_core.Ap[5] ),
    .A2(net1818));
 sg13g2_a21oi_1 _7775_ (.A1(net1820),
    .A2(_3370_),
    .Y(_3373_),
    .B1(_3372_));
 sg13g2_a22oi_1 _7776_ (.Y(_3374_),
    .B1(net1877),
    .B2(\z80.tv80s.i_tv80_core.R[5] ),
    .A2(net1879),
    .A1(\z80.tv80s.i_tv80_core.I[5] ));
 sg13g2_a21oi_1 _7777_ (.A1(net1859),
    .A2(_3374_),
    .Y(_3375_),
    .B1(net1848));
 sg13g2_o21ai_1 _7778_ (.B1(_3375_),
    .Y(_3376_),
    .A1(net1858),
    .A2(_3373_));
 sg13g2_a21oi_1 _7779_ (.A1(_2220_),
    .A2(net1847),
    .Y(_3377_),
    .B1(net1959));
 sg13g2_a22oi_1 _7780_ (.Y(_3378_),
    .B1(_3376_),
    .B2(_3377_),
    .A2(net1959),
    .A1(net277));
 sg13g2_inv_1 _7781_ (.Y(_0521_),
    .A(net278));
 sg13g2_xnor2_1 _7782_ (.Y(_3379_),
    .A(\z80.tv80s.i_tv80_core.ACC[6] ),
    .B(net1680));
 sg13g2_nand2b_1 _7783_ (.Y(_3380_),
    .B(net1905),
    .A_N(\z80.tv80s.i_tv80_core.ACC[6] ));
 sg13g2_o21ai_1 _7784_ (.B1(_3380_),
    .Y(_3381_),
    .A1(\z80.tv80s.i_tv80_core.Ap[6] ),
    .A2(net1818));
 sg13g2_a21oi_1 _7785_ (.A1(net1820),
    .A2(_3379_),
    .Y(_3382_),
    .B1(_3381_));
 sg13g2_a22oi_1 _7786_ (.Y(_3383_),
    .B1(net1877),
    .B2(\z80.tv80s.i_tv80_core.R[6] ),
    .A2(net1879),
    .A1(\z80.tv80s.i_tv80_core.I[6] ));
 sg13g2_a21oi_1 _7787_ (.A1(net1859),
    .A2(_3383_),
    .Y(_3384_),
    .B1(net1847));
 sg13g2_o21ai_1 _7788_ (.B1(_3384_),
    .Y(_3385_),
    .A1(net1859),
    .A2(_3382_));
 sg13g2_a21oi_1 _7789_ (.A1(_2271_),
    .A2(net1847),
    .Y(_3386_),
    .B1(net1962));
 sg13g2_a22oi_1 _7790_ (.Y(_3387_),
    .B1(_3385_),
    .B2(_3386_),
    .A2(net1959),
    .A1(net282));
 sg13g2_inv_1 _7791_ (.Y(_0522_),
    .A(net283));
 sg13g2_xnor2_1 _7792_ (.Y(_3388_),
    .A(\z80.tv80s.i_tv80_core.ACC[7] ),
    .B(net1680));
 sg13g2_nand2b_1 _7793_ (.Y(_3389_),
    .B(net1905),
    .A_N(\z80.tv80s.i_tv80_core.ACC[7] ));
 sg13g2_o21ai_1 _7794_ (.B1(_3389_),
    .Y(_3390_),
    .A1(\z80.tv80s.i_tv80_core.Ap[7] ),
    .A2(net1819));
 sg13g2_a21oi_1 _7795_ (.A1(net1821),
    .A2(_3388_),
    .Y(_3391_),
    .B1(_3390_));
 sg13g2_a22oi_1 _7796_ (.Y(_3392_),
    .B1(net1880),
    .B2(\z80.tv80s.i_tv80_core.I[7] ),
    .A2(\z80.tv80s.i_tv80_core.R[7] ),
    .A1(net2079));
 sg13g2_a21oi_1 _7797_ (.A1(net1860),
    .A2(_3392_),
    .Y(_3393_),
    .B1(net1848));
 sg13g2_o21ai_1 _7798_ (.B1(_3393_),
    .Y(_3394_),
    .A1(net1860),
    .A2(_3391_));
 sg13g2_a21oi_1 _7799_ (.A1(_2323_),
    .A2(net1848),
    .Y(_3395_),
    .B1(net1960));
 sg13g2_a22oi_1 _7800_ (.Y(_3396_),
    .B1(_3394_),
    .B2(_3395_),
    .A2(net1960),
    .A1(net249));
 sg13g2_inv_1 _7801_ (.Y(_0523_),
    .A(net250));
 sg13g2_o21ai_1 _7802_ (.B1(_3262_),
    .Y(_3397_),
    .A1(_2499_),
    .A2(_3260_));
 sg13g2_nand2b_1 _7803_ (.Y(_3398_),
    .B(net478),
    .A_N(\z80.tv80s.i_tv80_core.ts[2] ));
 sg13g2_a221oi_1 _7804_ (.B2(_0681_),
    .C1(\z80.tv80s.i_tv80_core.IntE ),
    .B1(_3258_),
    .A1(_1188_),
    .Y(_3399_),
    .A2(_1685_));
 sg13g2_o21ai_1 _7805_ (.B1(\z80.tv80s.i_tv80_core.ts[2] ),
    .Y(_3400_),
    .A1(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .A2(_2572_));
 sg13g2_o21ai_1 _7806_ (.B1(_3398_),
    .Y(_3401_),
    .A1(_3399_),
    .A2(_3400_));
 sg13g2_nand3b_1 _7807_ (.B(_3397_),
    .C(_3401_),
    .Y(_3402_),
    .A_N(_3265_));
 sg13g2_o21ai_1 _7808_ (.B1(_3402_),
    .Y(_0524_),
    .A1(net2227),
    .A2(_0806_));
 sg13g2_nand2_1 _7809_ (.Y(_3403_),
    .A(net1993),
    .B(_3094_));
 sg13g2_nand2_1 _7810_ (.Y(_3404_),
    .A(net230),
    .B(net1777));
 sg13g2_o21ai_1 _7811_ (.B1(_3404_),
    .Y(_0525_),
    .A1(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A2(net1777));
 sg13g2_nand2_1 _7812_ (.Y(_3405_),
    .A(net221),
    .B(net1777));
 sg13g2_o21ai_1 _7813_ (.B1(_3405_),
    .Y(_0526_),
    .A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(net1777));
 sg13g2_nand2_1 _7814_ (.Y(_3406_),
    .A(net215),
    .B(net1776));
 sg13g2_o21ai_1 _7815_ (.B1(_3406_),
    .Y(_0527_),
    .A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(net1776));
 sg13g2_nand2_1 _7816_ (.Y(_3407_),
    .A(net210),
    .B(net1776));
 sg13g2_o21ai_1 _7817_ (.B1(_3407_),
    .Y(_0528_),
    .A1(net2146),
    .A2(net1776));
 sg13g2_nand2_1 _7818_ (.Y(_3408_),
    .A(net213),
    .B(net1776));
 sg13g2_o21ai_1 _7819_ (.B1(_3408_),
    .Y(_0529_),
    .A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(net1776));
 sg13g2_nand2_1 _7820_ (.Y(_3409_),
    .A(net195),
    .B(net1776));
 sg13g2_o21ai_1 _7821_ (.B1(_3409_),
    .Y(_0530_),
    .A1(net2145),
    .A2(net1776));
 sg13g2_nand2_1 _7822_ (.Y(_3410_),
    .A(net217),
    .B(net1777));
 sg13g2_o21ai_1 _7823_ (.B1(_3410_),
    .Y(_0531_),
    .A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(net1777));
 sg13g2_nand2_1 _7824_ (.Y(_3411_),
    .A(net211),
    .B(net1780));
 sg13g2_o21ai_1 _7825_ (.B1(_3411_),
    .Y(_0532_),
    .A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(net1780));
 sg13g2_nand2_1 _7826_ (.Y(_3412_),
    .A(net205),
    .B(net1778));
 sg13g2_o21ai_1 _7827_ (.B1(_3412_),
    .Y(_0533_),
    .A1(net2151),
    .A2(net1778));
 sg13g2_nand2_1 _7828_ (.Y(_3413_),
    .A(net201),
    .B(net1778));
 sg13g2_o21ai_1 _7829_ (.B1(_3413_),
    .Y(_0534_),
    .A1(net2150),
    .A2(net1778));
 sg13g2_nand2_1 _7830_ (.Y(_3414_),
    .A(net235),
    .B(net1779));
 sg13g2_o21ai_1 _7831_ (.B1(_3414_),
    .Y(_0535_),
    .A1(net2147),
    .A2(net1779));
 sg13g2_nand2_1 _7832_ (.Y(_3415_),
    .A(net207),
    .B(net1779));
 sg13g2_o21ai_1 _7833_ (.B1(_3415_),
    .Y(_0536_),
    .A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(net1779));
 sg13g2_nand2_1 _7834_ (.Y(_3416_),
    .A(net223),
    .B(net1778));
 sg13g2_o21ai_1 _7835_ (.B1(_3416_),
    .Y(_0537_),
    .A1(\z80.tv80s.i_tv80_core.F[4] ),
    .A2(net1778));
 sg13g2_nand2_1 _7836_ (.Y(_3417_),
    .A(net196),
    .B(net1779));
 sg13g2_o21ai_1 _7837_ (.B1(_3417_),
    .Y(_0538_),
    .A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(net1779));
 sg13g2_nand2_1 _7838_ (.Y(_3418_),
    .A(net203),
    .B(net1780));
 sg13g2_o21ai_1 _7839_ (.B1(_3418_),
    .Y(_0539_),
    .A1(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(net1780));
 sg13g2_nand2_1 _7840_ (.Y(_3419_),
    .A(net198),
    .B(net1778));
 sg13g2_o21ai_1 _7841_ (.B1(_3419_),
    .Y(_0540_),
    .A1(\z80.tv80s.i_tv80_core.F[7] ),
    .A2(net1778));
 sg13g2_a21oi_1 _7842_ (.A1(net2123),
    .A2(\z80.tv80s.i_tv80_core.ts[4] ),
    .Y(_3420_),
    .B1(_0820_));
 sg13g2_nor2_1 _7843_ (.A(_1750_),
    .B(_3420_),
    .Y(_3421_));
 sg13g2_or2_1 _7844_ (.X(_3422_),
    .B(_3420_),
    .A(_1750_));
 sg13g2_nand2_1 _7845_ (.Y(_3423_),
    .A(net2142),
    .B(_2593_));
 sg13g2_nand2b_1 _7846_ (.Y(_3424_),
    .B(net2142),
    .A_N(net2051));
 sg13g2_o21ai_1 _7847_ (.B1(_3424_),
    .Y(_3425_),
    .A1(net2142),
    .A2(\z80.tv80s.i_tv80_core.SP[0] ));
 sg13g2_nand2b_1 _7848_ (.Y(_3426_),
    .B(_3423_),
    .A_N(_3425_));
 sg13g2_o21ai_1 _7849_ (.B1(_3426_),
    .Y(_3427_),
    .A1(net2051),
    .A2(_3423_));
 sg13g2_a21oi_1 _7850_ (.A1(\z80.tv80s.i_tv80_core.SP[0] ),
    .A2(net1772),
    .Y(_3428_),
    .B1(net1753));
 sg13g2_o21ai_1 _7851_ (.B1(_3428_),
    .Y(_3429_),
    .A1(net1772),
    .A2(_3427_));
 sg13g2_a21oi_1 _7852_ (.A1(net1753),
    .A2(_2593_),
    .Y(_3430_),
    .B1(net1909));
 sg13g2_nor2_2 _7853_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .B(_3062_),
    .Y(_3431_));
 sg13g2_and2_1 _7854_ (.A(_1767_),
    .B(_3431_),
    .X(_3432_));
 sg13g2_nand2_2 _7855_ (.Y(_3433_),
    .A(_1767_),
    .B(_3431_));
 sg13g2_a22oi_1 _7856_ (.Y(_3434_),
    .B1(_3429_),
    .B2(_3430_),
    .A2(net1909),
    .A1(\z80.tv80s.i_tv80_core.SP[0] ));
 sg13g2_a21oi_1 _7857_ (.A1(_1831_),
    .A2(net1851),
    .Y(_3435_),
    .B1(net1963));
 sg13g2_o21ai_1 _7858_ (.B1(_3435_),
    .Y(_3436_),
    .A1(net1851),
    .A2(_3434_));
 sg13g2_o21ai_1 _7859_ (.B1(_3436_),
    .Y(_0541_),
    .A1(_0660_),
    .A2(net1994));
 sg13g2_nor2_2 _7860_ (.A(net2138),
    .B(_1847_),
    .Y(_3437_));
 sg13g2_or3_2 _7861_ (.A(net2143),
    .B(_1836_),
    .C(_1846_),
    .X(_3438_));
 sg13g2_nand2_1 _7862_ (.Y(_3439_),
    .A(net2143),
    .B(_0172_));
 sg13g2_nand2_1 _7863_ (.Y(_3440_),
    .A(_3438_),
    .B(_3439_));
 sg13g2_nor2_1 _7864_ (.A(net2141),
    .B(\z80.tv80s.i_tv80_core.SP[1] ),
    .Y(_3441_));
 sg13g2_a21oi_1 _7865_ (.A1(net2141),
    .A2(_2650_),
    .Y(_3442_),
    .B1(_3441_));
 sg13g2_nand3_1 _7866_ (.B(_3439_),
    .C(_3442_),
    .A(_3438_),
    .Y(_3443_));
 sg13g2_a21oi_1 _7867_ (.A1(_3438_),
    .A2(_3439_),
    .Y(_3444_),
    .B1(_3442_));
 sg13g2_xor2_1 _7868_ (.B(_3442_),
    .A(_3440_),
    .X(_3445_));
 sg13g2_xnor2_1 _7869_ (.Y(_3446_),
    .A(_3426_),
    .B(_3445_));
 sg13g2_a21oi_1 _7870_ (.A1(\z80.tv80s.i_tv80_core.SP[1] ),
    .A2(net1772),
    .Y(_3447_),
    .B1(net1753));
 sg13g2_o21ai_1 _7871_ (.B1(_3447_),
    .Y(_3448_),
    .A1(net1772),
    .A2(_3446_));
 sg13g2_a21oi_1 _7872_ (.A1(net1753),
    .A2(_2650_),
    .Y(_3449_),
    .B1(net1907));
 sg13g2_a22oi_1 _7873_ (.Y(_3450_),
    .B1(_3448_),
    .B2(_3449_),
    .A2(net1907),
    .A1(\z80.tv80s.i_tv80_core.SP[1] ));
 sg13g2_o21ai_1 _7874_ (.B1(net1984),
    .Y(_3451_),
    .A1(_2005_),
    .A2(_3433_));
 sg13g2_a21oi_1 _7875_ (.A1(_3433_),
    .A2(_3450_),
    .Y(_3452_),
    .B1(_3451_));
 sg13g2_a21oi_1 _7876_ (.A1(_0659_),
    .A2(net1964),
    .Y(_0542_),
    .B1(_3452_));
 sg13g2_o21ai_1 _7877_ (.B1(_3438_),
    .Y(_3453_),
    .A1(_0682_),
    .A2(_0764_));
 sg13g2_mux2_1 _7878_ (.A0(\z80.tv80s.i_tv80_core.SP[2] ),
    .A1(_2673_),
    .S(net2141),
    .X(_3454_));
 sg13g2_nor2b_1 _7879_ (.A(_3453_),
    .B_N(_3454_),
    .Y(_3455_));
 sg13g2_xnor2_1 _7880_ (.Y(_3456_),
    .A(_3453_),
    .B(_3454_));
 sg13g2_o21ai_1 _7881_ (.B1(_3443_),
    .Y(_3457_),
    .A1(_3426_),
    .A2(_3444_));
 sg13g2_xnor2_1 _7882_ (.Y(_3458_),
    .A(_3456_),
    .B(_3457_));
 sg13g2_a21oi_1 _7883_ (.A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .A2(net1771),
    .Y(_3459_),
    .B1(net1753));
 sg13g2_o21ai_1 _7884_ (.B1(_3459_),
    .Y(_3460_),
    .A1(net1771),
    .A2(_3458_));
 sg13g2_o21ai_1 _7885_ (.B1(_3460_),
    .Y(_3461_),
    .A1(net1752),
    .A2(_2673_));
 sg13g2_a21oi_1 _7886_ (.A1(net1899),
    .A2(_3461_),
    .Y(_3462_),
    .B1(net1851));
 sg13g2_o21ai_1 _7887_ (.B1(_3462_),
    .Y(_3463_),
    .A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .A2(net1899));
 sg13g2_a21oi_1 _7888_ (.A1(_2050_),
    .A2(_3432_),
    .Y(_3464_),
    .B1(net1963));
 sg13g2_a22oi_1 _7889_ (.Y(_3465_),
    .B1(_3463_),
    .B2(_3464_),
    .A2(net1963),
    .A1(net252));
 sg13g2_inv_1 _7890_ (.Y(_0543_),
    .A(net253));
 sg13g2_a21oi_1 _7891_ (.A1(net2140),
    .A2(_0178_),
    .Y(_3466_),
    .B1(_3437_));
 sg13g2_nor2_1 _7892_ (.A(net2141),
    .B(\z80.tv80s.i_tv80_core.SP[3] ),
    .Y(_3467_));
 sg13g2_a21oi_1 _7893_ (.A1(net2141),
    .A2(_2700_),
    .Y(_3468_),
    .B1(_3467_));
 sg13g2_nand2_1 _7894_ (.Y(_3469_),
    .A(_3466_),
    .B(_3468_));
 sg13g2_xnor2_1 _7895_ (.Y(_3470_),
    .A(_3466_),
    .B(_3468_));
 sg13g2_a21oi_1 _7896_ (.A1(_3456_),
    .A2(_3457_),
    .Y(_3471_),
    .B1(_3455_));
 sg13g2_xor2_1 _7897_ (.B(_3471_),
    .A(_3470_),
    .X(_3472_));
 sg13g2_nand2_1 _7898_ (.Y(_3473_),
    .A(net1774),
    .B(_3472_));
 sg13g2_a21oi_1 _7899_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(net1771),
    .Y(_3474_),
    .B1(net1753));
 sg13g2_a22oi_1 _7900_ (.Y(_3475_),
    .B1(_3473_),
    .B2(_3474_),
    .A2(_2700_),
    .A1(net1754));
 sg13g2_nor2_1 _7901_ (.A(net1907),
    .B(_3475_),
    .Y(_3476_));
 sg13g2_o21ai_1 _7902_ (.B1(_3433_),
    .Y(_3477_),
    .A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(net1897));
 sg13g2_a21oi_1 _7903_ (.A1(_2101_),
    .A2(net1851),
    .Y(_3478_),
    .B1(net1961));
 sg13g2_o21ai_1 _7904_ (.B1(_3478_),
    .Y(_3479_),
    .A1(_3476_),
    .A2(_3477_));
 sg13g2_o21ai_1 _7905_ (.B1(_3479_),
    .Y(_0544_),
    .A1(_0658_),
    .A2(net1984));
 sg13g2_a21oi_1 _7906_ (.A1(net2138),
    .A2(_0181_),
    .Y(_3480_),
    .B1(_3437_));
 sg13g2_mux2_1 _7907_ (.A0(\z80.tv80s.i_tv80_core.SP[4] ),
    .A1(_2727_),
    .S(net2141),
    .X(_3481_));
 sg13g2_and2_1 _7908_ (.A(_3480_),
    .B(_3481_),
    .X(_3482_));
 sg13g2_xnor2_1 _7909_ (.Y(_3483_),
    .A(_3480_),
    .B(_3481_));
 sg13g2_inv_1 _7910_ (.Y(_3484_),
    .A(_3483_));
 sg13g2_o21ai_1 _7911_ (.B1(_3469_),
    .Y(_3485_),
    .A1(_3470_),
    .A2(_3471_));
 sg13g2_xnor2_1 _7912_ (.Y(_3486_),
    .A(_3484_),
    .B(_3485_));
 sg13g2_o21ai_1 _7913_ (.B1(net1752),
    .Y(_3487_),
    .A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(net1775));
 sg13g2_a21o_1 _7914_ (.A2(_3486_),
    .A1(net1774),
    .B1(_3487_),
    .X(_3488_));
 sg13g2_a21oi_1 _7915_ (.A1(net1753),
    .A2(_2727_),
    .Y(_3489_),
    .B1(net1910));
 sg13g2_a21oi_1 _7916_ (.A1(_3488_),
    .A2(_3489_),
    .Y(_3490_),
    .B1(net1851));
 sg13g2_o21ai_1 _7917_ (.B1(_3490_),
    .Y(_3491_),
    .A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(net1898));
 sg13g2_a21oi_1 _7918_ (.A1(_2147_),
    .A2(net1851),
    .Y(_3492_),
    .B1(net1962));
 sg13g2_a22oi_1 _7919_ (.Y(_3493_),
    .B1(_3491_),
    .B2(_3492_),
    .A2(net1964),
    .A1(net264));
 sg13g2_inv_1 _7920_ (.Y(_0545_),
    .A(net265));
 sg13g2_nand2_1 _7921_ (.Y(_3494_),
    .A(net191),
    .B(net1975));
 sg13g2_a21oi_1 _7922_ (.A1(net2140),
    .A2(_0184_),
    .Y(_3495_),
    .B1(_3437_));
 sg13g2_nor2_1 _7923_ (.A(net2140),
    .B(\z80.tv80s.i_tv80_core.SP[5] ),
    .Y(_3496_));
 sg13g2_a21oi_1 _7924_ (.A1(net2141),
    .A2(_2752_),
    .Y(_3497_),
    .B1(_3496_));
 sg13g2_nand2_1 _7925_ (.Y(_3498_),
    .A(_3495_),
    .B(_3497_));
 sg13g2_xnor2_1 _7926_ (.Y(_3499_),
    .A(_3495_),
    .B(_3497_));
 sg13g2_a21oi_1 _7927_ (.A1(_3484_),
    .A2(_3485_),
    .Y(_3500_),
    .B1(_3482_));
 sg13g2_xnor2_1 _7928_ (.Y(_3501_),
    .A(_3499_),
    .B(_3500_));
 sg13g2_o21ai_1 _7929_ (.B1(net1752),
    .Y(_3502_),
    .A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(net1774));
 sg13g2_a21o_1 _7930_ (.A2(_3501_),
    .A1(net1774),
    .B1(_3502_),
    .X(_3503_));
 sg13g2_a21oi_1 _7931_ (.A1(net1754),
    .A2(_2753_),
    .Y(_3504_),
    .B1(net1909));
 sg13g2_o21ai_1 _7932_ (.B1(_3433_),
    .Y(_3505_),
    .A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(net1898));
 sg13g2_a21oi_1 _7933_ (.A1(_3503_),
    .A2(_3504_),
    .Y(_3506_),
    .B1(_3505_));
 sg13g2_o21ai_1 _7934_ (.B1(net1985),
    .Y(_3507_),
    .A1(_2219_),
    .A2(_3433_));
 sg13g2_o21ai_1 _7935_ (.B1(_3494_),
    .Y(_0546_),
    .A1(_3506_),
    .A2(_3507_));
 sg13g2_nand2_1 _7936_ (.Y(_3508_),
    .A(net240),
    .B(net1964));
 sg13g2_a21o_1 _7937_ (.A2(_0187_),
    .A1(net2138),
    .B1(_3437_),
    .X(_3509_));
 sg13g2_nor2_1 _7938_ (.A(net2140),
    .B(\z80.tv80s.i_tv80_core.SP[6] ),
    .Y(_3510_));
 sg13g2_a21oi_1 _7939_ (.A1(net2140),
    .A2(_2780_),
    .Y(_3511_),
    .B1(_3510_));
 sg13g2_nand2b_1 _7940_ (.Y(_3512_),
    .B(_3511_),
    .A_N(_3509_));
 sg13g2_inv_1 _7941_ (.Y(_3513_),
    .A(_3512_));
 sg13g2_xnor2_1 _7942_ (.Y(_3514_),
    .A(_3509_),
    .B(_3511_));
 sg13g2_o21ai_1 _7943_ (.B1(_3498_),
    .Y(_3515_),
    .A1(_3499_),
    .A2(_3500_));
 sg13g2_xnor2_1 _7944_ (.Y(_3516_),
    .A(_3514_),
    .B(_3515_));
 sg13g2_o21ai_1 _7945_ (.B1(net1752),
    .Y(_3517_),
    .A1(\z80.tv80s.i_tv80_core.SP[6] ),
    .A2(net1774));
 sg13g2_a21o_1 _7946_ (.A2(_3516_),
    .A1(net1774),
    .B1(_3517_),
    .X(_3518_));
 sg13g2_a21oi_1 _7947_ (.A1(net1753),
    .A2(_2781_),
    .Y(_3519_),
    .B1(net1909));
 sg13g2_o21ai_1 _7948_ (.B1(_3433_),
    .Y(_3520_),
    .A1(\z80.tv80s.i_tv80_core.SP[6] ),
    .A2(net1898));
 sg13g2_a21oi_1 _7949_ (.A1(_3518_),
    .A2(_3519_),
    .Y(_3521_),
    .B1(_3520_));
 sg13g2_o21ai_1 _7950_ (.B1(net1984),
    .Y(_3522_),
    .A1(_2270_),
    .A2(_3433_));
 sg13g2_o21ai_1 _7951_ (.B1(_3508_),
    .Y(_0547_),
    .A1(_3521_),
    .A2(_3522_));
 sg13g2_a21oi_1 _7952_ (.A1(_3514_),
    .A2(_3515_),
    .Y(_3523_),
    .B1(_3513_));
 sg13g2_a21oi_1 _7953_ (.A1(net2138),
    .A2(_0190_),
    .Y(_3524_),
    .B1(_3437_));
 sg13g2_a21o_2 _7954_ (.A2(_0190_),
    .A1(net2138),
    .B1(_3437_),
    .X(_3525_));
 sg13g2_nor2_1 _7955_ (.A(net2138),
    .B(\z80.tv80s.i_tv80_core.SP[7] ),
    .Y(_3526_));
 sg13g2_a21oi_2 _7956_ (.B1(_3526_),
    .Y(_3527_),
    .A2(_2809_),
    .A1(net2139));
 sg13g2_nor2_1 _7957_ (.A(net1770),
    .B(_3527_),
    .Y(_3528_));
 sg13g2_xnor2_1 _7958_ (.Y(_3529_),
    .A(net1770),
    .B(_3527_));
 sg13g2_xnor2_1 _7959_ (.Y(_3530_),
    .A(_3523_),
    .B(_3529_));
 sg13g2_o21ai_1 _7960_ (.B1(net1750),
    .Y(_3531_),
    .A1(\z80.tv80s.i_tv80_core.SP[7] ),
    .A2(net1774));
 sg13g2_a21oi_1 _7961_ (.A1(net1774),
    .A2(_3530_),
    .Y(_3532_),
    .B1(_3531_));
 sg13g2_o21ai_1 _7962_ (.B1(net1898),
    .Y(_3533_),
    .A1(net1751),
    .A2(_2809_));
 sg13g2_a21oi_1 _7963_ (.A1(_0725_),
    .A2(net1910),
    .Y(_3534_),
    .B1(net1851));
 sg13g2_o21ai_1 _7964_ (.B1(_3534_),
    .Y(_3535_),
    .A1(_3532_),
    .A2(_3533_));
 sg13g2_a21oi_1 _7965_ (.A1(_2323_),
    .A2(net1851),
    .Y(_3536_),
    .B1(net1974));
 sg13g2_a22oi_1 _7966_ (.Y(_3537_),
    .B1(_3535_),
    .B2(_3536_),
    .A2(net1974),
    .A1(net266));
 sg13g2_inv_1 _7967_ (.Y(_0548_),
    .A(_3537_));
 sg13g2_mux2_1 _7968_ (.A0(\z80.tv80s.i_tv80_core.SP[8] ),
    .A1(_2836_),
    .S(net2138),
    .X(_3538_));
 sg13g2_xnor2_1 _7969_ (.Y(_3539_),
    .A(net1770),
    .B(_3538_));
 sg13g2_a221oi_1 _7970_ (.B2(_3527_),
    .C1(_3513_),
    .B1(net1770),
    .A1(_3514_),
    .Y(_3540_),
    .A2(_3515_));
 sg13g2_nor3_1 _7971_ (.A(_3528_),
    .B(_3539_),
    .C(_3540_),
    .Y(_3541_));
 sg13g2_o21ai_1 _7972_ (.B1(_3539_),
    .Y(_3542_),
    .A1(_3528_),
    .A2(_3540_));
 sg13g2_nand2b_2 _7973_ (.Y(_3543_),
    .B(_3542_),
    .A_N(_3541_));
 sg13g2_o21ai_1 _7974_ (.B1(net1751),
    .Y(_3544_),
    .A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .A2(net1773));
 sg13g2_a21o_1 _7975_ (.A2(_3543_),
    .A1(net1773),
    .B1(_3544_),
    .X(_3545_));
 sg13g2_a21oi_1 _7976_ (.A1(net1754),
    .A2(_2836_),
    .Y(_3546_),
    .B1(net1910));
 sg13g2_and2_1 _7977_ (.A(_2382_),
    .B(_3431_),
    .X(_3547_));
 sg13g2_a21oi_1 _7978_ (.A1(_3545_),
    .A2(_3546_),
    .Y(_3548_),
    .B1(net1850));
 sg13g2_o21ai_1 _7979_ (.B1(_3548_),
    .Y(_3549_),
    .A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .A2(net1898));
 sg13g2_a21oi_1 _7980_ (.A1(_1831_),
    .A2(net1849),
    .Y(_3550_),
    .B1(net1974));
 sg13g2_a22oi_1 _7981_ (.Y(_3551_),
    .B1(_3549_),
    .B2(_3550_),
    .A2(net1974),
    .A1(net242));
 sg13g2_inv_1 _7982_ (.Y(_0549_),
    .A(net243));
 sg13g2_a21o_1 _7983_ (.A2(_3538_),
    .A1(net1770),
    .B1(_3541_),
    .X(_3552_));
 sg13g2_nand2_1 _7984_ (.Y(_3553_),
    .A(_0682_),
    .B(\z80.tv80s.i_tv80_core.SP[9] ));
 sg13g2_nand2_1 _7985_ (.Y(_3554_),
    .A(net2137),
    .B(_2867_));
 sg13g2_a21oi_1 _7986_ (.A1(_3553_),
    .A2(_3554_),
    .Y(_3555_),
    .B1(_3525_));
 sg13g2_nand3_1 _7987_ (.B(_3553_),
    .C(_3554_),
    .A(_3525_),
    .Y(_3556_));
 sg13g2_nand2b_1 _7988_ (.Y(_3557_),
    .B(_3556_),
    .A_N(_3555_));
 sg13g2_xnor2_1 _7989_ (.Y(_3558_),
    .A(_3552_),
    .B(_3557_));
 sg13g2_nor2_1 _7990_ (.A(net1771),
    .B(_3558_),
    .Y(_3559_));
 sg13g2_o21ai_1 _7991_ (.B1(net1751),
    .Y(_3560_),
    .A1(\z80.tv80s.i_tv80_core.SP[9] ),
    .A2(net1773));
 sg13g2_a21oi_1 _7992_ (.A1(net1754),
    .A2(_2867_),
    .Y(_3561_),
    .B1(net1910));
 sg13g2_o21ai_1 _7993_ (.B1(_3561_),
    .Y(_3562_),
    .A1(_3559_),
    .A2(_3560_));
 sg13g2_o21ai_1 _7994_ (.B1(_3562_),
    .Y(_3563_),
    .A1(\z80.tv80s.i_tv80_core.SP[9] ),
    .A2(net1898));
 sg13g2_a21oi_1 _7995_ (.A1(_2005_),
    .A2(net1849),
    .Y(_3564_),
    .B1(net1962));
 sg13g2_o21ai_1 _7996_ (.B1(_3564_),
    .Y(_3565_),
    .A1(net1849),
    .A2(_3563_));
 sg13g2_o21ai_1 _7997_ (.B1(_3565_),
    .Y(_0550_),
    .A1(_0657_),
    .A2(net1984));
 sg13g2_nor2_1 _7998_ (.A(net2137),
    .B(\z80.tv80s.i_tv80_core.SP[10] ),
    .Y(_3566_));
 sg13g2_a21oi_2 _7999_ (.B1(_3566_),
    .Y(_3567_),
    .A2(_2902_),
    .A1(net2137));
 sg13g2_nand2_1 _8000_ (.Y(_3568_),
    .A(net1770),
    .B(_3567_));
 sg13g2_xnor2_1 _8001_ (.Y(_3569_),
    .A(net1769),
    .B(_3567_));
 sg13g2_a21oi_2 _8002_ (.B1(_3555_),
    .Y(_3570_),
    .A2(_3556_),
    .A1(_3552_));
 sg13g2_xor2_1 _8003_ (.B(_3570_),
    .A(_3569_),
    .X(_3571_));
 sg13g2_nor2_1 _8004_ (.A(net1771),
    .B(_3571_),
    .Y(_3572_));
 sg13g2_o21ai_1 _8005_ (.B1(net1750),
    .Y(_3573_),
    .A1(\z80.tv80s.i_tv80_core.SP[10] ),
    .A2(net1773));
 sg13g2_o21ai_1 _8006_ (.B1(net1900),
    .Y(_3574_),
    .A1(net1750),
    .A2(_2902_));
 sg13g2_inv_1 _8007_ (.Y(_3575_),
    .A(_3574_));
 sg13g2_o21ai_1 _8008_ (.B1(_3575_),
    .Y(_3576_),
    .A1(_3572_),
    .A2(_3573_));
 sg13g2_a21oi_1 _8009_ (.A1(_0701_),
    .A2(net1910),
    .Y(_3577_),
    .B1(_3547_));
 sg13g2_a221oi_1 _8010_ (.B2(_3577_),
    .C1(net1974),
    .B1(_3576_),
    .A1(_2050_),
    .Y(_3578_),
    .A2(net1849));
 sg13g2_a21o_1 _8011_ (.A2(net1974),
    .A1(net370),
    .B1(_3578_),
    .X(_0551_));
 sg13g2_nor2_1 _8012_ (.A(net2137),
    .B(\z80.tv80s.i_tv80_core.SP[11] ),
    .Y(_3579_));
 sg13g2_a21oi_1 _8013_ (.A1(net2137),
    .A2(_2924_),
    .Y(_3580_),
    .B1(_3579_));
 sg13g2_xnor2_1 _8014_ (.Y(_3581_),
    .A(_3525_),
    .B(_3580_));
 sg13g2_o21ai_1 _8015_ (.B1(_3568_),
    .Y(_3582_),
    .A1(_3569_),
    .A2(_3570_));
 sg13g2_xor2_1 _8016_ (.B(_3582_),
    .A(_3581_),
    .X(_3583_));
 sg13g2_nor2_1 _8017_ (.A(\z80.tv80s.i_tv80_core.SP[11] ),
    .B(net1773),
    .Y(_3584_));
 sg13g2_o21ai_1 _8018_ (.B1(net1750),
    .Y(_3585_),
    .A1(net1771),
    .A2(_3583_));
 sg13g2_a21oi_1 _8019_ (.A1(net1754),
    .A2(_2925_),
    .Y(_3586_),
    .B1(net1910));
 sg13g2_o21ai_1 _8020_ (.B1(_3586_),
    .Y(_3587_),
    .A1(_3584_),
    .A2(_3585_));
 sg13g2_o21ai_1 _8021_ (.B1(_3587_),
    .Y(_3588_),
    .A1(\z80.tv80s.i_tv80_core.SP[11] ),
    .A2(net1897));
 sg13g2_a21oi_1 _8022_ (.A1(_2101_),
    .A2(net1850),
    .Y(_3589_),
    .B1(net1961));
 sg13g2_o21ai_1 _8023_ (.B1(_3589_),
    .Y(_3590_),
    .A1(net1850),
    .A2(_3588_));
 sg13g2_o21ai_1 _8024_ (.B1(_3590_),
    .Y(_0552_),
    .A1(_0656_),
    .A2(net1984));
 sg13g2_nor2_1 _8025_ (.A(net2140),
    .B(\z80.tv80s.i_tv80_core.SP[12] ),
    .Y(_3591_));
 sg13g2_a21oi_1 _8026_ (.A1(net2140),
    .A2(_2959_),
    .Y(_3592_),
    .B1(_3591_));
 sg13g2_and2_1 _8027_ (.A(net1769),
    .B(_3592_),
    .X(_3593_));
 sg13g2_xnor2_1 _8028_ (.Y(_3594_),
    .A(net1769),
    .B(_3592_));
 sg13g2_inv_1 _8029_ (.Y(_3595_),
    .A(_3594_));
 sg13g2_o21ai_1 _8030_ (.B1(net1769),
    .Y(_3596_),
    .A1(_3567_),
    .A2(_3580_));
 sg13g2_nand2b_1 _8031_ (.Y(_3597_),
    .B(_3581_),
    .A_N(_3569_));
 sg13g2_o21ai_1 _8032_ (.B1(_3596_),
    .Y(_3598_),
    .A1(_3570_),
    .A2(_3597_));
 sg13g2_xnor2_1 _8033_ (.Y(_3599_),
    .A(_3594_),
    .B(_3598_));
 sg13g2_nor2_1 _8034_ (.A(net1771),
    .B(_3599_),
    .Y(_3600_));
 sg13g2_o21ai_1 _8035_ (.B1(net1750),
    .Y(_3601_),
    .A1(\z80.tv80s.i_tv80_core.SP[12] ),
    .A2(net1775));
 sg13g2_o21ai_1 _8036_ (.B1(net1900),
    .Y(_3602_),
    .A1(net1751),
    .A2(_2959_));
 sg13g2_inv_1 _8037_ (.Y(_3603_),
    .A(_3602_));
 sg13g2_o21ai_1 _8038_ (.B1(_3603_),
    .Y(_3604_),
    .A1(_3600_),
    .A2(_3601_));
 sg13g2_a21oi_1 _8039_ (.A1(_0710_),
    .A2(net1906),
    .Y(_3605_),
    .B1(net1849));
 sg13g2_a221oi_1 _8040_ (.B2(_3605_),
    .C1(net1961),
    .B1(_3604_),
    .A1(_2147_),
    .Y(_3606_),
    .A2(net1849));
 sg13g2_a21o_1 _8041_ (.A2(net1961),
    .A1(net346),
    .B1(_3606_),
    .X(_0553_));
 sg13g2_nand2_1 _8042_ (.Y(_3607_),
    .A(net200),
    .B(net1962));
 sg13g2_nor2_1 _8043_ (.A(net2139),
    .B(\z80.tv80s.i_tv80_core.SP[13] ),
    .Y(_3608_));
 sg13g2_a21oi_1 _8044_ (.A1(net2139),
    .A2(_2983_),
    .Y(_3609_),
    .B1(_3608_));
 sg13g2_xnor2_1 _8045_ (.Y(_3610_),
    .A(net1769),
    .B(_3609_));
 sg13g2_a21oi_1 _8046_ (.A1(_3595_),
    .A2(_3598_),
    .Y(_3611_),
    .B1(_3593_));
 sg13g2_xor2_1 _8047_ (.B(_3611_),
    .A(_3610_),
    .X(_3612_));
 sg13g2_mux2_1 _8048_ (.A0(\z80.tv80s.i_tv80_core.SP[13] ),
    .A1(_3612_),
    .S(net1773),
    .X(_3613_));
 sg13g2_o21ai_1 _8049_ (.B1(net1900),
    .Y(_3614_),
    .A1(net1751),
    .A2(_2983_));
 sg13g2_a21oi_1 _8050_ (.A1(net1751),
    .A2(_3613_),
    .Y(_3615_),
    .B1(_3614_));
 sg13g2_nor2_1 _8051_ (.A(\z80.tv80s.i_tv80_core.SP[13] ),
    .B(net1897),
    .Y(_3616_));
 sg13g2_nor3_1 _8052_ (.A(net1850),
    .B(_3615_),
    .C(_3616_),
    .Y(_3617_));
 sg13g2_a21o_1 _8053_ (.A2(net1850),
    .A1(_2220_),
    .B1(net1962),
    .X(_3618_));
 sg13g2_o21ai_1 _8054_ (.B1(_3607_),
    .Y(_0554_),
    .A1(_3617_),
    .A2(_3618_));
 sg13g2_nor2_1 _8055_ (.A(net2137),
    .B(\z80.tv80s.i_tv80_core.SP[14] ),
    .Y(_3619_));
 sg13g2_a21oi_1 _8056_ (.A1(net2139),
    .A2(_3016_),
    .Y(_3620_),
    .B1(_3619_));
 sg13g2_nand2_1 _8057_ (.Y(_3621_),
    .A(net1769),
    .B(_3620_));
 sg13g2_xnor2_1 _8058_ (.Y(_3622_),
    .A(net1769),
    .B(_3620_));
 sg13g2_nor2_1 _8059_ (.A(_3594_),
    .B(_3610_),
    .Y(_3623_));
 sg13g2_a221oi_1 _8060_ (.B2(_3598_),
    .C1(_3593_),
    .B1(_3623_),
    .A1(net1769),
    .Y(_3624_),
    .A2(_3609_));
 sg13g2_xor2_1 _8061_ (.B(_3624_),
    .A(_3622_),
    .X(_3625_));
 sg13g2_nor2_1 _8062_ (.A(net1771),
    .B(_3625_),
    .Y(_3626_));
 sg13g2_o21ai_1 _8063_ (.B1(net1750),
    .Y(_3627_),
    .A1(\z80.tv80s.i_tv80_core.SP[14] ),
    .A2(net1775));
 sg13g2_o21ai_1 _8064_ (.B1(net1900),
    .Y(_3628_),
    .A1(net1751),
    .A2(_3016_));
 sg13g2_inv_1 _8065_ (.Y(_3629_),
    .A(_3628_));
 sg13g2_o21ai_1 _8066_ (.B1(_3629_),
    .Y(_3630_),
    .A1(_3626_),
    .A2(_3627_));
 sg13g2_a21oi_1 _8067_ (.A1(_0718_),
    .A2(net1906),
    .Y(_3631_),
    .B1(net1850));
 sg13g2_a221oi_1 _8068_ (.B2(_3631_),
    .C1(net1962),
    .B1(_3630_),
    .A1(_2271_),
    .Y(_3632_),
    .A2(net1850));
 sg13g2_a21o_1 _8069_ (.A2(net1962),
    .A1(net349),
    .B1(_3632_),
    .X(_0555_));
 sg13g2_and2_1 _8070_ (.A(net517),
    .B(net1974),
    .X(_3633_));
 sg13g2_o21ai_1 _8071_ (.B1(_3621_),
    .Y(_3634_),
    .A1(_3622_),
    .A2(_3624_));
 sg13g2_nor2_1 _8072_ (.A(net2137),
    .B(\z80.tv80s.i_tv80_core.SP[15] ),
    .Y(_3635_));
 sg13g2_a21oi_1 _8073_ (.A1(net2137),
    .A2(_3040_),
    .Y(_3636_),
    .B1(_3635_));
 sg13g2_xnor2_1 _8074_ (.Y(_3637_),
    .A(_3525_),
    .B(_3636_));
 sg13g2_xnor2_1 _8075_ (.Y(_3638_),
    .A(_3634_),
    .B(_3637_));
 sg13g2_o21ai_1 _8076_ (.B1(net1750),
    .Y(_3639_),
    .A1(\z80.tv80s.i_tv80_core.SP[15] ),
    .A2(net1773));
 sg13g2_a21oi_1 _8077_ (.A1(net1773),
    .A2(_3638_),
    .Y(_3640_),
    .B1(_3639_));
 sg13g2_o21ai_1 _8078_ (.B1(net1900),
    .Y(_3641_),
    .A1(net1750),
    .A2(_3040_));
 sg13g2_a21oi_1 _8079_ (.A1(_0724_),
    .A2(net1910),
    .Y(_3642_),
    .B1(net1849));
 sg13g2_o21ai_1 _8080_ (.B1(_3642_),
    .Y(_3643_),
    .A1(_3640_),
    .A2(_3641_));
 sg13g2_a21oi_1 _8081_ (.A1(_2323_),
    .A2(net1849),
    .Y(_3644_),
    .B1(net1974));
 sg13g2_a21o_1 _8082_ (.A2(_3644_),
    .A1(_3643_),
    .B1(_3633_),
    .X(_0556_));
 sg13g2_nor2_1 _8083_ (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .B(_2473_),
    .Y(_3645_));
 sg13g2_nor2_1 _8084_ (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .B(_2373_),
    .Y(_3646_));
 sg13g2_o21ai_1 _8085_ (.B1(net1687),
    .Y(_3647_),
    .A1(_3645_),
    .A2(_3646_));
 sg13g2_nand4_1 _8086_ (.B(_1134_),
    .C(_1344_),
    .A(net1687),
    .Y(_3648_),
    .D(_3647_));
 sg13g2_inv_1 _8087_ (.Y(_3649_),
    .A(_3648_));
 sg13g2_nand4_1 _8088_ (.B(_1344_),
    .C(_2476_),
    .A(_1134_),
    .Y(_3650_),
    .D(_3647_));
 sg13g2_a22oi_1 _8089_ (.Y(_0557_),
    .B1(_3650_),
    .B2(_0655_),
    .A2(_3649_),
    .A1(_0687_));
 sg13g2_a22oi_1 _8090_ (.Y(_0558_),
    .B1(_3650_),
    .B2(_0683_),
    .A2(_3649_),
    .A1(_0686_));
 sg13g2_nand2_1 _8091_ (.Y(_3651_),
    .A(\z80.tv80s.i_tv80_core.ts[2] ),
    .B(_3650_));
 sg13g2_o21ai_1 _8092_ (.B1(_3651_),
    .Y(_0559_),
    .A1(net476),
    .A2(_3648_));
 sg13g2_nand2_1 _8093_ (.Y(_3652_),
    .A(net2142),
    .B(_3650_));
 sg13g2_o21ai_1 _8094_ (.B1(_3652_),
    .Y(_0560_),
    .A1(net516),
    .A2(_3648_));
 sg13g2_nand2_1 _8095_ (.Y(_3653_),
    .A(net545),
    .B(_3650_));
 sg13g2_o21ai_1 _8096_ (.B1(_3653_),
    .Y(_0561_),
    .A1(_0023_),
    .A2(_3648_));
 sg13g2_a22oi_1 _8097_ (.Y(_3654_),
    .B1(_3650_),
    .B2(net189),
    .A2(_3649_),
    .A1(\z80.tv80s.i_tv80_core.ts[4] ));
 sg13g2_inv_1 _8098_ (.Y(_0562_),
    .A(net190));
 sg13g2_nand2_1 _8099_ (.Y(_3655_),
    .A(\z80.tv80s.i_tv80_core.ts[6] ),
    .B(_3650_));
 sg13g2_o21ai_1 _8100_ (.B1(_3655_),
    .Y(_0563_),
    .A1(net183),
    .A2(_3648_));
 sg13g2_nor2_1 _8101_ (.A(\z80.tv80s.i_tv80_core.Halt_FF ),
    .B(_1592_),
    .Y(_3656_));
 sg13g2_nand3_1 _8102_ (.B(_2601_),
    .C(_3656_),
    .A(_2568_),
    .Y(_3657_));
 sg13g2_o21ai_1 _8103_ (.B1(_0833_),
    .Y(_3658_),
    .A1(net1726),
    .A2(_3657_));
 sg13g2_nand2_1 _8104_ (.Y(_3659_),
    .A(_0826_),
    .B(_3658_));
 sg13g2_inv_2 _8105_ (.Y(_3660_),
    .A(net1695));
 sg13g2_or3_1 _8106_ (.A(_0971_),
    .B(net1884),
    .C(_1431_),
    .X(_3661_));
 sg13g2_nand2_1 _8107_ (.Y(_3662_),
    .A(_0903_),
    .B(_1511_));
 sg13g2_nor3_2 _8108_ (.A(_1666_),
    .B(_3661_),
    .C(_3662_),
    .Y(_3663_));
 sg13g2_nand3_1 _8109_ (.B(_1245_),
    .C(_2352_),
    .A(_0931_),
    .Y(_3664_));
 sg13g2_a22oi_1 _8110_ (.Y(_3665_),
    .B1(_3664_),
    .B2(_0677_),
    .A2(net1922),
    .A1(_1011_));
 sg13g2_o21ai_1 _8111_ (.B1(_3665_),
    .Y(_3666_),
    .A1(net1942),
    .A2(_3663_));
 sg13g2_nand3_1 _8112_ (.B(_1147_),
    .C(_1241_),
    .A(_0975_),
    .Y(_3667_));
 sg13g2_or2_1 _8113_ (.X(_3668_),
    .B(_1173_),
    .A(_0997_));
 sg13g2_nand3_1 _8114_ (.B(_1233_),
    .C(_1234_),
    .A(_1177_),
    .Y(_3669_));
 sg13g2_nand4_1 _8115_ (.B(_0934_),
    .C(_2360_),
    .A(net1950),
    .Y(_3670_),
    .D(_2577_));
 sg13g2_nor4_1 _8116_ (.A(_0981_),
    .B(_0992_),
    .C(_1008_),
    .D(_3670_),
    .Y(_3671_));
 sg13g2_nand2b_1 _8117_ (.Y(_3672_),
    .B(_3671_),
    .A_N(_3664_));
 sg13g2_nor4_1 _8118_ (.A(_1016_),
    .B(_1161_),
    .C(_3669_),
    .D(_3672_),
    .Y(_3673_));
 sg13g2_nand2_1 _8119_ (.Y(_3674_),
    .A(_3663_),
    .B(_3673_));
 sg13g2_nor3_1 _8120_ (.A(_3667_),
    .B(_3668_),
    .C(_3674_),
    .Y(_3675_));
 sg13g2_o21ai_1 _8121_ (.B1(net2171),
    .Y(_3676_),
    .A1(_3666_),
    .A2(_3675_));
 sg13g2_nor4_2 _8122_ (.A(_0911_),
    .B(_0936_),
    .C(_1168_),
    .Y(_3677_),
    .D(_1172_));
 sg13g2_a221oi_1 _8123_ (.B2(net2131),
    .C1(net1884),
    .B1(_1011_),
    .A1(_0942_),
    .Y(_3678_),
    .A2(_0948_));
 sg13g2_nor4_1 _8124_ (.A(_0945_),
    .B(_0972_),
    .C(_1013_),
    .D(_1148_),
    .Y(_3679_));
 sg13g2_nor3_1 _8125_ (.A(_0933_),
    .B(_0941_),
    .C(_0944_),
    .Y(_3680_));
 sg13g2_nand4_1 _8126_ (.B(_3678_),
    .C(_3679_),
    .A(_1146_),
    .Y(_3681_),
    .D(_3680_));
 sg13g2_nor4_1 _8127_ (.A(_0926_),
    .B(_0964_),
    .C(_1244_),
    .D(_1259_),
    .Y(_3682_));
 sg13g2_nor4_1 _8128_ (.A(net2017),
    .B(_0887_),
    .C(_1526_),
    .D(_1527_),
    .Y(_3683_));
 sg13g2_nand4_1 _8129_ (.B(_1530_),
    .C(_3682_),
    .A(_1266_),
    .Y(_3684_),
    .D(_3683_));
 sg13g2_nor4_2 _8130_ (.A(_1524_),
    .B(_2480_),
    .C(_3681_),
    .Y(_3685_),
    .D(_3684_));
 sg13g2_or4_2 _8131_ (.A(_1524_),
    .B(_2480_),
    .C(_3681_),
    .D(_3684_),
    .X(_3686_));
 sg13g2_nor2b_2 _8132_ (.A(_2350_),
    .B_N(_3677_),
    .Y(_3687_));
 sg13g2_nand2b_1 _8133_ (.Y(_3688_),
    .B(_3677_),
    .A_N(_2350_));
 sg13g2_nand4_1 _8134_ (.B(_1523_),
    .C(_1530_),
    .A(_1176_),
    .Y(_3689_),
    .D(_2479_));
 sg13g2_nor3_1 _8135_ (.A(_1259_),
    .B(_1526_),
    .C(_1527_),
    .Y(_3690_));
 sg13g2_nor3_1 _8136_ (.A(_0926_),
    .B(_0932_),
    .C(_0981_),
    .Y(_3691_));
 sg13g2_nand4_1 _8137_ (.B(_1709_),
    .C(_3690_),
    .A(_1146_),
    .Y(_3692_),
    .D(_3691_));
 sg13g2_nor4_1 _8138_ (.A(_0941_),
    .B(_0944_),
    .C(_0945_),
    .D(_0972_),
    .Y(_3693_));
 sg13g2_nor4_1 _8139_ (.A(_0933_),
    .B(_0964_),
    .C(_1013_),
    .D(_1148_),
    .Y(_3694_));
 sg13g2_nand4_1 _8140_ (.B(_2478_),
    .C(_3693_),
    .A(_1243_),
    .Y(_3695_),
    .D(_3694_));
 sg13g2_nor4_2 _8141_ (.A(_2350_),
    .B(_3689_),
    .C(_3692_),
    .Y(_3696_),
    .D(_3695_));
 sg13g2_and4_2 _8142_ (.A(_1554_),
    .B(_2358_),
    .C(_3677_),
    .D(_3696_),
    .X(_3697_));
 sg13g2_a21oi_2 _8143_ (.B1(\z80.tv80s.i_tv80_core.BTR_r ),
    .Y(_3698_),
    .A2(_3687_),
    .A1(_3685_));
 sg13g2_a21oi_1 _8144_ (.A1(_0033_),
    .A2(_1138_),
    .Y(_3699_),
    .B1(net2025));
 sg13g2_nand2_1 _8145_ (.Y(_3700_),
    .A(net185),
    .B(net1900));
 sg13g2_o21ai_1 _8146_ (.B1(_3676_),
    .Y(_3701_),
    .A1(net1943),
    .A2(_1278_));
 sg13g2_nor3_1 _8147_ (.A(_3699_),
    .B(_3700_),
    .C(_3701_),
    .Y(_3702_));
 sg13g2_a22oi_1 _8148_ (.Y(_3703_),
    .B1(_3698_),
    .B2(_3702_),
    .A2(net1997),
    .A1(net1903));
 sg13g2_inv_1 _8149_ (.Y(_3704_),
    .A(net1714));
 sg13g2_o21ai_1 _8150_ (.B1(_3660_),
    .Y(_3705_),
    .A1(net1692),
    .A2(net1715));
 sg13g2_nor3_1 _8151_ (.A(_0169_),
    .B(_3686_),
    .C(_3688_),
    .Y(_3706_));
 sg13g2_nor2_1 _8152_ (.A(_3698_),
    .B(_3706_),
    .Y(_3707_));
 sg13g2_xnor2_1 _8153_ (.Y(_3708_),
    .A(_0194_),
    .B(_3707_));
 sg13g2_nor2_1 _8154_ (.A(net2136),
    .B(net1920),
    .Y(_3709_));
 sg13g2_nor2_1 _8155_ (.A(\z80.tv80s.i_tv80_core.PC[0] ),
    .B(net1872),
    .Y(_3710_));
 sg13g2_nor3_1 _8156_ (.A(net1758),
    .B(_3709_),
    .C(_3710_),
    .Y(_3711_));
 sg13g2_o21ai_1 _8157_ (.B1(net1841),
    .Y(_3712_),
    .A1(_2603_),
    .A2(_3711_));
 sg13g2_a21oi_1 _8158_ (.A1(_2594_),
    .A2(_3712_),
    .Y(_3713_),
    .B1(net1725));
 sg13g2_nor3_1 _8159_ (.A(_2585_),
    .B(_3703_),
    .C(_3713_),
    .Y(_3714_));
 sg13g2_a22oi_1 _8160_ (.Y(_3715_),
    .B1(_3714_),
    .B2(net1693),
    .A2(_3708_),
    .A1(_3703_));
 sg13g2_nor2_1 _8161_ (.A(net1696),
    .B(_3715_),
    .Y(_3716_));
 sg13g2_a21oi_1 _8162_ (.A1(_0735_),
    .A2(_3705_),
    .Y(_0564_),
    .B1(_3716_));
 sg13g2_nand2_1 _8163_ (.Y(_3717_),
    .A(net528),
    .B(_3705_));
 sg13g2_o21ai_1 _8164_ (.B1(\z80.tv80s.i_tv80_core.PC[0] ),
    .Y(_3718_),
    .A1(_3698_),
    .A2(_3706_));
 sg13g2_a21oi_2 _8165_ (.B1(_0798_),
    .Y(_3719_),
    .A2(_3687_),
    .A1(_3685_));
 sg13g2_o21ai_1 _8166_ (.B1(_0229_),
    .Y(_3720_),
    .A1(_3686_),
    .A2(_3688_));
 sg13g2_and3_1 _8167_ (.X(_3721_),
    .A(_0172_),
    .B(_3685_),
    .C(_3687_));
 sg13g2_nand3b_1 _8168_ (.B(_0196_),
    .C(_3720_),
    .Y(_3722_),
    .A_N(_3721_));
 sg13g2_o21ai_1 _8169_ (.B1(_0771_),
    .Y(_3723_),
    .A1(_3719_),
    .A2(_3721_));
 sg13g2_a21oi_1 _8170_ (.A1(_3722_),
    .A2(_3723_),
    .Y(_3724_),
    .B1(_3718_));
 sg13g2_nand3_1 _8171_ (.B(_3722_),
    .C(_3723_),
    .A(_3718_),
    .Y(_3725_));
 sg13g2_nor2_1 _8172_ (.A(net1703),
    .B(_3724_),
    .Y(_3726_));
 sg13g2_nand2_1 _8173_ (.Y(_3727_),
    .A(\z80.tv80s.i_tv80_core.PC[1] ),
    .B(net1920));
 sg13g2_a21oi_1 _8174_ (.A1(_2639_),
    .A2(_3727_),
    .Y(_3728_),
    .B1(net1782));
 sg13g2_a21oi_1 _8175_ (.A1(net2135),
    .A2(net1782),
    .Y(_3729_),
    .B1(_3728_));
 sg13g2_mux2_1 _8176_ (.A0(_2650_),
    .A1(_3729_),
    .S(net1840),
    .X(_3730_));
 sg13g2_nor2_1 _8177_ (.A(net1724),
    .B(_3730_),
    .Y(_3731_));
 sg13g2_a21oi_1 _8178_ (.A1(net2135),
    .A2(net1725),
    .Y(_3732_),
    .B1(_3731_));
 sg13g2_nor2_1 _8179_ (.A(net1716),
    .B(_3732_),
    .Y(_3733_));
 sg13g2_a22oi_1 _8180_ (.Y(_3734_),
    .B1(_3733_),
    .B2(net1693),
    .A2(_3726_),
    .A1(_3725_));
 sg13g2_o21ai_1 _8181_ (.B1(_3717_),
    .Y(_0565_),
    .A1(net1696),
    .A2(_3734_));
 sg13g2_nand2_1 _8182_ (.Y(_3735_),
    .A(net544),
    .B(_3705_));
 sg13g2_nor3_1 _8183_ (.A(_0741_),
    .B(_3719_),
    .C(_3721_),
    .Y(_3736_));
 sg13g2_a21o_1 _8184_ (.A2(_3697_),
    .A1(_0175_),
    .B1(_3719_),
    .X(_3737_));
 sg13g2_xnor2_1 _8185_ (.Y(_3738_),
    .A(\z80.tv80s.i_tv80_core.PC[2] ),
    .B(_3737_));
 sg13g2_o21ai_1 _8186_ (.B1(_3738_),
    .Y(_3739_),
    .A1(_3724_),
    .A2(_3736_));
 sg13g2_nor3_1 _8187_ (.A(_3724_),
    .B(_3736_),
    .C(_3738_),
    .Y(_3740_));
 sg13g2_nor2_1 _8188_ (.A(net1703),
    .B(_3740_),
    .Y(_3741_));
 sg13g2_nand2_1 _8189_ (.Y(_3742_),
    .A(\z80.tv80s.i_tv80_core.PC[2] ),
    .B(net1921));
 sg13g2_a21oi_1 _8190_ (.A1(_2665_),
    .A2(_3742_),
    .Y(_3743_),
    .B1(net1783));
 sg13g2_a21o_1 _8191_ (.A2(net1781),
    .A1(net2134),
    .B1(_3743_),
    .X(_3744_));
 sg13g2_a21oi_1 _8192_ (.A1(net1838),
    .A2(_3744_),
    .Y(_3745_),
    .B1(_2687_));
 sg13g2_mux2_1 _8193_ (.A0(_3745_),
    .A1(_0763_),
    .S(net1726),
    .X(_3746_));
 sg13g2_nor2_1 _8194_ (.A(net1716),
    .B(_3746_),
    .Y(_3747_));
 sg13g2_a22oi_1 _8195_ (.Y(_3748_),
    .B1(_3747_),
    .B2(net1693),
    .A2(_3741_),
    .A1(_3739_));
 sg13g2_o21ai_1 _8196_ (.B1(_3735_),
    .Y(_0566_),
    .A1(net1696),
    .A2(_3748_));
 sg13g2_nand2_1 _8197_ (.Y(_3749_),
    .A(net549),
    .B(_3705_));
 sg13g2_or2_1 _8198_ (.X(_3750_),
    .B(_3737_),
    .A(_0198_));
 sg13g2_a21oi_1 _8199_ (.A1(_0178_),
    .A2(_3697_),
    .Y(_3751_),
    .B1(_3719_));
 sg13g2_and2_1 _8200_ (.A(\z80.tv80s.i_tv80_core.PC[3] ),
    .B(_3751_),
    .X(_3752_));
 sg13g2_xnor2_1 _8201_ (.Y(_3753_),
    .A(\z80.tv80s.i_tv80_core.PC[3] ),
    .B(_3751_));
 sg13g2_a21oi_1 _8202_ (.A1(_3739_),
    .A2(_3750_),
    .Y(_3754_),
    .B1(_3753_));
 sg13g2_and3_1 _8203_ (.X(_3755_),
    .A(_3739_),
    .B(_3750_),
    .C(_3753_));
 sg13g2_nor3_1 _8204_ (.A(_3704_),
    .B(_3754_),
    .C(_3755_),
    .Y(_3756_));
 sg13g2_nand2_1 _8205_ (.Y(_3757_),
    .A(_0762_),
    .B(net1867));
 sg13g2_o21ai_1 _8206_ (.B1(_3757_),
    .Y(_3758_),
    .A1(\z80.tv80s.i_tv80_core.PC[3] ),
    .A2(net1867));
 sg13g2_o21ai_1 _8207_ (.B1(_2703_),
    .Y(_3759_),
    .A1(net1759),
    .A2(_3758_));
 sg13g2_a21oi_1 _8208_ (.A1(net1838),
    .A2(_3759_),
    .Y(_3760_),
    .B1(_2702_));
 sg13g2_nor2_1 _8209_ (.A(net1721),
    .B(_3760_),
    .Y(_3761_));
 sg13g2_a21oi_2 _8210_ (.B1(_3761_),
    .Y(_3762_),
    .A2(net1721),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sg13g2_nor2_1 _8211_ (.A(net1716),
    .B(_3762_),
    .Y(_3763_));
 sg13g2_a21oi_1 _8212_ (.A1(net1692),
    .A2(_3763_),
    .Y(_3764_),
    .B1(_3756_));
 sg13g2_o21ai_1 _8213_ (.B1(_3749_),
    .Y(_0567_),
    .A1(net1696),
    .A2(_3764_));
 sg13g2_nand2_1 _8214_ (.Y(_3765_),
    .A(net551),
    .B(_3705_));
 sg13g2_a21o_1 _8215_ (.A2(_3697_),
    .A1(_0181_),
    .B1(_3719_),
    .X(_3766_));
 sg13g2_xnor2_1 _8216_ (.Y(_3767_),
    .A(\z80.tv80s.i_tv80_core.PC[4] ),
    .B(_3766_));
 sg13g2_o21ai_1 _8217_ (.B1(_3767_),
    .Y(_3768_),
    .A1(_3752_),
    .A2(_3754_));
 sg13g2_nor3_1 _8218_ (.A(_3752_),
    .B(_3754_),
    .C(_3767_),
    .Y(_3769_));
 sg13g2_nor2_1 _8219_ (.A(_3704_),
    .B(_3769_),
    .Y(_3770_));
 sg13g2_nor2_1 _8220_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .B(net1921),
    .Y(_3771_));
 sg13g2_nor2_1 _8221_ (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .B(net1867),
    .Y(_3772_));
 sg13g2_nor3_1 _8222_ (.A(net1756),
    .B(_3771_),
    .C(_3772_),
    .Y(_3773_));
 sg13g2_o21ai_1 _8223_ (.B1(net1838),
    .Y(_3774_),
    .A1(_2719_),
    .A2(_3773_));
 sg13g2_a21oi_1 _8224_ (.A1(_2740_),
    .A2(_3774_),
    .Y(_3775_),
    .B1(net1721));
 sg13g2_a21oi_1 _8225_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net1726),
    .Y(_3776_),
    .B1(_3775_));
 sg13g2_nor2_1 _8226_ (.A(net1716),
    .B(_3776_),
    .Y(_3777_));
 sg13g2_a22oi_1 _8227_ (.Y(_3778_),
    .B1(_3777_),
    .B2(net1693),
    .A2(_3770_),
    .A1(_3768_));
 sg13g2_o21ai_1 _8228_ (.B1(_3765_),
    .Y(_0568_),
    .A1(net1696),
    .A2(_3778_));
 sg13g2_or2_1 _8229_ (.X(_3779_),
    .B(_3766_),
    .A(_0202_));
 sg13g2_nand2_1 _8230_ (.Y(_3780_),
    .A(_3768_),
    .B(_3779_));
 sg13g2_nand2_1 _8231_ (.Y(_3781_),
    .A(_0184_),
    .B(_3697_));
 sg13g2_and3_1 _8232_ (.X(_3782_),
    .A(\z80.tv80s.i_tv80_core.PC[5] ),
    .B(_3720_),
    .C(_3781_));
 sg13g2_a21oi_1 _8233_ (.A1(_3720_),
    .A2(_3781_),
    .Y(_3783_),
    .B1(\z80.tv80s.i_tv80_core.PC[5] ));
 sg13g2_nor2_1 _8234_ (.A(_3782_),
    .B(_3783_),
    .Y(_3784_));
 sg13g2_a21oi_1 _8235_ (.A1(_3780_),
    .A2(_3784_),
    .Y(_3785_),
    .B1(net1703));
 sg13g2_o21ai_1 _8236_ (.B1(_3785_),
    .Y(_3786_),
    .A1(_3780_),
    .A2(_3784_));
 sg13g2_nand2_1 _8237_ (.Y(_3787_),
    .A(\z80.tv80s.i_tv80_core.PC[5] ),
    .B(net1921));
 sg13g2_a21oi_1 _8238_ (.A1(_2755_),
    .A2(_3787_),
    .Y(_3788_),
    .B1(net1781));
 sg13g2_a21oi_1 _8239_ (.A1(net2133),
    .A2(net1781),
    .Y(_3789_),
    .B1(_3788_));
 sg13g2_mux2_1 _8240_ (.A0(_2752_),
    .A1(_3789_),
    .S(net1839),
    .X(_3790_));
 sg13g2_o21ai_1 _8241_ (.B1(_2767_),
    .Y(_3791_),
    .A1(net1726),
    .A2(_3790_));
 sg13g2_nand3_1 _8242_ (.B(_3704_),
    .C(_3791_),
    .A(net1693),
    .Y(_3792_));
 sg13g2_a21oi_1 _8243_ (.A1(_3786_),
    .A2(_3792_),
    .Y(_3793_),
    .B1(net1696));
 sg13g2_a21o_1 _8244_ (.A2(_3705_),
    .A1(net603),
    .B1(_3793_),
    .X(_0569_));
 sg13g2_a21oi_1 _8245_ (.A1(_3768_),
    .A2(_3779_),
    .Y(_3794_),
    .B1(_3783_));
 sg13g2_a21o_1 _8246_ (.A2(_3697_),
    .A1(_0187_),
    .B1(_3719_),
    .X(_3795_));
 sg13g2_xnor2_1 _8247_ (.Y(_3796_),
    .A(\z80.tv80s.i_tv80_core.PC[6] ),
    .B(_3795_));
 sg13g2_nor3_1 _8248_ (.A(_3782_),
    .B(_3794_),
    .C(_3796_),
    .Y(_3797_));
 sg13g2_o21ai_1 _8249_ (.B1(_3796_),
    .Y(_3798_),
    .A1(_3782_),
    .A2(_3794_));
 sg13g2_nand3b_1 _8250_ (.B(_3798_),
    .C(_3703_),
    .Y(_3799_),
    .A_N(_3797_));
 sg13g2_nand2_1 _8251_ (.Y(_3800_),
    .A(\z80.tv80s.i_tv80_core.PC[6] ),
    .B(net1921));
 sg13g2_a21oi_1 _8252_ (.A1(_2784_),
    .A2(_3800_),
    .Y(_3801_),
    .B1(net1782));
 sg13g2_o21ai_1 _8253_ (.B1(net1841),
    .Y(_3802_),
    .A1(_2783_),
    .A2(_3801_));
 sg13g2_a21oi_1 _8254_ (.A1(_2782_),
    .A2(_3802_),
    .Y(_3803_),
    .B1(net1724));
 sg13g2_or2_1 _8255_ (.X(_3804_),
    .B(_3803_),
    .A(_2772_));
 sg13g2_mux2_1 _8256_ (.A0(\z80.tv80s.i_tv80_core.PC[6] ),
    .A1(_3804_),
    .S(net1693),
    .X(_3805_));
 sg13g2_a21oi_1 _8257_ (.A1(net1703),
    .A2(_3805_),
    .Y(_3806_),
    .B1(net1697));
 sg13g2_a22oi_1 _8258_ (.Y(_0570_),
    .B1(_3799_),
    .B2(_3806_),
    .A2(net1697),
    .A1(_0749_));
 sg13g2_a21oi_1 _8259_ (.A1(_0190_),
    .A2(_3697_),
    .Y(_3807_),
    .B1(_3719_));
 sg13g2_a21o_2 _8260_ (.A2(_3697_),
    .A1(_0190_),
    .B1(_3719_),
    .X(_3808_));
 sg13g2_nor2_1 _8261_ (.A(_0751_),
    .B(_3808_),
    .Y(_3809_));
 sg13g2_xnor2_1 _8262_ (.Y(_3810_),
    .A(\z80.tv80s.i_tv80_core.PC[7] ),
    .B(net1846));
 sg13g2_nand2b_1 _8263_ (.Y(_3811_),
    .B(_0776_),
    .A_N(_3795_));
 sg13g2_nand3_1 _8264_ (.B(_3810_),
    .C(_3811_),
    .A(_3798_),
    .Y(_3812_));
 sg13g2_a21oi_1 _8265_ (.A1(_3798_),
    .A2(_3811_),
    .Y(_3813_),
    .B1(_3810_));
 sg13g2_nand2_1 _8266_ (.Y(_3814_),
    .A(_0751_),
    .B(net1920));
 sg13g2_o21ai_1 _8267_ (.B1(_3814_),
    .Y(_3815_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A2(net1920));
 sg13g2_o21ai_1 _8268_ (.B1(_2801_),
    .Y(_3816_),
    .A1(net1758),
    .A2(_3815_));
 sg13g2_a21oi_1 _8269_ (.A1(net1840),
    .A2(_3816_),
    .Y(_3817_),
    .B1(_2822_));
 sg13g2_o21ai_1 _8270_ (.B1(_2824_),
    .Y(_3818_),
    .A1(net1723),
    .A2(_3817_));
 sg13g2_a21oi_1 _8271_ (.A1(_0751_),
    .A2(net1687),
    .Y(_3819_),
    .B1(net1716));
 sg13g2_o21ai_1 _8272_ (.B1(_3819_),
    .Y(_3820_),
    .A1(net1687),
    .A2(_3818_));
 sg13g2_nor2_1 _8273_ (.A(net1703),
    .B(_3813_),
    .Y(_3821_));
 sg13g2_a21oi_1 _8274_ (.A1(_3812_),
    .A2(_3821_),
    .Y(_3822_),
    .B1(net1696));
 sg13g2_a22oi_1 _8275_ (.Y(_0571_),
    .B1(_3820_),
    .B2(_3822_),
    .A2(net1696),
    .A1(_0751_));
 sg13g2_xnor2_1 _8276_ (.Y(_3823_),
    .A(\z80.tv80s.i_tv80_core.PC[8] ),
    .B(net1846));
 sg13g2_inv_1 _8277_ (.Y(_3824_),
    .A(_3823_));
 sg13g2_o21ai_1 _8278_ (.B1(_3824_),
    .Y(_3825_),
    .A1(_3809_),
    .A2(_3813_));
 sg13g2_nor3_1 _8279_ (.A(_3809_),
    .B(_3813_),
    .C(_3824_),
    .Y(_3826_));
 sg13g2_nand2_1 _8280_ (.Y(_3827_),
    .A(\z80.tv80s.i_tv80_core.PC[8] ),
    .B(net1920));
 sg13g2_a21oi_1 _8281_ (.A1(_2839_),
    .A2(_3827_),
    .Y(_3828_),
    .B1(net1758));
 sg13g2_o21ai_1 _8282_ (.B1(net1840),
    .Y(_3829_),
    .A1(_2838_),
    .A2(_3828_));
 sg13g2_a21oi_1 _8283_ (.A1(_2837_),
    .A2(_3829_),
    .Y(_3830_),
    .B1(net1723));
 sg13g2_nor2_1 _8284_ (.A(_2857_),
    .B(_3830_),
    .Y(_3831_));
 sg13g2_nor2_1 _8285_ (.A(\z80.tv80s.i_tv80_core.PC[8] ),
    .B(net1692),
    .Y(_3832_));
 sg13g2_a21oi_1 _8286_ (.A1(net1692),
    .A2(_3831_),
    .Y(_3833_),
    .B1(_3832_));
 sg13g2_nand3b_1 _8287_ (.B(net1715),
    .C(_3825_),
    .Y(_3834_),
    .A_N(_3826_));
 sg13g2_a21oi_1 _8288_ (.A1(net1703),
    .A2(_3833_),
    .Y(_3835_),
    .B1(net1697));
 sg13g2_a22oi_1 _8289_ (.Y(_0572_),
    .B1(_3834_),
    .B2(_3835_),
    .A2(net1697),
    .A1(_0734_));
 sg13g2_nand2b_1 _8290_ (.Y(_3836_),
    .B(net1846),
    .A_N(_0171_));
 sg13g2_nand2_1 _8291_ (.Y(_3837_),
    .A(_3825_),
    .B(_3836_));
 sg13g2_nand2_1 _8292_ (.Y(_3838_),
    .A(_0740_),
    .B(_3808_));
 sg13g2_nand2_1 _8293_ (.Y(_3839_),
    .A(\z80.tv80s.i_tv80_core.PC[9] ),
    .B(net1846));
 sg13g2_nand2_1 _8294_ (.Y(_3840_),
    .A(_3838_),
    .B(_3839_));
 sg13g2_xor2_1 _8295_ (.B(_3840_),
    .A(_3837_),
    .X(_3841_));
 sg13g2_nor2_1 _8296_ (.A(_0740_),
    .B(net1870),
    .Y(_3842_));
 sg13g2_a21oi_1 _8297_ (.A1(\z80.tv80s.i_tv80_core.I[1] ),
    .A2(net1870),
    .Y(_3843_),
    .B1(_3842_));
 sg13g2_o21ai_1 _8298_ (.B1(_2869_),
    .Y(_3844_),
    .A1(net1757),
    .A2(_3843_));
 sg13g2_a21oi_1 _8299_ (.A1(net1836),
    .A2(_3844_),
    .Y(_3845_),
    .B1(_2868_));
 sg13g2_o21ai_1 _8300_ (.B1(_2885_),
    .Y(_3846_),
    .A1(net1722),
    .A2(_3845_));
 sg13g2_nand2_1 _8301_ (.Y(_3847_),
    .A(net1690),
    .B(_3846_));
 sg13g2_o21ai_1 _8302_ (.B1(_3847_),
    .Y(_3848_),
    .A1(_0740_),
    .A2(net1691));
 sg13g2_a21oi_1 _8303_ (.A1(net1715),
    .A2(_3841_),
    .Y(_3849_),
    .B1(net1695));
 sg13g2_o21ai_1 _8304_ (.B1(_3849_),
    .Y(_3850_),
    .A1(net1716),
    .A2(_3848_));
 sg13g2_o21ai_1 _8305_ (.B1(_3850_),
    .Y(_0573_),
    .A1(_0740_),
    .A2(_3660_));
 sg13g2_nand3_1 _8306_ (.B(_3836_),
    .C(_3839_),
    .A(_3825_),
    .Y(_3851_));
 sg13g2_xnor2_1 _8307_ (.Y(_3852_),
    .A(\z80.tv80s.i_tv80_core.PC[10] ),
    .B(net1845));
 sg13g2_inv_1 _8308_ (.Y(_3853_),
    .A(_3852_));
 sg13g2_nand3_1 _8309_ (.B(_3851_),
    .C(_3853_),
    .A(_3838_),
    .Y(_3854_));
 sg13g2_a21o_1 _8310_ (.A2(_3851_),
    .A1(_3838_),
    .B1(_3853_),
    .X(_3855_));
 sg13g2_nand3_1 _8311_ (.B(_3854_),
    .C(_3855_),
    .A(net1715),
    .Y(_3856_));
 sg13g2_nand2_1 _8312_ (.Y(_3857_),
    .A(\z80.tv80s.i_tv80_core.PC[10] ),
    .B(net1920));
 sg13g2_a21oi_1 _8313_ (.A1(_2890_),
    .A2(_3857_),
    .Y(_3858_),
    .B1(net1757));
 sg13g2_o21ai_1 _8314_ (.B1(net1836),
    .Y(_3859_),
    .A1(_2889_),
    .A2(_3858_));
 sg13g2_a21oi_1 _8315_ (.A1(_2913_),
    .A2(_3859_),
    .Y(_3860_),
    .B1(net1723));
 sg13g2_a21oi_1 _8316_ (.A1(net2049),
    .A2(net1723),
    .Y(_3861_),
    .B1(_3860_));
 sg13g2_nand2b_1 _8317_ (.Y(_3862_),
    .B(net1690),
    .A_N(_3861_));
 sg13g2_o21ai_1 _8318_ (.B1(_3862_),
    .Y(_3863_),
    .A1(_0744_),
    .A2(net1691));
 sg13g2_a21oi_1 _8319_ (.A1(net1703),
    .A2(_3863_),
    .Y(_3864_),
    .B1(net1695));
 sg13g2_a22oi_1 _8320_ (.Y(_0574_),
    .B1(_3856_),
    .B2(_3864_),
    .A2(net1695),
    .A1(_0744_));
 sg13g2_o21ai_1 _8321_ (.B1(_3854_),
    .Y(_3865_),
    .A1(_0177_),
    .A2(_3808_));
 sg13g2_xnor2_1 _8322_ (.Y(_3866_),
    .A(_0745_),
    .B(net1845));
 sg13g2_xnor2_1 _8323_ (.Y(_3867_),
    .A(_3865_),
    .B(_3866_));
 sg13g2_nor2_1 _8324_ (.A(_0745_),
    .B(net1869),
    .Y(_3868_));
 sg13g2_a21oi_1 _8325_ (.A1(\z80.tv80s.i_tv80_core.I[3] ),
    .A2(net1869),
    .Y(_3869_),
    .B1(_3868_));
 sg13g2_o21ai_1 _8326_ (.B1(_2927_),
    .Y(_3870_),
    .A1(net1757),
    .A2(_3869_));
 sg13g2_a21oi_1 _8327_ (.A1(net1835),
    .A2(_3870_),
    .Y(_3871_),
    .B1(_2926_));
 sg13g2_o21ai_1 _8328_ (.B1(_2940_),
    .Y(_3872_),
    .A1(net1722),
    .A2(_3871_));
 sg13g2_nand2_1 _8329_ (.Y(_3873_),
    .A(net1690),
    .B(_3872_));
 sg13g2_o21ai_1 _8330_ (.B1(_3873_),
    .Y(_3874_),
    .A1(_0745_),
    .A2(net1691));
 sg13g2_a21oi_1 _8331_ (.A1(net1715),
    .A2(_3867_),
    .Y(_3875_),
    .B1(net1698));
 sg13g2_o21ai_1 _8332_ (.B1(_3875_),
    .Y(_3876_),
    .A1(net1714),
    .A2(_3874_));
 sg13g2_o21ai_1 _8333_ (.B1(_3876_),
    .Y(_0575_),
    .A1(_0745_),
    .A2(_3660_));
 sg13g2_nand4_1 _8334_ (.B(_3851_),
    .C(_3853_),
    .A(_3838_),
    .Y(_3877_),
    .D(_3866_));
 sg13g2_o21ai_1 _8335_ (.B1(_0180_),
    .Y(_3878_),
    .A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .A2(_0177_));
 sg13g2_nand2_1 _8336_ (.Y(_3879_),
    .A(net1845),
    .B(_3878_));
 sg13g2_xnor2_1 _8337_ (.Y(_3880_),
    .A(\z80.tv80s.i_tv80_core.PC[12] ),
    .B(net1845));
 sg13g2_a21oi_2 _8338_ (.B1(_3880_),
    .Y(_3881_),
    .A2(_3879_),
    .A1(_3877_));
 sg13g2_nand3_1 _8339_ (.B(_3879_),
    .C(_3880_),
    .A(_3877_),
    .Y(_3882_));
 sg13g2_nand2b_1 _8340_ (.Y(_3883_),
    .B(_3882_),
    .A_N(_3881_));
 sg13g2_nor2_1 _8341_ (.A(_0746_),
    .B(net1866),
    .Y(_3884_));
 sg13g2_a21oi_1 _8342_ (.A1(\z80.tv80s.i_tv80_core.I[4] ),
    .A2(net1866),
    .Y(_3885_),
    .B1(_3884_));
 sg13g2_o21ai_1 _8343_ (.B1(_2946_),
    .Y(_3886_),
    .A1(net1756),
    .A2(_3885_));
 sg13g2_a21oi_1 _8344_ (.A1(net1835),
    .A2(_3886_),
    .Y(_3887_),
    .B1(_2970_));
 sg13g2_o21ai_1 _8345_ (.B1(_2972_),
    .Y(_3888_),
    .A1(net1722),
    .A2(_3887_));
 sg13g2_nand2_1 _8346_ (.Y(_3889_),
    .A(net1691),
    .B(_3888_));
 sg13g2_a21oi_1 _8347_ (.A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .A2(net1687),
    .Y(_3890_),
    .B1(net1714));
 sg13g2_a221oi_1 _8348_ (.B2(_3890_),
    .C1(net1698),
    .B1(_3889_),
    .A1(net1714),
    .Y(_3891_),
    .A2(_3883_));
 sg13g2_a21o_1 _8349_ (.A2(net1698),
    .A1(net574),
    .B1(_3891_),
    .X(_0576_));
 sg13g2_nand2_1 _8350_ (.Y(_3892_),
    .A(net543),
    .B(net1695));
 sg13g2_nor2_1 _8351_ (.A(_0183_),
    .B(_3808_),
    .Y(_3893_));
 sg13g2_xnor2_1 _8352_ (.Y(_3894_),
    .A(_0747_),
    .B(net1845));
 sg13g2_o21ai_1 _8353_ (.B1(_3894_),
    .Y(_3895_),
    .A1(_3881_),
    .A2(_3893_));
 sg13g2_or3_1 _8354_ (.A(_3881_),
    .B(_3893_),
    .C(_3894_),
    .X(_3896_));
 sg13g2_a21oi_1 _8355_ (.A1(_3895_),
    .A2(_3896_),
    .Y(_3897_),
    .B1(net1703));
 sg13g2_nor2_1 _8356_ (.A(_0747_),
    .B(net1869),
    .Y(_3898_));
 sg13g2_a21oi_1 _8357_ (.A1(\z80.tv80s.i_tv80_core.I[5] ),
    .A2(net1869),
    .Y(_3899_),
    .B1(_3898_));
 sg13g2_o21ai_1 _8358_ (.B1(_2986_),
    .Y(_3900_),
    .A1(net1757),
    .A2(_3899_));
 sg13g2_a21oi_1 _8359_ (.A1(net1835),
    .A2(_3900_),
    .Y(_3901_),
    .B1(_2985_));
 sg13g2_o21ai_1 _8360_ (.B1(_2999_),
    .Y(_3902_),
    .A1(net1722),
    .A2(_3901_));
 sg13g2_nand2_1 _8361_ (.Y(_3903_),
    .A(net1690),
    .B(_3902_));
 sg13g2_o21ai_1 _8362_ (.B1(_3903_),
    .Y(_3904_),
    .A1(_0747_),
    .A2(net1690));
 sg13g2_o21ai_1 _8363_ (.B1(_3660_),
    .Y(_3905_),
    .A1(net1714),
    .A2(_3904_));
 sg13g2_o21ai_1 _8364_ (.B1(_3892_),
    .Y(_0577_),
    .A1(_3897_),
    .A2(_3905_));
 sg13g2_nand2_1 _8365_ (.Y(_3906_),
    .A(_0767_),
    .B(net1845));
 sg13g2_xnor2_1 _8366_ (.Y(_3907_),
    .A(\z80.tv80s.i_tv80_core.PC[14] ),
    .B(net1845));
 sg13g2_a21oi_1 _8367_ (.A1(_3895_),
    .A2(_3906_),
    .Y(_3908_),
    .B1(_3907_));
 sg13g2_nand3_1 _8368_ (.B(_3906_),
    .C(_3907_),
    .A(_3895_),
    .Y(_3909_));
 sg13g2_nand2b_1 _8369_ (.Y(_3910_),
    .B(_3909_),
    .A_N(_3908_));
 sg13g2_nor2_1 _8370_ (.A(_0748_),
    .B(net1865),
    .Y(_3911_));
 sg13g2_a21oi_1 _8371_ (.A1(\z80.tv80s.i_tv80_core.I[6] ),
    .A2(net1865),
    .Y(_3912_),
    .B1(_3911_));
 sg13g2_o21ai_1 _8372_ (.B1(_3003_),
    .Y(_3913_),
    .A1(net1756),
    .A2(_3912_));
 sg13g2_a21oi_1 _8373_ (.A1(net1837),
    .A2(_3913_),
    .Y(_3914_),
    .B1(_3027_));
 sg13g2_o21ai_1 _8374_ (.B1(_3029_),
    .Y(_3915_),
    .A1(net1721),
    .A2(_3914_));
 sg13g2_nand2_1 _8375_ (.Y(_3916_),
    .A(net1690),
    .B(_3915_));
 sg13g2_a21oi_1 _8376_ (.A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .A2(net1687),
    .Y(_3917_),
    .B1(net1714));
 sg13g2_a221oi_1 _8377_ (.B2(_3917_),
    .C1(net1695),
    .B1(_3916_),
    .A1(net1714),
    .Y(_3918_),
    .A2(_3910_));
 sg13g2_a21o_1 _8378_ (.A2(net1695),
    .A1(net589),
    .B1(_3918_),
    .X(_0578_));
 sg13g2_nand4_1 _8379_ (.B(\z80.tv80s.i_tv80_core.PC[14] ),
    .C(_3808_),
    .A(\z80.tv80s.i_tv80_core.PC[13] ),
    .Y(_3919_),
    .D(_3881_));
 sg13g2_nand2_1 _8380_ (.Y(_3920_),
    .A(_0189_),
    .B(net1845));
 sg13g2_o21ai_1 _8381_ (.B1(_3919_),
    .Y(_3921_),
    .A1(_3908_),
    .A2(_3920_));
 sg13g2_xnor2_1 _8382_ (.Y(_3922_),
    .A(\z80.tv80s.i_tv80_core.PC[15] ),
    .B(_3921_));
 sg13g2_nor2_1 _8383_ (.A(_0750_),
    .B(net1865),
    .Y(_3923_));
 sg13g2_a21oi_1 _8384_ (.A1(\z80.tv80s.i_tv80_core.I[7] ),
    .A2(net1865),
    .Y(_3924_),
    .B1(_3923_));
 sg13g2_o21ai_1 _8385_ (.B1(_3043_),
    .Y(_3925_),
    .A1(net1756),
    .A2(_3924_));
 sg13g2_a21oi_1 _8386_ (.A1(net1837),
    .A2(_3925_),
    .Y(_3926_),
    .B1(_3042_));
 sg13g2_o21ai_1 _8387_ (.B1(_3056_),
    .Y(_3927_),
    .A1(net1721),
    .A2(_3926_));
 sg13g2_nand2_1 _8388_ (.Y(_3928_),
    .A(net1690),
    .B(_3927_));
 sg13g2_o21ai_1 _8389_ (.B1(_3928_),
    .Y(_3929_),
    .A1(_0750_),
    .A2(net1690));
 sg13g2_a21oi_1 _8390_ (.A1(net1714),
    .A2(_3922_),
    .Y(_3930_),
    .B1(net1695));
 sg13g2_o21ai_1 _8391_ (.B1(_3930_),
    .Y(_3931_),
    .A1(net1716),
    .A2(_3929_));
 sg13g2_o21ai_1 _8392_ (.B1(_3931_),
    .Y(_0579_),
    .A1(_0750_),
    .A2(_3660_));
 sg13g2_nand4_1 _8393_ (.B(net1995),
    .C(_1716_),
    .A(net1903),
    .Y(_3932_),
    .D(_2482_));
 sg13g2_mux2_1 _8394_ (.A0(_0020_),
    .A1(net532),
    .S(_3932_),
    .X(_0580_));
 sg13g2_and2_1 _8395_ (.A(net2106),
    .B(net2144),
    .X(_3933_));
 sg13g2_nand2_1 _8396_ (.Y(_3934_),
    .A(net2106),
    .B(net2144));
 sg13g2_or2_2 _8397_ (.X(_3935_),
    .B(_2596_),
    .A(net1997));
 sg13g2_nand3_1 _8398_ (.B(net1915),
    .C(net1792),
    .A(net2136),
    .Y(_3936_));
 sg13g2_o21ai_1 _8399_ (.B1(_3936_),
    .Y(_3937_),
    .A1(_3427_),
    .A2(net1916));
 sg13g2_nand2_1 _8400_ (.Y(_3938_),
    .A(net1901),
    .B(_3937_));
 sg13g2_nand2_1 _8401_ (.Y(_3939_),
    .A(net2114),
    .B(_1277_));
 sg13g2_a22oi_1 _8402_ (.Y(_3940_),
    .B1(_1673_),
    .B2(_3939_),
    .A2(_1200_),
    .A1(_1189_));
 sg13g2_nand2b_1 _8403_ (.Y(_3941_),
    .B(_0924_),
    .A_N(_3661_));
 sg13g2_o21ai_1 _8404_ (.B1(net2118),
    .Y(_3942_),
    .A1(_1677_),
    .A2(_3941_));
 sg13g2_nor2_1 _8405_ (.A(_1244_),
    .B(_2481_),
    .Y(_3943_));
 sg13g2_nor4_2 _8406_ (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(_0028_),
    .C(_0874_),
    .Y(_3944_),
    .D(_1018_));
 sg13g2_nand4_1 _8407_ (.B(_1233_),
    .C(_2352_),
    .A(_1015_),
    .Y(_3945_),
    .D(_3944_));
 sg13g2_nand3_1 _8408_ (.B(_2478_),
    .C(_2479_),
    .A(_1162_),
    .Y(_3946_));
 sg13g2_nor3_1 _8409_ (.A(_3941_),
    .B(_3945_),
    .C(_3946_),
    .Y(_3947_));
 sg13g2_nand4_1 _8410_ (.B(_1713_),
    .C(_3943_),
    .A(_0998_),
    .Y(_3948_),
    .D(_3947_));
 sg13g2_o21ai_1 _8411_ (.B1(_3942_),
    .Y(_3949_),
    .A1(_2598_),
    .A2(_3948_));
 sg13g2_a21oi_2 _8412_ (.B1(_3940_),
    .Y(_3950_),
    .A2(_3949_),
    .A1(net2168));
 sg13g2_nor2_1 _8413_ (.A(_0682_),
    .B(_3950_),
    .Y(_3951_));
 sg13g2_nand2b_2 _8414_ (.Y(_3952_),
    .B(net2143),
    .A_N(_3950_));
 sg13g2_nand3_1 _8415_ (.B(_0693_),
    .C(_2604_),
    .A(_0016_),
    .Y(_3953_));
 sg13g2_nand2_1 _8416_ (.Y(_3954_),
    .A(_0820_),
    .B(_3953_));
 sg13g2_a21oi_2 _8417_ (.B1(_3954_),
    .Y(_3955_),
    .A2(\z80.tv80s.i_tv80_core.IStatus[2] ),
    .A1(\z80.tv80s.i_tv80_core.IntCycle ));
 sg13g2_mux2_1 _8418_ (.A0(net2136),
    .A1(net5),
    .S(net1855),
    .X(_3956_));
 sg13g2_a21oi_1 _8419_ (.A1(net1912),
    .A2(_3956_),
    .Y(_3957_),
    .B1(net1755));
 sg13g2_o21ai_1 _8420_ (.B1(net1995),
    .Y(_3958_),
    .A1(_3424_),
    .A2(_3950_));
 sg13g2_a21oi_1 _8421_ (.A1(_3938_),
    .A2(_3957_),
    .Y(_3959_),
    .B1(_3958_));
 sg13g2_a21o_1 _8422_ (.A2(net1979),
    .A1(net2136),
    .B1(_3959_),
    .X(_0581_));
 sg13g2_nand3_1 _8423_ (.B(net1916),
    .C(net1793),
    .A(net2135),
    .Y(_3960_));
 sg13g2_o21ai_1 _8424_ (.B1(_3960_),
    .Y(_3961_),
    .A1(_3446_),
    .A2(net1916));
 sg13g2_nand2_1 _8425_ (.Y(_3962_),
    .A(net1901),
    .B(_3961_));
 sg13g2_mux2_1 _8426_ (.A0(net2135),
    .A1(net6),
    .S(net1855),
    .X(_3963_));
 sg13g2_a21oi_1 _8427_ (.A1(net1912),
    .A2(_3963_),
    .Y(_3964_),
    .B1(net1755));
 sg13g2_o21ai_1 _8428_ (.B1(net1995),
    .Y(_3965_),
    .A1(net2050),
    .A2(_3952_));
 sg13g2_a21oi_1 _8429_ (.A1(_3962_),
    .A2(_3964_),
    .Y(_3966_),
    .B1(_3965_));
 sg13g2_a21o_1 _8430_ (.A2(net1979),
    .A1(net2135),
    .B1(_3966_),
    .X(_0582_));
 sg13g2_nand3_1 _8431_ (.B(net1915),
    .C(net1792),
    .A(net2134),
    .Y(_3967_));
 sg13g2_o21ai_1 _8432_ (.B1(_3967_),
    .Y(_3968_),
    .A1(_3458_),
    .A2(net1915));
 sg13g2_nand2b_1 _8433_ (.Y(_3969_),
    .B(net1855),
    .A_N(net7));
 sg13g2_o21ai_1 _8434_ (.B1(_3969_),
    .Y(_3970_),
    .A1(net2134),
    .A2(net1855));
 sg13g2_a21oi_1 _8435_ (.A1(net1911),
    .A2(_3970_),
    .Y(_3971_),
    .B1(net1755));
 sg13g2_o21ai_1 _8436_ (.B1(_3971_),
    .Y(_3972_),
    .A1(net1909),
    .A2(_3968_));
 sg13g2_a21oi_1 _8437_ (.A1(net552),
    .A2(net1755),
    .Y(_3973_),
    .B1(net1976));
 sg13g2_a22oi_1 _8438_ (.Y(_0583_),
    .B1(_3972_),
    .B2(_3973_),
    .A2(net1975),
    .A1(_0763_));
 sg13g2_o21ai_1 _8439_ (.B1(net1915),
    .Y(_3974_),
    .A1(net2079),
    .A2(net1793));
 sg13g2_a21oi_1 _8440_ (.A1(_0762_),
    .A2(net1792),
    .Y(_3975_),
    .B1(_3974_));
 sg13g2_a21oi_1 _8441_ (.A1(_3472_),
    .A2(net1919),
    .Y(_3976_),
    .B1(_3975_));
 sg13g2_nor2_1 _8442_ (.A(net1909),
    .B(_3976_),
    .Y(_3977_));
 sg13g2_mux2_1 _8443_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A1(net8),
    .S(net1855),
    .X(_3978_));
 sg13g2_a21oi_1 _8444_ (.A1(net1911),
    .A2(_3978_),
    .Y(_3979_),
    .B1(_3977_));
 sg13g2_a21oi_1 _8445_ (.A1(net2048),
    .A2(net1755),
    .Y(_3980_),
    .B1(net1975));
 sg13g2_o21ai_1 _8446_ (.B1(_3980_),
    .Y(_3981_),
    .A1(net1755),
    .A2(_3979_));
 sg13g2_o21ai_1 _8447_ (.B1(_3981_),
    .Y(_3982_),
    .A1(net597),
    .A2(net1991));
 sg13g2_inv_1 _8448_ (.Y(_0584_),
    .A(_3982_));
 sg13g2_nand2_1 _8449_ (.Y(_3983_),
    .A(net556),
    .B(net1975));
 sg13g2_nand2_1 _8450_ (.Y(_3984_),
    .A(_3486_),
    .B(net1919));
 sg13g2_nor2_1 _8451_ (.A(net2021),
    .B(net1792),
    .Y(_3985_));
 sg13g2_a21oi_1 _8452_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net1793),
    .Y(_3986_),
    .B1(_3985_));
 sg13g2_a21oi_1 _8453_ (.A1(net1916),
    .A2(_3986_),
    .Y(_3987_),
    .B1(net1912));
 sg13g2_mux2_1 _8454_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A1(net9),
    .S(_3955_),
    .X(_3988_));
 sg13g2_a221oi_1 _8455_ (.B2(net1912),
    .C1(_3951_),
    .B1(_3988_),
    .A1(_3984_),
    .Y(_3989_),
    .A2(_3987_));
 sg13g2_o21ai_1 _8456_ (.B1(net1995),
    .Y(_3990_),
    .A1(net2047),
    .A2(_3952_));
 sg13g2_o21ai_1 _8457_ (.B1(_3983_),
    .Y(_0585_),
    .A1(_3989_),
    .A2(_3990_));
 sg13g2_nand2_1 _8458_ (.Y(_3991_),
    .A(net2133),
    .B(net1975));
 sg13g2_nand2_1 _8459_ (.Y(_3992_),
    .A(_3501_),
    .B(net1919));
 sg13g2_nand2b_1 _8460_ (.Y(_3993_),
    .B(net1792),
    .A_N(net2133));
 sg13g2_o21ai_1 _8461_ (.B1(_3993_),
    .Y(_3994_),
    .A1(net2063),
    .A2(net1792));
 sg13g2_a21oi_1 _8462_ (.A1(net1916),
    .A2(_3994_),
    .Y(_3995_),
    .B1(net1912));
 sg13g2_mux2_1 _8463_ (.A0(net2133),
    .A1(net10),
    .S(net1855),
    .X(_3996_));
 sg13g2_a221oi_1 _8464_ (.B2(net1912),
    .C1(_3951_),
    .B1(_3996_),
    .A1(_3992_),
    .Y(_3997_),
    .A2(_3995_));
 sg13g2_o21ai_1 _8465_ (.B1(net1995),
    .Y(_3998_),
    .A1(\z80.tv80s.di_reg[5] ),
    .A2(_3952_));
 sg13g2_o21ai_1 _8466_ (.B1(_3991_),
    .Y(_0586_),
    .A1(_3997_),
    .A2(_3998_));
 sg13g2_nand3_1 _8467_ (.B(net1915),
    .C(net1792),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .Y(_3999_));
 sg13g2_o21ai_1 _8468_ (.B1(_3999_),
    .Y(_4000_),
    .A1(_3516_),
    .A2(net1915));
 sg13g2_nand2_1 _8469_ (.Y(_4001_),
    .A(net1901),
    .B(_4000_));
 sg13g2_mux2_1 _8470_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A1(net11),
    .S(_3955_),
    .X(_4002_));
 sg13g2_a21oi_1 _8471_ (.A1(net1912),
    .A2(_4002_),
    .Y(_4003_),
    .B1(net1755));
 sg13g2_a221oi_1 _8472_ (.B2(_4003_),
    .C1(net1975),
    .B1(_4001_),
    .A1(_0719_),
    .Y(_4004_),
    .A2(_3951_));
 sg13g2_a21o_1 _8473_ (.A2(net1975),
    .A1(net573),
    .B1(_4004_),
    .X(_0587_));
 sg13g2_nand2_1 _8474_ (.Y(_4005_),
    .A(net584),
    .B(net1975));
 sg13g2_nand3_1 _8475_ (.B(net1915),
    .C(net1792),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .Y(_4006_));
 sg13g2_o21ai_1 _8476_ (.B1(_4006_),
    .Y(_4007_),
    .A1(_3530_),
    .A2(net1915));
 sg13g2_or2_1 _8477_ (.X(_4008_),
    .B(net1855),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sg13g2_a21oi_1 _8478_ (.A1(_0794_),
    .A2(net1855),
    .Y(_4009_),
    .B1(net1901));
 sg13g2_a221oi_1 _8479_ (.B2(_4009_),
    .C1(net1755),
    .B1(_4008_),
    .A1(net1901),
    .Y(_4010_),
    .A2(_4007_));
 sg13g2_o21ai_1 _8480_ (.B1(net1995),
    .Y(_4011_),
    .A1(net2044),
    .A2(_3952_));
 sg13g2_o21ai_1 _8481_ (.B1(_4005_),
    .Y(_0588_),
    .A1(_4010_),
    .A2(_4011_));
 sg13g2_nand3_1 _8482_ (.B(_1160_),
    .C(_3943_),
    .A(net2170),
    .Y(_4012_));
 sg13g2_nor2_1 _8483_ (.A(_2480_),
    .B(_4012_),
    .Y(_4013_));
 sg13g2_nand3_1 _8484_ (.B(_3677_),
    .C(_4013_),
    .A(_2599_),
    .Y(_4014_));
 sg13g2_o21ai_1 _8485_ (.B1(_1278_),
    .Y(_4015_),
    .A1(_3667_),
    .A2(_4014_));
 sg13g2_nand3_1 _8486_ (.B(net1889),
    .C(_4015_),
    .A(net2144),
    .Y(_4016_));
 sg13g2_inv_1 _8487_ (.Y(_4017_),
    .A(net1767));
 sg13g2_nand2b_1 _8488_ (.Y(_4018_),
    .B(net1911),
    .A_N(\z80.tv80s.i_tv80_core.TmpAddr[8] ));
 sg13g2_nand3_1 _8489_ (.B(net1918),
    .C(net1794),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .Y(_4019_));
 sg13g2_o21ai_1 _8490_ (.B1(_4019_),
    .Y(_4020_),
    .A1(_3543_),
    .A2(_3934_));
 sg13g2_o21ai_1 _8491_ (.B1(_4018_),
    .Y(_4021_),
    .A1(net1911),
    .A2(_4020_));
 sg13g2_o21ai_1 _8492_ (.B1(net1991),
    .Y(_4022_),
    .A1(net2051),
    .A2(net1767));
 sg13g2_a21oi_1 _8493_ (.A1(net1767),
    .A2(_4021_),
    .Y(_4023_),
    .B1(_4022_));
 sg13g2_a21o_1 _8494_ (.A2(net1979),
    .A1(net561),
    .B1(_4023_),
    .X(_0589_));
 sg13g2_nor2_1 _8495_ (.A(net557),
    .B(net1991),
    .Y(_4024_));
 sg13g2_and2_1 _8496_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .B(net1918),
    .X(_4025_));
 sg13g2_a221oi_1 _8497_ (.B2(_4025_),
    .C1(net1911),
    .B1(net1794),
    .A1(_3558_),
    .Y(_4026_),
    .A2(_3933_));
 sg13g2_o21ai_1 _8498_ (.B1(net1768),
    .Y(_4027_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .A2(net1902));
 sg13g2_nor2_1 _8499_ (.A(_4026_),
    .B(_4027_),
    .Y(_4028_));
 sg13g2_a21oi_1 _8500_ (.A1(net2050),
    .A2(_4017_),
    .Y(_4029_),
    .B1(_4028_));
 sg13g2_a21oi_1 _8501_ (.A1(net1990),
    .A2(_4029_),
    .Y(_0590_),
    .B1(_4024_));
 sg13g2_nand2_1 _8502_ (.Y(_4030_),
    .A(_3571_),
    .B(net1919));
 sg13g2_nand3_1 _8503_ (.B(net1918),
    .C(net1794),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .Y(_4031_));
 sg13g2_nand3_1 _8504_ (.B(_4030_),
    .C(_4031_),
    .A(net1903),
    .Y(_4032_));
 sg13g2_o21ai_1 _8505_ (.B1(_4032_),
    .Y(_4033_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(net1902));
 sg13g2_o21ai_1 _8506_ (.B1(net1990),
    .Y(_4034_),
    .A1(net2049),
    .A2(net1767));
 sg13g2_a21oi_1 _8507_ (.A1(net1767),
    .A2(_4033_),
    .Y(_4035_),
    .B1(_4034_));
 sg13g2_a21o_1 _8508_ (.A2(net1978),
    .A1(net534),
    .B1(_4035_),
    .X(_0591_));
 sg13g2_nand2_1 _8509_ (.Y(_4036_),
    .A(_3583_),
    .B(net1919));
 sg13g2_nand3_1 _8510_ (.B(net1918),
    .C(net1794),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .Y(_4037_));
 sg13g2_nand3_1 _8511_ (.B(_4036_),
    .C(_4037_),
    .A(net1902),
    .Y(_4038_));
 sg13g2_o21ai_1 _8512_ (.B1(_4038_),
    .Y(_4039_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2(net1902));
 sg13g2_o21ai_1 _8513_ (.B1(net1990),
    .Y(_4040_),
    .A1(net2048),
    .A2(net1767));
 sg13g2_a21oi_1 _8514_ (.A1(net1767),
    .A2(_4039_),
    .Y(_4041_),
    .B1(_4040_));
 sg13g2_a21o_1 _8515_ (.A2(net1978),
    .A1(net539),
    .B1(_4041_),
    .X(_0592_));
 sg13g2_nand2_1 _8516_ (.Y(_4042_),
    .A(_3599_),
    .B(net1919));
 sg13g2_nand3_1 _8517_ (.B(net1918),
    .C(net1794),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .Y(_4043_));
 sg13g2_nand3_1 _8518_ (.B(_4042_),
    .C(_4043_),
    .A(net1902),
    .Y(_4044_));
 sg13g2_o21ai_1 _8519_ (.B1(_4044_),
    .Y(_4045_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(net1902));
 sg13g2_o21ai_1 _8520_ (.B1(net1990),
    .Y(_4046_),
    .A1(net2047),
    .A2(net1768));
 sg13g2_a21oi_1 _8521_ (.A1(net1768),
    .A2(_4045_),
    .Y(_4047_),
    .B1(_4046_));
 sg13g2_a21o_1 _8522_ (.A2(net1977),
    .A1(net513),
    .B1(_4047_),
    .X(_0593_));
 sg13g2_nor2_1 _8523_ (.A(net535),
    .B(net1990),
    .Y(_4048_));
 sg13g2_and2_1 _8524_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .B(net1918),
    .X(_4049_));
 sg13g2_a221oi_1 _8525_ (.B2(_4049_),
    .C1(net1914),
    .B1(net1794),
    .A1(_3612_),
    .Y(_4050_),
    .A2(net1919));
 sg13g2_o21ai_1 _8526_ (.B1(net1767),
    .Y(_4051_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(net1902));
 sg13g2_nor2_1 _8527_ (.A(_4050_),
    .B(_4051_),
    .Y(_4052_));
 sg13g2_a21oi_1 _8528_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_4017_),
    .Y(_4053_),
    .B1(_4052_));
 sg13g2_a21oi_1 _8529_ (.A1(net1990),
    .A2(_4053_),
    .Y(_0594_),
    .B1(_4048_));
 sg13g2_nand2_1 _8530_ (.Y(_4054_),
    .A(net464),
    .B(net1977));
 sg13g2_nor2_1 _8531_ (.A(net464),
    .B(net1900),
    .Y(_4055_));
 sg13g2_and2_1 _8532_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .B(net1917),
    .X(_4056_));
 sg13g2_a221oi_1 _8533_ (.B2(_4056_),
    .C1(net1914),
    .B1(net1794),
    .A1(_3625_),
    .Y(_4057_),
    .A2(net1919));
 sg13g2_o21ai_1 _8534_ (.B1(net1768),
    .Y(_4058_),
    .A1(_4055_),
    .A2(_4057_));
 sg13g2_o21ai_1 _8535_ (.B1(_4058_),
    .Y(_4059_),
    .A1(net2045),
    .A2(net1768));
 sg13g2_o21ai_1 _8536_ (.B1(_4054_),
    .Y(_0595_),
    .A1(net1977),
    .A2(_4059_));
 sg13g2_nand3_1 _8537_ (.B(net1918),
    .C(net1794),
    .A(net507),
    .Y(_4060_));
 sg13g2_o21ai_1 _8538_ (.B1(_4060_),
    .Y(_4061_),
    .A1(_3638_),
    .A2(net1917));
 sg13g2_o21ai_1 _8539_ (.B1(net1768),
    .Y(_4062_),
    .A1(net507),
    .A2(net1902));
 sg13g2_inv_1 _8540_ (.Y(_4063_),
    .A(_4062_));
 sg13g2_o21ai_1 _8541_ (.B1(_4063_),
    .Y(_4064_),
    .A1(net1911),
    .A2(_4061_));
 sg13g2_a21oi_1 _8542_ (.A1(net2044),
    .A2(_4017_),
    .Y(_4065_),
    .B1(net1977));
 sg13g2_a22oi_1 _8543_ (.Y(_0596_),
    .B1(_4064_),
    .B2(_4065_),
    .A2(net1977),
    .A1(_0768_));
 sg13g2_nand2_1 _8544_ (.Y(_4066_),
    .A(_0236_),
    .B(_0237_));
 sg13g2_nor2_1 _8545_ (.A(_0236_),
    .B(_0237_),
    .Y(_4067_));
 sg13g2_nand2_1 _8546_ (.Y(_4068_),
    .A(_0805_),
    .B(_4067_));
 sg13g2_o21ai_1 _8547_ (.B1(net2104),
    .Y(_4069_),
    .A1(_0238_),
    .A2(_4066_));
 sg13g2_a21oi_1 _8548_ (.A1(_4066_),
    .A2(_4068_),
    .Y(_4070_),
    .B1(_4069_));
 sg13g2_and2_1 _8549_ (.A(_1134_),
    .B(_2496_),
    .X(_4071_));
 sg13g2_o21ai_1 _8550_ (.B1(_2498_),
    .Y(_4072_),
    .A1(net461),
    .A2(net1679));
 sg13g2_a21oi_1 _8551_ (.A1(_4070_),
    .A2(_4071_),
    .Y(_0597_),
    .B1(_4072_));
 sg13g2_nor3_1 _8552_ (.A(net2025),
    .B(_0804_),
    .C(_0237_),
    .Y(_4073_));
 sg13g2_a22oi_1 _8553_ (.Y(_4074_),
    .B1(_0805_),
    .B2(_4073_),
    .A2(net2124),
    .A1(net2025));
 sg13g2_or2_1 _8554_ (.X(_4075_),
    .B(_2495_),
    .A(_1338_));
 sg13g2_nor2_1 _8555_ (.A(_4074_),
    .B(_4075_),
    .Y(_4076_));
 sg13g2_mux2_1 _8556_ (.A0(net2121),
    .A1(_4076_),
    .S(_1135_),
    .X(_0598_));
 sg13g2_and4_1 _8557_ (.A(net2103),
    .B(_0804_),
    .C(_0237_),
    .D(_0805_),
    .X(_4077_));
 sg13g2_a21o_1 _8558_ (.A2(_2494_),
    .A1(_1074_),
    .B1(_4077_),
    .X(_4078_));
 sg13g2_nand3_1 _8559_ (.B(_2496_),
    .C(_4078_),
    .A(_1134_),
    .Y(_4079_));
 sg13g2_o21ai_1 _8560_ (.B1(_4079_),
    .Y(_0599_),
    .A1(_0679_),
    .A2(net1679));
 sg13g2_o21ai_1 _8561_ (.B1(_4069_),
    .Y(_4080_),
    .A1(net2103),
    .A2(net2110));
 sg13g2_nor2_1 _8562_ (.A(_4075_),
    .B(_4080_),
    .Y(_4081_));
 sg13g2_mux2_1 _8563_ (.A0(net2107),
    .A1(_4081_),
    .S(net1679),
    .X(_0600_));
 sg13g2_nand3_1 _8564_ (.B(_0238_),
    .C(_4067_),
    .A(net2103),
    .Y(_4082_));
 sg13g2_a21oi_1 _8565_ (.A1(_1340_),
    .A2(_4082_),
    .Y(_4083_),
    .B1(_4075_));
 sg13g2_mux2_1 _8566_ (.A0(net554),
    .A1(_4083_),
    .S(net1679),
    .X(_0601_));
 sg13g2_nor2_1 _8567_ (.A(net2103),
    .B(net627),
    .Y(_4084_));
 sg13g2_a221oi_1 _8568_ (.B2(_2494_),
    .C1(_1338_),
    .B1(_4084_),
    .A1(_0238_),
    .Y(_4085_),
    .A2(_4073_));
 sg13g2_nor2_1 _8569_ (.A(net2106),
    .B(net1679),
    .Y(_4086_));
 sg13g2_a21oi_2 _8570_ (.B1(_4086_),
    .Y(_0602_),
    .A2(_4085_),
    .A1(net1679));
 sg13g2_nand4_1 _8571_ (.B(_0804_),
    .C(net586),
    .A(net2103),
    .Y(_4087_),
    .D(_0238_));
 sg13g2_a21oi_1 _8572_ (.A1(_1353_),
    .A2(net587),
    .Y(_4088_),
    .B1(_4075_));
 sg13g2_nand2_1 _8573_ (.Y(_4089_),
    .A(net1679),
    .B(_4088_));
 sg13g2_o21ai_1 _8574_ (.B1(_4089_),
    .Y(_0603_),
    .A1(net2025),
    .A2(net1679));
 sg13g2_a21oi_1 _8575_ (.A1(net2105),
    .A2(net2166),
    .Y(_4090_),
    .B1(net1913));
 sg13g2_nor3_1 _8576_ (.A(net1997),
    .B(net1980),
    .C(_4090_),
    .Y(_4091_));
 sg13g2_nand3_1 _8577_ (.B(net484),
    .C(net1913),
    .A(\z80.tv80s.i_tv80_core.IntCycle ),
    .Y(_4092_));
 sg13g2_and2_2 _8578_ (.A(net1854),
    .B(_4092_),
    .X(_4093_));
 sg13g2_nand2_2 _8579_ (.Y(_4094_),
    .A(net1913),
    .B(_3953_));
 sg13g2_nand2_1 _8580_ (.Y(_4095_),
    .A(net5),
    .B(_4094_));
 sg13g2_nor2_1 _8581_ (.A(net2102),
    .B(net1854),
    .Y(_4096_));
 sg13g2_a21oi_1 _8582_ (.A1(_4093_),
    .A2(_4095_),
    .Y(_0604_),
    .B1(_4096_));
 sg13g2_nand2_1 _8583_ (.Y(_4097_),
    .A(net6),
    .B(_4094_));
 sg13g2_nor2_1 _8584_ (.A(net2097),
    .B(net1854),
    .Y(_4098_));
 sg13g2_a21oi_1 _8585_ (.A1(_4093_),
    .A2(_4097_),
    .Y(_0605_),
    .B1(_4098_));
 sg13g2_nand2_1 _8586_ (.Y(_4099_),
    .A(net7),
    .B(_4094_));
 sg13g2_nor2_1 _8587_ (.A(net2093),
    .B(net1854),
    .Y(_4100_));
 sg13g2_a21oi_1 _8588_ (.A1(_4093_),
    .A2(_4099_),
    .Y(_0606_),
    .B1(_4100_));
 sg13g2_nand2_1 _8589_ (.Y(_4101_),
    .A(net8),
    .B(_4094_));
 sg13g2_nor2_1 _8590_ (.A(net2079),
    .B(net1854),
    .Y(_4102_));
 sg13g2_a21oi_1 _8591_ (.A1(_4093_),
    .A2(_4101_),
    .Y(_0607_),
    .B1(_4102_));
 sg13g2_nand2_1 _8592_ (.Y(_4103_),
    .A(net9),
    .B(_4094_));
 sg13g2_nor2_1 _8593_ (.A(net2072),
    .B(net1854),
    .Y(_4104_));
 sg13g2_a21oi_1 _8594_ (.A1(_4093_),
    .A2(_4103_),
    .Y(_0608_),
    .B1(_4104_));
 sg13g2_nand2_1 _8595_ (.Y(_4105_),
    .A(net10),
    .B(_4094_));
 sg13g2_nor2_1 _8596_ (.A(net2069),
    .B(net1854),
    .Y(_4106_));
 sg13g2_a21oi_1 _8597_ (.A1(_4093_),
    .A2(_4105_),
    .Y(_0609_),
    .B1(_4106_));
 sg13g2_nand2_1 _8598_ (.Y(_4107_),
    .A(net11),
    .B(_4094_));
 sg13g2_nor2_1 _8599_ (.A(net2059),
    .B(_4091_),
    .Y(_4108_));
 sg13g2_a21oi_2 _8600_ (.B1(_4108_),
    .Y(_0610_),
    .A2(_4107_),
    .A1(_4093_));
 sg13g2_nand2_1 _8601_ (.Y(_4109_),
    .A(net12),
    .B(_4094_));
 sg13g2_nor2_1 _8602_ (.A(net2057),
    .B(net1854),
    .Y(_4110_));
 sg13g2_a21oi_2 _8603_ (.B1(_4110_),
    .Y(_0611_),
    .A2(_4109_),
    .A1(_4093_));
 sg13g2_o21ai_1 _8604_ (.B1(_1133_),
    .Y(_4111_),
    .A1(\z80.m1_n ),
    .A2(_0833_));
 sg13g2_nand2b_1 _8605_ (.Y(_4112_),
    .B(_1344_),
    .A_N(\z80.m1_n ));
 sg13g2_nand2_1 _8606_ (.Y(_4113_),
    .A(_1345_),
    .B(_4112_));
 sg13g2_o21ai_1 _8607_ (.B1(_4113_),
    .Y(_4114_),
    .A1(_2497_),
    .A2(_4111_));
 sg13g2_nor3_1 _8608_ (.A(\z80.m1_n ),
    .B(_0833_),
    .C(_1344_),
    .Y(_4115_));
 sg13g2_nor3_1 _8609_ (.A(net2183),
    .B(\z80.tv80s.i_tv80_core.ts[0] ),
    .C(_4115_),
    .Y(_4116_));
 sg13g2_a22oi_1 _8610_ (.Y(_0612_),
    .B1(_4114_),
    .B2(_4116_),
    .A2(net2182),
    .A1(_0654_));
 sg13g2_o21ai_1 _8611_ (.B1(_0834_),
    .Y(_4117_),
    .A1(_0837_),
    .A2(_0841_));
 sg13g2_nor3_1 _8612_ (.A(net2063),
    .B(_0843_),
    .C(_4117_),
    .Y(_4118_));
 sg13g2_a21o_1 _8613_ (.A2(_4117_),
    .A1(net499),
    .B1(_4118_),
    .X(_0613_));
 sg13g2_nor4_1 _8614_ (.A(net2060),
    .B(_0843_),
    .C(_1041_),
    .D(_4117_),
    .Y(_4119_));
 sg13g2_a21o_1 _8615_ (.A2(_4117_),
    .A1(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .B1(_4119_),
    .X(_0614_));
 sg13g2_nor2_1 _8616_ (.A(net1900),
    .B(_0837_),
    .Y(_4120_));
 sg13g2_nand2_1 _8617_ (.Y(_4121_),
    .A(_0826_),
    .B(_3700_));
 sg13g2_o21ai_1 _8618_ (.B1(net2053),
    .Y(_4122_),
    .A1(_4120_),
    .A2(_4121_));
 sg13g2_o21ai_1 _8619_ (.B1(_4122_),
    .Y(_0615_),
    .A1(net185),
    .A2(_0825_));
 sg13g2_nand3_1 _8620_ (.B(_0865_),
    .C(_1685_),
    .A(_0671_),
    .Y(_4123_));
 sg13g2_nor3_2 _8621_ (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .B(_2634_),
    .C(_4123_),
    .Y(_4124_));
 sg13g2_a21o_1 _8622_ (.A2(net1686),
    .A1(net448),
    .B1(_4124_),
    .X(_0616_));
 sg13g2_mux2_1 _8623_ (.A0(net5),
    .A1(net2051),
    .S(net1894),
    .X(_0617_));
 sg13g2_mux2_1 _8624_ (.A0(net6),
    .A1(net2050),
    .S(_0824_),
    .X(_0618_));
 sg13g2_mux2_1 _8625_ (.A0(net7),
    .A1(net2049),
    .S(_0824_),
    .X(_0619_));
 sg13g2_nor2_1 _8626_ (.A(net8),
    .B(net1894),
    .Y(_4125_));
 sg13g2_a21oi_1 _8627_ (.A1(_0705_),
    .A2(net1894),
    .Y(_0620_),
    .B1(_4125_));
 sg13g2_mux2_1 _8628_ (.A0(net9),
    .A1(net2047),
    .S(net1894),
    .X(_0621_));
 sg13g2_mux2_1 _8629_ (.A0(net10),
    .A1(net2046),
    .S(net1894),
    .X(_0622_));
 sg13g2_nor2_1 _8630_ (.A(net11),
    .B(net1894),
    .Y(_4126_));
 sg13g2_a21oi_1 _8631_ (.A1(_0719_),
    .A2(net1894),
    .Y(_0623_),
    .B1(_4126_));
 sg13g2_mux2_1 _8632_ (.A0(net12),
    .A1(net2043),
    .S(net1894),
    .X(_0624_));
 sg13g2_nand2_1 _8633_ (.Y(_4127_),
    .A(net466),
    .B(net1963));
 sg13g2_a21oi_1 _8634_ (.A1(net2102),
    .A2(net2166),
    .Y(_4128_),
    .B1(net1952));
 sg13g2_o21ai_1 _8635_ (.B1(_1268_),
    .Y(_4129_),
    .A1(net2023),
    .A2(_1548_));
 sg13g2_o21ai_1 _8636_ (.B1(_1298_),
    .Y(_4130_),
    .A1(net2023),
    .A2(_0931_));
 sg13g2_a21oi_1 _8637_ (.A1(net2110),
    .A2(net1935),
    .Y(_4131_),
    .B1(net2115));
 sg13g2_a21oi_2 _8638_ (.B1(_4131_),
    .Y(_4132_),
    .A2(net1935),
    .A1(net2115));
 sg13g2_a21oi_1 _8639_ (.A1(_1014_),
    .A2(_1647_),
    .Y(_4133_),
    .B1(net2112));
 sg13g2_a221oi_1 _8640_ (.B2(_1244_),
    .C1(_4133_),
    .B1(_4132_),
    .A1(net2118),
    .Y(_4134_),
    .A2(_4130_));
 sg13g2_nor3_1 _8641_ (.A(_0872_),
    .B(_0924_),
    .C(_1038_),
    .Y(_4135_));
 sg13g2_nor3_1 _8642_ (.A(_0034_),
    .B(net1883),
    .C(net1875),
    .Y(_4136_));
 sg13g2_nor3_1 _8643_ (.A(net2014),
    .B(net1934),
    .C(_1647_),
    .Y(_4137_));
 sg13g2_nor4_1 _8644_ (.A(_1621_),
    .B(_4135_),
    .C(_4136_),
    .D(_4137_),
    .Y(_4138_));
 sg13g2_nand3_1 _8645_ (.B(_4134_),
    .C(_4138_),
    .A(net1844),
    .Y(_4139_));
 sg13g2_nand3_1 _8646_ (.B(_4129_),
    .C(_4139_),
    .A(net2169),
    .Y(_4140_));
 sg13g2_xnor2_1 _8647_ (.Y(_4141_),
    .A(net2107),
    .B(net1936));
 sg13g2_nor2_1 _8648_ (.A(_1633_),
    .B(_4141_),
    .Y(_4142_));
 sg13g2_a221oi_1 _8649_ (.B2(net2081),
    .C1(_4142_),
    .B1(_1628_),
    .A1(net2116),
    .Y(_4143_),
    .A2(_0859_));
 sg13g2_and2_1 _8650_ (.A(_1570_),
    .B(_4143_),
    .X(_4144_));
 sg13g2_a21o_1 _8651_ (.A2(_4140_),
    .A1(_4128_),
    .B1(_4144_),
    .X(_4145_));
 sg13g2_nor2_1 _8652_ (.A(net1891),
    .B(_1229_),
    .Y(_4146_));
 sg13g2_or4_1 _8653_ (.A(_0902_),
    .B(_0921_),
    .C(_1148_),
    .D(_1496_),
    .X(_4147_));
 sg13g2_nor3_1 _8654_ (.A(_0930_),
    .B(_1264_),
    .C(_4147_),
    .Y(_4148_));
 sg13g2_nand4_1 _8655_ (.B(_1263_),
    .C(_1500_),
    .A(_0983_),
    .Y(_4149_),
    .D(_4148_));
 sg13g2_nor4_2 _8656_ (.A(_1242_),
    .B(_2369_),
    .C(_2483_),
    .Y(_4150_),
    .D(_4149_));
 sg13g2_and2_1 _8657_ (.A(net2111),
    .B(_4150_),
    .X(_4151_));
 sg13g2_a221oi_1 _8658_ (.B2(net1889),
    .C1(_4150_),
    .B1(_1148_),
    .A1(_0680_),
    .Y(_4152_),
    .A2(_0902_));
 sg13g2_nor3_1 _8659_ (.A(net2015),
    .B(_4151_),
    .C(_4152_),
    .Y(_4153_));
 sg13g2_or2_2 _8660_ (.X(_4154_),
    .B(_4153_),
    .A(_4146_));
 sg13g2_nor2b_1 _8661_ (.A(_4154_),
    .B_N(net1733),
    .Y(_4155_));
 sg13g2_o21ai_1 _8662_ (.B1(_4127_),
    .Y(_0625_),
    .A1(_2633_),
    .A2(_4155_));
 sg13g2_nand2_1 _8663_ (.Y(_4156_),
    .A(net527),
    .B(net1963));
 sg13g2_nor2_1 _8664_ (.A(_1635_),
    .B(_4154_),
    .Y(_4157_));
 sg13g2_o21ai_1 _8665_ (.B1(_4156_),
    .Y(_0626_),
    .A1(_2633_),
    .A2(_4157_));
 sg13g2_nand2_1 _8666_ (.Y(_4158_),
    .A(net276),
    .B(net1963));
 sg13g2_nor2_1 _8667_ (.A(_1657_),
    .B(_4154_),
    .Y(_4159_));
 sg13g2_o21ai_1 _8668_ (.B1(_4158_),
    .Y(_0627_),
    .A1(_2633_),
    .A2(_4159_));
 sg13g2_a21oi_1 _8669_ (.A1(net2089),
    .A2(net2058),
    .Y(_4160_),
    .B1(net1934));
 sg13g2_nand3_1 _8670_ (.B(_1260_),
    .C(_4160_),
    .A(_0870_),
    .Y(_4161_));
 sg13g2_nor4_1 _8671_ (.A(_0911_),
    .B(_0936_),
    .C(_1021_),
    .D(_4161_),
    .Y(_4162_));
 sg13g2_nand3_1 _8672_ (.B(_1711_),
    .C(_4162_),
    .A(_1495_),
    .Y(_4163_));
 sg13g2_nor3_1 _8673_ (.A(net2128),
    .B(net2111),
    .C(net1934),
    .Y(_4164_));
 sg13g2_o21ai_1 _8674_ (.B1(net2170),
    .Y(_4165_),
    .A1(_0934_),
    .A2(_4164_));
 sg13g2_a21oi_1 _8675_ (.A1(_0934_),
    .A2(_4163_),
    .Y(_4166_),
    .B1(_4165_));
 sg13g2_nor3_1 _8676_ (.A(net1891),
    .B(net1934),
    .C(_1633_),
    .Y(_4167_));
 sg13g2_or3_2 _8677_ (.A(_4146_),
    .B(_4166_),
    .C(_4167_),
    .X(_4168_));
 sg13g2_inv_1 _8678_ (.Y(_4169_),
    .A(_4168_));
 sg13g2_nor3_1 _8679_ (.A(_2633_),
    .B(_4154_),
    .C(_4169_),
    .Y(_4170_));
 sg13g2_a21o_1 _8680_ (.A2(net1963),
    .A1(net531),
    .B1(_4170_),
    .X(_0628_));
 sg13g2_nand2_1 _8681_ (.Y(_4171_),
    .A(net510),
    .B(net1963));
 sg13g2_o21ai_1 _8682_ (.B1(_0940_),
    .Y(_4172_),
    .A1(net2004),
    .A2(net1928));
 sg13g2_a221oi_1 _8683_ (.B2(_4172_),
    .C1(_1207_),
    .B1(_1184_),
    .A1(_0914_),
    .Y(_4173_),
    .A2(_1183_));
 sg13g2_nand4_1 _8684_ (.B(_1208_),
    .C(_1211_),
    .A(_1187_),
    .Y(_4174_),
    .D(_4173_));
 sg13g2_nor3_1 _8685_ (.A(_1221_),
    .B(_1227_),
    .C(_4174_),
    .Y(_4175_));
 sg13g2_nand2_1 _8686_ (.Y(_4176_),
    .A(_1179_),
    .B(_4175_));
 sg13g2_nor2_1 _8687_ (.A(net2111),
    .B(_0853_),
    .Y(_4177_));
 sg13g2_a22oi_1 _8688_ (.Y(_4178_),
    .B1(_4177_),
    .B2(_1180_),
    .A2(_4176_),
    .A1(net2130));
 sg13g2_nor2_1 _8689_ (.A(_0675_),
    .B(_4178_),
    .Y(_4179_));
 sg13g2_nor3_1 _8690_ (.A(net1876),
    .B(_1230_),
    .C(_1313_),
    .Y(_4180_));
 sg13g2_a21oi_1 _8691_ (.A1(_0884_),
    .A2(net1889),
    .Y(_4181_),
    .B1(_4180_));
 sg13g2_a221oi_1 _8692_ (.B2(_1630_),
    .C1(_1654_),
    .B1(_1425_),
    .A1(net2129),
    .Y(_4182_),
    .A2(_1107_));
 sg13g2_a21oi_2 _8693_ (.B1(net1892),
    .Y(_4183_),
    .A2(_4182_),
    .A1(_4181_));
 sg13g2_nand3_1 _8694_ (.B(_0926_),
    .C(_1425_),
    .A(net2080),
    .Y(_4184_));
 sg13g2_nor3_1 _8695_ (.A(_1594_),
    .B(_1615_),
    .C(_1646_),
    .Y(_4185_));
 sg13g2_nand4_1 _8696_ (.B(_1554_),
    .C(_4184_),
    .A(_1553_),
    .Y(_4186_),
    .D(_4185_));
 sg13g2_a21oi_1 _8697_ (.A1(_1243_),
    .A2(_1647_),
    .Y(_4187_),
    .B1(net1943));
 sg13g2_nor4_1 _8698_ (.A(_1268_),
    .B(_1621_),
    .C(_4186_),
    .D(_4187_),
    .Y(_4188_));
 sg13g2_nor3_1 _8699_ (.A(net2016),
    .B(_1618_),
    .C(_4188_),
    .Y(_4189_));
 sg13g2_nor4_2 _8700_ (.A(_4154_),
    .B(_4179_),
    .C(_4183_),
    .Y(_4190_),
    .D(_4189_));
 sg13g2_o21ai_1 _8701_ (.B1(_4171_),
    .Y(_0629_),
    .A1(_2633_),
    .A2(_4190_));
 sg13g2_nand2b_1 _8702_ (.Y(_4191_),
    .B(net2021),
    .A_N(_4123_));
 sg13g2_nand2_1 _8703_ (.Y(_4192_),
    .A(_1106_),
    .B(_1110_));
 sg13g2_nand3_1 _8704_ (.B(_1685_),
    .C(_4192_),
    .A(\z80.tv80s.i_tv80_core.F[6] ),
    .Y(_4193_));
 sg13g2_nand2b_1 _8705_ (.Y(_4194_),
    .B(_1688_),
    .A_N(net2147));
 sg13g2_nand4_1 _8706_ (.B(_4191_),
    .C(_4193_),
    .A(net2229),
    .Y(_4195_),
    .D(_4194_));
 sg13g2_o21ai_1 _8707_ (.B1(_4195_),
    .Y(_4196_),
    .A1(net2229),
    .A2(net566));
 sg13g2_inv_1 _8708_ (.Y(_0630_),
    .A(_4196_));
 sg13g2_nand4_1 _8709_ (.B(_1254_),
    .C(_1366_),
    .A(_0870_),
    .Y(_4197_),
    .D(_1531_));
 sg13g2_nor3_2 _8710_ (.A(_1715_),
    .B(_2483_),
    .C(_4197_),
    .Y(_4198_));
 sg13g2_a21o_1 _8711_ (.A2(net1971),
    .A1(net591),
    .B1(_4198_),
    .X(_0631_));
 sg13g2_nand2_1 _8712_ (.Y(_4199_),
    .A(net310),
    .B(net1972));
 sg13g2_nor2b_1 _8713_ (.A(_1112_),
    .B_N(_1229_),
    .Y(_4200_));
 sg13g2_nand2b_1 _8714_ (.Y(_4201_),
    .B(_4200_),
    .A_N(_0034_));
 sg13g2_nor2_1 _8715_ (.A(net2024),
    .B(net2129),
    .Y(_4202_));
 sg13g2_nand2_1 _8716_ (.Y(_4203_),
    .A(net2129),
    .B(_0034_));
 sg13g2_nand2b_1 _8717_ (.Y(_4204_),
    .B(_4203_),
    .A_N(_1840_));
 sg13g2_nand2_1 _8718_ (.Y(_4205_),
    .A(_1104_),
    .B(_1313_));
 sg13g2_a22oi_1 _8719_ (.Y(_4206_),
    .B1(_4202_),
    .B2(_1107_),
    .A2(_1839_),
    .A1(_0884_));
 sg13g2_nand3_1 _8720_ (.B(_1109_),
    .C(_4203_),
    .A(net2121),
    .Y(_4207_));
 sg13g2_a21oi_1 _8721_ (.A1(_1110_),
    .A2(_4205_),
    .Y(_4208_),
    .B1(_4204_));
 sg13g2_nor4_1 _8722_ (.A(net1892),
    .B(_1190_),
    .C(_1654_),
    .D(_4208_),
    .Y(_4209_));
 sg13g2_nand4_1 _8723_ (.B(_4206_),
    .C(_4207_),
    .A(_4201_),
    .Y(_4210_),
    .D(_4209_));
 sg13g2_and4_1 _8724_ (.A(_0951_),
    .B(_1234_),
    .C(_1262_),
    .D(_1669_),
    .X(_4211_));
 sg13g2_and3_2 _8725_ (.X(_4212_),
    .A(_1514_),
    .B(_2353_),
    .C(_4211_));
 sg13g2_nand4_1 _8726_ (.B(_1256_),
    .C(_1493_),
    .A(_1015_),
    .Y(_4213_),
    .D(_4212_));
 sg13g2_and2_1 _8727_ (.A(_1493_),
    .B(_4213_),
    .X(_4214_));
 sg13g2_nor3_1 _8728_ (.A(_1552_),
    .B(_4204_),
    .C(_4214_),
    .Y(_4215_));
 sg13g2_o21ai_1 _8729_ (.B1(_1069_),
    .Y(_4216_),
    .A1(_0034_),
    .A2(_4212_));
 sg13g2_o21ai_1 _8730_ (.B1(net2171),
    .Y(_4217_),
    .A1(_4215_),
    .A2(_4216_));
 sg13g2_nor2_2 _8731_ (.A(_1180_),
    .B(_1372_),
    .Y(_4218_));
 sg13g2_inv_1 _8732_ (.Y(_4219_),
    .A(_4218_));
 sg13g2_nand2_1 _8733_ (.Y(_4220_),
    .A(_1195_),
    .B(_1201_));
 sg13g2_nor2_1 _8734_ (.A(_4174_),
    .B(_4220_),
    .Y(_4221_));
 sg13g2_nor3_1 _8735_ (.A(_0932_),
    .B(_0950_),
    .C(_1174_),
    .Y(_4222_));
 sg13g2_nand3_1 _8736_ (.B(_2479_),
    .C(_4222_),
    .A(_1160_),
    .Y(_4223_));
 sg13g2_nor4_2 _8737_ (.A(_1159_),
    .B(_1227_),
    .C(_3668_),
    .Y(_4224_),
    .D(_4223_));
 sg13g2_nand2b_1 _8738_ (.Y(_4225_),
    .B(_4224_),
    .A_N(_4174_));
 sg13g2_nand3_1 _8739_ (.B(_4218_),
    .C(_4221_),
    .A(_4202_),
    .Y(_4226_));
 sg13g2_nand2_1 _8740_ (.Y(_4227_),
    .A(_0034_),
    .B(_0853_));
 sg13g2_a22oi_1 _8741_ (.Y(_4228_),
    .B1(_1837_),
    .B2(_0852_),
    .A2(_1245_),
    .A1(_0931_));
 sg13g2_a221oi_1 _8742_ (.B2(_0852_),
    .C1(_0955_),
    .B1(_1838_),
    .A1(net1949),
    .Y(_4229_),
    .A2(_0864_));
 sg13g2_o21ai_1 _8743_ (.B1(_4227_),
    .Y(_4230_),
    .A1(_4228_),
    .A2(_4229_));
 sg13g2_o21ai_1 _8744_ (.B1(_4230_),
    .Y(_4231_),
    .A1(_1840_),
    .A2(_4221_));
 sg13g2_nor2b_1 _8745_ (.A(_4231_),
    .B_N(_4226_),
    .Y(_4232_));
 sg13g2_o21ai_1 _8746_ (.B1(_4217_),
    .Y(_4233_),
    .A1(_0033_),
    .A2(_4232_));
 sg13g2_o21ai_1 _8747_ (.B1(_4210_),
    .Y(_4234_),
    .A1(net1954),
    .A2(_4233_));
 sg13g2_o21ai_1 _8748_ (.B1(net1875),
    .Y(_4235_),
    .A1(net2131),
    .A2(_1648_));
 sg13g2_nor2_1 _8749_ (.A(net2061),
    .B(_4212_),
    .Y(_4236_));
 sg13g2_nand2_1 _8750_ (.Y(_4237_),
    .A(net2066),
    .B(net1943));
 sg13g2_nor2_1 _8751_ (.A(_1014_),
    .B(_4237_),
    .Y(_4238_));
 sg13g2_nor3_1 _8752_ (.A(_1255_),
    .B(_4236_),
    .C(_4238_),
    .Y(_4239_));
 sg13g2_o21ai_1 _8753_ (.B1(_4239_),
    .Y(_4240_),
    .A1(_4214_),
    .A2(_4235_));
 sg13g2_a21o_1 _8754_ (.A2(net2061),
    .A1(net2122),
    .B1(_0885_),
    .X(_4241_));
 sg13g2_o21ai_1 _8755_ (.B1(_4241_),
    .Y(_4242_),
    .A1(_0860_),
    .A2(_4237_));
 sg13g2_a22oi_1 _8756_ (.Y(_4243_),
    .B1(_1110_),
    .B2(_4205_),
    .A2(net2061),
    .A1(net2129));
 sg13g2_nor2_1 _8757_ (.A(_1106_),
    .B(_1640_),
    .Y(_4244_));
 sg13g2_or4_1 _8758_ (.A(_4200_),
    .B(_4242_),
    .C(_4243_),
    .D(_4244_),
    .X(_4245_));
 sg13g2_a21oi_1 _8759_ (.A1(net2061),
    .A2(_4200_),
    .Y(_4246_),
    .B1(net1892));
 sg13g2_nand2_1 _8760_ (.Y(_4247_),
    .A(_0852_),
    .B(_1648_));
 sg13g2_o21ai_1 _8761_ (.B1(_4247_),
    .Y(_4248_),
    .A1(net2061),
    .A2(_0852_));
 sg13g2_o21ai_1 _8762_ (.B1(net2167),
    .Y(_4249_),
    .A1(_4218_),
    .A2(_4248_));
 sg13g2_a21oi_1 _8763_ (.A1(_1640_),
    .A2(_4218_),
    .Y(_4250_),
    .B1(_4249_));
 sg13g2_a22oi_1 _8764_ (.Y(_4251_),
    .B1(_4245_),
    .B2(_4246_),
    .A2(_4240_),
    .A1(net2171));
 sg13g2_nor2b_2 _8765_ (.A(_4250_),
    .B_N(_4251_),
    .Y(_4252_));
 sg13g2_nand4_1 _8766_ (.B(\z80.tv80s.i_tv80_core.ISet[1] ),
    .C(net1996),
    .A(net2110),
    .Y(_4253_),
    .D(_4252_));
 sg13g2_o21ai_1 _8767_ (.B1(_4199_),
    .Y(_0632_),
    .A1(_4234_),
    .A2(_4253_));
 sg13g2_nand2_1 _8768_ (.Y(_4254_),
    .A(net2042),
    .B(net1972));
 sg13g2_o21ai_1 _8769_ (.B1(_4254_),
    .Y(_0633_),
    .A1(net1686),
    .A2(_4234_));
 sg13g2_or4_1 _8770_ (.A(net2022),
    .B(net2129),
    .C(_4219_),
    .D(_4225_),
    .X(_4255_));
 sg13g2_nand2_1 _8771_ (.Y(_4256_),
    .A(net2021),
    .B(net2018));
 sg13g2_nand3_1 _8772_ (.B(net2120),
    .C(net1886),
    .A(net2057),
    .Y(_4257_));
 sg13g2_nand3_1 _8773_ (.B(_1575_),
    .C(_4257_),
    .A(_0852_),
    .Y(_4258_));
 sg13g2_a21oi_1 _8774_ (.A1(_0026_),
    .A2(_0853_),
    .Y(_4259_),
    .B1(_4218_));
 sg13g2_a22oi_1 _8775_ (.Y(_4260_),
    .B1(_4258_),
    .B2(_4259_),
    .A2(_4256_),
    .A1(_4225_));
 sg13g2_a21oi_1 _8776_ (.A1(_4255_),
    .A2(_4260_),
    .Y(_4261_),
    .B1(_0033_));
 sg13g2_nand2_1 _8777_ (.Y(_4262_),
    .A(net2130),
    .B(_0026_));
 sg13g2_nand2_1 _8778_ (.Y(_4263_),
    .A(_4256_),
    .B(_4262_));
 sg13g2_nor3_1 _8779_ (.A(_1552_),
    .B(_4213_),
    .C(_4263_),
    .Y(_4264_));
 sg13g2_o21ai_1 _8780_ (.B1(_4262_),
    .Y(_4265_),
    .A1(net2075),
    .A2(net1947));
 sg13g2_a21oi_1 _8781_ (.A1(net1875),
    .A2(_4265_),
    .Y(_4266_),
    .B1(_1493_));
 sg13g2_nor3_1 _8782_ (.A(net2021),
    .B(_0870_),
    .C(_1014_),
    .Y(_4267_));
 sg13g2_nor3_1 _8783_ (.A(_1011_),
    .B(_4266_),
    .C(_4267_),
    .Y(_4268_));
 sg13g2_o21ai_1 _8784_ (.B1(_4268_),
    .Y(_4269_),
    .A1(_0026_),
    .A2(_4212_));
 sg13g2_o21ai_1 _8785_ (.B1(net2171),
    .Y(_4270_),
    .A1(_4264_),
    .A2(_4269_));
 sg13g2_nor2_1 _8786_ (.A(net1954),
    .B(_4261_),
    .Y(_4271_));
 sg13g2_nand3_1 _8787_ (.B(net2121),
    .C(_0884_),
    .A(net2080),
    .Y(_4272_));
 sg13g2_a21o_1 _8788_ (.A2(_4272_),
    .A1(_1112_),
    .B1(_0026_),
    .X(_4273_));
 sg13g2_nand2_1 _8789_ (.Y(_4274_),
    .A(net2116),
    .B(_0026_));
 sg13g2_a22oi_1 _8790_ (.Y(_4275_),
    .B1(_3271_),
    .B2(_4274_),
    .A2(_0859_),
    .A1(net2023));
 sg13g2_a21oi_1 _8791_ (.A1(net2021),
    .A2(net1942),
    .Y(_4276_),
    .B1(_4275_));
 sg13g2_nor2_1 _8792_ (.A(_4205_),
    .B(_4263_),
    .Y(_4277_));
 sg13g2_nand3_1 _8793_ (.B(net1943),
    .C(_1190_),
    .A(net2075),
    .Y(_4278_));
 sg13g2_a21o_1 _8794_ (.A2(_4256_),
    .A1(_1107_),
    .B1(_1571_),
    .X(_4279_));
 sg13g2_o21ai_1 _8795_ (.B1(_4278_),
    .Y(_4280_),
    .A1(_1110_),
    .A2(_4265_));
 sg13g2_nor4_1 _8796_ (.A(_4276_),
    .B(_4277_),
    .C(_4279_),
    .D(_4280_),
    .Y(_4281_));
 sg13g2_a221oi_1 _8797_ (.B2(_4281_),
    .C1(net1686),
    .B1(_4273_),
    .A1(_4270_),
    .Y(_4282_),
    .A2(_4271_));
 sg13g2_a21o_1 _8798_ (.A2(net1967),
    .A1(net2037),
    .B1(_4282_),
    .X(_0634_));
 sg13g2_nand2_1 _8799_ (.Y(_4283_),
    .A(net267),
    .B(net1972));
 sg13g2_o21ai_1 _8800_ (.B1(_4283_),
    .Y(_0635_),
    .A1(net1686),
    .A2(_4252_));
 sg13g2_nor2b_1 _8801_ (.A(_4218_),
    .B_N(_4177_),
    .Y(_4284_));
 sg13g2_a21oi_1 _8802_ (.A1(net2130),
    .A2(_4218_),
    .Y(_4285_),
    .B1(_4284_));
 sg13g2_a21oi_1 _8803_ (.A1(net2171),
    .A2(_1257_),
    .Y(_4286_),
    .B1(net1954));
 sg13g2_o21ai_1 _8804_ (.B1(_4286_),
    .Y(_4287_),
    .A1(_0033_),
    .A2(_4285_));
 sg13g2_nand3b_1 _8805_ (.B(_4287_),
    .C(_1569_),
    .Y(_4288_),
    .A_N(net1686));
 sg13g2_o21ai_1 _8806_ (.B1(_4288_),
    .Y(_0636_),
    .A1(_0778_),
    .A2(net1996));
 sg13g2_nand4_1 _8807_ (.B(_1015_),
    .C(_1165_),
    .A(net1883),
    .Y(_4289_),
    .D(_1669_));
 sg13g2_nor3_1 _8808_ (.A(_1663_),
    .B(_1666_),
    .C(_4289_),
    .Y(_4290_));
 sg13g2_nand4_1 _8809_ (.B(_1262_),
    .C(_1263_),
    .A(_0951_),
    .Y(_4291_),
    .D(_1505_));
 sg13g2_nor2_1 _8810_ (.A(_1662_),
    .B(_4291_),
    .Y(_4292_));
 sg13g2_nand3_1 _8811_ (.B(_4290_),
    .C(_4292_),
    .A(_2353_),
    .Y(_4293_));
 sg13g2_nor4_1 _8812_ (.A(_1257_),
    .B(_1555_),
    .C(_1619_),
    .D(_1646_),
    .Y(_4294_));
 sg13g2_a21oi_1 _8813_ (.A1(_4293_),
    .A2(_4294_),
    .Y(_4295_),
    .B1(net2017));
 sg13g2_o21ai_1 _8814_ (.B1(_4295_),
    .Y(_4296_),
    .A1(_1549_),
    .A2(_4293_));
 sg13g2_nor2_1 _8815_ (.A(net1953),
    .B(_4179_),
    .Y(_4297_));
 sg13g2_a221oi_1 _8816_ (.B2(net1922),
    .C1(_1654_),
    .B1(_1109_),
    .A1(net2124),
    .Y(_4298_),
    .A2(_1107_));
 sg13g2_a221oi_1 _8817_ (.B2(_1572_),
    .C1(net1686),
    .B1(_4298_),
    .A1(_4296_),
    .Y(_4299_),
    .A2(_4297_));
 sg13g2_a21o_1 _8818_ (.A2(net1971),
    .A1(net2033),
    .B1(_4299_),
    .X(_0637_));
 sg13g2_nand2_1 _8819_ (.Y(_4300_),
    .A(net600),
    .B(net1965));
 sg13g2_nor2_1 _8820_ (.A(_1635_),
    .B(_1657_),
    .Y(_4301_));
 sg13g2_o21ai_1 _8821_ (.B1(net1985),
    .Y(_4302_),
    .A1(_4169_),
    .A2(_4301_));
 sg13g2_a21oi_2 _8822_ (.B1(_4168_),
    .Y(_4303_),
    .A2(_1657_),
    .A1(_1635_));
 sg13g2_inv_2 _8823_ (.Y(_4304_),
    .A(_4303_));
 sg13g2_mux2_1 _8824_ (.A0(_1910_),
    .A1(_2331_),
    .S(net1732),
    .X(_4305_));
 sg13g2_nand2_1 _8825_ (.Y(_4306_),
    .A(_4168_),
    .B(_4301_));
 sg13g2_nor2_2 _8826_ (.A(net1733),
    .B(_4306_),
    .Y(_4307_));
 sg13g2_nor2b_2 _8827_ (.A(_4306_),
    .B_N(net1733),
    .Y(_4308_));
 sg13g2_nand3_1 _8828_ (.B(_1657_),
    .C(_4169_),
    .A(_1635_),
    .Y(_4309_));
 sg13g2_nor2b_2 _8829_ (.A(_4309_),
    .B_N(net1733),
    .Y(_4310_));
 sg13g2_nor2_2 _8830_ (.A(net1733),
    .B(_4309_),
    .Y(_4311_));
 sg13g2_a22oi_1 _8831_ (.Y(_4312_),
    .B1(_4311_),
    .B2(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(_4308_),
    .A1(\z80.tv80s.i_tv80_core.SP[7] ));
 sg13g2_o21ai_1 _8832_ (.B1(_4312_),
    .Y(_4313_),
    .A1(_4304_),
    .A2(_4305_));
 sg13g2_a221oi_1 _8833_ (.B2(net2043),
    .C1(_4313_),
    .B1(_4310_),
    .A1(\z80.tv80s.i_tv80_core.SP[15] ),
    .Y(_4314_),
    .A2(_4307_));
 sg13g2_o21ai_1 _8834_ (.B1(_4300_),
    .Y(_0638_),
    .A1(_4302_),
    .A2(_4314_));
 sg13g2_nand2_1 _8835_ (.Y(_4315_),
    .A(net2030),
    .B(net1966));
 sg13g2_mux2_1 _8836_ (.A0(_1919_),
    .A1(_2278_),
    .S(net1732),
    .X(_4316_));
 sg13g2_a22oi_1 _8837_ (.Y(_4317_),
    .B1(_4311_),
    .B2(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_4310_),
    .A1(net2045));
 sg13g2_o21ai_1 _8838_ (.B1(_4317_),
    .Y(_4318_),
    .A1(_4304_),
    .A2(_4316_));
 sg13g2_a221oi_1 _8839_ (.B2(\z80.tv80s.i_tv80_core.SP[6] ),
    .C1(_4318_),
    .B1(_4308_),
    .A1(\z80.tv80s.i_tv80_core.SP[14] ),
    .Y(_4319_),
    .A2(_4307_));
 sg13g2_o21ai_1 _8840_ (.B1(_4315_),
    .Y(_0639_),
    .A1(_4302_),
    .A2(_4319_));
 sg13g2_nand2_1 _8841_ (.Y(_4320_),
    .A(net2029),
    .B(net1966));
 sg13g2_mux2_1 _8842_ (.A0(_1928_),
    .A1(_2227_),
    .S(net1732),
    .X(_4321_));
 sg13g2_a22oi_1 _8843_ (.Y(_4322_),
    .B1(_4311_),
    .B2(net2145),
    .A2(_4308_),
    .A1(\z80.tv80s.i_tv80_core.SP[5] ));
 sg13g2_o21ai_1 _8844_ (.B1(_4322_),
    .Y(_4323_),
    .A1(_4304_),
    .A2(_4321_));
 sg13g2_a221oi_1 _8845_ (.B2(net2046),
    .C1(_4323_),
    .B1(_4310_),
    .A1(\z80.tv80s.i_tv80_core.SP[13] ),
    .Y(_4324_),
    .A2(_4307_));
 sg13g2_o21ai_1 _8846_ (.B1(_4320_),
    .Y(_0640_),
    .A1(_4302_),
    .A2(_4324_));
 sg13g2_nand2_1 _8847_ (.Y(_4325_),
    .A(net598),
    .B(net1965));
 sg13g2_mux2_1 _8848_ (.A0(_1935_),
    .A1(_2159_),
    .S(net1732),
    .X(_4326_));
 sg13g2_a22oi_1 _8849_ (.Y(_4327_),
    .B1(_4308_),
    .B2(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(_4307_),
    .A1(\z80.tv80s.i_tv80_core.SP[12] ));
 sg13g2_o21ai_1 _8850_ (.B1(_4327_),
    .Y(_4328_),
    .A1(_4304_),
    .A2(_4326_));
 sg13g2_a221oi_1 _8851_ (.B2(\z80.tv80s.i_tv80_core.ACC[4] ),
    .C1(_4328_),
    .B1(_4311_),
    .A1(net2047),
    .Y(_4329_),
    .A2(_4310_));
 sg13g2_o21ai_1 _8852_ (.B1(_4325_),
    .Y(_0641_),
    .A1(_4302_),
    .A2(_4329_));
 sg13g2_nand2_1 _8853_ (.Y(_4330_),
    .A(net572),
    .B(net1966));
 sg13g2_mux2_1 _8854_ (.A0(_1867_),
    .A1(_2107_),
    .S(net1732),
    .X(_4331_));
 sg13g2_a22oi_1 _8855_ (.Y(_4332_),
    .B1(_4311_),
    .B2(net2146),
    .A2(_4308_),
    .A1(\z80.tv80s.i_tv80_core.SP[3] ));
 sg13g2_o21ai_1 _8856_ (.B1(_4332_),
    .Y(_4333_),
    .A1(_4304_),
    .A2(_4331_));
 sg13g2_a221oi_1 _8857_ (.B2(net2048),
    .C1(_4333_),
    .B1(_4310_),
    .A1(\z80.tv80s.i_tv80_core.SP[11] ),
    .Y(_4334_),
    .A2(_4307_));
 sg13g2_o21ai_1 _8858_ (.B1(_4330_),
    .Y(_0642_),
    .A1(_4302_),
    .A2(_4334_));
 sg13g2_nand2_1 _8859_ (.Y(_4335_),
    .A(net2028),
    .B(net1965));
 sg13g2_mux2_1 _8860_ (.A0(_1897_),
    .A1(_2056_),
    .S(net1732),
    .X(_4336_));
 sg13g2_a22oi_1 _8861_ (.Y(_4337_),
    .B1(_4311_),
    .B2(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_4308_),
    .A1(\z80.tv80s.i_tv80_core.SP[2] ));
 sg13g2_o21ai_1 _8862_ (.B1(_4337_),
    .Y(_4338_),
    .A1(_4304_),
    .A2(_4336_));
 sg13g2_a221oi_1 _8863_ (.B2(net2049),
    .C1(_4338_),
    .B1(_4310_),
    .A1(\z80.tv80s.i_tv80_core.SP[10] ),
    .Y(_4339_),
    .A2(_4307_));
 sg13g2_o21ai_1 _8864_ (.B1(_4335_),
    .Y(_0643_),
    .A1(_4302_),
    .A2(_4339_));
 sg13g2_o21ai_1 _8865_ (.B1(_4303_),
    .Y(_4340_),
    .A1(_1881_),
    .A2(net1732));
 sg13g2_a21oi_2 _8866_ (.B1(_4340_),
    .Y(_4341_),
    .A2(net1733),
    .A1(_2012_));
 sg13g2_a22oi_1 _8867_ (.Y(_4342_),
    .B1(_4311_),
    .B2(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_4307_),
    .A1(\z80.tv80s.i_tv80_core.SP[9] ));
 sg13g2_a221oi_1 _8868_ (.B2(net2050),
    .C1(_4341_),
    .B1(_4310_),
    .A1(\z80.tv80s.i_tv80_core.SP[1] ),
    .Y(_4343_),
    .A2(_4308_));
 sg13g2_a21oi_2 _8869_ (.B1(_4302_),
    .Y(_4344_),
    .A2(_4343_),
    .A1(_4342_));
 sg13g2_a21o_1 _8870_ (.A2(net1967),
    .A1(net2027),
    .B1(_4344_),
    .X(_0644_));
 sg13g2_o21ai_1 _8871_ (.B1(_4303_),
    .Y(_4345_),
    .A1(_1888_),
    .A2(net1732));
 sg13g2_a21oi_1 _8872_ (.A1(_1950_),
    .A2(net1733),
    .Y(_4346_),
    .B1(_4345_));
 sg13g2_a22oi_1 _8873_ (.Y(_4347_),
    .B1(_4311_),
    .B2(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A2(_4310_),
    .A1(net2051));
 sg13g2_a221oi_1 _8874_ (.B2(\z80.tv80s.i_tv80_core.SP[0] ),
    .C1(_4346_),
    .B1(_4308_),
    .A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .Y(_4348_),
    .A2(_4307_));
 sg13g2_a21o_2 _8875_ (.A2(_4348_),
    .A1(_4347_),
    .B1(_4302_),
    .X(_4349_));
 sg13g2_o21ai_1 _8876_ (.B1(_4349_),
    .Y(_0645_),
    .A1(_0782_),
    .A2(net1994));
 sg13g2_nand2_1 _8877_ (.Y(_4350_),
    .A(net567),
    .B(net1969));
 sg13g2_nor3_1 _8878_ (.A(_0982_),
    .B(_1016_),
    .C(_1019_),
    .Y(_4351_));
 sg13g2_and4_1 _8879_ (.A(_0991_),
    .B(_0996_),
    .C(_1248_),
    .D(_4351_),
    .X(_4352_));
 sg13g2_nor4_1 _8880_ (.A(_1010_),
    .B(_1150_),
    .C(_1544_),
    .D(_1668_),
    .Y(_4353_));
 sg13g2_nor2_1 _8881_ (.A(_0937_),
    .B(_1242_),
    .Y(_4354_));
 sg13g2_nand3_1 _8882_ (.B(_4353_),
    .C(_4354_),
    .A(_4352_),
    .Y(_4355_));
 sg13g2_a221oi_1 _8883_ (.B2(net1935),
    .C1(_1555_),
    .B1(_1646_),
    .A1(_0881_),
    .Y(_4356_),
    .A2(_1003_));
 sg13g2_nand4_1 _8884_ (.B(_1593_),
    .C(_4355_),
    .A(_1586_),
    .Y(_4357_),
    .D(_4356_));
 sg13g2_o21ai_1 _8885_ (.B1(net2170),
    .Y(_4358_),
    .A1(_4164_),
    .A2(_4355_));
 sg13g2_nand2b_1 _8886_ (.Y(_4359_),
    .B(_4357_),
    .A_N(_4358_));
 sg13g2_a21oi_1 _8887_ (.A1(net2014),
    .A2(net1934),
    .Y(_4360_),
    .B1(_1574_));
 sg13g2_nor2b_1 _8888_ (.A(net2115),
    .B_N(_4360_),
    .Y(_4361_));
 sg13g2_o21ai_1 _8889_ (.B1(net1935),
    .Y(_4362_),
    .A1(_1654_),
    .A2(_4361_));
 sg13g2_a221oi_1 _8890_ (.B2(net1876),
    .C1(net1891),
    .B1(_1578_),
    .A1(net2126),
    .Y(_4363_),
    .A2(_1107_));
 sg13g2_a221oi_1 _8891_ (.B2(_4363_),
    .C1(net2105),
    .B1(_4362_),
    .A1(net1891),
    .Y(_4364_),
    .A2(_4359_));
 sg13g2_nand3_1 _8892_ (.B(_1609_),
    .C(_4364_),
    .A(_1584_),
    .Y(_4365_));
 sg13g2_nand2_2 _8893_ (.Y(_4366_),
    .A(net1993),
    .B(_4365_));
 sg13g2_nor2_1 _8894_ (.A(net1797),
    .B(_2336_),
    .Y(_4367_));
 sg13g2_a22oi_1 _8895_ (.Y(_4368_),
    .B1(_1238_),
    .B2(_1577_),
    .A2(net1864),
    .A1(_0149_));
 sg13g2_o21ai_1 _8896_ (.B1(net2118),
    .Y(_4369_),
    .A1(_1174_),
    .A2(_1297_));
 sg13g2_a21oi_1 _8897_ (.A1(net2131),
    .A2(net1933),
    .Y(_4370_),
    .B1(_1292_));
 sg13g2_nor2_1 _8898_ (.A(_0149_),
    .B(_0864_),
    .Y(_4371_));
 sg13g2_a22oi_1 _8899_ (.Y(_4372_),
    .B1(_4371_),
    .B2(_0955_),
    .A2(_4370_),
    .A1(_0981_));
 sg13g2_o21ai_1 _8900_ (.B1(_4372_),
    .Y(_4373_),
    .A1(_1002_),
    .A2(_2473_));
 sg13g2_a21oi_1 _8901_ (.A1(net1882),
    .A2(_4132_),
    .Y(_4374_),
    .B1(_4373_));
 sg13g2_o21ai_1 _8902_ (.B1(net2127),
    .Y(_4375_),
    .A1(_0982_),
    .A2(_1264_));
 sg13g2_o21ai_1 _8903_ (.B1(_0886_),
    .Y(_4376_),
    .A1(_0915_),
    .A2(_1431_));
 sg13g2_nand4_1 _8904_ (.B(_4374_),
    .C(_4375_),
    .A(_4369_),
    .Y(_4377_),
    .D(_4376_));
 sg13g2_a221oi_1 _8905_ (.B2(_1268_),
    .C1(_4377_),
    .B1(_4368_),
    .A1(net1884),
    .Y(_4378_),
    .A2(_2580_));
 sg13g2_o21ai_1 _8906_ (.B1(_4128_),
    .Y(_4379_),
    .A1(net2015),
    .A2(_4378_));
 sg13g2_a21oi_1 _8907_ (.A1(_0859_),
    .A2(_4132_),
    .Y(_4380_),
    .B1(_1571_));
 sg13g2_a22oi_1 _8908_ (.Y(_4381_),
    .B1(_4131_),
    .B2(_4360_),
    .A2(_1578_),
    .A1(net2080));
 sg13g2_a21oi_1 _8909_ (.A1(_4380_),
    .A2(_4381_),
    .Y(_4382_),
    .B1(net2105));
 sg13g2_a22oi_1 _8910_ (.Y(_4383_),
    .B1(_4379_),
    .B2(_4382_),
    .A2(_0733_),
    .A1(net2105));
 sg13g2_inv_4 _8911_ (.A(net1730),
    .Y(_4384_));
 sg13g2_o21ai_1 _8912_ (.B1(net1786),
    .Y(_4385_),
    .A1(_0140_),
    .A2(net1814));
 sg13g2_a21oi_1 _8913_ (.A1(_0727_),
    .A2(net2010),
    .Y(_4386_),
    .B1(_4385_));
 sg13g2_nor2_1 _8914_ (.A(_0136_),
    .B(net1814),
    .Y(_4387_));
 sg13g2_o21ai_1 _8915_ (.B1(net1804),
    .Y(_4388_),
    .A1(_0135_),
    .A2(net2163));
 sg13g2_o21ai_1 _8916_ (.B1(net1799),
    .Y(_4389_),
    .A1(_4387_),
    .A2(_4388_));
 sg13g2_o21ai_1 _8917_ (.B1(net1730),
    .Y(_4390_),
    .A1(_4386_),
    .A2(_4389_));
 sg13g2_nand2_1 _8918_ (.Y(_4391_),
    .A(_1584_),
    .B(_1609_));
 sg13g2_a21oi_1 _8919_ (.A1(_1584_),
    .A2(_1609_),
    .Y(_4392_),
    .B1(_4364_));
 sg13g2_nand2b_2 _8920_ (.Y(_4393_),
    .B(_4391_),
    .A_N(_4364_));
 sg13g2_a221oi_1 _8921_ (.B2(_0728_),
    .C1(net1785),
    .B1(net1808),
    .A1(_0729_),
    .Y(_4394_),
    .A2(net2009));
 sg13g2_a221oi_1 _8922_ (.B2(_0731_),
    .C1(net1802),
    .B1(net1808),
    .A1(_0732_),
    .Y(_4395_),
    .A2(net2009));
 sg13g2_nor3_1 _8923_ (.A(_1963_),
    .B(_4394_),
    .C(_4395_),
    .Y(_4396_));
 sg13g2_nor2_1 _8924_ (.A(net1731),
    .B(_4396_),
    .Y(_4397_));
 sg13g2_o21ai_1 _8925_ (.B1(_4397_),
    .Y(_4398_),
    .A1(net1797),
    .A2(_2455_));
 sg13g2_o21ai_1 _8926_ (.B1(_4398_),
    .Y(_4399_),
    .A1(_4367_),
    .A2(_4390_));
 sg13g2_nand3_1 _8927_ (.B(_1609_),
    .C(_4364_),
    .A(_1583_),
    .Y(_4400_));
 sg13g2_nor2_2 _8928_ (.A(_4383_),
    .B(_4400_),
    .Y(_4401_));
 sg13g2_nand2b_2 _8929_ (.Y(_4402_),
    .B(_4364_),
    .A_N(_1609_));
 sg13g2_nor2_1 _8930_ (.A(_4384_),
    .B(_4402_),
    .Y(_4403_));
 sg13g2_nor3_2 _8931_ (.A(_1584_),
    .B(_4384_),
    .C(_4402_),
    .Y(_4404_));
 sg13g2_or2_1 _8932_ (.X(_4405_),
    .B(_4391_),
    .A(_4364_));
 sg13g2_nor2_2 _8933_ (.A(_4384_),
    .B(_4405_),
    .Y(_4406_));
 sg13g2_nor3_2 _8934_ (.A(_1583_),
    .B(_4383_),
    .C(_4402_),
    .Y(_4407_));
 sg13g2_nor2_2 _8935_ (.A(_4384_),
    .B(_4400_),
    .Y(_4408_));
 sg13g2_a22oi_1 _8936_ (.Y(_4409_),
    .B1(_4408_),
    .B2(\z80.tv80s.i_tv80_core.PC[7] ),
    .A2(_4407_),
    .A1(\z80.tv80s.i_tv80_core.F[7] ));
 sg13g2_nor2_2 _8937_ (.A(_4383_),
    .B(_4405_),
    .Y(_4410_));
 sg13g2_nor3_2 _8938_ (.A(_1584_),
    .B(net1730),
    .C(_4402_),
    .Y(_4411_));
 sg13g2_nand2_1 _8939_ (.Y(_4412_),
    .A(\z80.tv80s.i_tv80_core.SP[15] ),
    .B(_4411_));
 sg13g2_a22oi_1 _8940_ (.Y(_4413_),
    .B1(_4404_),
    .B2(\z80.tv80s.i_tv80_core.SP[7] ),
    .A2(_4401_),
    .A1(\z80.tv80s.i_tv80_core.PC[15] ));
 sg13g2_nand3_1 _8941_ (.B(_4412_),
    .C(_4413_),
    .A(_4409_),
    .Y(_4414_));
 sg13g2_a22oi_1 _8942_ (.Y(_4415_),
    .B1(_4410_),
    .B2(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(_4406_),
    .A1(net2043));
 sg13g2_o21ai_1 _8943_ (.B1(_4415_),
    .Y(_4416_),
    .A1(_4393_),
    .A2(_4399_));
 sg13g2_nor2_2 _8944_ (.A(_4414_),
    .B(_4416_),
    .Y(_4417_));
 sg13g2_o21ai_1 _8945_ (.B1(_4350_),
    .Y(_0646_),
    .A1(_4366_),
    .A2(_4417_));
 sg13g2_nand2_1 _8946_ (.Y(_4418_),
    .A(net578),
    .B(net1970));
 sg13g2_o21ai_1 _8947_ (.B1(net1786),
    .Y(_4419_),
    .A1(_0123_),
    .A2(net2165));
 sg13g2_a21oi_1 _8948_ (.A1(_0720_),
    .A2(net1809),
    .Y(_4420_),
    .B1(_4419_));
 sg13g2_nor2_1 _8949_ (.A(_0120_),
    .B(net1813),
    .Y(_4421_));
 sg13g2_o21ai_1 _8950_ (.B1(net1805),
    .Y(_4422_),
    .A1(_0119_),
    .A2(net2165));
 sg13g2_o21ai_1 _8951_ (.B1(net1800),
    .Y(_4423_),
    .A1(_4421_),
    .A2(_4422_));
 sg13g2_o21ai_1 _8952_ (.B1(net1730),
    .Y(_4424_),
    .A1(_4420_),
    .A2(_4423_));
 sg13g2_nor2_1 _8953_ (.A(_2240_),
    .B(_4424_),
    .Y(_4425_));
 sg13g2_a22oi_1 _8954_ (.Y(_4426_),
    .B1(net1807),
    .B2(_0722_),
    .A2(net2009),
    .A1(_0723_));
 sg13g2_nor2_1 _8955_ (.A(_0128_),
    .B(net1812),
    .Y(_4427_));
 sg13g2_o21ai_1 _8956_ (.B1(net1803),
    .Y(_4428_),
    .A1(_0127_),
    .A2(net2164));
 sg13g2_o21ai_1 _8957_ (.B1(net1797),
    .Y(_4429_),
    .A1(_4427_),
    .A2(_4428_));
 sg13g2_a21oi_2 _8958_ (.B1(_4429_),
    .Y(_4430_),
    .A2(_4426_),
    .A1(net1785));
 sg13g2_o21ai_1 _8959_ (.B1(_4384_),
    .Y(_4431_),
    .A1(net1798),
    .A2(_2445_));
 sg13g2_nor2_1 _8960_ (.A(_4393_),
    .B(_4425_),
    .Y(_4432_));
 sg13g2_o21ai_1 _8961_ (.B1(_4432_),
    .Y(_4433_),
    .A1(_4430_),
    .A2(_4431_));
 sg13g2_a22oi_1 _8962_ (.Y(_4434_),
    .B1(_4407_),
    .B2(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(_4404_),
    .A1(\z80.tv80s.i_tv80_core.SP[6] ));
 sg13g2_a22oi_1 _8963_ (.Y(_4435_),
    .B1(_4411_),
    .B2(\z80.tv80s.i_tv80_core.SP[14] ),
    .A2(_4408_),
    .A1(\z80.tv80s.i_tv80_core.PC[6] ));
 sg13g2_a22oi_1 _8964_ (.Y(_4436_),
    .B1(_4410_),
    .B2(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_4401_),
    .A1(\z80.tv80s.i_tv80_core.PC[14] ));
 sg13g2_nand4_1 _8965_ (.B(_4434_),
    .C(_4435_),
    .A(_4433_),
    .Y(_4437_),
    .D(_4436_));
 sg13g2_a21oi_2 _8966_ (.B1(_4437_),
    .Y(_4438_),
    .A2(_4406_),
    .A1(\z80.tv80s.di_reg[6] ));
 sg13g2_o21ai_1 _8967_ (.B1(_4418_),
    .Y(_0647_),
    .A1(_4366_),
    .A2(_4438_));
 sg13g2_nand2_1 _8968_ (.Y(_4439_),
    .A(net575),
    .B(net1970));
 sg13g2_o21ai_1 _8969_ (.B1(net1786),
    .Y(_4440_),
    .A1(_0108_),
    .A2(net1814));
 sg13g2_a21oi_1 _8970_ (.A1(_0714_),
    .A2(net2010),
    .Y(_4441_),
    .B1(_4440_));
 sg13g2_nor2_1 _8971_ (.A(_0104_),
    .B(net1814),
    .Y(_4442_));
 sg13g2_o21ai_1 _8972_ (.B1(net1804),
    .Y(_4443_),
    .A1(_0103_),
    .A2(net2163));
 sg13g2_o21ai_1 _8973_ (.B1(net1799),
    .Y(_4444_),
    .A1(_4442_),
    .A2(_4443_));
 sg13g2_o21ai_1 _8974_ (.B1(net1730),
    .Y(_4445_),
    .A1(_4441_),
    .A2(_4444_));
 sg13g2_nor2_1 _8975_ (.A(_2236_),
    .B(_4445_),
    .Y(_4446_));
 sg13g2_nor2_1 _8976_ (.A(_4393_),
    .B(_4446_),
    .Y(_4447_));
 sg13g2_o21ai_1 _8977_ (.B1(_4447_),
    .Y(_4448_),
    .A1(_2441_),
    .A2(net1731));
 sg13g2_a22oi_1 _8978_ (.Y(_4449_),
    .B1(_4410_),
    .B2(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2(_4404_),
    .A1(\z80.tv80s.i_tv80_core.SP[5] ));
 sg13g2_a22oi_1 _8979_ (.Y(_4450_),
    .B1(_4411_),
    .B2(\z80.tv80s.i_tv80_core.SP[13] ),
    .A2(_4406_),
    .A1(net2046));
 sg13g2_a22oi_1 _8980_ (.Y(_4451_),
    .B1(_4407_),
    .B2(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_4401_),
    .A1(\z80.tv80s.i_tv80_core.PC[13] ));
 sg13g2_nand4_1 _8981_ (.B(_4449_),
    .C(_4450_),
    .A(_4448_),
    .Y(_4452_),
    .D(_4451_));
 sg13g2_a21oi_2 _8982_ (.B1(_4452_),
    .Y(_4453_),
    .A2(_4408_),
    .A1(\z80.tv80s.i_tv80_core.PC[5] ));
 sg13g2_o21ai_1 _8983_ (.B1(_4439_),
    .Y(_0648_),
    .A1(_4366_),
    .A2(_4453_));
 sg13g2_nand2_1 _8984_ (.Y(_4454_),
    .A(net569),
    .B(net1970));
 sg13g2_o21ai_1 _8985_ (.B1(net1802),
    .Y(_4455_),
    .A1(_0095_),
    .A2(net2164));
 sg13g2_a21oi_1 _8986_ (.A1(_0712_),
    .A2(net1807),
    .Y(_4456_),
    .B1(_4455_));
 sg13g2_o21ai_1 _8987_ (.B1(net1785),
    .Y(_4457_),
    .A1(_0099_),
    .A2(net2164));
 sg13g2_a21oi_1 _8988_ (.A1(_0713_),
    .A2(net1807),
    .Y(_4458_),
    .B1(_4457_));
 sg13g2_nor3_1 _8989_ (.A(_1963_),
    .B(_4456_),
    .C(_4458_),
    .Y(_4459_));
 sg13g2_nor2_1 _8990_ (.A(net1731),
    .B(_4459_),
    .Y(_4460_));
 sg13g2_o21ai_1 _8991_ (.B1(_4460_),
    .Y(_4461_),
    .A1(net1797),
    .A2(_2423_));
 sg13g2_a21oi_2 _8992_ (.B1(_4393_),
    .Y(_4462_),
    .A2(net1730),
    .A1(_2173_));
 sg13g2_a22oi_1 _8993_ (.Y(_4463_),
    .B1(_4410_),
    .B2(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(_4407_),
    .A1(\z80.tv80s.i_tv80_core.F[4] ));
 sg13g2_a22oi_1 _8994_ (.Y(_4464_),
    .B1(_4411_),
    .B2(\z80.tv80s.i_tv80_core.SP[12] ),
    .A2(_4404_),
    .A1(\z80.tv80s.i_tv80_core.SP[4] ));
 sg13g2_a22oi_1 _8995_ (.Y(_4465_),
    .B1(_4406_),
    .B2(net2047),
    .A2(_4401_),
    .A1(\z80.tv80s.i_tv80_core.PC[12] ));
 sg13g2_nand3_1 _8996_ (.B(_4464_),
    .C(_4465_),
    .A(_4463_),
    .Y(_4466_));
 sg13g2_a221oi_1 _8997_ (.B2(_4462_),
    .C1(_4466_),
    .B1(_4461_),
    .A1(\z80.tv80s.i_tv80_core.PC[4] ),
    .Y(_4467_),
    .A2(_4408_));
 sg13g2_o21ai_1 _8998_ (.B1(_4454_),
    .Y(_0649_),
    .A1(_4366_),
    .A2(_4467_));
 sg13g2_nand2_1 _8999_ (.Y(_4468_),
    .A(net594),
    .B(net1970));
 sg13g2_nand2b_1 _9000_ (.Y(_4469_),
    .B(_1963_),
    .A_N(_2419_));
 sg13g2_o21ai_1 _9001_ (.B1(net1785),
    .Y(_4470_),
    .A1(_0083_),
    .A2(net2164));
 sg13g2_a21oi_1 _9002_ (.A1(_0709_),
    .A2(net1807),
    .Y(_4471_),
    .B1(_4470_));
 sg13g2_o21ai_1 _9003_ (.B1(net1802),
    .Y(_4472_),
    .A1(_0079_),
    .A2(net2164));
 sg13g2_o21ai_1 _9004_ (.B1(net1797),
    .Y(_4473_),
    .A1(_2421_),
    .A2(_4472_));
 sg13g2_nor2_1 _9005_ (.A(_4471_),
    .B(_4473_),
    .Y(_4474_));
 sg13g2_nor2_1 _9006_ (.A(net1731),
    .B(_4474_),
    .Y(_4475_));
 sg13g2_a221oi_1 _9007_ (.B2(_4475_),
    .C1(_4393_),
    .B1(_4469_),
    .A1(_2120_),
    .Y(_4476_),
    .A2(net1730));
 sg13g2_nand2_1 _9008_ (.Y(_4477_),
    .A(\z80.tv80s.i_tv80_core.SP[3] ),
    .B(_4404_));
 sg13g2_a22oi_1 _9009_ (.Y(_4478_),
    .B1(_4410_),
    .B2(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_4408_),
    .A1(\z80.tv80s.i_tv80_core.PC[3] ));
 sg13g2_a22oi_1 _9010_ (.Y(_4479_),
    .B1(_4411_),
    .B2(\z80.tv80s.i_tv80_core.SP[11] ),
    .A2(_4407_),
    .A1(\z80.tv80s.i_tv80_core.F[3] ));
 sg13g2_a221oi_1 _9011_ (.B2(net2048),
    .C1(_4476_),
    .B1(_4406_),
    .A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .Y(_4480_),
    .A2(_4401_));
 sg13g2_and4_2 _9012_ (.A(_4477_),
    .B(_4478_),
    .C(_4479_),
    .D(_4480_),
    .X(_4481_));
 sg13g2_o21ai_1 _9013_ (.B1(_4468_),
    .Y(_0650_),
    .A1(_4366_),
    .A2(_4481_));
 sg13g2_nand2_1 _9014_ (.Y(_4482_),
    .A(net542),
    .B(net1969));
 sg13g2_o21ai_1 _9015_ (.B1(net1786),
    .Y(_4483_),
    .A1(_0060_),
    .A2(net1813));
 sg13g2_a21oi_1 _9016_ (.A1(_0702_),
    .A2(net2010),
    .Y(_4484_),
    .B1(_4483_));
 sg13g2_nor2_1 _9017_ (.A(_0056_),
    .B(net1813),
    .Y(_4485_));
 sg13g2_o21ai_1 _9018_ (.B1(net1805),
    .Y(_4486_),
    .A1(_0055_),
    .A2(net2163));
 sg13g2_o21ai_1 _9019_ (.B1(net1799),
    .Y(_4487_),
    .A1(_4485_),
    .A2(_4486_));
 sg13g2_o21ai_1 _9020_ (.B1(net1730),
    .Y(_4488_),
    .A1(_4484_),
    .A2(_4487_));
 sg13g2_nor3_1 _9021_ (.A(_2406_),
    .B(_2411_),
    .C(net1731),
    .Y(_4489_));
 sg13g2_nor2_1 _9022_ (.A(_4393_),
    .B(_4489_),
    .Y(_4490_));
 sg13g2_o21ai_1 _9023_ (.B1(_4490_),
    .Y(_4491_),
    .A1(_2067_),
    .A2(_4488_));
 sg13g2_a22oi_1 _9024_ (.Y(_4492_),
    .B1(_4407_),
    .B2(\z80.tv80s.i_tv80_core.F[2] ),
    .A2(_4401_),
    .A1(\z80.tv80s.i_tv80_core.PC[10] ));
 sg13g2_a22oi_1 _9025_ (.Y(_4493_),
    .B1(_4411_),
    .B2(\z80.tv80s.i_tv80_core.SP[10] ),
    .A2(_4408_),
    .A1(\z80.tv80s.i_tv80_core.PC[2] ));
 sg13g2_a22oi_1 _9026_ (.Y(_4494_),
    .B1(_4406_),
    .B2(\z80.tv80s.di_reg[2] ),
    .A2(_4404_),
    .A1(\z80.tv80s.i_tv80_core.SP[2] ));
 sg13g2_nand4_1 _9027_ (.B(_4492_),
    .C(_4493_),
    .A(_4491_),
    .Y(_4495_),
    .D(_4494_));
 sg13g2_a21oi_2 _9028_ (.B1(_4495_),
    .Y(_4496_),
    .A2(_4410_),
    .A1(\z80.tv80s.i_tv80_core.ACC[2] ));
 sg13g2_o21ai_1 _9029_ (.B1(_4482_),
    .Y(_0651_),
    .A1(_4366_),
    .A2(_4496_));
 sg13g2_nand2_1 _9030_ (.Y(_4497_),
    .A(net562),
    .B(net1970));
 sg13g2_o21ai_1 _9031_ (.B1(net1785),
    .Y(_4498_),
    .A1(_0166_),
    .A2(net1812));
 sg13g2_a21oi_1 _9032_ (.A1(net2009),
    .A2(_0743_),
    .Y(_4499_),
    .B1(_4498_));
 sg13g2_o21ai_1 _9033_ (.B1(net1802),
    .Y(_4500_),
    .A1(_0162_),
    .A2(net1812));
 sg13g2_a21oi_1 _9034_ (.A1(net2009),
    .A2(_0742_),
    .Y(_4501_),
    .B1(_4500_));
 sg13g2_o21ai_1 _9035_ (.B1(net1797),
    .Y(_4502_),
    .A1(_4499_),
    .A2(_4501_));
 sg13g2_a21oi_2 _9036_ (.B1(net1731),
    .Y(_4503_),
    .A2(_4502_),
    .A1(_2399_));
 sg13g2_o21ai_1 _9037_ (.B1(net1804),
    .Y(_4504_),
    .A1(_0047_),
    .A2(net2163));
 sg13g2_a21oi_1 _9038_ (.A1(_0697_),
    .A2(net1809),
    .Y(_4505_),
    .B1(_4504_));
 sg13g2_o21ai_1 _9039_ (.B1(net1786),
    .Y(_4506_),
    .A1(_0051_),
    .A2(net2163));
 sg13g2_a21oi_1 _9040_ (.A1(_0698_),
    .A2(net1809),
    .Y(_4507_),
    .B1(_4506_));
 sg13g2_nor3_1 _9041_ (.A(_1963_),
    .B(_4505_),
    .C(_4507_),
    .Y(_4508_));
 sg13g2_nor2_2 _9042_ (.A(_2019_),
    .B(_4508_),
    .Y(_4509_));
 sg13g2_a21oi_2 _9043_ (.B1(_4503_),
    .Y(_4510_),
    .A2(_4509_),
    .A1(net1731));
 sg13g2_a22oi_1 _9044_ (.Y(_4511_),
    .B1(_4410_),
    .B2(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_4404_),
    .A1(\z80.tv80s.i_tv80_core.SP[1] ));
 sg13g2_a22oi_1 _9045_ (.Y(_4512_),
    .B1(_4408_),
    .B2(\z80.tv80s.i_tv80_core.PC[1] ),
    .A2(_4401_),
    .A1(\z80.tv80s.i_tv80_core.PC[9] ));
 sg13g2_a22oi_1 _9046_ (.Y(_4513_),
    .B1(_4407_),
    .B2(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_4406_),
    .A1(\z80.tv80s.di_reg[1] ));
 sg13g2_nand3_1 _9047_ (.B(_4512_),
    .C(_4513_),
    .A(_4511_),
    .Y(_4514_));
 sg13g2_a221oi_1 _9048_ (.B2(_4392_),
    .C1(_4514_),
    .B1(_4510_),
    .A1(\z80.tv80s.i_tv80_core.SP[9] ),
    .Y(_4515_),
    .A2(_4411_));
 sg13g2_o21ai_1 _9049_ (.B1(_4497_),
    .Y(_0652_),
    .A1(_4366_),
    .A2(_4515_));
 sg13g2_nand2_1 _9050_ (.Y(_4516_),
    .A(net582),
    .B(net1971));
 sg13g2_nor2_1 _9051_ (.A(_0154_),
    .B(net1812),
    .Y(_4517_));
 sg13g2_o21ai_1 _9052_ (.B1(net1803),
    .Y(_4518_),
    .A1(net2164),
    .A2(_0153_));
 sg13g2_a22oi_1 _9053_ (.Y(_4519_),
    .B1(net1808),
    .B2(_0738_),
    .A2(_0739_),
    .A1(net2010));
 sg13g2_a21oi_1 _9054_ (.A1(net1785),
    .A2(_4519_),
    .Y(_4520_),
    .B1(_1963_));
 sg13g2_o21ai_1 _9055_ (.B1(_4520_),
    .Y(_4521_),
    .A1(_4517_),
    .A2(_4518_));
 sg13g2_o21ai_1 _9056_ (.B1(_4521_),
    .Y(_4522_),
    .A1(net1798),
    .A2(_2387_));
 sg13g2_mux2_2 _9057_ (.A0(_1969_),
    .A1(_4522_),
    .S(_4384_),
    .X(_4523_));
 sg13g2_o21ai_1 _9058_ (.B1(_4403_),
    .Y(_4524_),
    .A1(\z80.tv80s.i_tv80_core.SP[0] ),
    .A2(_1584_));
 sg13g2_a22oi_1 _9059_ (.Y(_4525_),
    .B1(_4408_),
    .B2(\z80.tv80s.i_tv80_core.PC[0] ),
    .A2(_4407_),
    .A1(net2151));
 sg13g2_a22oi_1 _9060_ (.Y(_4526_),
    .B1(_4411_),
    .B2(\z80.tv80s.i_tv80_core.SP[8] ),
    .A2(_4406_),
    .A1(\z80.tv80s.di_reg[0] ));
 sg13g2_a22oi_1 _9061_ (.Y(_4527_),
    .B1(_4410_),
    .B2(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A2(_4401_),
    .A1(\z80.tv80s.i_tv80_core.PC[8] ));
 sg13g2_nand4_1 _9062_ (.B(_4525_),
    .C(_4526_),
    .A(_4524_),
    .Y(_4528_),
    .D(_4527_));
 sg13g2_a21oi_2 _9063_ (.B1(_4528_),
    .Y(_4529_),
    .A2(_4523_),
    .A1(_4392_));
 sg13g2_o21ai_1 _9064_ (.B1(_4516_),
    .Y(_0653_),
    .A1(_4366_),
    .A2(_4529_));
 sg13g2_dfrbp_1 _9065_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2198),
    .D(net564),
    .Q_N(_4618_),
    .Q(\z80.tv80s.i_tv80_core.R[0] ));
 sg13g2_dfrbp_1 _9066_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2198),
    .D(net504),
    .Q_N(_4617_),
    .Q(\z80.tv80s.i_tv80_core.R[1] ));
 sg13g2_dfrbp_1 _9067_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2194),
    .D(net541),
    .Q_N(_4616_),
    .Q(\z80.tv80s.i_tv80_core.R[2] ));
 sg13g2_dfrbp_1 _9068_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2194),
    .D(net538),
    .Q_N(_4615_),
    .Q(\z80.tv80s.i_tv80_core.R[3] ));
 sg13g2_dfrbp_1 _9069_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2189),
    .D(net522),
    .Q_N(_4614_),
    .Q(\z80.tv80s.i_tv80_core.R[4] ));
 sg13g2_dfrbp_1 _9070_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2194),
    .D(_0302_),
    .Q_N(_4613_),
    .Q(\z80.tv80s.i_tv80_core.R[5] ));
 sg13g2_dfrbp_1 _9071_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2194),
    .D(_0303_),
    .Q_N(_4612_),
    .Q(\z80.tv80s.i_tv80_core.R[6] ));
 sg13g2_dfrbp_1 _9072_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net59),
    .D(_0304_),
    .Q_N(_4611_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sg13g2_dfrbp_1 _9073_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net58),
    .D(_0305_),
    .Q_N(_4610_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sg13g2_dfrbp_1 _9074_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net57),
    .D(net194),
    .Q_N(_0150_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ));
 sg13g2_dfrbp_1 _9075_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net21),
    .D(net188),
    .Q_N(_0040_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ));
 sg13g2_dfrbp_1 _9076_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2219),
    .D(_0012_),
    .Q_N(_4619_),
    .Q(\z80.tv80s.i_tv80_core.mcycles[1] ));
 sg13g2_dfrbp_1 _9077_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2219),
    .D(_0013_),
    .Q_N(_4620_),
    .Q(\z80.tv80s.i_tv80_core.mcycles[2] ));
 sg13g2_dfrbp_1 _9078_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2221),
    .D(_0014_),
    .Q_N(_4621_),
    .Q(\z80.tv80s.i_tv80_core.mcycles[4] ));
 sg13g2_dfrbp_1 _9079_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2224),
    .D(_0015_),
    .Q_N(_4609_),
    .Q(\z80.tv80s.i_tv80_core.mcycles[5] ));
 sg13g2_dfrbp_1 _9080_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2205),
    .D(_0308_),
    .Q_N(_4608_),
    .Q(\z80.tv80s.i_tv80_core.PreserveC_r ));
 sg13g2_dfrbp_1 _9081_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2222),
    .D(net548),
    .Q_N(\z80.tv80s.i_tv80_core.ISet[0] ),
    .Q(_0239_));
 sg13g2_dfrbp_1 _9082_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2222),
    .D(_0000_),
    .Q_N(_4622_),
    .Q(\z80.tv80s.i_tv80_core.ISet[1] ));
 sg13g2_dfrbp_1 _9083_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2222),
    .D(_0001_),
    .Q_N(_0033_),
    .Q(\z80.tv80s.i_tv80_core.ISet[2] ));
 sg13g2_dfrbp_1 _9084_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2205),
    .D(_0002_),
    .Q_N(_4607_),
    .Q(\z80.tv80s.i_tv80_core.ISet[3] ));
 sg13g2_dfrbp_1 _9085_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net56),
    .D(_0309_),
    .Q_N(_0043_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ));
 sg13g2_dfrbp_1 _9086_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net55),
    .D(_0310_),
    .Q_N(_0051_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ));
 sg13g2_dfrbp_1 _9087_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net54),
    .D(_0311_),
    .Q_N(_0059_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ));
 sg13g2_dfrbp_1 _9088_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net53),
    .D(_0312_),
    .Q_N(_0075_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ));
 sg13g2_dfrbp_1 _9089_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net52),
    .D(_0313_),
    .Q_N(_0091_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ));
 sg13g2_dfrbp_1 _9090_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net51),
    .D(_0314_),
    .Q_N(_0107_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ));
 sg13g2_dfrbp_1 _9091_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net50),
    .D(_0315_),
    .Q_N(_0123_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ));
 sg13g2_dfrbp_1 _9092_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net49),
    .D(_0316_),
    .Q_N(_0139_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ));
 sg13g2_dfrbp_1 _9093_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net48),
    .D(_0317_),
    .Q_N(_0042_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ));
 sg13g2_dfrbp_1 _9094_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net47),
    .D(_0318_),
    .Q_N(_0050_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ));
 sg13g2_dfrbp_1 _9095_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net46),
    .D(_0319_),
    .Q_N(_0058_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ));
 sg13g2_dfrbp_1 _9096_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net45),
    .D(_0320_),
    .Q_N(_0074_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ));
 sg13g2_dfrbp_1 _9097_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net44),
    .D(_0321_),
    .Q_N(_0090_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ));
 sg13g2_dfrbp_1 _9098_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net43),
    .D(_0322_),
    .Q_N(_0106_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ));
 sg13g2_dfrbp_1 _9099_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net42),
    .D(_0323_),
    .Q_N(_0122_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ));
 sg13g2_dfrbp_1 _9100_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net41),
    .D(_0324_),
    .Q_N(_0138_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ));
 sg13g2_dfrbp_1 _9101_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net40),
    .D(_0325_),
    .Q_N(_0041_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ));
 sg13g2_dfrbp_1 _9102_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net39),
    .D(_0326_),
    .Q_N(_0049_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ));
 sg13g2_dfrbp_1 _9103_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net38),
    .D(_0327_),
    .Q_N(_0057_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ));
 sg13g2_dfrbp_1 _9104_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net37),
    .D(_0328_),
    .Q_N(_0073_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ));
 sg13g2_dfrbp_1 _9105_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net36),
    .D(_0329_),
    .Q_N(_0089_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ));
 sg13g2_dfrbp_1 _9106_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net35),
    .D(_0330_),
    .Q_N(_0105_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ));
 sg13g2_dfrbp_1 _9107_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net34),
    .D(_0331_),
    .Q_N(_0121_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ));
 sg13g2_dfrbp_1 _9108_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net33),
    .D(_0332_),
    .Q_N(_0137_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ));
 sg13g2_dfrbp_1 _9109_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net32),
    .D(_0333_),
    .Q_N(_0038_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ));
 sg13g2_dfrbp_1 _9110_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net31),
    .D(_0334_),
    .Q_N(_0048_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ));
 sg13g2_dfrbp_1 _9111_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net30),
    .D(_0335_),
    .Q_N(_0056_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ));
 sg13g2_dfrbp_1 _9112_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net29),
    .D(_0336_),
    .Q_N(_0072_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ));
 sg13g2_dfrbp_1 _9113_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net28),
    .D(_0337_),
    .Q_N(_0088_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ));
 sg13g2_dfrbp_1 _9114_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net27),
    .D(_0338_),
    .Q_N(_0104_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ));
 sg13g2_dfrbp_1 _9115_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net26),
    .D(_0339_),
    .Q_N(_0120_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ));
 sg13g2_dfrbp_1 _9116_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net25),
    .D(_0340_),
    .Q_N(_0136_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ));
 sg13g2_dfrbp_1 _9117_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2210),
    .D(_0341_),
    .Q_N(\z80.tv80s.wr_n ),
    .Q(_0240_));
 sg13g2_dfrbp_1 _9118_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2209),
    .D(_0342_),
    .Q_N(\z80.iorq_n ),
    .Q(_0241_));
 sg13g2_dfrbp_1 _9119_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2210),
    .D(_0343_),
    .Q_N(\z80.rd_n ),
    .Q(_0242_));
 sg13g2_dfrbp_1 _9120_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2210),
    .D(net327),
    .Q_N(\z80.mreq_n ),
    .Q(_0243_));
 sg13g2_dfrbp_1 _9121_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net18),
    .D(_0345_),
    .Q_N(_0157_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ));
 sg13g2_dfrbp_1 _9122_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net17),
    .D(_0346_),
    .Q_N(_0165_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ));
 sg13g2_dfrbp_1 _9123_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net16),
    .D(_0347_),
    .Q_N(_0067_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ));
 sg13g2_dfrbp_1 _9124_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net15),
    .D(_0348_),
    .Q_N(_0083_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ));
 sg13g2_dfrbp_1 _9125_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net14),
    .D(_0349_),
    .Q_N(_0099_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ));
 sg13g2_dfrbp_1 _9126_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net13),
    .D(_0350_),
    .Q_N(_0115_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ));
 sg13g2_dfrbp_1 _9127_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net182),
    .D(_0351_),
    .Q_N(_0131_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ));
 sg13g2_dfrbp_1 _9128_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net181),
    .D(_0352_),
    .Q_N(_0147_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ));
 sg13g2_dfrbp_1 _9129_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net180),
    .D(_0353_),
    .Q_N(_0044_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ));
 sg13g2_dfrbp_1 _9130_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net179),
    .D(_0354_),
    .Q_N(_0052_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ));
 sg13g2_dfrbp_1 _9131_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net178),
    .D(_0355_),
    .Q_N(_0060_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ));
 sg13g2_dfrbp_1 _9132_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net177),
    .D(_0356_),
    .Q_N(_0076_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ));
 sg13g2_dfrbp_1 _9133_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net176),
    .D(_0357_),
    .Q_N(_0092_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ));
 sg13g2_dfrbp_1 _9134_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net175),
    .D(_0358_),
    .Q_N(_0108_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ));
 sg13g2_dfrbp_1 _9135_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net174),
    .D(_0359_),
    .Q_N(_0124_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ));
 sg13g2_dfrbp_1 _9136_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net173),
    .D(_0360_),
    .Q_N(_0140_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ));
 sg13g2_dfrbp_1 _9137_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net172),
    .D(_0361_),
    .Q_N(_0156_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ));
 sg13g2_dfrbp_1 _9138_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net171),
    .D(_0362_),
    .Q_N(_0164_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ));
 sg13g2_dfrbp_1 _9139_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net170),
    .D(_0363_),
    .Q_N(_0066_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ));
 sg13g2_dfrbp_1 _9140_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net169),
    .D(_0364_),
    .Q_N(_0082_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ));
 sg13g2_dfrbp_1 _9141_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net168),
    .D(_0365_),
    .Q_N(_0098_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ));
 sg13g2_dfrbp_1 _9142_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net167),
    .D(_0366_),
    .Q_N(_0114_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ));
 sg13g2_dfrbp_1 _9143_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net166),
    .D(_0367_),
    .Q_N(_0130_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ));
 sg13g2_dfrbp_1 _9144_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net165),
    .D(_0368_),
    .Q_N(_0146_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ));
 sg13g2_dfrbp_1 _9145_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net164),
    .D(_0369_),
    .Q_N(_0036_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ));
 sg13g2_dfrbp_1 _9146_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net163),
    .D(_0370_),
    .Q_N(_0046_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ));
 sg13g2_dfrbp_1 _9147_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net162),
    .D(_0371_),
    .Q_N(_0054_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ));
 sg13g2_dfrbp_1 _9148_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net161),
    .D(_0372_),
    .Q_N(_0070_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ));
 sg13g2_dfrbp_1 _9149_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net160),
    .D(_0373_),
    .Q_N(_0086_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ));
 sg13g2_dfrbp_1 _9150_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net159),
    .D(_0374_),
    .Q_N(_0102_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ));
 sg13g2_dfrbp_1 _9151_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net158),
    .D(_0375_),
    .Q_N(_0118_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ));
 sg13g2_dfrbp_1 _9152_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net157),
    .D(_0376_),
    .Q_N(_0134_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ));
 sg13g2_dfrbp_1 _9153_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net156),
    .D(_0377_),
    .Q_N(_0151_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ));
 sg13g2_dfrbp_1 _9154_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net155),
    .D(_0378_),
    .Q_N(_0159_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ));
 sg13g2_dfrbp_1 _9155_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net154),
    .D(_0379_),
    .Q_N(_0061_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ));
 sg13g2_dfrbp_1 _9156_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net153),
    .D(_0380_),
    .Q_N(_0077_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ));
 sg13g2_dfrbp_1 _9157_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net152),
    .D(_0381_),
    .Q_N(_0093_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ));
 sg13g2_dfrbp_1 _9158_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net151),
    .D(_0382_),
    .Q_N(_0109_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ));
 sg13g2_dfrbp_1 _9159_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net150),
    .D(_0383_),
    .Q_N(_0125_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ));
 sg13g2_dfrbp_1 _9160_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net149),
    .D(_0384_),
    .Q_N(_0141_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ));
 sg13g2_dfrbp_1 _9161_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net148),
    .D(_0385_),
    .Q_N(_0152_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ));
 sg13g2_dfrbp_1 _9162_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net147),
    .D(_0386_),
    .Q_N(_0160_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ));
 sg13g2_dfrbp_1 _9163_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net146),
    .D(_0387_),
    .Q_N(_0062_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ));
 sg13g2_dfrbp_1 _9164_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net145),
    .D(_0388_),
    .Q_N(_0078_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ));
 sg13g2_dfrbp_1 _9165_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net144),
    .D(_0389_),
    .Q_N(_0094_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ));
 sg13g2_dfrbp_1 _9166_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net143),
    .D(_0390_),
    .Q_N(_0110_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ));
 sg13g2_dfrbp_1 _9167_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net142),
    .D(_0391_),
    .Q_N(_0126_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ));
 sg13g2_dfrbp_1 _9168_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net141),
    .D(_0392_),
    .Q_N(_0142_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ));
 sg13g2_dfrbp_1 _9169_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net140),
    .D(_0393_),
    .Q_N(_0037_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ));
 sg13g2_dfrbp_1 _9170_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net139),
    .D(_0394_),
    .Q_N(_0047_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ));
 sg13g2_dfrbp_1 _9171_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net138),
    .D(_0395_),
    .Q_N(_0055_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ));
 sg13g2_dfrbp_1 _9172_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net137),
    .D(_0396_),
    .Q_N(_0071_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ));
 sg13g2_dfrbp_1 _9173_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net136),
    .D(_0397_),
    .Q_N(_0087_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ));
 sg13g2_dfrbp_1 _9174_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net135),
    .D(_0398_),
    .Q_N(_0103_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ));
 sg13g2_dfrbp_1 _9175_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net134),
    .D(_0399_),
    .Q_N(_0119_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ));
 sg13g2_dfrbp_1 _9176_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net133),
    .D(_0400_),
    .Q_N(_0135_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ));
 sg13g2_dfrbp_1 _9177_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net132),
    .D(_0401_),
    .Q_N(_0154_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ));
 sg13g2_dfrbp_1 _9178_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net131),
    .D(_0402_),
    .Q_N(_0162_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ));
 sg13g2_dfrbp_1 _9179_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net130),
    .D(_0403_),
    .Q_N(_0064_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ));
 sg13g2_dfrbp_1 _9180_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net129),
    .D(_0404_),
    .Q_N(_0080_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ));
 sg13g2_dfrbp_1 _9181_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net128),
    .D(_0405_),
    .Q_N(_0096_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ));
 sg13g2_dfrbp_1 _9182_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net127),
    .D(_0406_),
    .Q_N(_0112_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ));
 sg13g2_dfrbp_1 _9183_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net126),
    .D(_0407_),
    .Q_N(_0128_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ));
 sg13g2_dfrbp_1 _9184_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net125),
    .D(_0408_),
    .Q_N(_0144_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ));
 sg13g2_dfrbp_1 _9185_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net124),
    .D(_0409_),
    .Q_N(_0155_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ));
 sg13g2_dfrbp_1 _9186_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net123),
    .D(_0410_),
    .Q_N(_0163_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ));
 sg13g2_dfrbp_1 _9187_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net122),
    .D(_0411_),
    .Q_N(_0065_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ));
 sg13g2_dfrbp_1 _9188_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net121),
    .D(_0412_),
    .Q_N(_0081_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ));
 sg13g2_dfrbp_1 _9189_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net120),
    .D(_0413_),
    .Q_N(_0097_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ));
 sg13g2_dfrbp_1 _9190_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net119),
    .D(_0414_),
    .Q_N(_0113_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ));
 sg13g2_dfrbp_1 _9191_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net118),
    .D(_0415_),
    .Q_N(_0129_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ));
 sg13g2_dfrbp_1 _9192_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net117),
    .D(_0416_),
    .Q_N(_0145_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ));
 sg13g2_dfrbp_1 _9193_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net116),
    .D(_0417_),
    .Q_N(_0158_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ));
 sg13g2_dfrbp_1 _9194_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net115),
    .D(_0418_),
    .Q_N(_0166_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ));
 sg13g2_dfrbp_1 _9195_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net114),
    .D(_0419_),
    .Q_N(_0068_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ));
 sg13g2_dfrbp_1 _9196_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net113),
    .D(_0420_),
    .Q_N(_0084_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ));
 sg13g2_dfrbp_1 _9197_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net112),
    .D(_0421_),
    .Q_N(_0100_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ));
 sg13g2_dfrbp_1 _9198_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net111),
    .D(_0422_),
    .Q_N(_0116_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ));
 sg13g2_dfrbp_1 _9199_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net110),
    .D(_0423_),
    .Q_N(_0132_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ));
 sg13g2_dfrbp_1 _9200_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net64),
    .D(_0424_),
    .Q_N(_0148_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ));
 sg13g2_dfrbp_1 _9201_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2224),
    .D(net345),
    .Q_N(_4623_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ));
 sg13g2_dfrbp_1 _9202_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2223),
    .D(_0006_),
    .Q_N(_4624_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ));
 sg13g2_dfrbp_1 _9203_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2223),
    .D(_0007_),
    .Q_N(_4625_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ));
 sg13g2_dfrbp_1 _9204_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2225),
    .D(_0008_),
    .Q_N(_4626_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ));
 sg13g2_dfrbp_1 _9205_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2223),
    .D(net489),
    .Q_N(_4627_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ));
 sg13g2_dfrbp_1 _9206_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2223),
    .D(_0010_),
    .Q_N(_4628_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ));
 sg13g2_dfrbp_1 _9207_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2223),
    .D(_0011_),
    .Q_N(_4606_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ));
 sg13g2_dfrbp_1 _9208_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net109),
    .D(_0425_),
    .Q_N(_0035_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ));
 sg13g2_dfrbp_1 _9209_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net108),
    .D(_0426_),
    .Q_N(_0045_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ));
 sg13g2_dfrbp_1 _9210_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net107),
    .D(_0427_),
    .Q_N(_0053_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ));
 sg13g2_dfrbp_1 _9211_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net106),
    .D(_0428_),
    .Q_N(_0069_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ));
 sg13g2_dfrbp_1 _9212_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net105),
    .D(_0429_),
    .Q_N(_0085_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ));
 sg13g2_dfrbp_1 _9213_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net104),
    .D(_0430_),
    .Q_N(_0101_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ));
 sg13g2_dfrbp_1 _9214_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net103),
    .D(_0431_),
    .Q_N(_0117_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ));
 sg13g2_dfrbp_1 _9215_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net66),
    .D(_0432_),
    .Q_N(_0133_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ));
 sg13g2_dfrbp_1 _9216_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2205),
    .D(_0003_),
    .Q_N(_4629_),
    .Q(\z80.tv80s.i_tv80_core.IStatus[1] ));
 sg13g2_dfrbp_1 _9217_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2205),
    .D(_0004_),
    .Q_N(_4605_),
    .Q(\z80.tv80s.i_tv80_core.IStatus[2] ));
 sg13g2_dfrbp_1 _9218_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net102),
    .D(_0433_),
    .Q_N(_0153_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ));
 sg13g2_dfrbp_1 _9219_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net101),
    .D(_0434_),
    .Q_N(_0161_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ));
 sg13g2_dfrbp_1 _9220_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net100),
    .D(_0435_),
    .Q_N(_0063_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ));
 sg13g2_dfrbp_1 _9221_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net99),
    .D(_0436_),
    .Q_N(_0079_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ));
 sg13g2_dfrbp_1 _9222_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net98),
    .D(_0437_),
    .Q_N(_0095_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ));
 sg13g2_dfrbp_1 _9223_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net97),
    .D(_0438_),
    .Q_N(_0111_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ));
 sg13g2_dfrbp_1 _9224_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net96),
    .D(_0439_),
    .Q_N(_0127_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ));
 sg13g2_dfrbp_1 _9225_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net95),
    .D(_0440_),
    .Q_N(_0143_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ));
 sg13g2_dfrbp_1 _9226_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2207),
    .D(net486),
    .Q_N(_0227_),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ));
 sg13g2_dfrbp_1 _9227_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2210),
    .D(net493),
    .Q_N(_0168_),
    .Q(\z80.tv80s.i_tv80_core.BusAck ));
 sg13g2_dfrbp_1 _9228_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2219),
    .D(net581),
    .Q_N(_0016_),
    .Q(\z80.tv80s.i_tv80_core.NMICycle ));
 sg13g2_dfrbp_1 _9229_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2209),
    .D(net472),
    .Q_N(_4604_),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ));
 sg13g2_dfrbp_1 _9230_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2220),
    .D(_0445_),
    .Q_N(_4603_),
    .Q(\z80.tv80s.i_tv80_core.BusReq_s ));
 sg13g2_dfrbp_1 _9231_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2220),
    .D(net227),
    .Q_N(_4630_),
    .Q(\z80.tv80s.i_tv80_core.NMI_s ));
 sg13g2_dfrbp_1 _9232_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2221),
    .D(_0017_),
    .Q_N(_4631_),
    .Q(_0236_));
 sg13g2_dfrbp_1 _9233_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2221),
    .D(_0018_),
    .Q_N(_4632_),
    .Q(_0237_));
 sg13g2_dfrbp_1 _9234_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2223),
    .D(_0019_),
    .Q_N(_4602_),
    .Q(_0238_));
 sg13g2_dfrbp_1 _9235_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2220),
    .D(_0447_),
    .Q_N(_4601_),
    .Q(\z80.tv80s.i_tv80_core.INT_s ));
 sg13g2_dfrbp_1 _9236_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2209),
    .D(_0448_),
    .Q_N(_4600_),
    .Q(\z80.tv80s.i_tv80_core.Oldnmi_n ));
 sg13g2_dfrbp_1 _9237_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2207),
    .D(_0449_),
    .Q_N(\z80.rfsh_n ),
    .Q(_0244_));
 sg13g2_dfrbp_1 _9238_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net92),
    .D(_0450_),
    .Q_N(_4599_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ));
 sg13g2_dfrbp_1 _9239_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net91),
    .D(_0451_),
    .Q_N(_4598_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ));
 sg13g2_dfrbp_1 _9240_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net89),
    .D(_0452_),
    .Q_N(_4597_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sg13g2_dfrbp_1 _9241_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net87),
    .D(_0453_),
    .Q_N(_4596_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sg13g2_dfrbp_1 _9242_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net86),
    .D(_0454_),
    .Q_N(_4595_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sg13g2_dfrbp_1 _9243_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net84),
    .D(_0455_),
    .Q_N(_4594_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[0] ));
 sg13g2_dfrbp_1 _9244_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net83),
    .D(_0456_),
    .Q_N(_4593_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[1] ));
 sg13g2_dfrbp_1 _9245_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net82),
    .D(_0457_),
    .Q_N(_4592_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[2] ));
 sg13g2_dfrbp_1 _9246_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net81),
    .D(net367),
    .Q_N(_4591_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[3] ));
 sg13g2_dfrbp_1 _9247_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net80),
    .D(net363),
    .Q_N(_4590_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[4] ));
 sg13g2_dfrbp_1 _9248_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net79),
    .D(net355),
    .Q_N(_4589_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[5] ));
 sg13g2_dfrbp_1 _9249_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net78),
    .D(net422),
    .Q_N(_4588_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[6] ));
 sg13g2_dfrbp_1 _9250_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net77),
    .D(net445),
    .Q_N(_4587_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[7] ));
 sg13g2_dfrbp_1 _9251_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net76),
    .D(net358),
    .Q_N(_4586_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[8] ));
 sg13g2_dfrbp_1 _9252_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net75),
    .D(_0464_),
    .Q_N(_4585_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[9] ));
 sg13g2_dfrbp_1 _9253_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net74),
    .D(net397),
    .Q_N(_4584_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[10] ));
 sg13g2_dfrbp_1 _9254_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net73),
    .D(_0466_),
    .Q_N(_4583_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[11] ));
 sg13g2_dfrbp_1 _9255_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net72),
    .D(net348),
    .Q_N(_4582_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[12] ));
 sg13g2_dfrbp_1 _9256_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net71),
    .D(net319),
    .Q_N(_4581_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[13] ));
 sg13g2_dfrbp_1 _9257_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net70),
    .D(_0469_),
    .Q_N(_4580_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[14] ));
 sg13g2_dfrbp_1 _9258_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net69),
    .D(net304),
    .Q_N(_4579_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[15] ));
 sg13g2_dfrbp_1 _9259_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net68),
    .D(_0471_),
    .Q_N(_4578_),
    .Q(\z80.tv80s.i_tv80_core.IncDecZ ));
 sg13g2_dfrbp_1 _9260_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2209),
    .D(net468),
    .Q_N(_0167_),
    .Q(\z80.tv80s.i_tv80_core.Halt_FF ));
 sg13g2_dfrbp_1 _9261_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2200),
    .D(net482),
    .Q_N(_4577_),
    .Q(\addr_bus[0] ));
 sg13g2_dfrbp_1 _9262_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2207),
    .D(_0474_),
    .Q_N(_4576_),
    .Q(\addr_bus[1] ));
 sg13g2_dfrbp_1 _9263_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2202),
    .D(_0475_),
    .Q_N(_4575_),
    .Q(\addr_bus[2] ));
 sg13g2_dfrbp_1 _9264_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2203),
    .D(_0476_),
    .Q_N(_4574_),
    .Q(\addr_bus[3] ));
 sg13g2_dfrbp_1 _9265_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2203),
    .D(_0477_),
    .Q_N(_4573_),
    .Q(\addr_bus[4] ));
 sg13g2_dfrbp_1 _9266_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2202),
    .D(_0478_),
    .Q_N(_4572_),
    .Q(\addr_bus[5] ));
 sg13g2_dfrbp_1 _9267_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2198),
    .D(net501),
    .Q_N(_4571_),
    .Q(\addr_bus[6] ));
 sg13g2_dfrbp_1 _9268_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net2206),
    .D(net458),
    .Q_N(_4570_),
    .Q(\addr_bus[7] ));
 sg13g2_dfrbp_1 _9269_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2198),
    .D(net480),
    .Q_N(_4569_),
    .Q(\addr_bus[8] ));
 sg13g2_dfrbp_1 _9270_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2207),
    .D(_0482_),
    .Q_N(_4568_),
    .Q(\addr_bus[9] ));
 sg13g2_dfrbp_1 _9271_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2208),
    .D(_0483_),
    .Q_N(_4567_),
    .Q(\addr_bus[10] ));
 sg13g2_dfrbp_1 _9272_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2208),
    .D(_0484_),
    .Q_N(_4566_),
    .Q(\addr_bus[11] ));
 sg13g2_dfrbp_1 _9273_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2207),
    .D(_0485_),
    .Q_N(_4565_),
    .Q(\addr_bus[12] ));
 sg13g2_dfrbp_1 _9274_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2208),
    .D(_0486_),
    .Q_N(_4564_),
    .Q(\addr_bus[13] ));
 sg13g2_dfrbp_1 _9275_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2208),
    .D(_0487_),
    .Q_N(_4563_),
    .Q(\addr_bus[14] ));
 sg13g2_dfrbp_1 _9276_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2208),
    .D(_0488_),
    .Q_N(_4562_),
    .Q(\addr_bus[15] ));
 sg13g2_dfrbp_1 _9277_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2204),
    .D(_0489_),
    .Q_N(\z80.tv80s.i_tv80_core.F[0] ),
    .Q(_0245_));
 sg13g2_dfrbp_1 _9278_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2192),
    .D(_0490_),
    .Q_N(\z80.tv80s.i_tv80_core.F[1] ),
    .Q(_0246_));
 sg13g2_dfrbp_1 _9279_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net2206),
    .D(net343),
    .Q_N(\z80.tv80s.i_tv80_core.F[2] ),
    .Q(_0247_));
 sg13g2_dfrbp_1 _9280_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2194),
    .D(_0492_),
    .Q_N(\z80.tv80s.i_tv80_core.F[3] ),
    .Q(_0248_));
 sg13g2_dfrbp_1 _9281_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2204),
    .D(_0493_),
    .Q_N(\z80.tv80s.i_tv80_core.F[4] ),
    .Q(_0249_));
 sg13g2_dfrbp_1 _9282_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2193),
    .D(_0494_),
    .Q_N(\z80.tv80s.i_tv80_core.F[5] ),
    .Q(_0250_));
 sg13g2_dfrbp_1 _9283_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2195),
    .D(_0495_),
    .Q_N(\z80.tv80s.i_tv80_core.F[6] ),
    .Q(_0251_));
 sg13g2_dfrbp_1 _9284_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2192),
    .D(_0496_),
    .Q_N(\z80.tv80s.i_tv80_core.F[7] ),
    .Q(_0252_));
 sg13g2_dfrbp_1 _9285_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2198),
    .D(_0497_),
    .Q_N(_4561_),
    .Q(\z80.tv80s.i_tv80_core.I[0] ));
 sg13g2_dfrbp_1 _9286_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2196),
    .D(net611),
    .Q_N(_4560_),
    .Q(\z80.tv80s.i_tv80_core.I[1] ));
 sg13g2_dfrbp_1 _9287_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2189),
    .D(net605),
    .Q_N(_4559_),
    .Q(\z80.tv80s.i_tv80_core.I[2] ));
 sg13g2_dfrbp_1 _9288_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2189),
    .D(_0500_),
    .Q_N(_4558_),
    .Q(\z80.tv80s.i_tv80_core.I[3] ));
 sg13g2_dfrbp_1 _9289_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2191),
    .D(net616),
    .Q_N(_4557_),
    .Q(\z80.tv80s.i_tv80_core.I[4] ));
 sg13g2_dfrbp_1 _9290_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2196),
    .D(_0502_),
    .Q_N(_4556_),
    .Q(\z80.tv80s.i_tv80_core.I[5] ));
 sg13g2_dfrbp_1 _9291_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2189),
    .D(net609),
    .Q_N(_4555_),
    .Q(\z80.tv80s.i_tv80_core.I[6] ));
 sg13g2_dfrbp_1 _9292_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2191),
    .D(net634),
    .Q_N(_4554_),
    .Q(\z80.tv80s.i_tv80_core.I[7] ));
 sg13g2_dfrbp_1 _9293_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2220),
    .D(net474),
    .Q_N(_0232_),
    .Q(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sg13g2_dfrbp_1 _9294_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2198),
    .D(_0506_),
    .Q_N(_4553_),
    .Q(\z80.tv80s.i_tv80_core.R[7] ));
 sg13g2_dfrbp_1 _9295_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2219),
    .D(_0507_),
    .Q_N(_0028_),
    .Q(\z80.tv80s.i_tv80_core.IntCycle ));
 sg13g2_dfrbp_1 _9296_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2203),
    .D(net506),
    .Q_N(_4552_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _9297_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2203),
    .D(_0509_),
    .Q_N(_4551_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _9298_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2203),
    .D(_0510_),
    .Q_N(_4550_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _9299_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2202),
    .D(_0511_),
    .Q_N(_4549_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _9300_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net2202),
    .D(_0512_),
    .Q_N(_4548_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _9301_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2202),
    .D(_0513_),
    .Q_N(_4547_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _9302_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net2202),
    .D(_0514_),
    .Q_N(_4546_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _9303_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2202),
    .D(_0515_),
    .Q_N(_4545_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _9304_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2193),
    .D(_0516_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[0] ),
    .Q(_0253_));
 sg13g2_dfrbp_1 _9305_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2190),
    .D(_0517_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[1] ),
    .Q(_0254_));
 sg13g2_dfrbp_1 _9306_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2190),
    .D(_0518_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[2] ),
    .Q(_0255_));
 sg13g2_dfrbp_1 _9307_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2191),
    .D(_0519_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[3] ),
    .Q(_0256_));
 sg13g2_dfrbp_1 _9308_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2190),
    .D(_0520_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[4] ),
    .Q(_0257_));
 sg13g2_dfrbp_1 _9309_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2189),
    .D(_0521_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[5] ),
    .Q(_0258_));
 sg13g2_dfrbp_1 _9310_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2189),
    .D(_0522_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[6] ),
    .Q(_0259_));
 sg13g2_dfrbp_1 _9311_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2193),
    .D(_0523_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[7] ),
    .Q(_0260_));
 sg13g2_dfrbp_1 _9312_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2220),
    .D(_0524_),
    .Q_N(_4544_),
    .Q(\z80.tv80s.i_tv80_core.IntE ));
 sg13g2_dfrbp_1 _9313_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2193),
    .D(net231),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[0] ),
    .Q(_0261_));
 sg13g2_dfrbp_1 _9314_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2190),
    .D(net222),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[1] ),
    .Q(_0262_));
 sg13g2_dfrbp_1 _9315_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2190),
    .D(net216),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[2] ),
    .Q(_0263_));
 sg13g2_dfrbp_1 _9316_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2190),
    .D(_0528_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[3] ),
    .Q(_0264_));
 sg13g2_dfrbp_1 _9317_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2190),
    .D(net214),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[4] ),
    .Q(_0265_));
 sg13g2_dfrbp_1 _9318_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2190),
    .D(_0530_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[5] ),
    .Q(_0266_));
 sg13g2_dfrbp_1 _9319_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2189),
    .D(net218),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[6] ),
    .Q(_0267_));
 sg13g2_dfrbp_1 _9320_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2193),
    .D(net212),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[7] ),
    .Q(_0268_));
 sg13g2_dfrbp_1 _9321_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2192),
    .D(_0533_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[0] ),
    .Q(_0269_));
 sg13g2_dfrbp_1 _9322_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2192),
    .D(net202),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[1] ),
    .Q(_0270_));
 sg13g2_dfrbp_1 _9323_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2192),
    .D(net236),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[2] ),
    .Q(_0271_));
 sg13g2_dfrbp_1 _9324_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2193),
    .D(net208),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[3] ),
    .Q(_0272_));
 sg13g2_dfrbp_1 _9325_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2192),
    .D(net224),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[4] ),
    .Q(_0273_));
 sg13g2_dfrbp_1 _9326_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2192),
    .D(net197),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[5] ),
    .Q(_0274_));
 sg13g2_dfrbp_1 _9327_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2194),
    .D(net204),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[6] ),
    .Q(_0275_));
 sg13g2_dfrbp_1 _9328_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2192),
    .D(net199),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[7] ),
    .Q(_0276_));
 sg13g2_dfrbp_1 _9329_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2199),
    .D(_0541_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[0] ),
    .Q(_0277_));
 sg13g2_dfrbp_1 _9330_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2198),
    .D(_0542_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[1] ),
    .Q(_0278_));
 sg13g2_dfrbp_1 _9331_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2198),
    .D(_0543_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[2] ),
    .Q(_0279_));
 sg13g2_dfrbp_1 _9332_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2196),
    .D(_0544_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[3] ),
    .Q(_0280_));
 sg13g2_dfrbp_1 _9333_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2196),
    .D(_0545_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[4] ),
    .Q(_0281_));
 sg13g2_dfrbp_1 _9334_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2199),
    .D(net192),
    .Q_N(\z80.tv80s.i_tv80_core.SP[5] ),
    .Q(_0282_));
 sg13g2_dfrbp_1 _9335_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2199),
    .D(_0547_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[6] ),
    .Q(_0283_));
 sg13g2_dfrbp_1 _9336_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2197),
    .D(_0548_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[7] ),
    .Q(_0284_));
 sg13g2_dfrbp_1 _9337_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2197),
    .D(_0549_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[8] ),
    .Q(_0285_));
 sg13g2_dfrbp_1 _9338_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2196),
    .D(_0550_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[9] ),
    .Q(_0286_));
 sg13g2_dfrbp_1 _9339_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2197),
    .D(_0551_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[10] ),
    .Q(_0287_));
 sg13g2_dfrbp_1 _9340_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2196),
    .D(_0552_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[11] ),
    .Q(_0288_));
 sg13g2_dfrbp_1 _9341_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2196),
    .D(_0553_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[12] ),
    .Q(_0289_));
 sg13g2_dfrbp_1 _9342_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2196),
    .D(_0554_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[13] ),
    .Q(_0290_));
 sg13g2_dfrbp_1 _9343_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2189),
    .D(_0555_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[14] ),
    .Q(_0291_));
 sg13g2_dfrbp_1 _9344_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2197),
    .D(_0556_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[15] ),
    .Q(_0292_));
 sg13g2_dfrbp_1 _9345_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2209),
    .D(net220),
    .Q_N(\z80.tv80s.i_tv80_core.ts[0] ),
    .Q(_0293_));
 sg13g2_dfrbp_1 _9346_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2209),
    .D(net470),
    .Q_N(_0032_),
    .Q(\z80.tv80s.i_tv80_core.ts[1] ));
 sg13g2_dfrbp_1 _9347_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2209),
    .D(net477),
    .Q_N(_0031_),
    .Q(\z80.tv80s.i_tv80_core.ts[2] ));
 sg13g2_dfrbp_1 _9348_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2206),
    .D(_0560_),
    .Q_N(_0023_),
    .Q(\z80.tv80s.i_tv80_core.ts[3] ));
 sg13g2_dfrbp_1 _9349_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2206),
    .D(net546),
    .Q_N(_4543_),
    .Q(\z80.tv80s.i_tv80_core.ts[4] ));
 sg13g2_dfrbp_1 _9350_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2205),
    .D(_0562_),
    .Q_N(_0030_),
    .Q(\z80.tv80s.i_tv80_core.ts[5] ));
 sg13g2_dfrbp_1 _9351_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2205),
    .D(net184),
    .Q_N(_0029_),
    .Q(\z80.tv80s.i_tv80_core.ts[6] ));
 sg13g2_dfrbp_1 _9352_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2217),
    .D(net519),
    .Q_N(_0194_),
    .Q(\z80.tv80s.i_tv80_core.PC[0] ));
 sg13g2_dfrbp_1 _9353_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2217),
    .D(net529),
    .Q_N(_0196_),
    .Q(\z80.tv80s.i_tv80_core.PC[1] ));
 sg13g2_dfrbp_1 _9354_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2217),
    .D(_0566_),
    .Q_N(_0198_),
    .Q(\z80.tv80s.i_tv80_core.PC[2] ));
 sg13g2_dfrbp_1 _9355_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2217),
    .D(_0567_),
    .Q_N(_0200_),
    .Q(\z80.tv80s.i_tv80_core.PC[3] ));
 sg13g2_dfrbp_1 _9356_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2217),
    .D(_0568_),
    .Q_N(_0202_),
    .Q(\z80.tv80s.i_tv80_core.PC[4] ));
 sg13g2_dfrbp_1 _9357_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2217),
    .D(_0569_),
    .Q_N(_4542_),
    .Q(\z80.tv80s.i_tv80_core.PC[5] ));
 sg13g2_dfrbp_1 _9358_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2217),
    .D(_0570_),
    .Q_N(_0205_),
    .Q(\z80.tv80s.i_tv80_core.PC[6] ));
 sg13g2_dfrbp_1 _9359_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2217),
    .D(net629),
    .Q_N(_0207_),
    .Q(\z80.tv80s.i_tv80_core.PC[7] ));
 sg13g2_dfrbp_1 _9360_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2216),
    .D(_0572_),
    .Q_N(_0171_),
    .Q(\z80.tv80s.i_tv80_core.PC[8] ));
 sg13g2_dfrbp_1 _9361_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2216),
    .D(_0573_),
    .Q_N(_0174_),
    .Q(\z80.tv80s.i_tv80_core.PC[9] ));
 sg13g2_dfrbp_1 _9362_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2216),
    .D(_0574_),
    .Q_N(_0177_),
    .Q(\z80.tv80s.i_tv80_core.PC[10] ));
 sg13g2_dfrbp_1 _9363_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2215),
    .D(_0575_),
    .Q_N(_0180_),
    .Q(\z80.tv80s.i_tv80_core.PC[11] ));
 sg13g2_dfrbp_1 _9364_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2215),
    .D(_0576_),
    .Q_N(_0183_),
    .Q(\z80.tv80s.i_tv80_core.PC[12] ));
 sg13g2_dfrbp_1 _9365_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2216),
    .D(_0577_),
    .Q_N(_0186_),
    .Q(\z80.tv80s.i_tv80_core.PC[13] ));
 sg13g2_dfrbp_1 _9366_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2216),
    .D(_0578_),
    .Q_N(_0189_),
    .Q(\z80.tv80s.i_tv80_core.PC[14] ));
 sg13g2_dfrbp_1 _9367_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2216),
    .D(_0579_),
    .Q_N(_0192_),
    .Q(\z80.tv80s.i_tv80_core.PC[15] ));
 sg13g2_dfrbp_1 _9368_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2215),
    .D(net533),
    .Q_N(_0020_),
    .Q(\z80.tv80s.i_tv80_core.Alternate ));
 sg13g2_dfrbp_1 _9369_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2218),
    .D(_0581_),
    .Q_N(_0193_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[0] ));
 sg13g2_dfrbp_1 _9370_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2213),
    .D(_0582_),
    .Q_N(_0195_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[1] ));
 sg13g2_dfrbp_1 _9371_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2213),
    .D(net553),
    .Q_N(_0197_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[2] ));
 sg13g2_dfrbp_1 _9372_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2213),
    .D(_0584_),
    .Q_N(_0199_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sg13g2_dfrbp_1 _9373_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2213),
    .D(_0585_),
    .Q_N(_0201_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sg13g2_dfrbp_1 _9374_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2213),
    .D(net607),
    .Q_N(_0203_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sg13g2_dfrbp_1 _9375_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2214),
    .D(_0587_),
    .Q_N(_0204_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sg13g2_dfrbp_1 _9376_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2213),
    .D(_0588_),
    .Q_N(_0206_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sg13g2_dfrbp_1 _9377_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2215),
    .D(_0589_),
    .Q_N(_0170_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[8] ));
 sg13g2_dfrbp_1 _9378_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2215),
    .D(_0590_),
    .Q_N(_0173_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[9] ));
 sg13g2_dfrbp_1 _9379_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2215),
    .D(_0591_),
    .Q_N(_0176_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[10] ));
 sg13g2_dfrbp_1 _9380_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2215),
    .D(_0592_),
    .Q_N(_0179_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[11] ));
 sg13g2_dfrbp_1 _9381_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2214),
    .D(net514),
    .Q_N(_0182_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[12] ));
 sg13g2_dfrbp_1 _9382_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2215),
    .D(net536),
    .Q_N(_0185_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[13] ));
 sg13g2_dfrbp_1 _9383_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2214),
    .D(_0595_),
    .Q_N(_0188_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[14] ));
 sg13g2_dfrbp_1 _9384_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2214),
    .D(net508),
    .Q_N(_0191_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[15] ));
 sg13g2_dfrbp_1 _9385_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2219),
    .D(net462),
    .Q_N(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .Q(_0294_));
 sg13g2_dfrbp_1 _9386_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2223),
    .D(_0598_),
    .Q_N(_0234_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sg13g2_dfrbp_1 _9387_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2223),
    .D(_0599_),
    .Q_N(_0021_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sg13g2_dfrbp_1 _9388_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2221),
    .D(_0600_),
    .Q_N(_0022_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sg13g2_dfrbp_1 _9389_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2221),
    .D(net555),
    .Q_N(_0025_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ));
 sg13g2_dfrbp_1 _9390_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2222),
    .D(_0602_),
    .Q_N(_0231_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sg13g2_dfrbp_1 _9391_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2221),
    .D(_0603_),
    .Q_N(_0230_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sg13g2_dfrbp_1 _9392_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2222),
    .D(_0604_),
    .Q_N(_0149_),
    .Q(\z80.tv80s.i_tv80_core.IR[0] ));
 sg13g2_dfrbp_1 _9393_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2219),
    .D(_0605_),
    .Q_N(_0024_),
    .Q(\z80.tv80s.i_tv80_core.IR[1] ));
 sg13g2_dfrbp_1 _9394_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2222),
    .D(_0606_),
    .Q_N(_0027_),
    .Q(\z80.tv80s.i_tv80_core.IR[2] ));
 sg13g2_dfrbp_1 _9395_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2219),
    .D(_0607_),
    .Q_N(_0034_),
    .Q(\z80.tv80s.i_tv80_core.IR[3] ));
 sg13g2_dfrbp_1 _9396_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2219),
    .D(_0608_),
    .Q_N(_0026_),
    .Q(\z80.tv80s.i_tv80_core.IR[4] ));
 sg13g2_dfrbp_1 _9397_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2209),
    .D(_0609_),
    .Q_N(_0235_),
    .Q(\z80.tv80s.i_tv80_core.IR[5] ));
 sg13g2_dfrbp_1 _9398_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2224),
    .D(_0610_),
    .Q_N(_4541_),
    .Q(\z80.tv80s.i_tv80_core.IR[6] ));
 sg13g2_dfrbp_1 _9399_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2224),
    .D(_0611_),
    .Q_N(_0233_),
    .Q(\z80.tv80s.i_tv80_core.IR[7] ));
 sg13g2_dfrbp_1 _9400_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2210),
    .D(net334),
    .Q_N(\z80.m1_n ),
    .Q(_0295_));
 sg13g2_dfrbp_1 _9401_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2222),
    .D(_0613_),
    .Q_N(_4540_),
    .Q(\z80.tv80s.i_tv80_core.XY_State[0] ));
 sg13g2_dfrbp_1 _9402_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2205),
    .D(net624),
    .Q_N(_0039_),
    .Q(\z80.tv80s.i_tv80_core.XY_State[1] ));
 sg13g2_dfrbp_1 _9403_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2213),
    .D(net186),
    .Q_N(_4539_),
    .Q(\z80.tv80s.i_tv80_core.XY_Ind ));
 sg13g2_dfrbp_1 _9404_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2218),
    .D(net449),
    .Q_N(_0229_),
    .Q(\z80.tv80s.i_tv80_core.BTR_r ));
 sg13g2_dfrbp_1 _9405_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2213),
    .D(_0617_),
    .Q_N(_0169_),
    .Q(\z80.tv80s.di_reg[0] ));
 sg13g2_dfrbp_1 _9406_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2199),
    .D(_0618_),
    .Q_N(_0172_),
    .Q(\z80.tv80s.di_reg[1] ));
 sg13g2_dfrbp_1 _9407_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2199),
    .D(_0619_),
    .Q_N(_0175_),
    .Q(\z80.tv80s.di_reg[2] ));
 sg13g2_dfrbp_1 _9408_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2200),
    .D(_0620_),
    .Q_N(_0178_),
    .Q(\z80.tv80s.di_reg[3] ));
 sg13g2_dfrbp_1 _9409_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2199),
    .D(_0621_),
    .Q_N(_0181_),
    .Q(\z80.tv80s.di_reg[4] ));
 sg13g2_dfrbp_1 _9410_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2200),
    .D(_0622_),
    .Q_N(_0184_),
    .Q(\z80.tv80s.di_reg[5] ));
 sg13g2_dfrbp_1 _9411_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2199),
    .D(_0623_),
    .Q_N(_0187_),
    .Q(\z80.tv80s.di_reg[6] ));
 sg13g2_dfrbp_1 _9412_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2199),
    .D(_0624_),
    .Q_N(_0190_),
    .Q(\z80.tv80s.di_reg[7] ));
 sg13g2_dfrbp_1 _9413_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2200),
    .D(_0625_),
    .Q_N(_4538_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ));
 sg13g2_dfrbp_1 _9414_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2200),
    .D(_0626_),
    .Q_N(_4537_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ));
 sg13g2_dfrbp_1 _9415_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2194),
    .D(_0627_),
    .Q_N(_4536_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ));
 sg13g2_dfrbp_1 _9416_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2194),
    .D(_0628_),
    .Q_N(_4535_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ));
 sg13g2_dfrbp_1 _9417_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2195),
    .D(_0629_),
    .Q_N(_0228_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ));
 sg13g2_dfrbp_1 _9418_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2222),
    .D(_0630_),
    .Q_N(_4534_),
    .Q(\z80.tv80s.i_tv80_core.No_BTR ));
 sg13g2_dfrbp_1 _9419_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2205),
    .D(_0631_),
    .Q_N(_4533_),
    .Q(\z80.tv80s.i_tv80_core.Arith16_r ));
 sg13g2_dfrbp_1 _9420_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2207),
    .D(net311),
    .Q_N(_4532_),
    .Q(\z80.tv80s.i_tv80_core.Z16_r ));
 sg13g2_dfrbp_1 _9421_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2207),
    .D(_0633_),
    .Q_N(_4531_),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ));
 sg13g2_dfrbp_1 _9422_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2202),
    .D(_0634_),
    .Q_N(_0225_),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ));
 sg13g2_dfrbp_1 _9423_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2207),
    .D(_0635_),
    .Q_N(_0226_),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ));
 sg13g2_dfrbp_1 _9424_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2203),
    .D(_0636_),
    .Q_N(_4530_),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sg13g2_dfrbp_1 _9425_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net2206),
    .D(_0637_),
    .Q_N(_0208_),
    .Q(\z80.tv80s.i_tv80_core.Save_ALU_r ));
 sg13g2_dfrbp_1 _9426_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net60),
    .D(_0638_),
    .Q_N(_0210_),
    .Q(\z80.tv80s.i_tv80_core.BusA[7] ));
 sg13g2_dfrbp_1 _9427_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net24),
    .D(_0639_),
    .Q_N(_0216_),
    .Q(\z80.tv80s.i_tv80_core.BusA[6] ));
 sg13g2_dfrbp_1 _9428_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net22),
    .D(_0640_),
    .Q_N(_0215_),
    .Q(\z80.tv80s.i_tv80_core.BusA[5] ));
 sg13g2_dfrbp_1 _9429_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net19),
    .D(_0641_),
    .Q_N(_0214_),
    .Q(\z80.tv80s.i_tv80_core.BusA[4] ));
 sg13g2_dfrbp_1 _9430_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net93),
    .D(_0642_),
    .Q_N(_0213_),
    .Q(\z80.tv80s.i_tv80_core.BusA[3] ));
 sg13g2_dfrbp_1 _9431_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net88),
    .D(_0643_),
    .Q_N(_0211_),
    .Q(\z80.tv80s.i_tv80_core.BusA[2] ));
 sg13g2_dfrbp_1 _9432_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net67),
    .D(_0644_),
    .Q_N(_0209_),
    .Q(\z80.tv80s.i_tv80_core.BusA[1] ));
 sg13g2_dfrbp_1 _9433_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net63),
    .D(_0645_),
    .Q_N(_0212_),
    .Q(\z80.tv80s.i_tv80_core.BusA[0] ));
 sg13g2_dfrbp_1 _9434_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net61),
    .D(_0646_),
    .Q_N(_0224_),
    .Q(\z80.tv80s.i_tv80_core.BusB[7] ));
 sg13g2_dfrbp_1 _9435_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net23),
    .D(net579),
    .Q_N(_0223_),
    .Q(\z80.tv80s.i_tv80_core.BusB[6] ));
 sg13g2_dfrbp_1 _9436_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net94),
    .D(_0648_),
    .Q_N(_0222_),
    .Q(\z80.tv80s.i_tv80_core.BusB[5] ));
 sg13g2_dfrbp_1 _9437_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net85),
    .D(_0649_),
    .Q_N(_0221_),
    .Q(\z80.tv80s.i_tv80_core.BusB[4] ));
 sg13g2_dfrbp_1 _9438_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net62),
    .D(_0650_),
    .Q_N(_0220_),
    .Q(\z80.tv80s.i_tv80_core.BusB[3] ));
 sg13g2_dfrbp_1 _9439_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net20),
    .D(_0651_),
    .Q_N(_0219_),
    .Q(\z80.tv80s.i_tv80_core.BusB[2] ));
 sg13g2_dfrbp_1 _9440_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net65),
    .D(_0652_),
    .Q_N(_0218_),
    .Q(\z80.tv80s.i_tv80_core.BusB[1] ));
 sg13g2_dfrbp_1 _9441_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net90),
    .D(_0653_),
    .Q_N(_0217_),
    .Q(\z80.tv80s.i_tv80_core.BusB[0] ));
 sg13g2_tiehi _9125__14 (.L_HI(net14));
 sg13g2_tiehi _9124__15 (.L_HI(net15));
 sg13g2_tiehi _9123__16 (.L_HI(net16));
 sg13g2_tiehi _9122__17 (.L_HI(net17));
 sg13g2_tiehi _9121__18 (.L_HI(net18));
 sg13g2_tiehi _9429__19 (.L_HI(net19));
 sg13g2_tiehi _9439__20 (.L_HI(net20));
 sg13g2_tiehi _9075__21 (.L_HI(net21));
 sg13g2_tiehi _9428__22 (.L_HI(net22));
 sg13g2_tiehi _9435__23 (.L_HI(net23));
 sg13g2_tiehi _9427__24 (.L_HI(net24));
 sg13g2_tiehi _9116__25 (.L_HI(net25));
 sg13g2_tiehi _9115__26 (.L_HI(net26));
 sg13g2_tiehi _9114__27 (.L_HI(net27));
 sg13g2_tiehi _9113__28 (.L_HI(net28));
 sg13g2_tiehi _9112__29 (.L_HI(net29));
 sg13g2_tiehi _9111__30 (.L_HI(net30));
 sg13g2_tiehi _9110__31 (.L_HI(net31));
 sg13g2_tiehi _9109__32 (.L_HI(net32));
 sg13g2_tiehi _9108__33 (.L_HI(net33));
 sg13g2_tiehi _9107__34 (.L_HI(net34));
 sg13g2_tiehi _9106__35 (.L_HI(net35));
 sg13g2_tiehi _9105__36 (.L_HI(net36));
 sg13g2_tiehi _9104__37 (.L_HI(net37));
 sg13g2_tiehi _9103__38 (.L_HI(net38));
 sg13g2_tiehi _9102__39 (.L_HI(net39));
 sg13g2_tiehi _9101__40 (.L_HI(net40));
 sg13g2_tiehi _9100__41 (.L_HI(net41));
 sg13g2_tiehi _9099__42 (.L_HI(net42));
 sg13g2_tiehi _9098__43 (.L_HI(net43));
 sg13g2_tiehi _9097__44 (.L_HI(net44));
 sg13g2_tiehi _9096__45 (.L_HI(net45));
 sg13g2_tiehi _9095__46 (.L_HI(net46));
 sg13g2_tiehi _9094__47 (.L_HI(net47));
 sg13g2_tiehi _9093__48 (.L_HI(net48));
 sg13g2_tiehi _9092__49 (.L_HI(net49));
 sg13g2_tiehi _9091__50 (.L_HI(net50));
 sg13g2_tiehi _9090__51 (.L_HI(net51));
 sg13g2_tiehi _9089__52 (.L_HI(net52));
 sg13g2_tiehi _9088__53 (.L_HI(net53));
 sg13g2_tiehi _9087__54 (.L_HI(net54));
 sg13g2_tiehi _9086__55 (.L_HI(net55));
 sg13g2_tiehi _9085__56 (.L_HI(net56));
 sg13g2_tiehi _9074__57 (.L_HI(net57));
 sg13g2_tiehi _9073__58 (.L_HI(net58));
 sg13g2_tiehi _9072__59 (.L_HI(net59));
 sg13g2_tiehi _9426__60 (.L_HI(net60));
 sg13g2_tiehi _9434__61 (.L_HI(net61));
 sg13g2_tiehi _9438__62 (.L_HI(net62));
 sg13g2_tiehi _9433__63 (.L_HI(net63));
 sg13g2_tiehi _9200__64 (.L_HI(net64));
 sg13g2_tiehi _9440__65 (.L_HI(net65));
 sg13g2_tiehi _9215__66 (.L_HI(net66));
 sg13g2_tiehi _9432__67 (.L_HI(net67));
 sg13g2_tiehi _9259__68 (.L_HI(net68));
 sg13g2_tiehi _9258__69 (.L_HI(net69));
 sg13g2_tiehi _9257__70 (.L_HI(net70));
 sg13g2_tiehi _9256__71 (.L_HI(net71));
 sg13g2_tiehi _9255__72 (.L_HI(net72));
 sg13g2_tiehi _9254__73 (.L_HI(net73));
 sg13g2_tiehi _9253__74 (.L_HI(net74));
 sg13g2_tiehi _9252__75 (.L_HI(net75));
 sg13g2_tiehi _9251__76 (.L_HI(net76));
 sg13g2_tiehi _9250__77 (.L_HI(net77));
 sg13g2_tiehi _9249__78 (.L_HI(net78));
 sg13g2_tiehi _9248__79 (.L_HI(net79));
 sg13g2_tiehi _9247__80 (.L_HI(net80));
 sg13g2_tiehi _9246__81 (.L_HI(net81));
 sg13g2_tiehi _9245__82 (.L_HI(net82));
 sg13g2_tiehi _9244__83 (.L_HI(net83));
 sg13g2_tiehi _9243__84 (.L_HI(net84));
 sg13g2_tiehi _9437__85 (.L_HI(net85));
 sg13g2_tiehi _9242__86 (.L_HI(net86));
 sg13g2_tiehi _9241__87 (.L_HI(net87));
 sg13g2_tiehi _9431__88 (.L_HI(net88));
 sg13g2_tiehi _9240__89 (.L_HI(net89));
 sg13g2_tiehi _9441__90 (.L_HI(net90));
 sg13g2_tiehi _9239__91 (.L_HI(net91));
 sg13g2_tiehi _9238__92 (.L_HI(net92));
 sg13g2_tiehi _9430__93 (.L_HI(net93));
 sg13g2_tiehi _9436__94 (.L_HI(net94));
 sg13g2_tiehi _9225__95 (.L_HI(net95));
 sg13g2_tiehi _9224__96 (.L_HI(net96));
 sg13g2_tiehi _9223__97 (.L_HI(net97));
 sg13g2_tiehi _9222__98 (.L_HI(net98));
 sg13g2_tiehi _9221__99 (.L_HI(net99));
 sg13g2_tiehi _9220__100 (.L_HI(net100));
 sg13g2_tiehi _9219__101 (.L_HI(net101));
 sg13g2_tiehi _9218__102 (.L_HI(net102));
 sg13g2_tiehi _9214__103 (.L_HI(net103));
 sg13g2_tiehi _9213__104 (.L_HI(net104));
 sg13g2_tiehi _9212__105 (.L_HI(net105));
 sg13g2_tiehi _9211__106 (.L_HI(net106));
 sg13g2_tiehi _9210__107 (.L_HI(net107));
 sg13g2_tiehi _9209__108 (.L_HI(net108));
 sg13g2_tiehi _9208__109 (.L_HI(net109));
 sg13g2_tiehi _9199__110 (.L_HI(net110));
 sg13g2_tiehi _9198__111 (.L_HI(net111));
 sg13g2_tiehi _9197__112 (.L_HI(net112));
 sg13g2_tiehi _9196__113 (.L_HI(net113));
 sg13g2_tiehi _9195__114 (.L_HI(net114));
 sg13g2_tiehi _9194__115 (.L_HI(net115));
 sg13g2_tiehi _9193__116 (.L_HI(net116));
 sg13g2_tiehi _9192__117 (.L_HI(net117));
 sg13g2_tiehi _9191__118 (.L_HI(net118));
 sg13g2_tiehi _9190__119 (.L_HI(net119));
 sg13g2_tiehi _9189__120 (.L_HI(net120));
 sg13g2_tiehi _9188__121 (.L_HI(net121));
 sg13g2_tiehi _9187__122 (.L_HI(net122));
 sg13g2_tiehi _9186__123 (.L_HI(net123));
 sg13g2_tiehi _9185__124 (.L_HI(net124));
 sg13g2_tiehi _9184__125 (.L_HI(net125));
 sg13g2_tiehi _9183__126 (.L_HI(net126));
 sg13g2_tiehi _9182__127 (.L_HI(net127));
 sg13g2_tiehi _9181__128 (.L_HI(net128));
 sg13g2_tiehi _9180__129 (.L_HI(net129));
 sg13g2_tiehi _9179__130 (.L_HI(net130));
 sg13g2_tiehi _9178__131 (.L_HI(net131));
 sg13g2_tiehi _9177__132 (.L_HI(net132));
 sg13g2_tiehi _9176__133 (.L_HI(net133));
 sg13g2_tiehi _9175__134 (.L_HI(net134));
 sg13g2_tiehi _9174__135 (.L_HI(net135));
 sg13g2_tiehi _9173__136 (.L_HI(net136));
 sg13g2_tiehi _9172__137 (.L_HI(net137));
 sg13g2_tiehi _9171__138 (.L_HI(net138));
 sg13g2_tiehi _9170__139 (.L_HI(net139));
 sg13g2_tiehi _9169__140 (.L_HI(net140));
 sg13g2_tiehi _9168__141 (.L_HI(net141));
 sg13g2_tiehi _9167__142 (.L_HI(net142));
 sg13g2_tiehi _9166__143 (.L_HI(net143));
 sg13g2_tiehi _9165__144 (.L_HI(net144));
 sg13g2_tiehi _9164__145 (.L_HI(net145));
 sg13g2_tiehi _9163__146 (.L_HI(net146));
 sg13g2_tiehi _9162__147 (.L_HI(net147));
 sg13g2_tiehi _9161__148 (.L_HI(net148));
 sg13g2_tiehi _9160__149 (.L_HI(net149));
 sg13g2_tiehi _9159__150 (.L_HI(net150));
 sg13g2_tiehi _9158__151 (.L_HI(net151));
 sg13g2_tiehi _9157__152 (.L_HI(net152));
 sg13g2_tiehi _9156__153 (.L_HI(net153));
 sg13g2_tiehi _9155__154 (.L_HI(net154));
 sg13g2_tiehi _9154__155 (.L_HI(net155));
 sg13g2_tiehi _9153__156 (.L_HI(net156));
 sg13g2_tiehi _9152__157 (.L_HI(net157));
 sg13g2_tiehi _9151__158 (.L_HI(net158));
 sg13g2_tiehi _9150__159 (.L_HI(net159));
 sg13g2_tiehi _9149__160 (.L_HI(net160));
 sg13g2_tiehi _9148__161 (.L_HI(net161));
 sg13g2_tiehi _9147__162 (.L_HI(net162));
 sg13g2_tiehi _9146__163 (.L_HI(net163));
 sg13g2_tiehi _9145__164 (.L_HI(net164));
 sg13g2_tiehi _9144__165 (.L_HI(net165));
 sg13g2_tiehi _9143__166 (.L_HI(net166));
 sg13g2_tiehi _9142__167 (.L_HI(net167));
 sg13g2_tiehi _9141__168 (.L_HI(net168));
 sg13g2_tiehi _9140__169 (.L_HI(net169));
 sg13g2_tiehi _9139__170 (.L_HI(net170));
 sg13g2_tiehi _9138__171 (.L_HI(net171));
 sg13g2_tiehi _9137__172 (.L_HI(net172));
 sg13g2_tiehi _9136__173 (.L_HI(net173));
 sg13g2_tiehi _9135__174 (.L_HI(net174));
 sg13g2_tiehi _9134__175 (.L_HI(net175));
 sg13g2_tiehi _9133__176 (.L_HI(net176));
 sg13g2_tiehi _9132__177 (.L_HI(net177));
 sg13g2_tiehi _9131__178 (.L_HI(net178));
 sg13g2_tiehi _9130__179 (.L_HI(net179));
 sg13g2_tiehi _9129__180 (.L_HI(net180));
 sg13g2_tiehi _9128__181 (.L_HI(net181));
 sg13g2_tiehi _9127__182 (.L_HI(net182));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _9612_ (.A(net1766),
    .X(uio_oe[0]));
 sg13g2_buf_1 _9613_ (.A(net1766),
    .X(uio_oe[1]));
 sg13g2_buf_1 _9614_ (.A(net1766),
    .X(uio_oe[2]));
 sg13g2_buf_1 _9615_ (.A(net1766),
    .X(uio_oe[3]));
 sg13g2_buf_1 _9616_ (.A(net1766),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9617_ (.A(net1766),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9618_ (.A(net1766),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9619_ (.A(net1766),
    .X(uio_oe[7]));
 sg13g2_buf_4 fanout1679 (.X(net1679),
    .A(_1135_));
 sg13g2_buf_4 fanout1680 (.X(net1680),
    .A(_3105_));
 sg13g2_buf_2 fanout1681 (.A(net1683),
    .X(net1681));
 sg13g2_buf_1 fanout1682 (.A(net1683),
    .X(net1682));
 sg13g2_buf_4 fanout1683 (.X(net1683),
    .A(_2636_));
 sg13g2_buf_2 fanout1684 (.A(_2635_),
    .X(net1684));
 sg13g2_buf_4 fanout1685 (.X(net1685),
    .A(_2635_));
 sg13g2_buf_4 fanout1686 (.X(net1686),
    .A(_2634_));
 sg13g2_buf_8 fanout1687 (.A(_1131_),
    .X(net1687));
 sg13g2_buf_2 fanout1688 (.A(net1694),
    .X(net1688));
 sg13g2_buf_4 fanout1689 (.X(net1689),
    .A(net1694));
 sg13g2_buf_2 fanout1690 (.A(net1691),
    .X(net1690));
 sg13g2_buf_1 fanout1691 (.A(net1692),
    .X(net1691));
 sg13g2_buf_1 fanout1692 (.A(net1693),
    .X(net1692));
 sg13g2_buf_2 fanout1693 (.A(net1694),
    .X(net1693));
 sg13g2_buf_4 fanout1694 (.X(net1694),
    .A(_1130_));
 sg13g2_buf_2 fanout1695 (.A(net1698),
    .X(net1695));
 sg13g2_buf_2 fanout1696 (.A(net1698),
    .X(net1696));
 sg13g2_buf_1 fanout1697 (.A(net1698),
    .X(net1697));
 sg13g2_buf_2 fanout1698 (.A(_3659_),
    .X(net1698));
 sg13g2_buf_2 fanout1699 (.A(net1700),
    .X(net1699));
 sg13g2_buf_2 fanout1700 (.A(_2615_),
    .X(net1700));
 sg13g2_buf_2 fanout1701 (.A(net1702),
    .X(net1701));
 sg13g2_buf_2 fanout1702 (.A(_1335_),
    .X(net1702));
 sg13g2_buf_2 fanout1703 (.A(_3704_),
    .X(net1703));
 sg13g2_buf_2 fanout1704 (.A(net1705),
    .X(net1704));
 sg13g2_buf_4 fanout1705 (.X(net1705),
    .A(_2614_));
 sg13g2_buf_2 fanout1706 (.A(net1707),
    .X(net1706));
 sg13g2_buf_2 fanout1707 (.A(_2613_),
    .X(net1707));
 sg13g2_buf_2 fanout1708 (.A(net1709),
    .X(net1708));
 sg13g2_buf_4 fanout1709 (.X(net1709),
    .A(_2610_));
 sg13g2_buf_2 fanout1710 (.A(net1713),
    .X(net1710));
 sg13g2_buf_2 fanout1711 (.A(net1713),
    .X(net1711));
 sg13g2_buf_2 fanout1712 (.A(net1713),
    .X(net1712));
 sg13g2_buf_2 fanout1713 (.A(_2607_),
    .X(net1713));
 sg13g2_buf_2 fanout1714 (.A(net1715),
    .X(net1714));
 sg13g2_buf_2 fanout1715 (.A(net1716),
    .X(net1715));
 sg13g2_buf_2 fanout1716 (.A(_3703_),
    .X(net1716));
 sg13g2_buf_2 fanout1717 (.A(net1718),
    .X(net1717));
 sg13g2_buf_1 fanout1718 (.A(net1719),
    .X(net1718));
 sg13g2_buf_1 fanout1719 (.A(net1720),
    .X(net1719));
 sg13g2_buf_1 fanout1720 (.A(_2584_),
    .X(net1720));
 sg13g2_buf_2 fanout1721 (.A(net1727),
    .X(net1721));
 sg13g2_buf_2 fanout1722 (.A(net1723),
    .X(net1722));
 sg13g2_buf_2 fanout1723 (.A(net1727),
    .X(net1723));
 sg13g2_buf_2 fanout1724 (.A(net1726),
    .X(net1724));
 sg13g2_buf_1 fanout1725 (.A(net1727),
    .X(net1725));
 sg13g2_buf_2 fanout1726 (.A(net1727),
    .X(net1726));
 sg13g2_buf_2 fanout1727 (.A(_2584_),
    .X(net1727));
 sg13g2_buf_4 fanout1728 (.X(net1728),
    .A(_2467_));
 sg13g2_buf_4 fanout1729 (.X(net1729),
    .A(_2462_));
 sg13g2_buf_4 fanout1730 (.X(net1730),
    .A(net1731));
 sg13g2_buf_4 fanout1731 (.X(net1731),
    .A(_4383_));
 sg13g2_buf_4 fanout1732 (.X(net1732),
    .A(net1733));
 sg13g2_buf_4 fanout1733 (.X(net1733),
    .A(_4145_));
 sg13g2_buf_4 fanout1734 (.X(net1734),
    .A(net1735));
 sg13g2_buf_4 fanout1735 (.X(net1735),
    .A(_1862_));
 sg13g2_buf_4 fanout1736 (.X(net1736),
    .A(_1861_));
 sg13g2_buf_4 fanout1737 (.X(net1737),
    .A(_1861_));
 sg13g2_buf_4 fanout1738 (.X(net1738),
    .A(net1739));
 sg13g2_buf_4 fanout1739 (.X(net1739),
    .A(_1860_));
 sg13g2_buf_4 fanout1740 (.X(net1740),
    .A(net1741));
 sg13g2_buf_4 fanout1741 (.X(net1741),
    .A(_1858_));
 sg13g2_buf_4 fanout1742 (.X(net1742),
    .A(net1743));
 sg13g2_buf_4 fanout1743 (.X(net1743),
    .A(_1855_));
 sg13g2_buf_4 fanout1744 (.X(net1744),
    .A(net1745));
 sg13g2_buf_4 fanout1745 (.X(net1745),
    .A(_1851_));
 sg13g2_buf_4 fanout1746 (.X(net1746),
    .A(net1747));
 sg13g2_buf_4 fanout1747 (.X(net1747),
    .A(_1849_));
 sg13g2_buf_4 fanout1748 (.X(net1748),
    .A(_1749_));
 sg13g2_buf_4 fanout1749 (.X(net1749),
    .A(_1749_));
 sg13g2_buf_2 fanout1750 (.A(net1751),
    .X(net1750));
 sg13g2_buf_2 fanout1751 (.A(net1752),
    .X(net1751));
 sg13g2_buf_2 fanout1752 (.A(_1518_),
    .X(net1752));
 sg13g2_buf_2 fanout1753 (.A(net1754),
    .X(net1753));
 sg13g2_buf_4 fanout1754 (.X(net1754),
    .A(_1517_));
 sg13g2_buf_2 fanout1755 (.A(_3951_),
    .X(net1755));
 sg13g2_buf_2 fanout1756 (.A(net1759),
    .X(net1756));
 sg13g2_buf_2 fanout1757 (.A(net1759),
    .X(net1757));
 sg13g2_buf_2 fanout1758 (.A(net1759),
    .X(net1758));
 sg13g2_buf_2 fanout1759 (.A(_2628_),
    .X(net1759));
 sg13g2_buf_2 fanout1760 (.A(net1763),
    .X(net1760));
 sg13g2_buf_1 fanout1761 (.A(net1763),
    .X(net1761));
 sg13g2_buf_2 fanout1762 (.A(net1763),
    .X(net1762));
 sg13g2_buf_2 fanout1763 (.A(_2619_),
    .X(net1763));
 sg13g2_buf_4 fanout1764 (.X(net1764),
    .A(_1734_));
 sg13g2_buf_2 fanout1765 (.A(_1733_),
    .X(net1765));
 sg13g2_buf_2 fanout1766 (.A(doe),
    .X(net1766));
 sg13g2_buf_2 fanout1767 (.A(net1768),
    .X(net1767));
 sg13g2_buf_2 fanout1768 (.A(_4016_),
    .X(net1768));
 sg13g2_buf_2 fanout1769 (.A(net1770),
    .X(net1769));
 sg13g2_buf_2 fanout1770 (.A(_3524_),
    .X(net1770));
 sg13g2_buf_2 fanout1771 (.A(_3422_),
    .X(net1771));
 sg13g2_buf_1 fanout1772 (.A(_3422_),
    .X(net1772));
 sg13g2_buf_2 fanout1773 (.A(net1775),
    .X(net1773));
 sg13g2_buf_2 fanout1774 (.A(net1775),
    .X(net1774));
 sg13g2_buf_2 fanout1775 (.A(_3421_),
    .X(net1775));
 sg13g2_buf_2 fanout1776 (.A(net1777),
    .X(net1776));
 sg13g2_buf_2 fanout1777 (.A(_3403_),
    .X(net1777));
 sg13g2_buf_2 fanout1778 (.A(net1780),
    .X(net1778));
 sg13g2_buf_2 fanout1779 (.A(net1780),
    .X(net1779));
 sg13g2_buf_2 fanout1780 (.A(_3403_),
    .X(net1780));
 sg13g2_buf_2 fanout1781 (.A(net1783),
    .X(net1781));
 sg13g2_buf_2 fanout1782 (.A(net1783),
    .X(net1782));
 sg13g2_buf_2 fanout1783 (.A(net1784),
    .X(net1783));
 sg13g2_buf_4 fanout1784 (.X(net1784),
    .A(_2602_));
 sg13g2_buf_4 fanout1785 (.X(net1785),
    .A(net1786));
 sg13g2_buf_4 fanout1786 (.X(net1786),
    .A(_1960_));
 sg13g2_buf_2 fanout1787 (.A(_1775_),
    .X(net1787));
 sg13g2_buf_2 fanout1788 (.A(_1775_),
    .X(net1788));
 sg13g2_buf_2 fanout1789 (.A(_1772_),
    .X(net1789));
 sg13g2_buf_4 fanout1790 (.X(net1790),
    .A(_1771_));
 sg13g2_buf_2 fanout1791 (.A(_1771_),
    .X(net1791));
 sg13g2_buf_2 fanout1792 (.A(net1793),
    .X(net1792));
 sg13g2_buf_1 fanout1793 (.A(_3935_),
    .X(net1793));
 sg13g2_buf_2 fanout1794 (.A(_3935_),
    .X(net1794));
 sg13g2_buf_2 fanout1795 (.A(net1796),
    .X(net1795));
 sg13g2_buf_2 fanout1796 (.A(_3081_),
    .X(net1796));
 sg13g2_buf_4 fanout1797 (.X(net1797),
    .A(net1801));
 sg13g2_buf_2 fanout1798 (.A(net1801),
    .X(net1798));
 sg13g2_buf_4 fanout1799 (.X(net1799),
    .A(net1801));
 sg13g2_buf_2 fanout1800 (.A(net1801),
    .X(net1800));
 sg13g2_buf_2 fanout1801 (.A(_1962_),
    .X(net1801));
 sg13g2_buf_4 fanout1802 (.X(net1802),
    .A(net1803));
 sg13g2_buf_4 fanout1803 (.X(net1803),
    .A(net1806));
 sg13g2_buf_4 fanout1804 (.X(net1804),
    .A(net1806));
 sg13g2_buf_4 fanout1805 (.X(net1805),
    .A(net1806));
 sg13g2_buf_2 fanout1806 (.A(_1961_),
    .X(net1806));
 sg13g2_buf_4 fanout1807 (.X(net1807),
    .A(net1808));
 sg13g2_buf_4 fanout1808 (.X(net1808),
    .A(net1811));
 sg13g2_buf_4 fanout1809 (.X(net1809),
    .A(net1810));
 sg13g2_buf_4 fanout1810 (.X(net1810),
    .A(net1811));
 sg13g2_buf_2 fanout1811 (.A(_1957_),
    .X(net1811));
 sg13g2_buf_4 fanout1812 (.X(net1812),
    .A(_1956_));
 sg13g2_buf_4 fanout1813 (.X(net1813),
    .A(net1814));
 sg13g2_buf_4 fanout1814 (.X(net1814),
    .A(_1956_));
 sg13g2_buf_2 fanout1815 (.A(net1816),
    .X(net1815));
 sg13g2_buf_2 fanout1816 (.A(net1817),
    .X(net1816));
 sg13g2_buf_2 fanout1817 (.A(_1848_),
    .X(net1817));
 sg13g2_buf_4 fanout1818 (.X(net1818),
    .A(_3095_));
 sg13g2_buf_2 fanout1819 (.A(_3095_),
    .X(net1819));
 sg13g2_buf_2 fanout1820 (.A(_3092_),
    .X(net1820));
 sg13g2_buf_1 fanout1821 (.A(_3092_),
    .X(net1821));
 sg13g2_buf_4 fanout1822 (.X(net1822),
    .A(net1823));
 sg13g2_buf_4 fanout1823 (.X(net1823),
    .A(_1847_));
 sg13g2_buf_4 fanout1824 (.X(net1824),
    .A(_1727_));
 sg13g2_buf_2 fanout1825 (.A(net1826),
    .X(net1825));
 sg13g2_buf_2 fanout1826 (.A(net1827),
    .X(net1826));
 sg13g2_buf_4 fanout1827 (.X(net1827),
    .A(_1720_));
 sg13g2_buf_2 fanout1828 (.A(net1830),
    .X(net1828));
 sg13g2_buf_2 fanout1829 (.A(net1830),
    .X(net1829));
 sg13g2_buf_4 fanout1830 (.X(net1830),
    .A(_1718_));
 sg13g2_buf_2 fanout1831 (.A(net1834),
    .X(net1831));
 sg13g2_buf_2 fanout1832 (.A(net1834),
    .X(net1832));
 sg13g2_buf_2 fanout1833 (.A(net1834),
    .X(net1833));
 sg13g2_buf_2 fanout1834 (.A(_1718_),
    .X(net1834));
 sg13g2_buf_2 fanout1835 (.A(net1836),
    .X(net1835));
 sg13g2_buf_2 fanout1836 (.A(_1536_),
    .X(net1836));
 sg13g2_buf_2 fanout1837 (.A(_1536_),
    .X(net1837));
 sg13g2_buf_2 fanout1838 (.A(net1842),
    .X(net1838));
 sg13g2_buf_2 fanout1839 (.A(net1842),
    .X(net1839));
 sg13g2_buf_2 fanout1840 (.A(net1842),
    .X(net1840));
 sg13g2_buf_2 fanout1841 (.A(net1842),
    .X(net1841));
 sg13g2_buf_1 fanout1842 (.A(_1536_),
    .X(net1842));
 sg13g2_buf_4 fanout1843 (.X(net1843),
    .A(_1267_));
 sg13g2_buf_1 fanout1844 (.A(_1267_),
    .X(net1844));
 sg13g2_buf_2 fanout1845 (.A(_3807_),
    .X(net1845));
 sg13g2_buf_1 fanout1846 (.A(_3807_),
    .X(net1846));
 sg13g2_buf_2 fanout1847 (.A(net1848),
    .X(net1847));
 sg13g2_buf_2 fanout1848 (.A(_3328_),
    .X(net1848));
 sg13g2_buf_2 fanout1849 (.A(net1850),
    .X(net1849));
 sg13g2_buf_2 fanout1850 (.A(_3547_),
    .X(net1850));
 sg13g2_buf_4 fanout1851 (.X(net1851),
    .A(_3432_));
 sg13g2_buf_2 fanout1852 (.A(_3273_),
    .X(net1852));
 sg13g2_buf_2 fanout1853 (.A(_3270_),
    .X(net1853));
 sg13g2_buf_2 fanout1854 (.A(_4091_),
    .X(net1854));
 sg13g2_buf_2 fanout1855 (.A(_3955_),
    .X(net1855));
 sg13g2_buf_2 fanout1856 (.A(net1857),
    .X(net1856));
 sg13g2_buf_2 fanout1857 (.A(_3272_),
    .X(net1857));
 sg13g2_buf_2 fanout1858 (.A(net1859),
    .X(net1858));
 sg13g2_buf_2 fanout1859 (.A(net1861),
    .X(net1859));
 sg13g2_buf_2 fanout1860 (.A(net1861),
    .X(net1860));
 sg13g2_buf_2 fanout1861 (.A(_3108_),
    .X(net1861));
 sg13g2_buf_2 fanout1862 (.A(_1463_),
    .X(net1862));
 sg13g2_buf_2 fanout1863 (.A(_1804_),
    .X(net1863));
 sg13g2_buf_4 fanout1864 (.X(net1864),
    .A(_1047_));
 sg13g2_buf_2 fanout1865 (.A(net1868),
    .X(net1865));
 sg13g2_buf_1 fanout1866 (.A(net1868),
    .X(net1866));
 sg13g2_buf_2 fanout1867 (.A(net1868),
    .X(net1867));
 sg13g2_buf_2 fanout1868 (.A(_2605_),
    .X(net1868));
 sg13g2_buf_2 fanout1869 (.A(net1871),
    .X(net1869));
 sg13g2_buf_1 fanout1870 (.A(net1871),
    .X(net1870));
 sg13g2_buf_1 fanout1871 (.A(net1872),
    .X(net1871));
 sg13g2_buf_2 fanout1872 (.A(_2605_),
    .X(net1872));
 sg13g2_buf_2 fanout1873 (.A(_1788_),
    .X(net1873));
 sg13g2_buf_2 fanout1874 (.A(_1779_),
    .X(net1874));
 sg13g2_buf_4 fanout1875 (.X(net1875),
    .A(net1876));
 sg13g2_buf_2 fanout1876 (.A(_1046_),
    .X(net1876));
 sg13g2_buf_4 fanout1877 (.X(net1877),
    .A(_1040_));
 sg13g2_buf_1 fanout1878 (.A(_1040_),
    .X(net1878));
 sg13g2_buf_4 fanout1879 (.X(net1879),
    .A(net1880));
 sg13g2_buf_2 fanout1880 (.A(_1033_),
    .X(net1880));
 sg13g2_buf_4 fanout1881 (.X(net1881),
    .A(_1020_));
 sg13g2_buf_4 fanout1882 (.X(net1882),
    .A(_1013_));
 sg13g2_buf_4 fanout1883 (.X(net1883),
    .A(_1009_));
 sg13g2_buf_4 fanout1884 (.X(net1884),
    .A(_1005_));
 sg13g2_buf_4 fanout1885 (.X(net1885),
    .A(_0955_));
 sg13g2_buf_4 fanout1886 (.X(net1886),
    .A(net1887));
 sg13g2_buf_4 fanout1887 (.X(net1887),
    .A(_0954_));
 sg13g2_buf_4 fanout1888 (.X(net1888),
    .A(_0918_));
 sg13g2_buf_4 fanout1889 (.X(net1889),
    .A(_0886_));
 sg13g2_buf_4 fanout1890 (.X(net1890),
    .A(_0866_));
 sg13g2_buf_2 fanout1891 (.A(net1893),
    .X(net1891));
 sg13g2_buf_4 fanout1892 (.X(net1892),
    .A(net1893));
 sg13g2_buf_1 fanout1893 (.A(_0846_),
    .X(net1893));
 sg13g2_buf_2 fanout1894 (.A(_0824_),
    .X(net1894));
 sg13g2_buf_2 fanout1895 (.A(net1896),
    .X(net1895));
 sg13g2_buf_2 fanout1896 (.A(net1904),
    .X(net1896));
 sg13g2_buf_4 fanout1897 (.X(net1897),
    .A(net1899));
 sg13g2_buf_2 fanout1898 (.A(net1899),
    .X(net1898));
 sg13g2_buf_2 fanout1899 (.A(net1904),
    .X(net1899));
 sg13g2_buf_4 fanout1900 (.X(net1900),
    .A(net1904));
 sg13g2_buf_2 fanout1901 (.A(net1904),
    .X(net1901));
 sg13g2_buf_2 fanout1902 (.A(net1903),
    .X(net1902));
 sg13g2_buf_2 fanout1903 (.A(net1904),
    .X(net1903));
 sg13g2_buf_2 fanout1904 (.A(_0809_),
    .X(net1904));
 sg13g2_buf_2 fanout1905 (.A(net1908),
    .X(net1905));
 sg13g2_buf_2 fanout1906 (.A(net1907),
    .X(net1906));
 sg13g2_buf_2 fanout1907 (.A(net1908),
    .X(net1907));
 sg13g2_buf_4 fanout1908 (.X(net1908),
    .A(_0808_));
 sg13g2_buf_2 fanout1909 (.A(net1910),
    .X(net1909));
 sg13g2_buf_2 fanout1910 (.A(net1911),
    .X(net1910));
 sg13g2_buf_4 fanout1911 (.X(net1911),
    .A(net1914));
 sg13g2_buf_2 fanout1912 (.A(net1913),
    .X(net1912));
 sg13g2_buf_4 fanout1913 (.X(net1913),
    .A(net1914));
 sg13g2_buf_2 fanout1914 (.A(_0808_),
    .X(net1914));
 sg13g2_buf_2 fanout1915 (.A(net1917),
    .X(net1915));
 sg13g2_buf_1 fanout1916 (.A(net1917),
    .X(net1916));
 sg13g2_buf_2 fanout1917 (.A(net1918),
    .X(net1917));
 sg13g2_buf_2 fanout1918 (.A(_3934_),
    .X(net1918));
 sg13g2_buf_2 fanout1919 (.A(_3933_),
    .X(net1919));
 sg13g2_buf_2 fanout1920 (.A(net1921),
    .X(net1920));
 sg13g2_buf_4 fanout1921 (.X(net1921),
    .A(_2606_));
 sg13g2_buf_4 fanout1922 (.X(net1922),
    .A(_1312_));
 sg13g2_buf_2 fanout1923 (.A(net1924),
    .X(net1923));
 sg13g2_buf_2 fanout1924 (.A(net1927),
    .X(net1924));
 sg13g2_buf_2 fanout1925 (.A(net1926),
    .X(net1925));
 sg13g2_buf_2 fanout1926 (.A(net1927),
    .X(net1926));
 sg13g2_buf_2 fanout1927 (.A(_1139_),
    .X(net1927));
 sg13g2_buf_4 fanout1928 (.X(net1928),
    .A(_0963_));
 sg13g2_buf_4 fanout1929 (.X(net1929),
    .A(_0938_));
 sg13g2_buf_2 fanout1930 (.A(_0938_),
    .X(net1930));
 sg13g2_buf_4 fanout1931 (.X(net1931),
    .A(net1932));
 sg13g2_buf_4 fanout1932 (.X(net1932),
    .A(_0905_));
 sg13g2_buf_4 fanout1933 (.X(net1933),
    .A(net1934));
 sg13g2_buf_4 fanout1934 (.X(net1934),
    .A(_0898_));
 sg13g2_buf_4 fanout1935 (.X(net1935),
    .A(net1936));
 sg13g2_buf_4 fanout1936 (.X(net1936),
    .A(_0897_));
 sg13g2_buf_4 fanout1937 (.X(net1937),
    .A(net1938));
 sg13g2_buf_2 fanout1938 (.A(net1939),
    .X(net1938));
 sg13g2_buf_4 fanout1939 (.X(net1939),
    .A(_0893_));
 sg13g2_buf_2 fanout1940 (.A(_0892_),
    .X(net1940));
 sg13g2_buf_2 fanout1941 (.A(_0892_),
    .X(net1941));
 sg13g2_buf_4 fanout1942 (.X(net1942),
    .A(_0869_));
 sg13g2_buf_4 fanout1943 (.X(net1943),
    .A(_0869_));
 sg13g2_buf_4 fanout1944 (.X(net1944),
    .A(net1945));
 sg13g2_buf_4 fanout1945 (.X(net1945),
    .A(_0867_));
 sg13g2_buf_2 fanout1946 (.A(_0862_),
    .X(net1946));
 sg13g2_buf_2 fanout1947 (.A(_0862_),
    .X(net1947));
 sg13g2_buf_4 fanout1948 (.X(net1948),
    .A(_0856_));
 sg13g2_buf_4 fanout1949 (.X(net1949),
    .A(_0848_));
 sg13g2_buf_2 fanout1950 (.A(_0848_),
    .X(net1950));
 sg13g2_buf_4 fanout1951 (.X(net1951),
    .A(_0847_));
 sg13g2_buf_2 fanout1952 (.A(net1953),
    .X(net1952));
 sg13g2_buf_2 fanout1953 (.A(net1954),
    .X(net1953));
 sg13g2_buf_4 fanout1954 (.X(net1954),
    .A(_0845_));
 sg13g2_buf_4 fanout1955 (.X(net1955),
    .A(net1956));
 sg13g2_buf_4 fanout1956 (.X(net1956),
    .A(_0839_));
 sg13g2_buf_4 fanout1957 (.X(net1957),
    .A(_0829_));
 sg13g2_buf_4 fanout1958 (.X(net1958),
    .A(_0829_));
 sg13g2_buf_2 fanout1959 (.A(net1960),
    .X(net1959));
 sg13g2_buf_2 fanout1960 (.A(net1973),
    .X(net1960));
 sg13g2_buf_2 fanout1961 (.A(net1962),
    .X(net1961));
 sg13g2_buf_2 fanout1962 (.A(net1964),
    .X(net1962));
 sg13g2_buf_2 fanout1963 (.A(net1964),
    .X(net1963));
 sg13g2_buf_2 fanout1964 (.A(net1973),
    .X(net1964));
 sg13g2_buf_2 fanout1965 (.A(net1966),
    .X(net1965));
 sg13g2_buf_2 fanout1966 (.A(net1969),
    .X(net1966));
 sg13g2_buf_2 fanout1967 (.A(net1969),
    .X(net1967));
 sg13g2_buf_1 fanout1968 (.A(net1969),
    .X(net1968));
 sg13g2_buf_2 fanout1969 (.A(net1973),
    .X(net1969));
 sg13g2_buf_2 fanout1970 (.A(net1972),
    .X(net1970));
 sg13g2_buf_1 fanout1971 (.A(net1972),
    .X(net1971));
 sg13g2_buf_2 fanout1972 (.A(net1973),
    .X(net1972));
 sg13g2_buf_2 fanout1973 (.A(_0823_),
    .X(net1973));
 sg13g2_buf_2 fanout1974 (.A(net1976),
    .X(net1974));
 sg13g2_buf_4 fanout1975 (.X(net1975),
    .A(net1976));
 sg13g2_buf_2 fanout1976 (.A(net1982),
    .X(net1976));
 sg13g2_buf_2 fanout1977 (.A(net1979),
    .X(net1977));
 sg13g2_buf_1 fanout1978 (.A(net1979),
    .X(net1978));
 sg13g2_buf_2 fanout1979 (.A(net1982),
    .X(net1979));
 sg13g2_buf_4 fanout1980 (.X(net1980),
    .A(net1982));
 sg13g2_buf_2 fanout1981 (.A(net1982),
    .X(net1981));
 sg13g2_buf_2 fanout1982 (.A(_0823_),
    .X(net1982));
 sg13g2_buf_2 fanout1983 (.A(net1985),
    .X(net1983));
 sg13g2_buf_4 fanout1984 (.X(net1984),
    .A(net1985));
 sg13g2_buf_4 fanout1985 (.X(net1985),
    .A(_0822_));
 sg13g2_buf_2 fanout1986 (.A(net1987),
    .X(net1986));
 sg13g2_buf_2 fanout1987 (.A(net1992),
    .X(net1987));
 sg13g2_buf_4 fanout1988 (.X(net1988),
    .A(net1992));
 sg13g2_buf_1 fanout1989 (.A(net1992),
    .X(net1989));
 sg13g2_buf_2 fanout1990 (.A(net1991),
    .X(net1990));
 sg13g2_buf_2 fanout1991 (.A(net1992),
    .X(net1991));
 sg13g2_buf_2 fanout1992 (.A(_0822_),
    .X(net1992));
 sg13g2_buf_4 fanout1993 (.X(net1993),
    .A(net1994));
 sg13g2_buf_4 fanout1994 (.X(net1994),
    .A(net1996));
 sg13g2_buf_2 fanout1995 (.A(net1996),
    .X(net1995));
 sg13g2_buf_4 fanout1996 (.X(net1996),
    .A(_0822_));
 sg13g2_buf_4 fanout1997 (.X(net1997),
    .A(_0821_));
 sg13g2_buf_2 fanout1998 (.A(net1999),
    .X(net1998));
 sg13g2_buf_4 fanout1999 (.X(net1999),
    .A(net2000));
 sg13g2_buf_4 fanout2000 (.X(net2000),
    .A(net2001));
 sg13g2_buf_4 fanout2001 (.X(net2001),
    .A(_0814_));
 sg13g2_buf_4 fanout2002 (.X(net2002),
    .A(_0813_));
 sg13g2_buf_4 fanout2003 (.X(net2003),
    .A(net2004));
 sg13g2_buf_4 fanout2004 (.X(net2004),
    .A(_0812_));
 sg13g2_buf_4 fanout2005 (.X(net2005),
    .A(_0810_));
 sg13g2_buf_4 fanout2006 (.X(net2006),
    .A(_0761_));
 sg13g2_buf_4 fanout2007 (.X(net2007),
    .A(_0761_));
 sg13g2_buf_4 fanout2008 (.X(net2008),
    .A(_0760_));
 sg13g2_buf_4 fanout2009 (.X(net2009),
    .A(_0736_));
 sg13g2_buf_2 fanout2010 (.A(_0736_),
    .X(net2010));
 sg13g2_buf_2 fanout2011 (.A(net2013),
    .X(net2011));
 sg13g2_buf_1 fanout2012 (.A(net2013),
    .X(net2012));
 sg13g2_buf_2 fanout2013 (.A(_0689_),
    .X(net2013));
 sg13g2_buf_4 fanout2014 (.X(net2014),
    .A(_0679_));
 sg13g2_buf_4 fanout2015 (.X(net2015),
    .A(net2017));
 sg13g2_buf_1 fanout2016 (.A(net2017),
    .X(net2016));
 sg13g2_buf_8 fanout2017 (.A(_0676_),
    .X(net2017));
 sg13g2_buf_4 fanout2018 (.X(net2018),
    .A(net2019));
 sg13g2_buf_4 fanout2019 (.X(net2019),
    .A(net2020));
 sg13g2_buf_4 fanout2020 (.X(net2020),
    .A(_0674_));
 sg13g2_buf_4 fanout2021 (.X(net2021),
    .A(_0673_));
 sg13g2_buf_2 fanout2022 (.A(_0673_),
    .X(net2022));
 sg13g2_buf_4 fanout2023 (.X(net2023),
    .A(net2024));
 sg13g2_buf_8 fanout2024 (.A(_0672_),
    .X(net2024));
 sg13g2_buf_4 fanout2025 (.X(net2025),
    .A(_0668_));
 sg13g2_buf_1 fanout2026 (.A(_0668_),
    .X(net2026));
 sg13g2_buf_2 fanout2027 (.A(net635),
    .X(net2027));
 sg13g2_buf_4 fanout2028 (.X(net2028),
    .A(net601));
 sg13g2_buf_4 fanout2029 (.X(net2029),
    .A(net602));
 sg13g2_buf_2 fanout2030 (.A(net2031),
    .X(net2030));
 sg13g2_buf_2 fanout2031 (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(net2031));
 sg13g2_buf_2 fanout2032 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net2032));
 sg13g2_buf_2 fanout2033 (.A(net593),
    .X(net2033));
 sg13g2_buf_2 fanout2034 (.A(net2035),
    .X(net2034));
 sg13g2_buf_2 fanout2035 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(net2035));
 sg13g2_buf_2 fanout2036 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .X(net2036));
 sg13g2_buf_4 fanout2037 (.X(net2037),
    .A(net2039));
 sg13g2_buf_2 fanout2038 (.A(net2039),
    .X(net2038));
 sg13g2_buf_2 fanout2039 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .X(net2039));
 sg13g2_buf_2 fanout2040 (.A(net2041),
    .X(net2040));
 sg13g2_buf_2 fanout2041 (.A(net2042),
    .X(net2041));
 sg13g2_buf_2 fanout2042 (.A(net559),
    .X(net2042));
 sg13g2_buf_4 fanout2043 (.X(net2043),
    .A(net612));
 sg13g2_buf_2 fanout2044 (.A(\z80.tv80s.di_reg[7] ),
    .X(net2044));
 sg13g2_buf_4 fanout2045 (.X(net2045),
    .A(\z80.tv80s.di_reg[6] ));
 sg13g2_buf_4 fanout2046 (.X(net2046),
    .A(\z80.tv80s.di_reg[5] ));
 sg13g2_buf_4 fanout2047 (.X(net2047),
    .A(\z80.tv80s.di_reg[4] ));
 sg13g2_buf_4 fanout2048 (.X(net2048),
    .A(\z80.tv80s.di_reg[3] ));
 sg13g2_buf_4 fanout2049 (.X(net2049),
    .A(\z80.tv80s.di_reg[2] ));
 sg13g2_buf_4 fanout2050 (.X(net2050),
    .A(\z80.tv80s.di_reg[1] ));
 sg13g2_buf_4 fanout2051 (.X(net2051),
    .A(\z80.tv80s.di_reg[0] ));
 sg13g2_buf_4 fanout2052 (.X(net2052),
    .A(net2053));
 sg13g2_buf_4 fanout2053 (.X(net2053),
    .A(\z80.tv80s.i_tv80_core.XY_Ind ));
 sg13g2_buf_1 fanout2054 (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(net2054));
 sg13g2_buf_4 fanout2055 (.X(net2055),
    .A(net2057));
 sg13g2_buf_1 fanout2056 (.A(net2057),
    .X(net2056));
 sg13g2_buf_2 fanout2057 (.A(net630),
    .X(net2057));
 sg13g2_buf_4 fanout2058 (.X(net2058),
    .A(\z80.tv80s.i_tv80_core.IR[6] ));
 sg13g2_buf_4 fanout2059 (.X(net2059),
    .A(net626));
 sg13g2_buf_2 fanout2060 (.A(net623),
    .X(net2060));
 sg13g2_buf_4 fanout2061 (.X(net2061),
    .A(_0235_));
 sg13g2_buf_2 fanout2062 (.A(net2063),
    .X(net2062));
 sg13g2_buf_4 fanout2063 (.X(net2063),
    .A(net2069));
 sg13g2_buf_4 fanout2064 (.X(net2064),
    .A(net2065));
 sg13g2_buf_2 fanout2065 (.A(net2066),
    .X(net2065));
 sg13g2_buf_2 fanout2066 (.A(net2067),
    .X(net2066));
 sg13g2_buf_2 fanout2067 (.A(net2068),
    .X(net2067));
 sg13g2_buf_4 fanout2068 (.X(net2068),
    .A(net2069));
 sg13g2_buf_2 fanout2069 (.A(net568),
    .X(net2069));
 sg13g2_buf_4 fanout2070 (.X(net2070),
    .A(net2071));
 sg13g2_buf_1 fanout2071 (.A(net2072),
    .X(net2071));
 sg13g2_buf_2 fanout2072 (.A(net585),
    .X(net2072));
 sg13g2_buf_4 fanout2073 (.X(net2073),
    .A(net2074));
 sg13g2_buf_2 fanout2074 (.A(net2075),
    .X(net2074));
 sg13g2_buf_4 fanout2075 (.X(net2075),
    .A(\z80.tv80s.i_tv80_core.IR[4] ));
 sg13g2_buf_4 fanout2076 (.X(net2076),
    .A(net2079));
 sg13g2_buf_2 fanout2077 (.A(net2078),
    .X(net2077));
 sg13g2_buf_2 fanout2078 (.A(net2079),
    .X(net2078));
 sg13g2_buf_4 fanout2079 (.X(net2079),
    .A(net617));
 sg13g2_buf_4 fanout2080 (.X(net2080),
    .A(net2081));
 sg13g2_buf_2 fanout2081 (.A(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(net2081));
 sg13g2_buf_4 fanout2082 (.X(net2082),
    .A(net2087));
 sg13g2_buf_4 fanout2083 (.X(net2083),
    .A(net2085));
 sg13g2_buf_1 fanout2084 (.A(net2085),
    .X(net2084));
 sg13g2_buf_1 fanout2085 (.A(net2086),
    .X(net2085));
 sg13g2_buf_2 fanout2086 (.A(net2087),
    .X(net2086));
 sg13g2_buf_2 fanout2087 (.A(net2088),
    .X(net2087));
 sg13g2_buf_4 fanout2088 (.X(net2088),
    .A(\z80.tv80s.i_tv80_core.IR[3] ));
 sg13g2_buf_2 fanout2089 (.A(net2092),
    .X(net2089));
 sg13g2_buf_2 fanout2090 (.A(net2091),
    .X(net2090));
 sg13g2_buf_4 fanout2091 (.X(net2091),
    .A(net2092));
 sg13g2_buf_2 fanout2092 (.A(net2093),
    .X(net2092));
 sg13g2_buf_4 fanout2093 (.X(net2093),
    .A(net571));
 sg13g2_buf_2 fanout2094 (.A(net2095),
    .X(net2094));
 sg13g2_buf_2 fanout2095 (.A(net2096),
    .X(net2095));
 sg13g2_buf_2 fanout2096 (.A(net2097),
    .X(net2096));
 sg13g2_buf_4 fanout2097 (.X(net2097),
    .A(net570));
 sg13g2_buf_2 fanout2098 (.A(net2100),
    .X(net2098));
 sg13g2_buf_2 fanout2099 (.A(net2100),
    .X(net2099));
 sg13g2_buf_1 fanout2100 (.A(net2101),
    .X(net2100));
 sg13g2_buf_2 fanout2101 (.A(net2102),
    .X(net2101));
 sg13g2_buf_4 fanout2102 (.X(net2102),
    .A(net565));
 sg13g2_buf_2 fanout2103 (.A(net2104),
    .X(net2103));
 sg13g2_buf_2 fanout2104 (.A(net2105),
    .X(net2104));
 sg13g2_buf_4 fanout2105 (.X(net2105),
    .A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sg13g2_buf_4 fanout2106 (.X(net2106),
    .A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sg13g2_buf_4 fanout2107 (.X(net2107),
    .A(net599));
 sg13g2_buf_2 fanout2108 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(net2108));
 sg13g2_buf_4 fanout2109 (.X(net2109),
    .A(net2110));
 sg13g2_buf_4 fanout2110 (.X(net2110),
    .A(net577));
 sg13g2_buf_4 fanout2111 (.X(net2111),
    .A(_0234_));
 sg13g2_buf_1 fanout2112 (.A(net2113),
    .X(net2112));
 sg13g2_buf_4 fanout2113 (.X(net2113),
    .A(_0234_));
 sg13g2_buf_2 fanout2114 (.A(net2117),
    .X(net2114));
 sg13g2_buf_1 fanout2115 (.A(net2117),
    .X(net2115));
 sg13g2_buf_2 fanout2116 (.A(net2117),
    .X(net2116));
 sg13g2_buf_2 fanout2117 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .X(net2117));
 sg13g2_buf_2 fanout2118 (.A(net2119),
    .X(net2118));
 sg13g2_buf_2 fanout2119 (.A(net2122),
    .X(net2119));
 sg13g2_buf_2 fanout2120 (.A(net2121),
    .X(net2120));
 sg13g2_buf_4 fanout2121 (.X(net2121),
    .A(net2122));
 sg13g2_buf_1 fanout2122 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .X(net2122));
 sg13g2_buf_4 fanout2123 (.X(net2123),
    .A(net2132));
 sg13g2_buf_4 fanout2124 (.X(net2124),
    .A(net2125));
 sg13g2_buf_2 fanout2125 (.A(net2126),
    .X(net2125));
 sg13g2_buf_4 fanout2126 (.X(net2126),
    .A(net2132));
 sg13g2_buf_2 fanout2127 (.A(net2130),
    .X(net2127));
 sg13g2_buf_2 fanout2128 (.A(net2130),
    .X(net2128));
 sg13g2_buf_2 fanout2129 (.A(net2130),
    .X(net2129));
 sg13g2_buf_4 fanout2130 (.X(net2130),
    .A(net2131));
 sg13g2_buf_4 fanout2131 (.X(net2131),
    .A(net2132));
 sg13g2_buf_2 fanout2132 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .X(net2132));
 sg13g2_buf_2 fanout2133 (.A(net606),
    .X(net2133));
 sg13g2_buf_2 fanout2134 (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .X(net2134));
 sg13g2_buf_4 fanout2135 (.X(net2135),
    .A(net595));
 sg13g2_buf_4 fanout2136 (.X(net2136),
    .A(net588));
 sg13g2_buf_2 fanout2137 (.A(net2139),
    .X(net2137));
 sg13g2_buf_2 fanout2138 (.A(net2139),
    .X(net2138));
 sg13g2_buf_2 fanout2139 (.A(net2140),
    .X(net2139));
 sg13g2_buf_2 fanout2140 (.A(net2141),
    .X(net2140));
 sg13g2_buf_2 fanout2141 (.A(net2143),
    .X(net2141));
 sg13g2_buf_2 fanout2142 (.A(net2143),
    .X(net2142));
 sg13g2_buf_2 fanout2143 (.A(net2144),
    .X(net2143));
 sg13g2_buf_4 fanout2144 (.X(net2144),
    .A(\z80.tv80s.i_tv80_core.ts[3] ));
 sg13g2_buf_4 fanout2145 (.X(net2145),
    .A(\z80.tv80s.i_tv80_core.ACC[5] ));
 sg13g2_buf_4 fanout2146 (.X(net2146),
    .A(\z80.tv80s.i_tv80_core.ACC[3] ));
 sg13g2_buf_4 fanout2147 (.X(net2147),
    .A(\z80.tv80s.i_tv80_core.F[2] ));
 sg13g2_buf_2 fanout2148 (.A(net2149),
    .X(net2148));
 sg13g2_buf_2 fanout2149 (.A(net2150),
    .X(net2149));
 sg13g2_buf_2 fanout2150 (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .X(net2150));
 sg13g2_buf_8 fanout2151 (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .X(net2151));
 sg13g2_buf_2 fanout2152 (.A(net2153),
    .X(net2152));
 sg13g2_buf_2 fanout2153 (.A(net2154),
    .X(net2153));
 sg13g2_buf_2 fanout2154 (.A(net2162),
    .X(net2154));
 sg13g2_buf_2 fanout2155 (.A(net2156),
    .X(net2155));
 sg13g2_buf_2 fanout2156 (.A(net2162),
    .X(net2156));
 sg13g2_buf_4 fanout2157 (.X(net2157),
    .A(net2161));
 sg13g2_buf_4 fanout2158 (.X(net2158),
    .A(net2159));
 sg13g2_buf_2 fanout2159 (.A(net2160),
    .X(net2159));
 sg13g2_buf_4 fanout2160 (.X(net2160),
    .A(net2161));
 sg13g2_buf_2 fanout2161 (.A(net2162),
    .X(net2161));
 sg13g2_buf_2 fanout2162 (.A(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .X(net2162));
 sg13g2_buf_4 fanout2163 (.X(net2163),
    .A(net2165));
 sg13g2_buf_4 fanout2164 (.X(net2164),
    .A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sg13g2_buf_2 fanout2165 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .X(net2165));
 sg13g2_buf_2 fanout2166 (.A(net620),
    .X(net2166));
 sg13g2_buf_2 fanout2167 (.A(\z80.tv80s.i_tv80_core.ISet[2] ),
    .X(net2167));
 sg13g2_buf_4 fanout2168 (.X(net2168),
    .A(net636));
 sg13g2_buf_2 fanout2169 (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(net2169));
 sg13g2_buf_2 fanout2170 (.A(net2171),
    .X(net2170));
 sg13g2_buf_4 fanout2171 (.X(net2171),
    .A(\z80.tv80s.i_tv80_core.ISet[0] ));
 sg13g2_buf_4 fanout2172 (.X(net2172),
    .A(net547));
 sg13g2_buf_4 fanout2173 (.X(net2173),
    .A(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sg13g2_buf_4 fanout2174 (.X(net2174),
    .A(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sg13g2_buf_4 fanout2175 (.X(net2175),
    .A(net2176));
 sg13g2_buf_4 fanout2176 (.X(net2176),
    .A(net2180));
 sg13g2_buf_4 fanout2177 (.X(net2177),
    .A(net2180));
 sg13g2_buf_4 fanout2178 (.X(net2178),
    .A(net2179));
 sg13g2_buf_4 fanout2179 (.X(net2179),
    .A(net2180));
 sg13g2_buf_4 fanout2180 (.X(net2180),
    .A(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sg13g2_buf_2 fanout2181 (.A(net2183),
    .X(net2181));
 sg13g2_buf_1 fanout2182 (.A(net2183),
    .X(net2182));
 sg13g2_buf_2 fanout2183 (.A(_0685_),
    .X(net2183));
 sg13g2_buf_2 fanout2184 (.A(net2185),
    .X(net2184));
 sg13g2_buf_2 fanout2185 (.A(ui_in[7]),
    .X(net2185));
 sg13g2_buf_2 fanout2186 (.A(net2188),
    .X(net2186));
 sg13g2_buf_1 fanout2187 (.A(net2188),
    .X(net2187));
 sg13g2_buf_2 fanout2188 (.A(ui_in[6]),
    .X(net2188));
 sg13g2_buf_4 fanout2189 (.X(net2189),
    .A(net2191));
 sg13g2_buf_4 fanout2190 (.X(net2190),
    .A(net2201));
 sg13g2_buf_2 fanout2191 (.A(net2201),
    .X(net2191));
 sg13g2_buf_4 fanout2192 (.X(net2192),
    .A(net2193));
 sg13g2_buf_4 fanout2193 (.X(net2193),
    .A(net2195));
 sg13g2_buf_4 fanout2194 (.X(net2194),
    .A(net2195));
 sg13g2_buf_2 fanout2195 (.A(net2201),
    .X(net2195));
 sg13g2_buf_4 fanout2196 (.X(net2196),
    .A(net2201));
 sg13g2_buf_2 fanout2197 (.A(net2201),
    .X(net2197));
 sg13g2_buf_4 fanout2198 (.X(net2198),
    .A(net2200));
 sg13g2_buf_4 fanout2199 (.X(net2199),
    .A(net2200));
 sg13g2_buf_4 fanout2200 (.X(net2200),
    .A(net2201));
 sg13g2_buf_4 fanout2201 (.X(net2201),
    .A(net2212));
 sg13g2_buf_4 fanout2202 (.X(net2202),
    .A(net2204));
 sg13g2_buf_4 fanout2203 (.X(net2203),
    .A(net2204));
 sg13g2_buf_4 fanout2204 (.X(net2204),
    .A(net2212));
 sg13g2_buf_4 fanout2205 (.X(net2205),
    .A(net2206));
 sg13g2_buf_4 fanout2206 (.X(net2206),
    .A(net2212));
 sg13g2_buf_4 fanout2207 (.X(net2207),
    .A(net2211));
 sg13g2_buf_2 fanout2208 (.A(net2211),
    .X(net2208));
 sg13g2_buf_4 fanout2209 (.X(net2209),
    .A(net2211));
 sg13g2_buf_2 fanout2210 (.A(net2211),
    .X(net2210));
 sg13g2_buf_1 fanout2211 (.A(net2212),
    .X(net2211));
 sg13g2_buf_2 fanout2212 (.A(net2226),
    .X(net2212));
 sg13g2_buf_4 fanout2213 (.X(net2213),
    .A(net2214));
 sg13g2_buf_4 fanout2214 (.X(net2214),
    .A(net2226));
 sg13g2_buf_4 fanout2215 (.X(net2215),
    .A(net2218));
 sg13g2_buf_4 fanout2216 (.X(net2216),
    .A(net2218));
 sg13g2_buf_4 fanout2217 (.X(net2217),
    .A(net2218));
 sg13g2_buf_2 fanout2218 (.A(net2226),
    .X(net2218));
 sg13g2_buf_4 fanout2219 (.X(net2219),
    .A(net2221));
 sg13g2_buf_2 fanout2220 (.A(net2221),
    .X(net2220));
 sg13g2_buf_4 fanout2221 (.X(net2221),
    .A(net2225));
 sg13g2_buf_4 fanout2222 (.X(net2222),
    .A(net2225));
 sg13g2_buf_4 fanout2223 (.X(net2223),
    .A(net2224));
 sg13g2_buf_4 fanout2224 (.X(net2224),
    .A(net2225));
 sg13g2_buf_2 fanout2225 (.A(net2226),
    .X(net2225));
 sg13g2_buf_2 fanout2226 (.A(rst_n),
    .X(net2226));
 sg13g2_buf_2 fanout2227 (.A(net2229),
    .X(net2227));
 sg13g2_buf_1 fanout2228 (.A(net2229),
    .X(net2228));
 sg13g2_buf_2 fanout2229 (.A(ena),
    .X(net2229));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[0]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[3]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[4]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[5]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[6]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[7]),
    .X(net12));
 sg13g2_tiehi _9126__13 (.L_HI(net13));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_62_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_11_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_59_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_61_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_63_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_64_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_65_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_9_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_13_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_24_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_8_clk));
 sg13g2_inv_2 clkload30 (.A(clknet_leaf_23_clk));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_51_clk));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_58_clk));
 sg13g2_inv_2 clkload35 (.A(clknet_leaf_54_clk));
 sg13g2_inv_1 clkload36 (.A(clknet_leaf_57_clk));
 sg13g2_inv_4 clkload37 (.A(clknet_leaf_44_clk));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_46_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_47_clk));
 sg13g2_inv_4 clkload40 (.A(clknet_leaf_40_clk));
 sg13g2_inv_8 clkload41 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload42 (.A(clknet_leaf_26_clk));
 sg13g2_inv_8 clkload43 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload44 (.A(clknet_leaf_53_clk));
 sg13g2_inv_2 clkload45 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload46 (.A(clknet_leaf_31_clk));
 sg13g2_inv_2 clkload47 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload48 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload49 (.A(clknet_leaf_37_clk));
 sg13g2_inv_8 clkload50 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload51 (.A(clknet_leaf_33_clk));
 sg13g2_inv_8 clkload52 (.A(clknet_leaf_34_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0030_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0563_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0231_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0615_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold5 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0307_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold7 (.A(\z80.tv80s.i_tv80_core.ts[5] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold8 (.A(_3654_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0282_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0546_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold11 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0306_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0266_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0274_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0538_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0276_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0540_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0290_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0270_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0534_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0275_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0539_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0269_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0248_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0272_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0536_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0250_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0264_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0268_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0532_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0265_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0529_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0263_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0527_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0267_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0531_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0029_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0557_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0262_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0526_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0273_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0537_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold43 (.A(\z80.tv80s.i_tv80_core.Oldnmi_n ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold44 (.A(_2504_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0446_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0240_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0278_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0261_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0525_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0256_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold51 (.A(_3360_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold52 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0271_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0535_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold55 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold56 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold57 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0283_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold59 (.A(\addr_bus[9] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0285_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold61 (.A(_3551_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold62 (.A(\addr_bus[1] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold63 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold64 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold65 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0252_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0260_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold68 (.A(_3396_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0245_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0279_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold71 (.A(_3465_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold72 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold73 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold74 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold75 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold76 (.A(\z80.tv80s.i_tv80_core.ISet[3] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold77 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold78 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold79 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold80 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold81 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0281_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold83 (.A(_3493_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0284_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold85 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold86 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold87 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold88 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold89 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold90 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold91 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold92 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold93 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold94 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0258_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold96 (.A(_3378_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold97 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold98 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold99 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0259_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold101 (.A(_3387_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold102 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold103 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold104 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold105 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold106 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold107 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold108 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold109 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold110 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold111 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold112 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold113 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold114 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold115 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold116 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold117 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold118 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold119 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold120 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold121 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[15] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0470_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold123 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold124 (.A(\addr_bus[13] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold125 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold126 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0286_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold128 (.A(\z80.tv80s.i_tv80_core.Z16_r ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0632_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold130 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold131 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold132 (.A(\addr_bus[12] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0254_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold134 (.A(_3342_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0249_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold136 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[13] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0468_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold138 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold139 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold140 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0288_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0246_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold143 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0243_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0344_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold146 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[14] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold147 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold148 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[2] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold149 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold150 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0295_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0612_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0251_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0255_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold155 (.A(_3351_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0280_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0253_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold158 (.A(_3333_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0277_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0247_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0491_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold162 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0005_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0289_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold165 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[12] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0467_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0291_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold168 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0244_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold170 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold171 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold172 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[5] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0460_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold174 (.A(\addr_bus[15] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold175 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[8] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0463_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold177 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold178 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold179 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold180 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[4] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0459_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold182 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold183 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold184 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[3] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0458_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold186 (.A(\addr_bus[11] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold187 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[9] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0287_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold189 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold190 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold191 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold192 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold193 (.A(\addr_bus[2] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold194 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold195 (.A(\addr_bus[3] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold196 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold197 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold198 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0257_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold200 (.A(_3369_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold201 (.A(\addr_bus[5] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold202 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold203 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold204 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold205 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold206 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold207 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold208 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold209 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold210 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold211 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold212 (.A(\addr_bus[14] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold213 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold214 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[10] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0465_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold216 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold217 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[11] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold218 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold219 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold220 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold221 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold222 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold223 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold224 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold225 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold226 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold227 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold228 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold229 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold230 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold231 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold232 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold233 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold234 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold235 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold236 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold237 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold238 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold239 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[6] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0461_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold241 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold242 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold243 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold244 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold245 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold246 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold247 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold248 (.A(\z80.tv80s.i_tv80_core.INT_s ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold249 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold250 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold251 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold252 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[1] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold253 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold254 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold255 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold256 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold257 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold258 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold259 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold260 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold261 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold262 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[7] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0462_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold264 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold265 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold266 (.A(\z80.tv80s.i_tv80_core.BTR_r ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0616_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold268 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold269 (.A(\addr_bus[10] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold270 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold271 (.A(\addr_bus[4] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold272 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold273 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold274 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold275 (.A(\addr_bus[7] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0480_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0241_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0242_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0294_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0597_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold281 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold282 (.A(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold283 (.A(uio_out[4]),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold284 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0167_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0472_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold287 (.A(\z80.tv80s.i_tv80_core.ts[0] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0558_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0227_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0444_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0232_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0505_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold293 (.A(uio_out[7]),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0032_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0559_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold296 (.A(\z80.tv80s.i_tv80_core.IntE ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold297 (.A(\addr_bus[8] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0481_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold299 (.A(\addr_bus[0] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0473_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold301 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold302 (.A(\z80.tv80s.i_tv80_core.IStatus[2] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold303 (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0441_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold305 (.A(uio_out[6]),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold306 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0009_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold308 (.A(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold309 (.A(\z80.tv80s.i_tv80_core.BusAck ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold310 (.A(_2477_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0442_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold312 (.A(\z80.tv80s.i_tv80_core.IncDecZ ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold313 (.A(uio_out[1]),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold314 (.A(uio_out[3]),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold315 (.A(uio_out[5]),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold316 (.A(uio_out[2]),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold317 (.A(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold318 (.A(\addr_bus[6] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0479_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold320 (.A(\z80.tv80s.i_tv80_core.R[1] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold321 (.A(_1470_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0298_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold323 (.A(uio_out[0]),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0508_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold325 (.A(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0596_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold327 (.A(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold328 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold329 (.A(\z80.tv80s.i_tv80_core.R[7] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold330 (.A(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold331 (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0593_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold333 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0031_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0292_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold336 (.A(\z80.tv80s.i_tv80_core.PC[0] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0564_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold338 (.A(\z80.tv80s.i_tv80_core.R[4] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold339 (.A(_1480_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0301_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold341 (.A(\z80.tv80s.i_tv80_core.R[6] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold342 (.A(_1486_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold343 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold344 (.A(\z80.tv80s.i_tv80_core.ISet[1] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold345 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold346 (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0565_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold348 (.A(\z80.tv80s.i_tv80_core.PreserveC_r ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold349 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold350 (.A(\z80.tv80s.i_tv80_core.Alternate ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0580_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold352 (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold353 (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0594_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold355 (.A(\z80.tv80s.i_tv80_core.R[3] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0300_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold357 (.A(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold358 (.A(\z80.tv80s.i_tv80_core.R[2] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0299_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold360 (.A(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold361 (.A(\z80.tv80s.i_tv80_core.PC[13] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold362 (.A(\z80.tv80s.i_tv80_core.PC[2] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold363 (.A(\z80.tv80s.i_tv80_core.ts[4] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0561_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold365 (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0296_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold367 (.A(\z80.tv80s.i_tv80_core.PC[3] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold368 (.A(\z80.tv80s.i_tv80_core.R[5] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold369 (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold370 (.A(\z80.tv80s.di_reg[2] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0583_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold372 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0601_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold374 (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold375 (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold376 (.A(\z80.tv80s.i_tv80_core.BusReq_s ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold377 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold378 (.A(\z80.tv80s.i_tv80_core.PC[9] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold379 (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold380 (.A(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold381 (.A(\z80.tv80s.i_tv80_core.R[0] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0297_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold383 (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold384 (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold385 (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold386 (.A(\z80.tv80s.i_tv80_core.IR[5] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold387 (.A(\z80.tv80s.i_tv80_core.BusB[4] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold388 (.A(\z80.tv80s.i_tv80_core.IR[1] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold389 (.A(\z80.tv80s.i_tv80_core.IR[2] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold390 (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold391 (.A(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold392 (.A(\z80.tv80s.i_tv80_core.PC[12] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold393 (.A(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold394 (.A(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold395 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold396 (.A(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0647_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold398 (.A(\z80.tv80s.i_tv80_core.NMI_s ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0443_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold400 (.A(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold401 (.A(\z80.tv80s.i_tv80_core.PC[11] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold402 (.A(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold403 (.A(\z80.tv80s.i_tv80_core.IR[4] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0237_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold405 (.A(_4087_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold406 (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold407 (.A(\z80.tv80s.i_tv80_core.PC[14] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold408 (.A(\z80.tv80s.i_tv80_core.PC[15] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold409 (.A(\z80.tv80s.i_tv80_core.Arith16_r ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold410 (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold411 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold412 (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold413 (.A(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold414 (.A(\z80.tv80s.i_tv80_core.IntCycle ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold415 (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold416 (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold417 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold418 (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold419 (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold420 (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold421 (.A(\z80.tv80s.i_tv80_core.PC[5] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold422 (.A(\z80.tv80s.i_tv80_core.I[2] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0499_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold424 (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0586_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold426 (.A(\z80.tv80s.i_tv80_core.I[6] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0503_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold428 (.A(\z80.tv80s.i_tv80_core.I[1] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0498_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold430 (.A(\z80.tv80s.di_reg[7] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold431 (.A(\z80.tv80s.i_tv80_core.I[5] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold432 (.A(\z80.tv80s.i_tv80_core.I[0] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold433 (.A(\z80.tv80s.i_tv80_core.I[4] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0501_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold435 (.A(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold436 (.A(\z80.tv80s.i_tv80_core.I[3] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold437 (.A(\z80.tv80s.i_tv80_core.PC[8] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold438 (.A(\z80.tv80s.i_tv80_core.ISet[2] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold439 (.A(_1421_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold440 (.A(\z80.tv80s.i_tv80_core.PC[10] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0235_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0614_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold443 (.A(\z80.tv80s.i_tv80_core.BusReq_s ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold444 (.A(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold445 (.A(_0025_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold446 (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0571_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold448 (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold449 (.A(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold450 (.A(\z80.tv80s.i_tv80_core.PC[6] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold451 (.A(\z80.tv80s.i_tv80_core.I[7] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0504_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold453 (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold454 (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(net636));
 sg13g2_antennanp ANTENNA_1 (.A(_0611_));
 sg13g2_antennanp ANTENNA_2 (.A(_3084_));
 sg13g2_antennanp ANTENNA_3 (.A(_3084_));
 sg13g2_antennanp ANTENNA_4 (.A(_3084_));
 sg13g2_antennanp ANTENNA_5 (.A(_0611_));
 sg13g2_antennanp ANTENNA_6 (.A(_0611_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_fill_2 FILLER_3_196 ();
 sg13g2_fill_1 FILLER_3_202 ();
 sg13g2_fill_2 FILLER_3_212 ();
 sg13g2_decap_8 FILLER_3_223 ();
 sg13g2_decap_8 FILLER_3_230 ();
 sg13g2_decap_8 FILLER_3_237 ();
 sg13g2_decap_8 FILLER_3_244 ();
 sg13g2_decap_8 FILLER_3_260 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_288 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_309 ();
 sg13g2_fill_2 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_fill_2 FILLER_4_185 ();
 sg13g2_fill_1 FILLER_4_187 ();
 sg13g2_decap_4 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_229 ();
 sg13g2_decap_4 FILLER_4_236 ();
 sg13g2_fill_2 FILLER_4_240 ();
 sg13g2_fill_2 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_fill_2 FILLER_4_281 ();
 sg13g2_fill_1 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_decap_8 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_4_415 ();
 sg13g2_decap_8 FILLER_4_422 ();
 sg13g2_decap_8 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_4_436 ();
 sg13g2_decap_8 FILLER_4_443 ();
 sg13g2_decap_8 FILLER_4_450 ();
 sg13g2_decap_8 FILLER_4_457 ();
 sg13g2_decap_8 FILLER_4_464 ();
 sg13g2_decap_8 FILLER_4_471 ();
 sg13g2_decap_8 FILLER_4_478 ();
 sg13g2_decap_8 FILLER_4_485 ();
 sg13g2_decap_8 FILLER_4_492 ();
 sg13g2_decap_8 FILLER_4_499 ();
 sg13g2_decap_8 FILLER_4_506 ();
 sg13g2_decap_8 FILLER_4_513 ();
 sg13g2_decap_8 FILLER_4_520 ();
 sg13g2_decap_8 FILLER_4_527 ();
 sg13g2_decap_8 FILLER_4_534 ();
 sg13g2_decap_8 FILLER_4_541 ();
 sg13g2_decap_8 FILLER_4_548 ();
 sg13g2_decap_8 FILLER_4_555 ();
 sg13g2_decap_8 FILLER_4_562 ();
 sg13g2_decap_8 FILLER_4_569 ();
 sg13g2_decap_8 FILLER_4_576 ();
 sg13g2_decap_8 FILLER_4_583 ();
 sg13g2_decap_8 FILLER_4_590 ();
 sg13g2_decap_8 FILLER_4_597 ();
 sg13g2_decap_8 FILLER_4_604 ();
 sg13g2_decap_8 FILLER_4_611 ();
 sg13g2_decap_8 FILLER_4_618 ();
 sg13g2_decap_8 FILLER_4_625 ();
 sg13g2_decap_8 FILLER_4_632 ();
 sg13g2_decap_8 FILLER_4_639 ();
 sg13g2_decap_8 FILLER_4_646 ();
 sg13g2_decap_8 FILLER_4_653 ();
 sg13g2_decap_8 FILLER_4_660 ();
 sg13g2_decap_8 FILLER_4_667 ();
 sg13g2_decap_8 FILLER_4_674 ();
 sg13g2_decap_8 FILLER_4_681 ();
 sg13g2_decap_8 FILLER_4_688 ();
 sg13g2_decap_8 FILLER_4_695 ();
 sg13g2_decap_8 FILLER_4_702 ();
 sg13g2_decap_8 FILLER_4_709 ();
 sg13g2_decap_8 FILLER_4_716 ();
 sg13g2_decap_8 FILLER_4_723 ();
 sg13g2_decap_8 FILLER_4_730 ();
 sg13g2_decap_8 FILLER_4_737 ();
 sg13g2_decap_8 FILLER_4_744 ();
 sg13g2_decap_8 FILLER_4_751 ();
 sg13g2_decap_8 FILLER_4_758 ();
 sg13g2_decap_8 FILLER_4_765 ();
 sg13g2_decap_8 FILLER_4_772 ();
 sg13g2_decap_8 FILLER_4_779 ();
 sg13g2_decap_8 FILLER_4_786 ();
 sg13g2_decap_8 FILLER_4_793 ();
 sg13g2_decap_8 FILLER_4_800 ();
 sg13g2_decap_8 FILLER_4_807 ();
 sg13g2_decap_8 FILLER_4_814 ();
 sg13g2_decap_8 FILLER_4_821 ();
 sg13g2_decap_8 FILLER_4_828 ();
 sg13g2_decap_8 FILLER_4_835 ();
 sg13g2_decap_8 FILLER_4_842 ();
 sg13g2_decap_8 FILLER_4_849 ();
 sg13g2_decap_4 FILLER_4_856 ();
 sg13g2_fill_2 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_fill_1 FILLER_5_161 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_fill_1 FILLER_5_270 ();
 sg13g2_fill_1 FILLER_5_297 ();
 sg13g2_fill_2 FILLER_5_327 ();
 sg13g2_decap_4 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_fill_1 FILLER_5_391 ();
 sg13g2_fill_2 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_5_415 ();
 sg13g2_fill_2 FILLER_5_436 ();
 sg13g2_fill_1 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_fill_1 FILLER_5_466 ();
 sg13g2_decap_8 FILLER_5_477 ();
 sg13g2_decap_4 FILLER_5_484 ();
 sg13g2_fill_1 FILLER_5_488 ();
 sg13g2_decap_8 FILLER_5_493 ();
 sg13g2_decap_8 FILLER_5_500 ();
 sg13g2_fill_2 FILLER_5_507 ();
 sg13g2_fill_1 FILLER_5_509 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_decap_8 FILLER_5_536 ();
 sg13g2_decap_8 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_550 ();
 sg13g2_decap_8 FILLER_5_557 ();
 sg13g2_decap_8 FILLER_5_564 ();
 sg13g2_decap_8 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_8 FILLER_5_599 ();
 sg13g2_decap_8 FILLER_5_606 ();
 sg13g2_decap_8 FILLER_5_613 ();
 sg13g2_decap_8 FILLER_5_620 ();
 sg13g2_decap_8 FILLER_5_627 ();
 sg13g2_decap_8 FILLER_5_634 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_decap_8 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_655 ();
 sg13g2_decap_8 FILLER_5_662 ();
 sg13g2_decap_8 FILLER_5_669 ();
 sg13g2_decap_8 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_683 ();
 sg13g2_decap_8 FILLER_5_690 ();
 sg13g2_decap_8 FILLER_5_697 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_725 ();
 sg13g2_decap_8 FILLER_5_732 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_4 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_128 ();
 sg13g2_decap_8 FILLER_6_138 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_fill_1 FILLER_6_172 ();
 sg13g2_decap_4 FILLER_6_229 ();
 sg13g2_fill_2 FILLER_6_252 ();
 sg13g2_fill_2 FILLER_6_267 ();
 sg13g2_fill_1 FILLER_6_269 ();
 sg13g2_fill_1 FILLER_6_293 ();
 sg13g2_decap_4 FILLER_6_304 ();
 sg13g2_fill_1 FILLER_6_334 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_fill_2 FILLER_6_382 ();
 sg13g2_fill_2 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_fill_2 FILLER_6_491 ();
 sg13g2_fill_1 FILLER_6_529 ();
 sg13g2_decap_8 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_599 ();
 sg13g2_decap_8 FILLER_6_606 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_4 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_112 ();
 sg13g2_fill_1 FILLER_7_195 ();
 sg13g2_fill_2 FILLER_7_240 ();
 sg13g2_fill_1 FILLER_7_242 ();
 sg13g2_decap_4 FILLER_7_295 ();
 sg13g2_fill_2 FILLER_7_299 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_4 FILLER_7_337 ();
 sg13g2_fill_2 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_fill_2 FILLER_7_367 ();
 sg13g2_fill_1 FILLER_7_369 ();
 sg13g2_fill_2 FILLER_7_405 ();
 sg13g2_fill_1 FILLER_7_407 ();
 sg13g2_fill_2 FILLER_7_418 ();
 sg13g2_decap_4 FILLER_7_460 ();
 sg13g2_fill_1 FILLER_7_464 ();
 sg13g2_fill_1 FILLER_7_479 ();
 sg13g2_fill_2 FILLER_7_516 ();
 sg13g2_fill_1 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_545 ();
 sg13g2_decap_8 FILLER_7_552 ();
 sg13g2_decap_8 FILLER_7_559 ();
 sg13g2_decap_8 FILLER_7_566 ();
 sg13g2_decap_8 FILLER_7_573 ();
 sg13g2_decap_8 FILLER_7_580 ();
 sg13g2_decap_8 FILLER_7_587 ();
 sg13g2_decap_8 FILLER_7_594 ();
 sg13g2_decap_8 FILLER_7_601 ();
 sg13g2_decap_8 FILLER_7_608 ();
 sg13g2_decap_8 FILLER_7_615 ();
 sg13g2_decap_8 FILLER_7_622 ();
 sg13g2_decap_8 FILLER_7_629 ();
 sg13g2_decap_8 FILLER_7_636 ();
 sg13g2_decap_8 FILLER_7_643 ();
 sg13g2_decap_8 FILLER_7_650 ();
 sg13g2_decap_8 FILLER_7_657 ();
 sg13g2_decap_8 FILLER_7_664 ();
 sg13g2_decap_8 FILLER_7_671 ();
 sg13g2_decap_8 FILLER_7_678 ();
 sg13g2_decap_8 FILLER_7_685 ();
 sg13g2_decap_8 FILLER_7_692 ();
 sg13g2_decap_8 FILLER_7_699 ();
 sg13g2_decap_8 FILLER_7_706 ();
 sg13g2_decap_8 FILLER_7_713 ();
 sg13g2_decap_8 FILLER_7_720 ();
 sg13g2_decap_8 FILLER_7_727 ();
 sg13g2_decap_8 FILLER_7_734 ();
 sg13g2_decap_8 FILLER_7_741 ();
 sg13g2_decap_8 FILLER_7_748 ();
 sg13g2_decap_8 FILLER_7_755 ();
 sg13g2_decap_8 FILLER_7_762 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_8 FILLER_7_804 ();
 sg13g2_decap_8 FILLER_7_811 ();
 sg13g2_decap_8 FILLER_7_818 ();
 sg13g2_decap_8 FILLER_7_825 ();
 sg13g2_decap_8 FILLER_7_832 ();
 sg13g2_decap_8 FILLER_7_839 ();
 sg13g2_decap_8 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_853 ();
 sg13g2_fill_2 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_decap_4 FILLER_8_210 ();
 sg13g2_fill_2 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_fill_1 FILLER_8_234 ();
 sg13g2_decap_4 FILLER_8_270 ();
 sg13g2_fill_2 FILLER_8_274 ();
 sg13g2_fill_1 FILLER_8_290 ();
 sg13g2_decap_4 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_363 ();
 sg13g2_fill_1 FILLER_8_365 ();
 sg13g2_fill_2 FILLER_8_452 ();
 sg13g2_fill_2 FILLER_8_512 ();
 sg13g2_fill_1 FILLER_8_514 ();
 sg13g2_fill_2 FILLER_8_543 ();
 sg13g2_fill_1 FILLER_8_545 ();
 sg13g2_fill_2 FILLER_8_556 ();
 sg13g2_fill_1 FILLER_8_558 ();
 sg13g2_decap_8 FILLER_8_577 ();
 sg13g2_decap_8 FILLER_8_584 ();
 sg13g2_decap_8 FILLER_8_591 ();
 sg13g2_decap_8 FILLER_8_598 ();
 sg13g2_decap_8 FILLER_8_605 ();
 sg13g2_decap_8 FILLER_8_612 ();
 sg13g2_decap_8 FILLER_8_619 ();
 sg13g2_decap_8 FILLER_8_626 ();
 sg13g2_decap_8 FILLER_8_633 ();
 sg13g2_decap_8 FILLER_8_640 ();
 sg13g2_decap_8 FILLER_8_647 ();
 sg13g2_decap_8 FILLER_8_654 ();
 sg13g2_decap_8 FILLER_8_661 ();
 sg13g2_decap_8 FILLER_8_668 ();
 sg13g2_decap_8 FILLER_8_675 ();
 sg13g2_decap_8 FILLER_8_682 ();
 sg13g2_decap_8 FILLER_8_689 ();
 sg13g2_decap_8 FILLER_8_696 ();
 sg13g2_decap_8 FILLER_8_703 ();
 sg13g2_decap_8 FILLER_8_710 ();
 sg13g2_decap_8 FILLER_8_717 ();
 sg13g2_decap_8 FILLER_8_724 ();
 sg13g2_decap_8 FILLER_8_731 ();
 sg13g2_decap_8 FILLER_8_738 ();
 sg13g2_decap_8 FILLER_8_745 ();
 sg13g2_decap_8 FILLER_8_752 ();
 sg13g2_decap_8 FILLER_8_759 ();
 sg13g2_decap_8 FILLER_8_766 ();
 sg13g2_decap_8 FILLER_8_773 ();
 sg13g2_decap_8 FILLER_8_780 ();
 sg13g2_decap_8 FILLER_8_787 ();
 sg13g2_decap_8 FILLER_8_794 ();
 sg13g2_decap_8 FILLER_8_801 ();
 sg13g2_decap_8 FILLER_8_808 ();
 sg13g2_decap_8 FILLER_8_815 ();
 sg13g2_decap_8 FILLER_8_822 ();
 sg13g2_decap_8 FILLER_8_829 ();
 sg13g2_decap_8 FILLER_8_836 ();
 sg13g2_decap_8 FILLER_8_843 ();
 sg13g2_decap_8 FILLER_8_850 ();
 sg13g2_decap_4 FILLER_8_857 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_4 FILLER_9_91 ();
 sg13g2_fill_2 FILLER_9_104 ();
 sg13g2_fill_1 FILLER_9_106 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_180 ();
 sg13g2_fill_2 FILLER_9_187 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_fill_1 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_240 ();
 sg13g2_fill_2 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_263 ();
 sg13g2_decap_4 FILLER_9_290 ();
 sg13g2_fill_2 FILLER_9_366 ();
 sg13g2_fill_2 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_406 ();
 sg13g2_fill_2 FILLER_9_426 ();
 sg13g2_fill_1 FILLER_9_428 ();
 sg13g2_fill_2 FILLER_9_469 ();
 sg13g2_fill_2 FILLER_9_515 ();
 sg13g2_fill_1 FILLER_9_517 ();
 sg13g2_fill_2 FILLER_9_544 ();
 sg13g2_fill_1 FILLER_9_546 ();
 sg13g2_fill_1 FILLER_9_573 ();
 sg13g2_decap_8 FILLER_9_584 ();
 sg13g2_decap_8 FILLER_9_591 ();
 sg13g2_fill_2 FILLER_9_598 ();
 sg13g2_fill_1 FILLER_9_600 ();
 sg13g2_decap_8 FILLER_9_611 ();
 sg13g2_decap_8 FILLER_9_618 ();
 sg13g2_decap_8 FILLER_9_625 ();
 sg13g2_decap_8 FILLER_9_632 ();
 sg13g2_decap_8 FILLER_9_639 ();
 sg13g2_decap_8 FILLER_9_646 ();
 sg13g2_decap_8 FILLER_9_653 ();
 sg13g2_decap_8 FILLER_9_660 ();
 sg13g2_decap_8 FILLER_9_667 ();
 sg13g2_decap_8 FILLER_9_674 ();
 sg13g2_decap_8 FILLER_9_681 ();
 sg13g2_decap_8 FILLER_9_688 ();
 sg13g2_decap_8 FILLER_9_695 ();
 sg13g2_decap_8 FILLER_9_702 ();
 sg13g2_decap_8 FILLER_9_709 ();
 sg13g2_decap_8 FILLER_9_716 ();
 sg13g2_decap_8 FILLER_9_723 ();
 sg13g2_decap_8 FILLER_9_730 ();
 sg13g2_decap_8 FILLER_9_737 ();
 sg13g2_decap_8 FILLER_9_744 ();
 sg13g2_decap_8 FILLER_9_751 ();
 sg13g2_decap_8 FILLER_9_758 ();
 sg13g2_decap_8 FILLER_9_765 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_decap_8 FILLER_9_779 ();
 sg13g2_decap_8 FILLER_9_786 ();
 sg13g2_decap_8 FILLER_9_793 ();
 sg13g2_decap_8 FILLER_9_800 ();
 sg13g2_decap_8 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_8 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_9_835 ();
 sg13g2_decap_8 FILLER_9_842 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_decap_4 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_fill_2 FILLER_10_84 ();
 sg13g2_fill_1 FILLER_10_86 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_4 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_167 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_219 ();
 sg13g2_fill_1 FILLER_10_226 ();
 sg13g2_decap_4 FILLER_10_286 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_342 ();
 sg13g2_fill_1 FILLER_10_344 ();
 sg13g2_fill_1 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_430 ();
 sg13g2_fill_2 FILLER_10_446 ();
 sg13g2_fill_1 FILLER_10_457 ();
 sg13g2_decap_4 FILLER_10_548 ();
 sg13g2_fill_1 FILLER_10_552 ();
 sg13g2_fill_2 FILLER_10_583 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_669 ();
 sg13g2_decap_8 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_683 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_4 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_fill_1 FILLER_11_70 ();
 sg13g2_fill_2 FILLER_11_107 ();
 sg13g2_fill_2 FILLER_11_145 ();
 sg13g2_decap_4 FILLER_11_153 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_192 ();
 sg13g2_fill_2 FILLER_11_229 ();
 sg13g2_decap_4 FILLER_11_239 ();
 sg13g2_fill_1 FILLER_11_250 ();
 sg13g2_fill_2 FILLER_11_285 ();
 sg13g2_fill_2 FILLER_11_300 ();
 sg13g2_fill_2 FILLER_11_346 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_4 FILLER_11_375 ();
 sg13g2_decap_4 FILLER_11_383 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_fill_2 FILLER_11_398 ();
 sg13g2_decap_8 FILLER_11_426 ();
 sg13g2_decap_4 FILLER_11_485 ();
 sg13g2_fill_1 FILLER_11_489 ();
 sg13g2_fill_2 FILLER_11_520 ();
 sg13g2_fill_1 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_549 ();
 sg13g2_fill_2 FILLER_11_556 ();
 sg13g2_fill_2 FILLER_11_566 ();
 sg13g2_decap_8 FILLER_11_578 ();
 sg13g2_decap_8 FILLER_11_585 ();
 sg13g2_fill_2 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_608 ();
 sg13g2_decap_4 FILLER_11_615 ();
 sg13g2_decap_8 FILLER_11_629 ();
 sg13g2_decap_8 FILLER_11_636 ();
 sg13g2_decap_8 FILLER_11_643 ();
 sg13g2_decap_8 FILLER_11_650 ();
 sg13g2_decap_8 FILLER_11_657 ();
 sg13g2_decap_8 FILLER_11_664 ();
 sg13g2_decap_8 FILLER_11_671 ();
 sg13g2_decap_8 FILLER_11_678 ();
 sg13g2_decap_8 FILLER_11_685 ();
 sg13g2_decap_8 FILLER_11_692 ();
 sg13g2_decap_8 FILLER_11_699 ();
 sg13g2_decap_8 FILLER_11_706 ();
 sg13g2_decap_8 FILLER_11_713 ();
 sg13g2_decap_8 FILLER_11_720 ();
 sg13g2_decap_8 FILLER_11_727 ();
 sg13g2_decap_8 FILLER_11_734 ();
 sg13g2_decap_8 FILLER_11_741 ();
 sg13g2_decap_8 FILLER_11_748 ();
 sg13g2_decap_8 FILLER_11_755 ();
 sg13g2_decap_8 FILLER_11_762 ();
 sg13g2_decap_8 FILLER_11_769 ();
 sg13g2_decap_8 FILLER_11_776 ();
 sg13g2_decap_8 FILLER_11_783 ();
 sg13g2_decap_8 FILLER_11_790 ();
 sg13g2_decap_8 FILLER_11_797 ();
 sg13g2_decap_8 FILLER_11_804 ();
 sg13g2_decap_8 FILLER_11_811 ();
 sg13g2_decap_8 FILLER_11_818 ();
 sg13g2_decap_8 FILLER_11_825 ();
 sg13g2_decap_8 FILLER_11_832 ();
 sg13g2_decap_8 FILLER_11_839 ();
 sg13g2_decap_8 FILLER_11_846 ();
 sg13g2_decap_8 FILLER_11_853 ();
 sg13g2_fill_2 FILLER_11_860 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_1 FILLER_12_85 ();
 sg13g2_fill_2 FILLER_12_122 ();
 sg13g2_fill_1 FILLER_12_124 ();
 sg13g2_fill_2 FILLER_12_138 ();
 sg13g2_fill_1 FILLER_12_161 ();
 sg13g2_fill_1 FILLER_12_166 ();
 sg13g2_decap_8 FILLER_12_197 ();
 sg13g2_decap_4 FILLER_12_235 ();
 sg13g2_fill_2 FILLER_12_239 ();
 sg13g2_fill_1 FILLER_12_249 ();
 sg13g2_fill_2 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_fill_2 FILLER_12_408 ();
 sg13g2_fill_2 FILLER_12_414 ();
 sg13g2_fill_1 FILLER_12_416 ();
 sg13g2_fill_2 FILLER_12_441 ();
 sg13g2_decap_4 FILLER_12_447 ();
 sg13g2_fill_2 FILLER_12_451 ();
 sg13g2_fill_1 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_fill_2 FILLER_12_490 ();
 sg13g2_fill_1 FILLER_12_492 ();
 sg13g2_decap_4 FILLER_12_504 ();
 sg13g2_fill_1 FILLER_12_544 ();
 sg13g2_fill_1 FILLER_12_551 ();
 sg13g2_decap_8 FILLER_12_650 ();
 sg13g2_decap_8 FILLER_12_657 ();
 sg13g2_decap_8 FILLER_12_664 ();
 sg13g2_decap_8 FILLER_12_671 ();
 sg13g2_decap_8 FILLER_12_678 ();
 sg13g2_decap_8 FILLER_12_685 ();
 sg13g2_decap_8 FILLER_12_692 ();
 sg13g2_decap_8 FILLER_12_699 ();
 sg13g2_decap_8 FILLER_12_706 ();
 sg13g2_decap_8 FILLER_12_713 ();
 sg13g2_decap_8 FILLER_12_720 ();
 sg13g2_decap_8 FILLER_12_727 ();
 sg13g2_decap_8 FILLER_12_734 ();
 sg13g2_decap_8 FILLER_12_741 ();
 sg13g2_decap_8 FILLER_12_748 ();
 sg13g2_decap_8 FILLER_12_755 ();
 sg13g2_decap_8 FILLER_12_762 ();
 sg13g2_decap_8 FILLER_12_769 ();
 sg13g2_decap_8 FILLER_12_776 ();
 sg13g2_decap_8 FILLER_12_783 ();
 sg13g2_decap_8 FILLER_12_790 ();
 sg13g2_decap_8 FILLER_12_797 ();
 sg13g2_decap_8 FILLER_12_804 ();
 sg13g2_decap_8 FILLER_12_811 ();
 sg13g2_decap_8 FILLER_12_818 ();
 sg13g2_decap_8 FILLER_12_825 ();
 sg13g2_decap_8 FILLER_12_832 ();
 sg13g2_decap_8 FILLER_12_839 ();
 sg13g2_decap_8 FILLER_12_846 ();
 sg13g2_decap_8 FILLER_12_853 ();
 sg13g2_fill_2 FILLER_12_860 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_fill_2 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_105 ();
 sg13g2_fill_1 FILLER_13_115 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_160 ();
 sg13g2_decap_4 FILLER_13_189 ();
 sg13g2_fill_2 FILLER_13_193 ();
 sg13g2_decap_4 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_decap_4 FILLER_13_293 ();
 sg13g2_fill_1 FILLER_13_297 ();
 sg13g2_decap_4 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_318 ();
 sg13g2_fill_2 FILLER_13_333 ();
 sg13g2_fill_2 FILLER_13_352 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_decap_4 FILLER_13_407 ();
 sg13g2_fill_2 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_475 ();
 sg13g2_fill_2 FILLER_13_482 ();
 sg13g2_fill_1 FILLER_13_484 ();
 sg13g2_fill_2 FILLER_13_507 ();
 sg13g2_fill_1 FILLER_13_509 ();
 sg13g2_fill_2 FILLER_13_537 ();
 sg13g2_decap_4 FILLER_13_547 ();
 sg13g2_fill_2 FILLER_13_561 ();
 sg13g2_fill_2 FILLER_13_578 ();
 sg13g2_decap_8 FILLER_13_649 ();
 sg13g2_decap_8 FILLER_13_656 ();
 sg13g2_decap_8 FILLER_13_663 ();
 sg13g2_decap_8 FILLER_13_670 ();
 sg13g2_decap_8 FILLER_13_677 ();
 sg13g2_decap_8 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_691 ();
 sg13g2_decap_8 FILLER_13_698 ();
 sg13g2_decap_8 FILLER_13_705 ();
 sg13g2_decap_8 FILLER_13_712 ();
 sg13g2_decap_8 FILLER_13_719 ();
 sg13g2_decap_8 FILLER_13_726 ();
 sg13g2_decap_8 FILLER_13_733 ();
 sg13g2_decap_8 FILLER_13_740 ();
 sg13g2_decap_8 FILLER_13_747 ();
 sg13g2_decap_8 FILLER_13_754 ();
 sg13g2_decap_8 FILLER_13_761 ();
 sg13g2_decap_8 FILLER_13_768 ();
 sg13g2_decap_8 FILLER_13_775 ();
 sg13g2_decap_8 FILLER_13_782 ();
 sg13g2_decap_8 FILLER_13_789 ();
 sg13g2_decap_8 FILLER_13_796 ();
 sg13g2_decap_8 FILLER_13_803 ();
 sg13g2_decap_8 FILLER_13_810 ();
 sg13g2_decap_8 FILLER_13_817 ();
 sg13g2_decap_8 FILLER_13_824 ();
 sg13g2_decap_8 FILLER_13_831 ();
 sg13g2_decap_8 FILLER_13_838 ();
 sg13g2_decap_8 FILLER_13_845 ();
 sg13g2_decap_8 FILLER_13_852 ();
 sg13g2_fill_2 FILLER_13_859 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_4 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_60 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_fill_2 FILLER_14_173 ();
 sg13g2_decap_8 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_fill_1 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_decap_4 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_4 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_277 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_fill_1 FILLER_14_325 ();
 sg13g2_fill_2 FILLER_14_352 ();
 sg13g2_fill_1 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_fill_1 FILLER_14_380 ();
 sg13g2_fill_1 FILLER_14_442 ();
 sg13g2_decap_8 FILLER_14_481 ();
 sg13g2_fill_2 FILLER_14_496 ();
 sg13g2_decap_4 FILLER_14_503 ();
 sg13g2_decap_8 FILLER_14_534 ();
 sg13g2_fill_1 FILLER_14_541 ();
 sg13g2_fill_2 FILLER_14_597 ();
 sg13g2_decap_4 FILLER_14_625 ();
 sg13g2_fill_1 FILLER_14_629 ();
 sg13g2_decap_8 FILLER_14_656 ();
 sg13g2_decap_8 FILLER_14_663 ();
 sg13g2_decap_8 FILLER_14_670 ();
 sg13g2_decap_8 FILLER_14_677 ();
 sg13g2_decap_8 FILLER_14_684 ();
 sg13g2_decap_8 FILLER_14_691 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_decap_8 FILLER_14_705 ();
 sg13g2_decap_8 FILLER_14_712 ();
 sg13g2_decap_8 FILLER_14_719 ();
 sg13g2_decap_8 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_733 ();
 sg13g2_decap_8 FILLER_14_740 ();
 sg13g2_decap_8 FILLER_14_747 ();
 sg13g2_decap_8 FILLER_14_754 ();
 sg13g2_decap_8 FILLER_14_761 ();
 sg13g2_decap_8 FILLER_14_768 ();
 sg13g2_decap_8 FILLER_14_775 ();
 sg13g2_decap_8 FILLER_14_782 ();
 sg13g2_decap_8 FILLER_14_789 ();
 sg13g2_decap_8 FILLER_14_796 ();
 sg13g2_decap_8 FILLER_14_803 ();
 sg13g2_decap_8 FILLER_14_810 ();
 sg13g2_decap_8 FILLER_14_817 ();
 sg13g2_decap_8 FILLER_14_824 ();
 sg13g2_decap_8 FILLER_14_831 ();
 sg13g2_decap_8 FILLER_14_838 ();
 sg13g2_decap_8 FILLER_14_845 ();
 sg13g2_decap_8 FILLER_14_852 ();
 sg13g2_fill_2 FILLER_14_859 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_83 ();
 sg13g2_fill_2 FILLER_15_95 ();
 sg13g2_fill_1 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_191 ();
 sg13g2_fill_2 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_212 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_fill_2 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_fill_2 FILLER_15_403 ();
 sg13g2_fill_1 FILLER_15_409 ();
 sg13g2_decap_4 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_4 FILLER_15_471 ();
 sg13g2_decap_8 FILLER_15_484 ();
 sg13g2_fill_1 FILLER_15_491 ();
 sg13g2_fill_2 FILLER_15_520 ();
 sg13g2_fill_2 FILLER_15_540 ();
 sg13g2_fill_1 FILLER_15_542 ();
 sg13g2_decap_4 FILLER_15_569 ();
 sg13g2_fill_2 FILLER_15_573 ();
 sg13g2_decap_4 FILLER_15_592 ();
 sg13g2_fill_2 FILLER_15_596 ();
 sg13g2_fill_2 FILLER_15_621 ();
 sg13g2_fill_1 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_647 ();
 sg13g2_decap_8 FILLER_15_654 ();
 sg13g2_decap_8 FILLER_15_661 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_decap_8 FILLER_15_675 ();
 sg13g2_decap_8 FILLER_15_682 ();
 sg13g2_decap_8 FILLER_15_689 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_710 ();
 sg13g2_decap_8 FILLER_15_717 ();
 sg13g2_decap_8 FILLER_15_724 ();
 sg13g2_decap_8 FILLER_15_731 ();
 sg13g2_decap_8 FILLER_15_738 ();
 sg13g2_decap_8 FILLER_15_745 ();
 sg13g2_decap_8 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_759 ();
 sg13g2_decap_8 FILLER_15_766 ();
 sg13g2_decap_8 FILLER_15_773 ();
 sg13g2_decap_8 FILLER_15_780 ();
 sg13g2_decap_8 FILLER_15_787 ();
 sg13g2_decap_8 FILLER_15_794 ();
 sg13g2_decap_8 FILLER_15_801 ();
 sg13g2_decap_8 FILLER_15_808 ();
 sg13g2_decap_8 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_822 ();
 sg13g2_decap_8 FILLER_15_829 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_8 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_4 FILLER_15_857 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_160 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_fill_2 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_258 ();
 sg13g2_fill_2 FILLER_16_284 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_321 ();
 sg13g2_fill_2 FILLER_16_346 ();
 sg13g2_fill_1 FILLER_16_366 ();
 sg13g2_fill_1 FILLER_16_385 ();
 sg13g2_fill_2 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_392 ();
 sg13g2_fill_2 FILLER_16_448 ();
 sg13g2_fill_2 FILLER_16_480 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_fill_2 FILLER_16_521 ();
 sg13g2_fill_1 FILLER_16_523 ();
 sg13g2_fill_2 FILLER_16_550 ();
 sg13g2_decap_8 FILLER_16_570 ();
 sg13g2_fill_2 FILLER_16_577 ();
 sg13g2_decap_8 FILLER_16_589 ();
 sg13g2_fill_1 FILLER_16_596 ();
 sg13g2_fill_2 FILLER_16_649 ();
 sg13g2_decap_8 FILLER_16_660 ();
 sg13g2_decap_8 FILLER_16_667 ();
 sg13g2_decap_8 FILLER_16_674 ();
 sg13g2_decap_8 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_688 ();
 sg13g2_decap_8 FILLER_16_695 ();
 sg13g2_decap_8 FILLER_16_702 ();
 sg13g2_decap_8 FILLER_16_709 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_737 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_decap_8 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_814 ();
 sg13g2_decap_8 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_46 ();
 sg13g2_fill_2 FILLER_17_92 ();
 sg13g2_fill_1 FILLER_17_94 ();
 sg13g2_fill_2 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_fill_2 FILLER_17_157 ();
 sg13g2_fill_1 FILLER_17_159 ();
 sg13g2_fill_2 FILLER_17_164 ();
 sg13g2_fill_2 FILLER_17_184 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_204 ();
 sg13g2_fill_2 FILLER_17_220 ();
 sg13g2_decap_4 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_236 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_fill_1 FILLER_17_311 ();
 sg13g2_fill_2 FILLER_17_333 ();
 sg13g2_fill_2 FILLER_17_364 ();
 sg13g2_fill_1 FILLER_17_395 ();
 sg13g2_fill_2 FILLER_17_422 ();
 sg13g2_fill_1 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_17_430 ();
 sg13g2_fill_2 FILLER_17_437 ();
 sg13g2_fill_1 FILLER_17_439 ();
 sg13g2_fill_2 FILLER_17_462 ();
 sg13g2_fill_1 FILLER_17_464 ();
 sg13g2_decap_4 FILLER_17_473 ();
 sg13g2_fill_2 FILLER_17_485 ();
 sg13g2_fill_1 FILLER_17_487 ();
 sg13g2_fill_1 FILLER_17_506 ();
 sg13g2_decap_4 FILLER_17_521 ();
 sg13g2_fill_2 FILLER_17_525 ();
 sg13g2_fill_2 FILLER_17_536 ();
 sg13g2_fill_1 FILLER_17_538 ();
 sg13g2_decap_8 FILLER_17_544 ();
 sg13g2_decap_4 FILLER_17_597 ();
 sg13g2_fill_1 FILLER_17_601 ();
 sg13g2_decap_8 FILLER_17_620 ();
 sg13g2_decap_4 FILLER_17_627 ();
 sg13g2_fill_1 FILLER_17_631 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_46 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_180 ();
 sg13g2_fill_2 FILLER_18_212 ();
 sg13g2_fill_1 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_279 ();
 sg13g2_decap_4 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_fill_2 FILLER_18_383 ();
 sg13g2_fill_1 FILLER_18_385 ();
 sg13g2_fill_1 FILLER_18_433 ();
 sg13g2_fill_2 FILLER_18_440 ();
 sg13g2_fill_2 FILLER_18_448 ();
 sg13g2_fill_1 FILLER_18_450 ();
 sg13g2_fill_2 FILLER_18_459 ();
 sg13g2_fill_1 FILLER_18_461 ();
 sg13g2_decap_4 FILLER_18_493 ();
 sg13g2_decap_4 FILLER_18_515 ();
 sg13g2_fill_2 FILLER_18_519 ();
 sg13g2_fill_2 FILLER_18_542 ();
 sg13g2_fill_1 FILLER_18_544 ();
 sg13g2_fill_1 FILLER_18_565 ();
 sg13g2_decap_4 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_677 ();
 sg13g2_decap_8 FILLER_18_684 ();
 sg13g2_decap_8 FILLER_18_691 ();
 sg13g2_decap_8 FILLER_18_698 ();
 sg13g2_decap_8 FILLER_18_705 ();
 sg13g2_decap_8 FILLER_18_712 ();
 sg13g2_decap_8 FILLER_18_719 ();
 sg13g2_decap_8 FILLER_18_726 ();
 sg13g2_decap_8 FILLER_18_733 ();
 sg13g2_decap_8 FILLER_18_740 ();
 sg13g2_decap_8 FILLER_18_747 ();
 sg13g2_decap_8 FILLER_18_754 ();
 sg13g2_decap_8 FILLER_18_761 ();
 sg13g2_decap_8 FILLER_18_768 ();
 sg13g2_decap_8 FILLER_18_775 ();
 sg13g2_decap_8 FILLER_18_782 ();
 sg13g2_decap_8 FILLER_18_789 ();
 sg13g2_decap_8 FILLER_18_796 ();
 sg13g2_decap_8 FILLER_18_803 ();
 sg13g2_decap_8 FILLER_18_810 ();
 sg13g2_decap_8 FILLER_18_817 ();
 sg13g2_decap_8 FILLER_18_824 ();
 sg13g2_decap_8 FILLER_18_831 ();
 sg13g2_decap_8 FILLER_18_838 ();
 sg13g2_decap_8 FILLER_18_845 ();
 sg13g2_decap_8 FILLER_18_852 ();
 sg13g2_fill_2 FILLER_18_859 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_39 ();
 sg13g2_fill_1 FILLER_19_67 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_243 ();
 sg13g2_decap_4 FILLER_19_298 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_330 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_fill_2 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_389 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_decap_4 FILLER_19_450 ();
 sg13g2_fill_1 FILLER_19_454 ();
 sg13g2_fill_1 FILLER_19_463 ();
 sg13g2_fill_2 FILLER_19_499 ();
 sg13g2_fill_1 FILLER_19_501 ();
 sg13g2_fill_2 FILLER_19_510 ();
 sg13g2_fill_1 FILLER_19_512 ();
 sg13g2_fill_1 FILLER_19_526 ();
 sg13g2_fill_1 FILLER_19_533 ();
 sg13g2_fill_2 FILLER_19_565 ();
 sg13g2_fill_1 FILLER_19_567 ();
 sg13g2_fill_1 FILLER_19_589 ();
 sg13g2_decap_8 FILLER_19_682 ();
 sg13g2_decap_8 FILLER_19_689 ();
 sg13g2_decap_8 FILLER_19_696 ();
 sg13g2_decap_8 FILLER_19_703 ();
 sg13g2_decap_8 FILLER_19_710 ();
 sg13g2_decap_8 FILLER_19_717 ();
 sg13g2_decap_8 FILLER_19_724 ();
 sg13g2_decap_8 FILLER_19_731 ();
 sg13g2_decap_8 FILLER_19_738 ();
 sg13g2_decap_8 FILLER_19_745 ();
 sg13g2_decap_8 FILLER_19_752 ();
 sg13g2_decap_8 FILLER_19_759 ();
 sg13g2_decap_8 FILLER_19_766 ();
 sg13g2_decap_8 FILLER_19_773 ();
 sg13g2_decap_8 FILLER_19_780 ();
 sg13g2_decap_8 FILLER_19_787 ();
 sg13g2_decap_8 FILLER_19_794 ();
 sg13g2_decap_8 FILLER_19_801 ();
 sg13g2_decap_8 FILLER_19_808 ();
 sg13g2_decap_8 FILLER_19_815 ();
 sg13g2_decap_8 FILLER_19_822 ();
 sg13g2_decap_8 FILLER_19_829 ();
 sg13g2_decap_8 FILLER_19_836 ();
 sg13g2_decap_8 FILLER_19_843 ();
 sg13g2_decap_8 FILLER_19_850 ();
 sg13g2_decap_4 FILLER_19_857 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_4 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_83 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_fill_2 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_345 ();
 sg13g2_decap_4 FILLER_20_387 ();
 sg13g2_decap_4 FILLER_20_457 ();
 sg13g2_decap_8 FILLER_20_479 ();
 sg13g2_decap_4 FILLER_20_486 ();
 sg13g2_fill_1 FILLER_20_490 ();
 sg13g2_fill_2 FILLER_20_513 ();
 sg13g2_fill_1 FILLER_20_515 ();
 sg13g2_decap_4 FILLER_20_522 ();
 sg13g2_fill_2 FILLER_20_539 ();
 sg13g2_fill_2 FILLER_20_545 ();
 sg13g2_fill_2 FILLER_20_578 ();
 sg13g2_fill_2 FILLER_20_590 ();
 sg13g2_fill_2 FILLER_20_624 ();
 sg13g2_fill_2 FILLER_20_645 ();
 sg13g2_fill_1 FILLER_20_647 ();
 sg13g2_decap_8 FILLER_20_678 ();
 sg13g2_decap_8 FILLER_20_685 ();
 sg13g2_decap_8 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_699 ();
 sg13g2_decap_8 FILLER_20_706 ();
 sg13g2_decap_8 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_720 ();
 sg13g2_decap_8 FILLER_20_727 ();
 sg13g2_decap_8 FILLER_20_734 ();
 sg13g2_decap_8 FILLER_20_741 ();
 sg13g2_decap_8 FILLER_20_748 ();
 sg13g2_decap_8 FILLER_20_755 ();
 sg13g2_decap_8 FILLER_20_762 ();
 sg13g2_decap_8 FILLER_20_769 ();
 sg13g2_decap_8 FILLER_20_776 ();
 sg13g2_decap_8 FILLER_20_783 ();
 sg13g2_decap_8 FILLER_20_790 ();
 sg13g2_decap_8 FILLER_20_797 ();
 sg13g2_decap_8 FILLER_20_804 ();
 sg13g2_decap_8 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_818 ();
 sg13g2_decap_8 FILLER_20_825 ();
 sg13g2_decap_8 FILLER_20_832 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_214 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_2 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_4 FILLER_21_312 ();
 sg13g2_decap_4 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_fill_2 FILLER_21_431 ();
 sg13g2_fill_1 FILLER_21_433 ();
 sg13g2_decap_4 FILLER_21_438 ();
 sg13g2_fill_2 FILLER_21_446 ();
 sg13g2_decap_4 FILLER_21_456 ();
 sg13g2_fill_1 FILLER_21_460 ();
 sg13g2_fill_2 FILLER_21_512 ();
 sg13g2_fill_1 FILLER_21_514 ();
 sg13g2_fill_2 FILLER_21_550 ();
 sg13g2_fill_1 FILLER_21_552 ();
 sg13g2_decap_8 FILLER_21_671 ();
 sg13g2_decap_8 FILLER_21_678 ();
 sg13g2_decap_8 FILLER_21_685 ();
 sg13g2_decap_8 FILLER_21_692 ();
 sg13g2_decap_8 FILLER_21_699 ();
 sg13g2_decap_8 FILLER_21_706 ();
 sg13g2_decap_8 FILLER_21_713 ();
 sg13g2_decap_8 FILLER_21_720 ();
 sg13g2_decap_8 FILLER_21_727 ();
 sg13g2_decap_8 FILLER_21_734 ();
 sg13g2_decap_8 FILLER_21_741 ();
 sg13g2_decap_8 FILLER_21_748 ();
 sg13g2_decap_8 FILLER_21_755 ();
 sg13g2_decap_8 FILLER_21_762 ();
 sg13g2_decap_8 FILLER_21_769 ();
 sg13g2_decap_8 FILLER_21_776 ();
 sg13g2_decap_8 FILLER_21_783 ();
 sg13g2_decap_8 FILLER_21_790 ();
 sg13g2_decap_8 FILLER_21_797 ();
 sg13g2_decap_8 FILLER_21_804 ();
 sg13g2_decap_8 FILLER_21_811 ();
 sg13g2_decap_8 FILLER_21_818 ();
 sg13g2_decap_8 FILLER_21_825 ();
 sg13g2_decap_8 FILLER_21_832 ();
 sg13g2_decap_8 FILLER_21_839 ();
 sg13g2_decap_8 FILLER_21_846 ();
 sg13g2_decap_8 FILLER_21_853 ();
 sg13g2_fill_2 FILLER_21_860 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_62 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_fill_2 FILLER_22_92 ();
 sg13g2_fill_1 FILLER_22_94 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_122 ();
 sg13g2_decap_4 FILLER_22_129 ();
 sg13g2_fill_1 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_145 ();
 sg13g2_fill_1 FILLER_22_156 ();
 sg13g2_decap_4 FILLER_22_175 ();
 sg13g2_fill_1 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_fill_1 FILLER_22_216 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_fill_2 FILLER_22_414 ();
 sg13g2_fill_2 FILLER_22_471 ();
 sg13g2_decap_4 FILLER_22_538 ();
 sg13g2_fill_2 FILLER_22_542 ();
 sg13g2_decap_8 FILLER_22_570 ();
 sg13g2_decap_4 FILLER_22_577 ();
 sg13g2_fill_1 FILLER_22_599 ();
 sg13g2_fill_1 FILLER_22_619 ();
 sg13g2_fill_2 FILLER_22_633 ();
 sg13g2_decap_8 FILLER_22_663 ();
 sg13g2_decap_8 FILLER_22_670 ();
 sg13g2_decap_8 FILLER_22_677 ();
 sg13g2_decap_8 FILLER_22_684 ();
 sg13g2_decap_8 FILLER_22_691 ();
 sg13g2_decap_8 FILLER_22_698 ();
 sg13g2_decap_8 FILLER_22_705 ();
 sg13g2_decap_8 FILLER_22_712 ();
 sg13g2_decap_8 FILLER_22_719 ();
 sg13g2_decap_8 FILLER_22_726 ();
 sg13g2_decap_8 FILLER_22_733 ();
 sg13g2_decap_8 FILLER_22_740 ();
 sg13g2_decap_8 FILLER_22_747 ();
 sg13g2_decap_8 FILLER_22_754 ();
 sg13g2_decap_8 FILLER_22_761 ();
 sg13g2_decap_8 FILLER_22_768 ();
 sg13g2_decap_8 FILLER_22_775 ();
 sg13g2_decap_8 FILLER_22_782 ();
 sg13g2_decap_8 FILLER_22_789 ();
 sg13g2_decap_8 FILLER_22_796 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_decap_8 FILLER_22_810 ();
 sg13g2_decap_8 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_decap_8 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_838 ();
 sg13g2_decap_8 FILLER_22_845 ();
 sg13g2_decap_8 FILLER_22_852 ();
 sg13g2_fill_2 FILLER_22_859 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_fill_2 FILLER_23_160 ();
 sg13g2_fill_1 FILLER_23_162 ();
 sg13g2_fill_1 FILLER_23_188 ();
 sg13g2_fill_2 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_fill_2 FILLER_23_202 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_fill_2 FILLER_23_228 ();
 sg13g2_fill_1 FILLER_23_230 ();
 sg13g2_decap_4 FILLER_23_250 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_decap_4 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_441 ();
 sg13g2_fill_1 FILLER_23_443 ();
 sg13g2_decap_8 FILLER_23_456 ();
 sg13g2_decap_4 FILLER_23_463 ();
 sg13g2_fill_1 FILLER_23_467 ();
 sg13g2_fill_1 FILLER_23_476 ();
 sg13g2_fill_1 FILLER_23_513 ();
 sg13g2_fill_1 FILLER_23_526 ();
 sg13g2_fill_2 FILLER_23_548 ();
 sg13g2_decap_4 FILLER_23_571 ();
 sg13g2_fill_2 FILLER_23_575 ();
 sg13g2_fill_2 FILLER_23_592 ();
 sg13g2_fill_1 FILLER_23_594 ();
 sg13g2_fill_2 FILLER_23_637 ();
 sg13g2_fill_1 FILLER_23_639 ();
 sg13g2_decap_8 FILLER_23_666 ();
 sg13g2_decap_8 FILLER_23_673 ();
 sg13g2_decap_8 FILLER_23_680 ();
 sg13g2_decap_8 FILLER_23_687 ();
 sg13g2_decap_8 FILLER_23_694 ();
 sg13g2_decap_8 FILLER_23_701 ();
 sg13g2_decap_8 FILLER_23_708 ();
 sg13g2_decap_8 FILLER_23_715 ();
 sg13g2_decap_8 FILLER_23_722 ();
 sg13g2_decap_8 FILLER_23_729 ();
 sg13g2_decap_8 FILLER_23_736 ();
 sg13g2_decap_8 FILLER_23_743 ();
 sg13g2_decap_8 FILLER_23_750 ();
 sg13g2_decap_8 FILLER_23_757 ();
 sg13g2_decap_8 FILLER_23_764 ();
 sg13g2_decap_8 FILLER_23_771 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_decap_8 FILLER_23_785 ();
 sg13g2_decap_8 FILLER_23_792 ();
 sg13g2_decap_8 FILLER_23_799 ();
 sg13g2_decap_8 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_813 ();
 sg13g2_decap_8 FILLER_23_820 ();
 sg13g2_decap_8 FILLER_23_827 ();
 sg13g2_decap_8 FILLER_23_834 ();
 sg13g2_decap_8 FILLER_23_841 ();
 sg13g2_decap_8 FILLER_23_848 ();
 sg13g2_decap_8 FILLER_23_855 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_94 ();
 sg13g2_fill_2 FILLER_24_110 ();
 sg13g2_decap_4 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_decap_8 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_262 ();
 sg13g2_decap_8 FILLER_24_269 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_302 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_310 ();
 sg13g2_fill_1 FILLER_24_324 ();
 sg13g2_decap_4 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_decap_4 FILLER_24_455 ();
 sg13g2_fill_1 FILLER_24_459 ();
 sg13g2_fill_2 FILLER_24_486 ();
 sg13g2_fill_2 FILLER_24_510 ();
 sg13g2_fill_1 FILLER_24_512 ();
 sg13g2_decap_4 FILLER_24_542 ();
 sg13g2_fill_1 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_570 ();
 sg13g2_fill_1 FILLER_24_587 ();
 sg13g2_decap_8 FILLER_24_667 ();
 sg13g2_decap_8 FILLER_24_674 ();
 sg13g2_decap_8 FILLER_24_681 ();
 sg13g2_decap_8 FILLER_24_688 ();
 sg13g2_decap_8 FILLER_24_695 ();
 sg13g2_decap_8 FILLER_24_702 ();
 sg13g2_decap_8 FILLER_24_709 ();
 sg13g2_decap_8 FILLER_24_716 ();
 sg13g2_decap_8 FILLER_24_723 ();
 sg13g2_decap_8 FILLER_24_730 ();
 sg13g2_decap_8 FILLER_24_737 ();
 sg13g2_decap_8 FILLER_24_744 ();
 sg13g2_decap_8 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_758 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_8 FILLER_24_772 ();
 sg13g2_decap_8 FILLER_24_779 ();
 sg13g2_decap_8 FILLER_24_786 ();
 sg13g2_decap_8 FILLER_24_793 ();
 sg13g2_decap_8 FILLER_24_800 ();
 sg13g2_decap_8 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_814 ();
 sg13g2_decap_8 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_decap_8 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_842 ();
 sg13g2_decap_8 FILLER_24_849 ();
 sg13g2_decap_4 FILLER_24_856 ();
 sg13g2_fill_2 FILLER_24_860 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_fill_2 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_79 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_decap_4 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_184 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_4 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_218 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_387 ();
 sg13g2_fill_2 FILLER_25_416 ();
 sg13g2_fill_1 FILLER_25_418 ();
 sg13g2_fill_2 FILLER_25_429 ();
 sg13g2_fill_1 FILLER_25_431 ();
 sg13g2_fill_2 FILLER_25_445 ();
 sg13g2_fill_1 FILLER_25_464 ();
 sg13g2_fill_2 FILLER_25_470 ();
 sg13g2_fill_1 FILLER_25_472 ();
 sg13g2_decap_4 FILLER_25_538 ();
 sg13g2_fill_1 FILLER_25_542 ();
 sg13g2_decap_4 FILLER_25_551 ();
 sg13g2_decap_8 FILLER_25_579 ();
 sg13g2_fill_1 FILLER_25_591 ();
 sg13g2_fill_1 FILLER_25_621 ();
 sg13g2_decap_8 FILLER_25_662 ();
 sg13g2_decap_8 FILLER_25_669 ();
 sg13g2_decap_8 FILLER_25_676 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_8 FILLER_25_690 ();
 sg13g2_decap_8 FILLER_25_697 ();
 sg13g2_decap_8 FILLER_25_704 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_8 FILLER_25_718 ();
 sg13g2_decap_8 FILLER_25_725 ();
 sg13g2_decap_8 FILLER_25_732 ();
 sg13g2_decap_8 FILLER_25_739 ();
 sg13g2_decap_8 FILLER_25_746 ();
 sg13g2_decap_8 FILLER_25_753 ();
 sg13g2_decap_8 FILLER_25_760 ();
 sg13g2_decap_8 FILLER_25_767 ();
 sg13g2_decap_8 FILLER_25_774 ();
 sg13g2_decap_8 FILLER_25_781 ();
 sg13g2_decap_8 FILLER_25_788 ();
 sg13g2_decap_8 FILLER_25_795 ();
 sg13g2_decap_8 FILLER_25_802 ();
 sg13g2_decap_8 FILLER_25_809 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_823 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_4 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_90 ();
 sg13g2_fill_1 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_decap_4 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_fill_2 FILLER_26_369 ();
 sg13g2_fill_2 FILLER_26_485 ();
 sg13g2_decap_8 FILLER_26_556 ();
 sg13g2_decap_8 FILLER_26_568 ();
 sg13g2_fill_1 FILLER_26_575 ();
 sg13g2_decap_4 FILLER_26_612 ();
 sg13g2_fill_2 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_654 ();
 sg13g2_decap_8 FILLER_26_661 ();
 sg13g2_decap_8 FILLER_26_668 ();
 sg13g2_decap_8 FILLER_26_675 ();
 sg13g2_decap_8 FILLER_26_682 ();
 sg13g2_decap_8 FILLER_26_689 ();
 sg13g2_decap_8 FILLER_26_696 ();
 sg13g2_decap_8 FILLER_26_703 ();
 sg13g2_decap_8 FILLER_26_710 ();
 sg13g2_decap_8 FILLER_26_717 ();
 sg13g2_decap_8 FILLER_26_724 ();
 sg13g2_decap_8 FILLER_26_731 ();
 sg13g2_decap_8 FILLER_26_738 ();
 sg13g2_decap_8 FILLER_26_745 ();
 sg13g2_decap_8 FILLER_26_752 ();
 sg13g2_decap_8 FILLER_26_759 ();
 sg13g2_decap_8 FILLER_26_766 ();
 sg13g2_decap_8 FILLER_26_773 ();
 sg13g2_decap_8 FILLER_26_780 ();
 sg13g2_decap_8 FILLER_26_787 ();
 sg13g2_decap_8 FILLER_26_794 ();
 sg13g2_decap_8 FILLER_26_801 ();
 sg13g2_decap_8 FILLER_26_808 ();
 sg13g2_decap_8 FILLER_26_815 ();
 sg13g2_decap_8 FILLER_26_822 ();
 sg13g2_decap_8 FILLER_26_829 ();
 sg13g2_decap_8 FILLER_26_836 ();
 sg13g2_decap_8 FILLER_26_843 ();
 sg13g2_decap_8 FILLER_26_850 ();
 sg13g2_decap_4 FILLER_26_857 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_93 ();
 sg13g2_fill_2 FILLER_27_130 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_decap_4 FILLER_27_272 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_fill_1 FILLER_27_388 ();
 sg13g2_decap_4 FILLER_27_417 ();
 sg13g2_fill_2 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_431 ();
 sg13g2_fill_1 FILLER_27_433 ();
 sg13g2_fill_1 FILLER_27_460 ();
 sg13g2_fill_2 FILLER_27_469 ();
 sg13g2_fill_1 FILLER_27_471 ();
 sg13g2_fill_2 FILLER_27_477 ();
 sg13g2_fill_1 FILLER_27_479 ();
 sg13g2_fill_2 FILLER_27_499 ();
 sg13g2_fill_1 FILLER_27_519 ();
 sg13g2_fill_2 FILLER_27_525 ();
 sg13g2_decap_4 FILLER_27_559 ();
 sg13g2_fill_1 FILLER_27_563 ();
 sg13g2_fill_1 FILLER_27_594 ();
 sg13g2_decap_8 FILLER_27_631 ();
 sg13g2_fill_2 FILLER_27_638 ();
 sg13g2_decap_8 FILLER_27_649 ();
 sg13g2_decap_8 FILLER_27_656 ();
 sg13g2_decap_8 FILLER_27_663 ();
 sg13g2_decap_8 FILLER_27_670 ();
 sg13g2_decap_8 FILLER_27_677 ();
 sg13g2_decap_8 FILLER_27_684 ();
 sg13g2_decap_8 FILLER_27_691 ();
 sg13g2_decap_8 FILLER_27_698 ();
 sg13g2_decap_8 FILLER_27_705 ();
 sg13g2_decap_8 FILLER_27_712 ();
 sg13g2_decap_8 FILLER_27_719 ();
 sg13g2_decap_8 FILLER_27_726 ();
 sg13g2_decap_8 FILLER_27_733 ();
 sg13g2_decap_8 FILLER_27_740 ();
 sg13g2_decap_8 FILLER_27_747 ();
 sg13g2_decap_8 FILLER_27_754 ();
 sg13g2_decap_8 FILLER_27_761 ();
 sg13g2_decap_8 FILLER_27_768 ();
 sg13g2_decap_8 FILLER_27_775 ();
 sg13g2_decap_8 FILLER_27_782 ();
 sg13g2_decap_8 FILLER_27_789 ();
 sg13g2_decap_8 FILLER_27_796 ();
 sg13g2_decap_8 FILLER_27_803 ();
 sg13g2_decap_8 FILLER_27_810 ();
 sg13g2_decap_8 FILLER_27_817 ();
 sg13g2_decap_8 FILLER_27_824 ();
 sg13g2_decap_8 FILLER_27_831 ();
 sg13g2_decap_8 FILLER_27_838 ();
 sg13g2_decap_8 FILLER_27_845 ();
 sg13g2_decap_8 FILLER_27_852 ();
 sg13g2_fill_2 FILLER_27_859 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_159 ();
 sg13g2_decap_4 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_fill_2 FILLER_28_252 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_decap_4 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_356 ();
 sg13g2_decap_4 FILLER_28_395 ();
 sg13g2_fill_2 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_405 ();
 sg13g2_fill_1 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_28_477 ();
 sg13g2_fill_1 FILLER_28_479 ();
 sg13g2_fill_2 FILLER_28_515 ();
 sg13g2_fill_2 FILLER_28_522 ();
 sg13g2_fill_1 FILLER_28_568 ();
 sg13g2_decap_8 FILLER_28_590 ();
 sg13g2_fill_2 FILLER_28_601 ();
 sg13g2_decap_4 FILLER_28_612 ();
 sg13g2_decap_8 FILLER_28_620 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_decap_8 FILLER_28_634 ();
 sg13g2_decap_8 FILLER_28_641 ();
 sg13g2_decap_8 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_655 ();
 sg13g2_decap_8 FILLER_28_662 ();
 sg13g2_decap_8 FILLER_28_669 ();
 sg13g2_decap_8 FILLER_28_676 ();
 sg13g2_decap_8 FILLER_28_683 ();
 sg13g2_decap_8 FILLER_28_690 ();
 sg13g2_decap_8 FILLER_28_697 ();
 sg13g2_decap_8 FILLER_28_704 ();
 sg13g2_decap_8 FILLER_28_711 ();
 sg13g2_decap_8 FILLER_28_718 ();
 sg13g2_decap_8 FILLER_28_725 ();
 sg13g2_decap_8 FILLER_28_732 ();
 sg13g2_decap_8 FILLER_28_739 ();
 sg13g2_decap_8 FILLER_28_746 ();
 sg13g2_decap_8 FILLER_28_753 ();
 sg13g2_decap_8 FILLER_28_760 ();
 sg13g2_decap_8 FILLER_28_767 ();
 sg13g2_decap_8 FILLER_28_774 ();
 sg13g2_decap_8 FILLER_28_781 ();
 sg13g2_decap_8 FILLER_28_788 ();
 sg13g2_decap_8 FILLER_28_795 ();
 sg13g2_decap_8 FILLER_28_802 ();
 sg13g2_decap_8 FILLER_28_809 ();
 sg13g2_decap_8 FILLER_28_816 ();
 sg13g2_decap_8 FILLER_28_823 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_decap_4 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_decap_4 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_decap_4 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_decap_4 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_321 ();
 sg13g2_fill_2 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_fill_2 FILLER_29_458 ();
 sg13g2_fill_1 FILLER_29_460 ();
 sg13g2_fill_2 FILLER_29_477 ();
 sg13g2_fill_2 FILLER_29_520 ();
 sg13g2_fill_2 FILLER_29_559 ();
 sg13g2_decap_8 FILLER_29_587 ();
 sg13g2_decap_8 FILLER_29_594 ();
 sg13g2_decap_8 FILLER_29_611 ();
 sg13g2_decap_8 FILLER_29_618 ();
 sg13g2_decap_8 FILLER_29_625 ();
 sg13g2_decap_8 FILLER_29_632 ();
 sg13g2_decap_8 FILLER_29_639 ();
 sg13g2_decap_8 FILLER_29_646 ();
 sg13g2_decap_8 FILLER_29_653 ();
 sg13g2_decap_8 FILLER_29_660 ();
 sg13g2_decap_8 FILLER_29_667 ();
 sg13g2_decap_8 FILLER_29_674 ();
 sg13g2_decap_8 FILLER_29_681 ();
 sg13g2_decap_8 FILLER_29_688 ();
 sg13g2_decap_8 FILLER_29_695 ();
 sg13g2_decap_8 FILLER_29_702 ();
 sg13g2_decap_8 FILLER_29_709 ();
 sg13g2_decap_8 FILLER_29_716 ();
 sg13g2_decap_8 FILLER_29_723 ();
 sg13g2_decap_8 FILLER_29_730 ();
 sg13g2_decap_8 FILLER_29_737 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_decap_8 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_758 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_8 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_8 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_828 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_842 ();
 sg13g2_decap_8 FILLER_29_849 ();
 sg13g2_decap_4 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_decap_4 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_decap_4 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_decap_4 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_409 ();
 sg13g2_fill_1 FILLER_30_416 ();
 sg13g2_decap_8 FILLER_30_458 ();
 sg13g2_fill_2 FILLER_30_509 ();
 sg13g2_fill_1 FILLER_30_552 ();
 sg13g2_decap_4 FILLER_30_579 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_fill_2 FILLER_31_256 ();
 sg13g2_decap_4 FILLER_31_273 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_decap_4 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_fill_2 FILLER_31_403 ();
 sg13g2_fill_1 FILLER_31_419 ();
 sg13g2_decap_8 FILLER_31_458 ();
 sg13g2_fill_1 FILLER_31_469 ();
 sg13g2_fill_1 FILLER_31_480 ();
 sg13g2_fill_1 FILLER_31_530 ();
 sg13g2_fill_2 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_603 ();
 sg13g2_decap_8 FILLER_31_610 ();
 sg13g2_decap_8 FILLER_31_617 ();
 sg13g2_decap_8 FILLER_31_624 ();
 sg13g2_decap_8 FILLER_31_631 ();
 sg13g2_decap_4 FILLER_31_638 ();
 sg13g2_decap_8 FILLER_31_668 ();
 sg13g2_decap_8 FILLER_31_675 ();
 sg13g2_decap_8 FILLER_31_682 ();
 sg13g2_decap_8 FILLER_31_689 ();
 sg13g2_decap_8 FILLER_31_696 ();
 sg13g2_decap_8 FILLER_31_703 ();
 sg13g2_decap_8 FILLER_31_710 ();
 sg13g2_decap_8 FILLER_31_717 ();
 sg13g2_decap_8 FILLER_31_724 ();
 sg13g2_decap_8 FILLER_31_731 ();
 sg13g2_decap_8 FILLER_31_738 ();
 sg13g2_decap_8 FILLER_31_745 ();
 sg13g2_decap_8 FILLER_31_752 ();
 sg13g2_decap_8 FILLER_31_759 ();
 sg13g2_decap_8 FILLER_31_766 ();
 sg13g2_decap_8 FILLER_31_773 ();
 sg13g2_decap_8 FILLER_31_780 ();
 sg13g2_decap_8 FILLER_31_787 ();
 sg13g2_decap_8 FILLER_31_794 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_decap_8 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_4 FILLER_31_857 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_4 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_decap_4 FILLER_32_202 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_decap_4 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_decap_4 FILLER_32_325 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_decap_4 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_decap_4 FILLER_32_397 ();
 sg13g2_fill_2 FILLER_32_411 ();
 sg13g2_fill_2 FILLER_32_443 ();
 sg13g2_fill_2 FILLER_32_457 ();
 sg13g2_decap_4 FILLER_32_483 ();
 sg13g2_fill_1 FILLER_32_487 ();
 sg13g2_decap_4 FILLER_32_508 ();
 sg13g2_fill_1 FILLER_32_512 ();
 sg13g2_fill_2 FILLER_32_558 ();
 sg13g2_decap_8 FILLER_32_603 ();
 sg13g2_decap_4 FILLER_32_610 ();
 sg13g2_fill_1 FILLER_32_614 ();
 sg13g2_decap_4 FILLER_32_622 ();
 sg13g2_fill_1 FILLER_32_626 ();
 sg13g2_decap_8 FILLER_32_653 ();
 sg13g2_fill_2 FILLER_32_660 ();
 sg13g2_fill_1 FILLER_32_662 ();
 sg13g2_fill_2 FILLER_32_667 ();
 sg13g2_fill_1 FILLER_32_669 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_8 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_4 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_144 ();
 sg13g2_fill_2 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_decap_8 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_2 FILLER_33_395 ();
 sg13g2_decap_4 FILLER_33_418 ();
 sg13g2_fill_1 FILLER_33_439 ();
 sg13g2_fill_1 FILLER_33_449 ();
 sg13g2_decap_4 FILLER_33_471 ();
 sg13g2_fill_1 FILLER_33_475 ();
 sg13g2_fill_1 FILLER_33_479 ();
 sg13g2_decap_8 FILLER_33_485 ();
 sg13g2_decap_4 FILLER_33_492 ();
 sg13g2_fill_2 FILLER_33_496 ();
 sg13g2_decap_4 FILLER_33_516 ();
 sg13g2_fill_2 FILLER_33_520 ();
 sg13g2_decap_8 FILLER_33_527 ();
 sg13g2_fill_2 FILLER_33_534 ();
 sg13g2_fill_1 FILLER_33_545 ();
 sg13g2_fill_2 FILLER_33_563 ();
 sg13g2_decap_4 FILLER_33_588 ();
 sg13g2_fill_1 FILLER_33_605 ();
 sg13g2_fill_1 FILLER_33_632 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_fill_2 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_685 ();
 sg13g2_decap_8 FILLER_33_692 ();
 sg13g2_decap_8 FILLER_33_699 ();
 sg13g2_decap_8 FILLER_33_706 ();
 sg13g2_decap_8 FILLER_33_713 ();
 sg13g2_decap_8 FILLER_33_720 ();
 sg13g2_decap_8 FILLER_33_727 ();
 sg13g2_decap_8 FILLER_33_734 ();
 sg13g2_decap_8 FILLER_33_741 ();
 sg13g2_decap_8 FILLER_33_748 ();
 sg13g2_decap_8 FILLER_33_755 ();
 sg13g2_decap_8 FILLER_33_762 ();
 sg13g2_decap_8 FILLER_33_769 ();
 sg13g2_decap_8 FILLER_33_776 ();
 sg13g2_decap_8 FILLER_33_783 ();
 sg13g2_decap_8 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_797 ();
 sg13g2_decap_8 FILLER_33_804 ();
 sg13g2_decap_8 FILLER_33_811 ();
 sg13g2_decap_8 FILLER_33_818 ();
 sg13g2_decap_8 FILLER_33_825 ();
 sg13g2_decap_8 FILLER_33_832 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_decap_8 FILLER_33_846 ();
 sg13g2_decap_8 FILLER_33_853 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_decap_4 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_4 FILLER_34_386 ();
 sg13g2_fill_2 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_8 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_411 ();
 sg13g2_decap_4 FILLER_34_417 ();
 sg13g2_fill_2 FILLER_34_424 ();
 sg13g2_fill_1 FILLER_34_426 ();
 sg13g2_decap_4 FILLER_34_441 ();
 sg13g2_fill_2 FILLER_34_445 ();
 sg13g2_fill_2 FILLER_34_474 ();
 sg13g2_fill_1 FILLER_34_480 ();
 sg13g2_fill_1 FILLER_34_507 ();
 sg13g2_fill_2 FILLER_34_526 ();
 sg13g2_fill_1 FILLER_34_528 ();
 sg13g2_fill_1 FILLER_34_542 ();
 sg13g2_decap_8 FILLER_34_548 ();
 sg13g2_decap_4 FILLER_34_564 ();
 sg13g2_decap_4 FILLER_34_573 ();
 sg13g2_fill_2 FILLER_34_587 ();
 sg13g2_fill_2 FILLER_34_611 ();
 sg13g2_fill_1 FILLER_34_613 ();
 sg13g2_fill_2 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_647 ();
 sg13g2_decap_4 FILLER_34_654 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_fill_2 FILLER_34_700 ();
 sg13g2_fill_1 FILLER_34_702 ();
 sg13g2_decap_8 FILLER_34_706 ();
 sg13g2_decap_8 FILLER_34_713 ();
 sg13g2_decap_8 FILLER_34_720 ();
 sg13g2_decap_8 FILLER_34_727 ();
 sg13g2_decap_8 FILLER_34_734 ();
 sg13g2_decap_8 FILLER_34_741 ();
 sg13g2_decap_8 FILLER_34_748 ();
 sg13g2_decap_8 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_762 ();
 sg13g2_decap_8 FILLER_34_769 ();
 sg13g2_decap_8 FILLER_34_776 ();
 sg13g2_decap_8 FILLER_34_783 ();
 sg13g2_decap_8 FILLER_34_790 ();
 sg13g2_decap_8 FILLER_34_797 ();
 sg13g2_decap_8 FILLER_34_804 ();
 sg13g2_decap_8 FILLER_34_811 ();
 sg13g2_decap_8 FILLER_34_818 ();
 sg13g2_decap_8 FILLER_34_825 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_fill_2 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_105 ();
 sg13g2_fill_1 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_fill_2 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_decap_4 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_decap_4 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_350 ();
 sg13g2_decap_4 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_4 FILLER_35_412 ();
 sg13g2_fill_2 FILLER_35_416 ();
 sg13g2_decap_4 FILLER_35_435 ();
 sg13g2_fill_2 FILLER_35_448 ();
 sg13g2_fill_1 FILLER_35_450 ();
 sg13g2_fill_2 FILLER_35_455 ();
 sg13g2_decap_4 FILLER_35_467 ();
 sg13g2_fill_1 FILLER_35_475 ();
 sg13g2_fill_1 FILLER_35_485 ();
 sg13g2_decap_4 FILLER_35_490 ();
 sg13g2_fill_1 FILLER_35_494 ();
 sg13g2_fill_1 FILLER_35_500 ();
 sg13g2_fill_2 FILLER_35_514 ();
 sg13g2_fill_1 FILLER_35_556 ();
 sg13g2_fill_2 FILLER_35_570 ();
 sg13g2_fill_1 FILLER_35_572 ();
 sg13g2_fill_2 FILLER_35_602 ();
 sg13g2_fill_2 FILLER_35_608 ();
 sg13g2_decap_4 FILLER_35_646 ();
 sg13g2_decap_4 FILLER_35_654 ();
 sg13g2_fill_2 FILLER_35_681 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_88 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_292 ();
 sg13g2_fill_1 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_decap_4 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_340 ();
 sg13g2_decap_4 FILLER_36_356 ();
 sg13g2_fill_1 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_386 ();
 sg13g2_fill_1 FILLER_36_409 ();
 sg13g2_decap_8 FILLER_36_437 ();
 sg13g2_decap_4 FILLER_36_444 ();
 sg13g2_fill_1 FILLER_36_448 ();
 sg13g2_fill_2 FILLER_36_465 ();
 sg13g2_fill_2 FILLER_36_485 ();
 sg13g2_decap_4 FILLER_36_518 ();
 sg13g2_fill_2 FILLER_36_540 ();
 sg13g2_fill_1 FILLER_36_542 ();
 sg13g2_fill_2 FILLER_36_567 ();
 sg13g2_fill_1 FILLER_36_569 ();
 sg13g2_decap_8 FILLER_36_591 ();
 sg13g2_fill_2 FILLER_36_626 ();
 sg13g2_fill_1 FILLER_36_628 ();
 sg13g2_decap_4 FILLER_36_642 ();
 sg13g2_fill_2 FILLER_36_646 ();
 sg13g2_fill_1 FILLER_36_651 ();
 sg13g2_fill_1 FILLER_36_657 ();
 sg13g2_fill_2 FILLER_36_683 ();
 sg13g2_fill_1 FILLER_36_685 ();
 sg13g2_decap_8 FILLER_36_695 ();
 sg13g2_decap_8 FILLER_36_721 ();
 sg13g2_decap_8 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_742 ();
 sg13g2_decap_8 FILLER_36_749 ();
 sg13g2_decap_8 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_decap_8 FILLER_36_770 ();
 sg13g2_decap_8 FILLER_36_777 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_decap_8 FILLER_36_791 ();
 sg13g2_decap_8 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_812 ();
 sg13g2_decap_8 FILLER_36_819 ();
 sg13g2_decap_8 FILLER_36_826 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_decap_8 FILLER_36_854 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_65 ();
 sg13g2_fill_2 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_decap_4 FILLER_37_298 ();
 sg13g2_decap_4 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_decap_4 FILLER_37_395 ();
 sg13g2_fill_1 FILLER_37_399 ();
 sg13g2_decap_4 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_429 ();
 sg13g2_fill_2 FILLER_37_436 ();
 sg13g2_fill_1 FILLER_37_438 ();
 sg13g2_fill_2 FILLER_37_461 ();
 sg13g2_decap_8 FILLER_37_491 ();
 sg13g2_fill_2 FILLER_37_498 ();
 sg13g2_fill_1 FILLER_37_500 ();
 sg13g2_fill_1 FILLER_37_516 ();
 sg13g2_decap_8 FILLER_37_529 ();
 sg13g2_fill_1 FILLER_37_536 ();
 sg13g2_fill_1 FILLER_37_542 ();
 sg13g2_fill_1 FILLER_37_566 ();
 sg13g2_decap_8 FILLER_37_586 ();
 sg13g2_fill_2 FILLER_37_593 ();
 sg13g2_decap_8 FILLER_37_600 ();
 sg13g2_fill_2 FILLER_37_607 ();
 sg13g2_fill_1 FILLER_37_628 ();
 sg13g2_fill_1 FILLER_37_690 ();
 sg13g2_decap_8 FILLER_37_717 ();
 sg13g2_decap_8 FILLER_37_724 ();
 sg13g2_decap_8 FILLER_37_731 ();
 sg13g2_decap_8 FILLER_37_738 ();
 sg13g2_decap_8 FILLER_37_745 ();
 sg13g2_decap_8 FILLER_37_752 ();
 sg13g2_decap_8 FILLER_37_759 ();
 sg13g2_decap_8 FILLER_37_766 ();
 sg13g2_decap_8 FILLER_37_773 ();
 sg13g2_decap_8 FILLER_37_780 ();
 sg13g2_decap_8 FILLER_37_787 ();
 sg13g2_decap_8 FILLER_37_794 ();
 sg13g2_decap_8 FILLER_37_801 ();
 sg13g2_decap_8 FILLER_37_808 ();
 sg13g2_decap_8 FILLER_37_815 ();
 sg13g2_decap_8 FILLER_37_822 ();
 sg13g2_decap_8 FILLER_37_829 ();
 sg13g2_decap_8 FILLER_37_836 ();
 sg13g2_decap_8 FILLER_37_843 ();
 sg13g2_decap_8 FILLER_37_850 ();
 sg13g2_decap_4 FILLER_37_857 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_101 ();
 sg13g2_fill_1 FILLER_38_111 ();
 sg13g2_decap_4 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_240 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_269 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_4 FILLER_38_292 ();
 sg13g2_decap_4 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_decap_4 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_315 ();
 sg13g2_fill_2 FILLER_38_335 ();
 sg13g2_fill_1 FILLER_38_337 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_fill_2 FILLER_38_354 ();
 sg13g2_fill_1 FILLER_38_376 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_fill_2 FILLER_38_391 ();
 sg13g2_fill_1 FILLER_38_393 ();
 sg13g2_decap_4 FILLER_38_413 ();
 sg13g2_fill_2 FILLER_38_417 ();
 sg13g2_decap_4 FILLER_38_430 ();
 sg13g2_fill_1 FILLER_38_434 ();
 sg13g2_fill_1 FILLER_38_440 ();
 sg13g2_decap_8 FILLER_38_463 ();
 sg13g2_fill_2 FILLER_38_479 ();
 sg13g2_decap_8 FILLER_38_486 ();
 sg13g2_decap_8 FILLER_38_493 ();
 sg13g2_fill_1 FILLER_38_500 ();
 sg13g2_decap_4 FILLER_38_519 ();
 sg13g2_fill_1 FILLER_38_523 ();
 sg13g2_decap_8 FILLER_38_528 ();
 sg13g2_fill_1 FILLER_38_535 ();
 sg13g2_fill_1 FILLER_38_563 ();
 sg13g2_fill_1 FILLER_38_576 ();
 sg13g2_fill_2 FILLER_38_587 ();
 sg13g2_fill_1 FILLER_38_589 ();
 sg13g2_fill_2 FILLER_38_596 ();
 sg13g2_fill_1 FILLER_38_598 ();
 sg13g2_fill_1 FILLER_38_604 ();
 sg13g2_fill_2 FILLER_38_626 ();
 sg13g2_fill_1 FILLER_38_628 ();
 sg13g2_decap_4 FILLER_38_639 ();
 sg13g2_fill_2 FILLER_38_643 ();
 sg13g2_fill_1 FILLER_38_668 ();
 sg13g2_fill_2 FILLER_38_677 ();
 sg13g2_decap_4 FILLER_38_696 ();
 sg13g2_fill_2 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_4 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_39 ();
 sg13g2_fill_2 FILLER_39_76 ();
 sg13g2_fill_1 FILLER_39_78 ();
 sg13g2_decap_4 FILLER_39_96 ();
 sg13g2_fill_1 FILLER_39_108 ();
 sg13g2_decap_8 FILLER_39_135 ();
 sg13g2_decap_4 FILLER_39_178 ();
 sg13g2_fill_2 FILLER_39_191 ();
 sg13g2_fill_1 FILLER_39_193 ();
 sg13g2_decap_8 FILLER_39_199 ();
 sg13g2_fill_1 FILLER_39_206 ();
 sg13g2_fill_1 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_262 ();
 sg13g2_fill_1 FILLER_39_264 ();
 sg13g2_fill_1 FILLER_39_273 ();
 sg13g2_fill_1 FILLER_39_296 ();
 sg13g2_decap_8 FILLER_39_318 ();
 sg13g2_decap_4 FILLER_39_338 ();
 sg13g2_fill_2 FILLER_39_342 ();
 sg13g2_decap_4 FILLER_39_352 ();
 sg13g2_fill_2 FILLER_39_356 ();
 sg13g2_decap_8 FILLER_39_376 ();
 sg13g2_fill_1 FILLER_39_383 ();
 sg13g2_fill_1 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_39_408 ();
 sg13g2_decap_4 FILLER_39_415 ();
 sg13g2_fill_1 FILLER_39_419 ();
 sg13g2_decap_8 FILLER_39_433 ();
 sg13g2_decap_8 FILLER_39_454 ();
 sg13g2_decap_4 FILLER_39_466 ();
 sg13g2_fill_2 FILLER_39_470 ();
 sg13g2_decap_4 FILLER_39_491 ();
 sg13g2_fill_1 FILLER_39_495 ();
 sg13g2_decap_4 FILLER_39_515 ();
 sg13g2_fill_1 FILLER_39_519 ();
 sg13g2_fill_2 FILLER_39_548 ();
 sg13g2_fill_2 FILLER_39_555 ();
 sg13g2_decap_8 FILLER_39_566 ();
 sg13g2_decap_4 FILLER_39_573 ();
 sg13g2_fill_2 FILLER_39_577 ();
 sg13g2_fill_2 FILLER_39_583 ();
 sg13g2_fill_2 FILLER_39_589 ();
 sg13g2_fill_1 FILLER_39_591 ();
 sg13g2_decap_4 FILLER_39_618 ();
 sg13g2_fill_2 FILLER_39_627 ();
 sg13g2_fill_1 FILLER_39_669 ();
 sg13g2_fill_1 FILLER_39_684 ();
 sg13g2_decap_8 FILLER_39_710 ();
 sg13g2_decap_8 FILLER_39_717 ();
 sg13g2_decap_8 FILLER_39_724 ();
 sg13g2_decap_8 FILLER_39_731 ();
 sg13g2_decap_8 FILLER_39_738 ();
 sg13g2_decap_8 FILLER_39_745 ();
 sg13g2_decap_8 FILLER_39_752 ();
 sg13g2_decap_8 FILLER_39_759 ();
 sg13g2_decap_8 FILLER_39_766 ();
 sg13g2_decap_8 FILLER_39_773 ();
 sg13g2_decap_8 FILLER_39_780 ();
 sg13g2_decap_8 FILLER_39_787 ();
 sg13g2_decap_8 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_801 ();
 sg13g2_decap_8 FILLER_39_808 ();
 sg13g2_decap_8 FILLER_39_815 ();
 sg13g2_decap_8 FILLER_39_822 ();
 sg13g2_decap_8 FILLER_39_829 ();
 sg13g2_decap_8 FILLER_39_836 ();
 sg13g2_decap_8 FILLER_39_843 ();
 sg13g2_decap_8 FILLER_39_850 ();
 sg13g2_decap_4 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_4 FILLER_40_28 ();
 sg13g2_fill_2 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_98 ();
 sg13g2_decap_4 FILLER_40_131 ();
 sg13g2_fill_2 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_152 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_fill_1 FILLER_40_215 ();
 sg13g2_fill_1 FILLER_40_222 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_fill_1 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_263 ();
 sg13g2_decap_8 FILLER_40_270 ();
 sg13g2_decap_8 FILLER_40_277 ();
 sg13g2_fill_2 FILLER_40_284 ();
 sg13g2_fill_1 FILLER_40_286 ();
 sg13g2_decap_8 FILLER_40_298 ();
 sg13g2_fill_1 FILLER_40_334 ();
 sg13g2_fill_2 FILLER_40_349 ();
 sg13g2_fill_2 FILLER_40_380 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_decap_4 FILLER_40_413 ();
 sg13g2_decap_4 FILLER_40_434 ();
 sg13g2_decap_4 FILLER_40_444 ();
 sg13g2_fill_2 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_498 ();
 sg13g2_fill_2 FILLER_40_505 ();
 sg13g2_decap_8 FILLER_40_512 ();
 sg13g2_decap_4 FILLER_40_519 ();
 sg13g2_fill_1 FILLER_40_523 ();
 sg13g2_fill_1 FILLER_40_558 ();
 sg13g2_fill_2 FILLER_40_572 ();
 sg13g2_decap_8 FILLER_40_605 ();
 sg13g2_decap_4 FILLER_40_612 ();
 sg13g2_fill_2 FILLER_40_624 ();
 sg13g2_fill_1 FILLER_40_630 ();
 sg13g2_decap_4 FILLER_40_641 ();
 sg13g2_fill_2 FILLER_40_645 ();
 sg13g2_fill_2 FILLER_40_653 ();
 sg13g2_fill_2 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_decap_8 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_847 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_192 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_fill_2 FILLER_41_238 ();
 sg13g2_decap_4 FILLER_41_272 ();
 sg13g2_decap_4 FILLER_41_304 ();
 sg13g2_fill_1 FILLER_41_317 ();
 sg13g2_decap_4 FILLER_41_322 ();
 sg13g2_fill_2 FILLER_41_326 ();
 sg13g2_decap_8 FILLER_41_338 ();
 sg13g2_decap_8 FILLER_41_345 ();
 sg13g2_fill_2 FILLER_41_360 ();
 sg13g2_fill_1 FILLER_41_362 ();
 sg13g2_fill_2 FILLER_41_377 ();
 sg13g2_fill_2 FILLER_41_387 ();
 sg13g2_fill_1 FILLER_41_389 ();
 sg13g2_fill_2 FILLER_41_402 ();
 sg13g2_fill_1 FILLER_41_404 ();
 sg13g2_decap_8 FILLER_41_416 ();
 sg13g2_decap_4 FILLER_41_423 ();
 sg13g2_fill_1 FILLER_41_427 ();
 sg13g2_decap_4 FILLER_41_446 ();
 sg13g2_fill_2 FILLER_41_450 ();
 sg13g2_fill_2 FILLER_41_474 ();
 sg13g2_decap_4 FILLER_41_489 ();
 sg13g2_fill_1 FILLER_41_493 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_fill_2 FILLER_41_504 ();
 sg13g2_fill_1 FILLER_41_506 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_decap_4 FILLER_41_539 ();
 sg13g2_fill_1 FILLER_41_543 ();
 sg13g2_fill_1 FILLER_41_553 ();
 sg13g2_fill_2 FILLER_41_584 ();
 sg13g2_fill_1 FILLER_41_591 ();
 sg13g2_decap_4 FILLER_41_610 ();
 sg13g2_fill_1 FILLER_41_614 ();
 sg13g2_fill_2 FILLER_41_623 ();
 sg13g2_fill_1 FILLER_41_625 ();
 sg13g2_fill_1 FILLER_41_661 ();
 sg13g2_fill_2 FILLER_41_676 ();
 sg13g2_fill_1 FILLER_41_691 ();
 sg13g2_decap_4 FILLER_41_712 ();
 sg13g2_fill_2 FILLER_41_716 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_fill_2 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_63 ();
 sg13g2_fill_1 FILLER_42_65 ();
 sg13g2_fill_1 FILLER_42_149 ();
 sg13g2_decap_4 FILLER_42_174 ();
 sg13g2_fill_2 FILLER_42_178 ();
 sg13g2_decap_4 FILLER_42_228 ();
 sg13g2_decap_8 FILLER_42_237 ();
 sg13g2_decap_4 FILLER_42_244 ();
 sg13g2_fill_2 FILLER_42_248 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_4 FILLER_42_382 ();
 sg13g2_fill_2 FILLER_42_386 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_445 ();
 sg13g2_fill_1 FILLER_42_459 ();
 sg13g2_fill_2 FILLER_42_479 ();
 sg13g2_fill_1 FILLER_42_497 ();
 sg13g2_decap_4 FILLER_42_509 ();
 sg13g2_decap_8 FILLER_42_524 ();
 sg13g2_decap_4 FILLER_42_568 ();
 sg13g2_fill_1 FILLER_42_572 ();
 sg13g2_decap_8 FILLER_42_578 ();
 sg13g2_fill_1 FILLER_42_585 ();
 sg13g2_decap_8 FILLER_42_591 ();
 sg13g2_fill_2 FILLER_42_598 ();
 sg13g2_fill_1 FILLER_42_600 ();
 sg13g2_fill_2 FILLER_42_609 ();
 sg13g2_fill_2 FILLER_42_637 ();
 sg13g2_fill_1 FILLER_42_639 ();
 sg13g2_decap_4 FILLER_42_653 ();
 sg13g2_fill_2 FILLER_42_675 ();
 sg13g2_fill_1 FILLER_42_683 ();
 sg13g2_fill_1 FILLER_42_701 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_826 ();
 sg13g2_decap_8 FILLER_42_833 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_fill_2 FILLER_43_42 ();
 sg13g2_fill_2 FILLER_43_79 ();
 sg13g2_fill_1 FILLER_43_81 ();
 sg13g2_fill_2 FILLER_43_102 ();
 sg13g2_fill_2 FILLER_43_114 ();
 sg13g2_fill_2 FILLER_43_121 ();
 sg13g2_fill_1 FILLER_43_123 ();
 sg13g2_fill_1 FILLER_43_139 ();
 sg13g2_fill_1 FILLER_43_172 ();
 sg13g2_decap_4 FILLER_43_189 ();
 sg13g2_fill_1 FILLER_43_193 ();
 sg13g2_fill_2 FILLER_43_208 ();
 sg13g2_fill_2 FILLER_43_250 ();
 sg13g2_fill_1 FILLER_43_252 ();
 sg13g2_fill_2 FILLER_43_263 ();
 sg13g2_fill_1 FILLER_43_265 ();
 sg13g2_decap_4 FILLER_43_271 ();
 sg13g2_fill_1 FILLER_43_275 ();
 sg13g2_decap_8 FILLER_43_314 ();
 sg13g2_decap_4 FILLER_43_321 ();
 sg13g2_fill_1 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_352 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_fill_1 FILLER_43_422 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_fill_1 FILLER_43_430 ();
 sg13g2_fill_2 FILLER_43_461 ();
 sg13g2_fill_1 FILLER_43_475 ();
 sg13g2_decap_8 FILLER_43_517 ();
 sg13g2_fill_1 FILLER_43_524 ();
 sg13g2_fill_2 FILLER_43_536 ();
 sg13g2_decap_8 FILLER_43_541 ();
 sg13g2_decap_4 FILLER_43_557 ();
 sg13g2_fill_2 FILLER_43_561 ();
 sg13g2_decap_4 FILLER_43_567 ();
 sg13g2_fill_1 FILLER_43_571 ();
 sg13g2_fill_1 FILLER_43_599 ();
 sg13g2_fill_2 FILLER_43_605 ();
 sg13g2_fill_1 FILLER_43_607 ();
 sg13g2_fill_1 FILLER_43_622 ();
 sg13g2_fill_2 FILLER_43_647 ();
 sg13g2_fill_1 FILLER_43_649 ();
 sg13g2_decap_8 FILLER_43_663 ();
 sg13g2_decap_4 FILLER_43_670 ();
 sg13g2_fill_1 FILLER_43_674 ();
 sg13g2_decap_8 FILLER_43_729 ();
 sg13g2_decap_8 FILLER_43_736 ();
 sg13g2_decap_8 FILLER_43_743 ();
 sg13g2_decap_8 FILLER_43_750 ();
 sg13g2_decap_8 FILLER_43_757 ();
 sg13g2_decap_8 FILLER_43_764 ();
 sg13g2_decap_8 FILLER_43_771 ();
 sg13g2_decap_8 FILLER_43_778 ();
 sg13g2_decap_8 FILLER_43_785 ();
 sg13g2_decap_8 FILLER_43_792 ();
 sg13g2_decap_8 FILLER_43_799 ();
 sg13g2_decap_8 FILLER_43_806 ();
 sg13g2_decap_8 FILLER_43_813 ();
 sg13g2_decap_8 FILLER_43_820 ();
 sg13g2_decap_8 FILLER_43_827 ();
 sg13g2_decap_8 FILLER_43_834 ();
 sg13g2_decap_8 FILLER_43_841 ();
 sg13g2_decap_8 FILLER_43_848 ();
 sg13g2_decap_8 FILLER_43_855 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_4 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_53 ();
 sg13g2_fill_2 FILLER_44_85 ();
 sg13g2_fill_1 FILLER_44_87 ();
 sg13g2_fill_1 FILLER_44_103 ();
 sg13g2_fill_2 FILLER_44_159 ();
 sg13g2_fill_1 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_173 ();
 sg13g2_fill_2 FILLER_44_233 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_fill_2 FILLER_44_250 ();
 sg13g2_decap_8 FILLER_44_283 ();
 sg13g2_decap_4 FILLER_44_290 ();
 sg13g2_decap_8 FILLER_44_299 ();
 sg13g2_fill_1 FILLER_44_306 ();
 sg13g2_decap_4 FILLER_44_345 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_374 ();
 sg13g2_decap_8 FILLER_44_381 ();
 sg13g2_fill_2 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_437 ();
 sg13g2_fill_1 FILLER_44_444 ();
 sg13g2_decap_8 FILLER_44_453 ();
 sg13g2_fill_2 FILLER_44_460 ();
 sg13g2_fill_2 FILLER_44_467 ();
 sg13g2_fill_1 FILLER_44_469 ();
 sg13g2_decap_4 FILLER_44_479 ();
 sg13g2_decap_4 FILLER_44_493 ();
 sg13g2_decap_8 FILLER_44_502 ();
 sg13g2_fill_1 FILLER_44_509 ();
 sg13g2_fill_2 FILLER_44_521 ();
 sg13g2_fill_2 FILLER_44_569 ();
 sg13g2_fill_1 FILLER_44_571 ();
 sg13g2_decap_4 FILLER_44_592 ();
 sg13g2_fill_1 FILLER_44_606 ();
 sg13g2_fill_1 FILLER_44_616 ();
 sg13g2_fill_1 FILLER_44_623 ();
 sg13g2_fill_1 FILLER_44_644 ();
 sg13g2_decap_4 FILLER_44_672 ();
 sg13g2_fill_1 FILLER_44_676 ();
 sg13g2_fill_2 FILLER_44_694 ();
 sg13g2_fill_1 FILLER_44_696 ();
 sg13g2_fill_1 FILLER_44_702 ();
 sg13g2_decap_8 FILLER_44_729 ();
 sg13g2_decap_8 FILLER_44_736 ();
 sg13g2_decap_8 FILLER_44_743 ();
 sg13g2_decap_8 FILLER_44_750 ();
 sg13g2_decap_8 FILLER_44_757 ();
 sg13g2_decap_8 FILLER_44_764 ();
 sg13g2_decap_8 FILLER_44_771 ();
 sg13g2_decap_8 FILLER_44_778 ();
 sg13g2_decap_8 FILLER_44_785 ();
 sg13g2_decap_8 FILLER_44_792 ();
 sg13g2_decap_8 FILLER_44_799 ();
 sg13g2_decap_8 FILLER_44_806 ();
 sg13g2_decap_8 FILLER_44_813 ();
 sg13g2_decap_8 FILLER_44_820 ();
 sg13g2_decap_8 FILLER_44_827 ();
 sg13g2_decap_8 FILLER_44_834 ();
 sg13g2_decap_8 FILLER_44_841 ();
 sg13g2_decap_8 FILLER_44_848 ();
 sg13g2_decap_8 FILLER_44_855 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_fill_1 FILLER_45_42 ();
 sg13g2_fill_1 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_108 ();
 sg13g2_fill_2 FILLER_45_132 ();
 sg13g2_fill_1 FILLER_45_158 ();
 sg13g2_fill_2 FILLER_45_168 ();
 sg13g2_fill_1 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_194 ();
 sg13g2_fill_1 FILLER_45_231 ();
 sg13g2_fill_2 FILLER_45_258 ();
 sg13g2_fill_2 FILLER_45_275 ();
 sg13g2_fill_1 FILLER_45_285 ();
 sg13g2_decap_4 FILLER_45_291 ();
 sg13g2_decap_4 FILLER_45_331 ();
 sg13g2_fill_1 FILLER_45_350 ();
 sg13g2_fill_1 FILLER_45_356 ();
 sg13g2_fill_1 FILLER_45_367 ();
 sg13g2_fill_1 FILLER_45_425 ();
 sg13g2_fill_2 FILLER_45_443 ();
 sg13g2_fill_1 FILLER_45_445 ();
 sg13g2_decap_8 FILLER_45_452 ();
 sg13g2_fill_2 FILLER_45_459 ();
 sg13g2_decap_8 FILLER_45_515 ();
 sg13g2_fill_2 FILLER_45_522 ();
 sg13g2_fill_1 FILLER_45_524 ();
 sg13g2_decap_8 FILLER_45_536 ();
 sg13g2_fill_1 FILLER_45_543 ();
 sg13g2_fill_1 FILLER_45_549 ();
 sg13g2_fill_2 FILLER_45_571 ();
 sg13g2_fill_1 FILLER_45_597 ();
 sg13g2_decap_4 FILLER_45_601 ();
 sg13g2_fill_2 FILLER_45_605 ();
 sg13g2_fill_2 FILLER_45_623 ();
 sg13g2_decap_8 FILLER_45_643 ();
 sg13g2_fill_2 FILLER_45_650 ();
 sg13g2_fill_2 FILLER_45_677 ();
 sg13g2_fill_2 FILLER_45_684 ();
 sg13g2_fill_1 FILLER_45_693 ();
 sg13g2_decap_8 FILLER_45_737 ();
 sg13g2_decap_8 FILLER_45_744 ();
 sg13g2_decap_8 FILLER_45_751 ();
 sg13g2_decap_8 FILLER_45_758 ();
 sg13g2_decap_8 FILLER_45_765 ();
 sg13g2_decap_8 FILLER_45_772 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_8 FILLER_45_786 ();
 sg13g2_decap_8 FILLER_45_793 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_decap_8 FILLER_45_807 ();
 sg13g2_decap_8 FILLER_45_814 ();
 sg13g2_decap_8 FILLER_45_821 ();
 sg13g2_decap_8 FILLER_45_828 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_4 FILLER_45_856 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_4 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_39 ();
 sg13g2_fill_1 FILLER_46_171 ();
 sg13g2_decap_4 FILLER_46_204 ();
 sg13g2_fill_1 FILLER_46_219 ();
 sg13g2_fill_2 FILLER_46_266 ();
 sg13g2_decap_4 FILLER_46_279 ();
 sg13g2_fill_1 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_319 ();
 sg13g2_decap_8 FILLER_46_330 ();
 sg13g2_fill_2 FILLER_46_337 ();
 sg13g2_decap_8 FILLER_46_368 ();
 sg13g2_fill_1 FILLER_46_375 ();
 sg13g2_fill_2 FILLER_46_412 ();
 sg13g2_fill_1 FILLER_46_435 ();
 sg13g2_decap_8 FILLER_46_451 ();
 sg13g2_decap_8 FILLER_46_458 ();
 sg13g2_fill_2 FILLER_46_485 ();
 sg13g2_decap_4 FILLER_46_492 ();
 sg13g2_fill_2 FILLER_46_496 ();
 sg13g2_decap_4 FILLER_46_502 ();
 sg13g2_fill_2 FILLER_46_544 ();
 sg13g2_fill_2 FILLER_46_556 ();
 sg13g2_fill_1 FILLER_46_558 ();
 sg13g2_decap_8 FILLER_46_589 ();
 sg13g2_fill_2 FILLER_46_596 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_fill_2 FILLER_46_616 ();
 sg13g2_fill_1 FILLER_46_618 ();
 sg13g2_fill_1 FILLER_46_624 ();
 sg13g2_decap_8 FILLER_46_652 ();
 sg13g2_fill_1 FILLER_46_659 ();
 sg13g2_fill_2 FILLER_46_679 ();
 sg13g2_fill_1 FILLER_46_690 ();
 sg13g2_decap_8 FILLER_46_737 ();
 sg13g2_decap_8 FILLER_46_744 ();
 sg13g2_decap_8 FILLER_46_751 ();
 sg13g2_decap_8 FILLER_46_758 ();
 sg13g2_decap_8 FILLER_46_765 ();
 sg13g2_decap_8 FILLER_46_772 ();
 sg13g2_decap_8 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_793 ();
 sg13g2_decap_8 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_decap_8 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_835 ();
 sg13g2_decap_8 FILLER_46_842 ();
 sg13g2_decap_8 FILLER_46_849 ();
 sg13g2_decap_4 FILLER_46_856 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_fill_1 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_77 ();
 sg13g2_fill_2 FILLER_47_98 ();
 sg13g2_fill_1 FILLER_47_142 ();
 sg13g2_fill_1 FILLER_47_185 ();
 sg13g2_fill_2 FILLER_47_204 ();
 sg13g2_fill_2 FILLER_47_227 ();
 sg13g2_fill_1 FILLER_47_229 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_fill_1 FILLER_47_285 ();
 sg13g2_fill_2 FILLER_47_310 ();
 sg13g2_fill_1 FILLER_47_312 ();
 sg13g2_decap_4 FILLER_47_343 ();
 sg13g2_fill_1 FILLER_47_347 ();
 sg13g2_decap_4 FILLER_47_353 ();
 sg13g2_fill_2 FILLER_47_357 ();
 sg13g2_fill_2 FILLER_47_388 ();
 sg13g2_fill_1 FILLER_47_414 ();
 sg13g2_fill_2 FILLER_47_425 ();
 sg13g2_fill_2 FILLER_47_437 ();
 sg13g2_fill_1 FILLER_47_439 ();
 sg13g2_fill_1 FILLER_47_445 ();
 sg13g2_decap_8 FILLER_47_460 ();
 sg13g2_decap_8 FILLER_47_467 ();
 sg13g2_fill_1 FILLER_47_474 ();
 sg13g2_decap_4 FILLER_47_485 ();
 sg13g2_fill_2 FILLER_47_489 ();
 sg13g2_decap_4 FILLER_47_496 ();
 sg13g2_decap_4 FILLER_47_524 ();
 sg13g2_fill_2 FILLER_47_532 ();
 sg13g2_fill_1 FILLER_47_534 ();
 sg13g2_fill_1 FILLER_47_559 ();
 sg13g2_decap_8 FILLER_47_580 ();
 sg13g2_fill_2 FILLER_47_587 ();
 sg13g2_fill_2 FILLER_47_688 ();
 sg13g2_fill_2 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_fill_1 FILLER_48_75 ();
 sg13g2_fill_2 FILLER_48_137 ();
 sg13g2_fill_1 FILLER_48_165 ();
 sg13g2_fill_2 FILLER_48_190 ();
 sg13g2_fill_1 FILLER_48_224 ();
 sg13g2_fill_1 FILLER_48_238 ();
 sg13g2_fill_1 FILLER_48_254 ();
 sg13g2_fill_1 FILLER_48_296 ();
 sg13g2_fill_2 FILLER_48_301 ();
 sg13g2_fill_1 FILLER_48_322 ();
 sg13g2_decap_4 FILLER_48_332 ();
 sg13g2_fill_2 FILLER_48_341 ();
 sg13g2_decap_4 FILLER_48_372 ();
 sg13g2_fill_2 FILLER_48_391 ();
 sg13g2_fill_1 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_430 ();
 sg13g2_fill_2 FILLER_48_471 ();
 sg13g2_fill_1 FILLER_48_473 ();
 sg13g2_decap_4 FILLER_48_489 ();
 sg13g2_fill_2 FILLER_48_493 ();
 sg13g2_fill_2 FILLER_48_515 ();
 sg13g2_fill_1 FILLER_48_517 ();
 sg13g2_fill_2 FILLER_48_538 ();
 sg13g2_fill_1 FILLER_48_591 ();
 sg13g2_fill_2 FILLER_48_616 ();
 sg13g2_fill_1 FILLER_48_618 ();
 sg13g2_fill_2 FILLER_48_660 ();
 sg13g2_fill_1 FILLER_48_667 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_fill_2 FILLER_48_686 ();
 sg13g2_fill_2 FILLER_48_698 ();
 sg13g2_fill_2 FILLER_48_706 ();
 sg13g2_decap_4 FILLER_48_718 ();
 sg13g2_decap_8 FILLER_48_733 ();
 sg13g2_decap_8 FILLER_48_740 ();
 sg13g2_decap_8 FILLER_48_747 ();
 sg13g2_fill_2 FILLER_48_754 ();
 sg13g2_fill_1 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_decap_8 FILLER_48_787 ();
 sg13g2_decap_8 FILLER_48_794 ();
 sg13g2_decap_8 FILLER_48_801 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_4 FILLER_48_857 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_fill_2 FILLER_49_49 ();
 sg13g2_fill_2 FILLER_49_82 ();
 sg13g2_fill_1 FILLER_49_122 ();
 sg13g2_fill_1 FILLER_49_128 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_158 ();
 sg13g2_fill_2 FILLER_49_221 ();
 sg13g2_fill_1 FILLER_49_263 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_fill_2 FILLER_49_303 ();
 sg13g2_fill_2 FILLER_49_313 ();
 sg13g2_fill_2 FILLER_49_346 ();
 sg13g2_fill_1 FILLER_49_348 ();
 sg13g2_fill_1 FILLER_49_446 ();
 sg13g2_fill_2 FILLER_49_452 ();
 sg13g2_decap_4 FILLER_49_475 ();
 sg13g2_fill_1 FILLER_49_495 ();
 sg13g2_decap_8 FILLER_49_506 ();
 sg13g2_decap_4 FILLER_49_513 ();
 sg13g2_fill_2 FILLER_49_517 ();
 sg13g2_fill_2 FILLER_49_533 ();
 sg13g2_decap_4 FILLER_49_542 ();
 sg13g2_fill_2 FILLER_49_580 ();
 sg13g2_fill_1 FILLER_49_582 ();
 sg13g2_decap_4 FILLER_49_615 ();
 sg13g2_decap_8 FILLER_49_627 ();
 sg13g2_decap_4 FILLER_49_646 ();
 sg13g2_fill_2 FILLER_49_650 ();
 sg13g2_fill_1 FILLER_49_673 ();
 sg13g2_decap_8 FILLER_49_683 ();
 sg13g2_fill_2 FILLER_49_690 ();
 sg13g2_fill_1 FILLER_49_692 ();
 sg13g2_decap_4 FILLER_49_717 ();
 sg13g2_fill_2 FILLER_49_745 ();
 sg13g2_fill_1 FILLER_49_747 ();
 sg13g2_fill_1 FILLER_49_760 ();
 sg13g2_fill_2 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_789 ();
 sg13g2_decap_8 FILLER_49_796 ();
 sg13g2_decap_8 FILLER_49_803 ();
 sg13g2_decap_8 FILLER_49_810 ();
 sg13g2_decap_8 FILLER_49_817 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_831 ();
 sg13g2_decap_8 FILLER_49_838 ();
 sg13g2_decap_8 FILLER_49_845 ();
 sg13g2_decap_8 FILLER_49_852 ();
 sg13g2_fill_2 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_fill_2 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_109 ();
 sg13g2_fill_1 FILLER_50_111 ();
 sg13g2_fill_2 FILLER_50_123 ();
 sg13g2_fill_1 FILLER_50_125 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_fill_1 FILLER_50_155 ();
 sg13g2_fill_1 FILLER_50_178 ();
 sg13g2_fill_2 FILLER_50_187 ();
 sg13g2_fill_2 FILLER_50_307 ();
 sg13g2_decap_8 FILLER_50_327 ();
 sg13g2_decap_8 FILLER_50_334 ();
 sg13g2_fill_2 FILLER_50_341 ();
 sg13g2_fill_1 FILLER_50_343 ();
 sg13g2_fill_2 FILLER_50_374 ();
 sg13g2_fill_1 FILLER_50_376 ();
 sg13g2_fill_2 FILLER_50_381 ();
 sg13g2_fill_2 FILLER_50_391 ();
 sg13g2_fill_1 FILLER_50_403 ();
 sg13g2_fill_2 FILLER_50_409 ();
 sg13g2_fill_1 FILLER_50_411 ();
 sg13g2_decap_8 FILLER_50_426 ();
 sg13g2_decap_4 FILLER_50_433 ();
 sg13g2_fill_1 FILLER_50_437 ();
 sg13g2_decap_4 FILLER_50_455 ();
 sg13g2_fill_2 FILLER_50_459 ();
 sg13g2_fill_2 FILLER_50_492 ();
 sg13g2_decap_4 FILLER_50_552 ();
 sg13g2_fill_1 FILLER_50_556 ();
 sg13g2_fill_1 FILLER_50_561 ();
 sg13g2_fill_2 FILLER_50_581 ();
 sg13g2_fill_1 FILLER_50_583 ();
 sg13g2_fill_1 FILLER_50_600 ();
 sg13g2_fill_1 FILLER_50_610 ();
 sg13g2_fill_2 FILLER_50_622 ();
 sg13g2_fill_1 FILLER_50_624 ();
 sg13g2_decap_4 FILLER_50_634 ();
 sg13g2_fill_2 FILLER_50_638 ();
 sg13g2_decap_8 FILLER_50_656 ();
 sg13g2_decap_4 FILLER_50_663 ();
 sg13g2_fill_1 FILLER_50_667 ();
 sg13g2_decap_4 FILLER_50_691 ();
 sg13g2_fill_1 FILLER_50_695 ();
 sg13g2_decap_4 FILLER_50_713 ();
 sg13g2_fill_2 FILLER_50_717 ();
 sg13g2_fill_2 FILLER_50_729 ();
 sg13g2_fill_1 FILLER_50_731 ();
 sg13g2_decap_4 FILLER_50_759 ();
 sg13g2_fill_1 FILLER_50_763 ();
 sg13g2_fill_1 FILLER_50_775 ();
 sg13g2_decap_8 FILLER_50_793 ();
 sg13g2_decap_8 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_807 ();
 sg13g2_decap_8 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_821 ();
 sg13g2_decap_8 FILLER_50_828 ();
 sg13g2_decap_8 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_842 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_75 ();
 sg13g2_fill_2 FILLER_51_90 ();
 sg13g2_fill_2 FILLER_51_100 ();
 sg13g2_fill_2 FILLER_51_123 ();
 sg13g2_fill_1 FILLER_51_125 ();
 sg13g2_fill_2 FILLER_51_153 ();
 sg13g2_fill_1 FILLER_51_155 ();
 sg13g2_fill_1 FILLER_51_231 ();
 sg13g2_fill_1 FILLER_51_286 ();
 sg13g2_fill_1 FILLER_51_297 ();
 sg13g2_fill_1 FILLER_51_317 ();
 sg13g2_fill_1 FILLER_51_328 ();
 sg13g2_decap_8 FILLER_51_338 ();
 sg13g2_fill_1 FILLER_51_345 ();
 sg13g2_fill_2 FILLER_51_368 ();
 sg13g2_fill_1 FILLER_51_370 ();
 sg13g2_fill_1 FILLER_51_384 ();
 sg13g2_fill_1 FILLER_51_405 ();
 sg13g2_decap_4 FILLER_51_459 ();
 sg13g2_decap_8 FILLER_51_471 ();
 sg13g2_fill_2 FILLER_51_478 ();
 sg13g2_decap_4 FILLER_51_509 ();
 sg13g2_fill_1 FILLER_51_513 ();
 sg13g2_fill_1 FILLER_51_540 ();
 sg13g2_fill_2 FILLER_51_546 ();
 sg13g2_fill_2 FILLER_51_557 ();
 sg13g2_fill_1 FILLER_51_559 ();
 sg13g2_fill_2 FILLER_51_571 ();
 sg13g2_fill_2 FILLER_51_590 ();
 sg13g2_decap_8 FILLER_51_606 ();
 sg13g2_fill_1 FILLER_51_613 ();
 sg13g2_decap_4 FILLER_51_632 ();
 sg13g2_fill_1 FILLER_51_636 ();
 sg13g2_fill_1 FILLER_51_647 ();
 sg13g2_decap_4 FILLER_51_664 ();
 sg13g2_fill_2 FILLER_51_668 ();
 sg13g2_fill_1 FILLER_51_691 ();
 sg13g2_fill_1 FILLER_51_696 ();
 sg13g2_fill_2 FILLER_51_711 ();
 sg13g2_fill_1 FILLER_51_713 ();
 sg13g2_fill_1 FILLER_51_736 ();
 sg13g2_fill_2 FILLER_51_761 ();
 sg13g2_decap_4 FILLER_51_785 ();
 sg13g2_fill_1 FILLER_51_789 ();
 sg13g2_decap_8 FILLER_51_805 ();
 sg13g2_fill_1 FILLER_51_812 ();
 sg13g2_fill_2 FILLER_51_822 ();
 sg13g2_fill_1 FILLER_51_824 ();
 sg13g2_decap_8 FILLER_51_833 ();
 sg13g2_decap_8 FILLER_51_840 ();
 sg13g2_decap_8 FILLER_51_847 ();
 sg13g2_decap_8 FILLER_51_854 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_4 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_42 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_2 FILLER_52_94 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_fill_2 FILLER_52_164 ();
 sg13g2_fill_2 FILLER_52_174 ();
 sg13g2_fill_1 FILLER_52_200 ();
 sg13g2_decap_4 FILLER_52_247 ();
 sg13g2_fill_1 FILLER_52_256 ();
 sg13g2_decap_8 FILLER_52_267 ();
 sg13g2_fill_2 FILLER_52_274 ();
 sg13g2_fill_1 FILLER_52_276 ();
 sg13g2_decap_4 FILLER_52_315 ();
 sg13g2_decap_8 FILLER_52_345 ();
 sg13g2_decap_4 FILLER_52_367 ();
 sg13g2_fill_2 FILLER_52_371 ();
 sg13g2_fill_1 FILLER_52_393 ();
 sg13g2_fill_2 FILLER_52_399 ();
 sg13g2_fill_1 FILLER_52_401 ();
 sg13g2_decap_8 FILLER_52_424 ();
 sg13g2_fill_1 FILLER_52_431 ();
 sg13g2_decap_4 FILLER_52_446 ();
 sg13g2_decap_8 FILLER_52_498 ();
 sg13g2_fill_2 FILLER_52_505 ();
 sg13g2_decap_8 FILLER_52_522 ();
 sg13g2_decap_8 FILLER_52_529 ();
 sg13g2_decap_8 FILLER_52_536 ();
 sg13g2_decap_8 FILLER_52_553 ();
 sg13g2_fill_2 FILLER_52_560 ();
 sg13g2_decap_4 FILLER_52_567 ();
 sg13g2_fill_2 FILLER_52_616 ();
 sg13g2_fill_2 FILLER_52_641 ();
 sg13g2_decap_4 FILLER_52_652 ();
 sg13g2_fill_1 FILLER_52_656 ();
 sg13g2_fill_2 FILLER_52_662 ();
 sg13g2_fill_1 FILLER_52_675 ();
 sg13g2_fill_2 FILLER_52_696 ();
 sg13g2_fill_1 FILLER_52_698 ();
 sg13g2_decap_8 FILLER_52_715 ();
 sg13g2_fill_2 FILLER_52_762 ();
 sg13g2_fill_1 FILLER_52_764 ();
 sg13g2_decap_4 FILLER_52_777 ();
 sg13g2_fill_2 FILLER_52_781 ();
 sg13g2_decap_4 FILLER_52_801 ();
 sg13g2_fill_2 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_848 ();
 sg13g2_decap_8 FILLER_52_855 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_18 ();
 sg13g2_fill_1 FILLER_53_111 ();
 sg13g2_fill_2 FILLER_53_121 ();
 sg13g2_fill_2 FILLER_53_137 ();
 sg13g2_decap_4 FILLER_53_156 ();
 sg13g2_fill_1 FILLER_53_186 ();
 sg13g2_fill_1 FILLER_53_208 ();
 sg13g2_fill_1 FILLER_53_215 ();
 sg13g2_fill_2 FILLER_53_257 ();
 sg13g2_decap_4 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_fill_2 FILLER_53_315 ();
 sg13g2_fill_2 FILLER_53_326 ();
 sg13g2_decap_4 FILLER_53_333 ();
 sg13g2_fill_1 FILLER_53_337 ();
 sg13g2_decap_4 FILLER_53_416 ();
 sg13g2_fill_2 FILLER_53_431 ();
 sg13g2_fill_1 FILLER_53_433 ();
 sg13g2_fill_1 FILLER_53_443 ();
 sg13g2_decap_4 FILLER_53_476 ();
 sg13g2_fill_1 FILLER_53_480 ();
 sg13g2_decap_4 FILLER_53_485 ();
 sg13g2_decap_4 FILLER_53_516 ();
 sg13g2_decap_8 FILLER_53_540 ();
 sg13g2_fill_1 FILLER_53_547 ();
 sg13g2_fill_2 FILLER_53_560 ();
 sg13g2_fill_1 FILLER_53_562 ();
 sg13g2_fill_1 FILLER_53_584 ();
 sg13g2_fill_1 FILLER_53_590 ();
 sg13g2_fill_2 FILLER_53_610 ();
 sg13g2_fill_2 FILLER_53_630 ();
 sg13g2_fill_1 FILLER_53_632 ();
 sg13g2_fill_2 FILLER_53_638 ();
 sg13g2_fill_1 FILLER_53_640 ();
 sg13g2_fill_1 FILLER_53_661 ();
 sg13g2_fill_1 FILLER_53_671 ();
 sg13g2_decap_4 FILLER_53_687 ();
 sg13g2_fill_1 FILLER_53_731 ();
 sg13g2_decap_4 FILLER_53_759 ();
 sg13g2_fill_2 FILLER_53_763 ();
 sg13g2_decap_4 FILLER_53_770 ();
 sg13g2_decap_8 FILLER_53_786 ();
 sg13g2_fill_1 FILLER_53_793 ();
 sg13g2_decap_8 FILLER_53_832 ();
 sg13g2_decap_4 FILLER_53_839 ();
 sg13g2_decap_8 FILLER_53_851 ();
 sg13g2_decap_4 FILLER_53_858 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_75 ();
 sg13g2_fill_2 FILLER_54_85 ();
 sg13g2_fill_1 FILLER_54_87 ();
 sg13g2_fill_1 FILLER_54_101 ();
 sg13g2_fill_2 FILLER_54_112 ();
 sg13g2_fill_1 FILLER_54_119 ();
 sg13g2_fill_2 FILLER_54_130 ();
 sg13g2_fill_1 FILLER_54_132 ();
 sg13g2_fill_1 FILLER_54_145 ();
 sg13g2_fill_2 FILLER_54_188 ();
 sg13g2_fill_2 FILLER_54_224 ();
 sg13g2_fill_1 FILLER_54_248 ();
 sg13g2_decap_8 FILLER_54_281 ();
 sg13g2_decap_8 FILLER_54_288 ();
 sg13g2_decap_4 FILLER_54_295 ();
 sg13g2_fill_1 FILLER_54_299 ();
 sg13g2_decap_8 FILLER_54_314 ();
 sg13g2_fill_1 FILLER_54_325 ();
 sg13g2_fill_1 FILLER_54_334 ();
 sg13g2_decap_8 FILLER_54_339 ();
 sg13g2_decap_4 FILLER_54_346 ();
 sg13g2_fill_2 FILLER_54_350 ();
 sg13g2_decap_4 FILLER_54_371 ();
 sg13g2_fill_2 FILLER_54_378 ();
 sg13g2_decap_4 FILLER_54_420 ();
 sg13g2_decap_4 FILLER_54_438 ();
 sg13g2_fill_1 FILLER_54_442 ();
 sg13g2_decap_4 FILLER_54_488 ();
 sg13g2_fill_1 FILLER_54_497 ();
 sg13g2_decap_8 FILLER_54_507 ();
 sg13g2_fill_2 FILLER_54_514 ();
 sg13g2_fill_1 FILLER_54_540 ();
 sg13g2_decap_8 FILLER_54_566 ();
 sg13g2_decap_4 FILLER_54_578 ();
 sg13g2_fill_1 FILLER_54_582 ();
 sg13g2_decap_4 FILLER_54_587 ();
 sg13g2_decap_4 FILLER_54_602 ();
 sg13g2_fill_2 FILLER_54_606 ();
 sg13g2_decap_4 FILLER_54_628 ();
 sg13g2_fill_1 FILLER_54_641 ();
 sg13g2_decap_8 FILLER_54_654 ();
 sg13g2_decap_8 FILLER_54_661 ();
 sg13g2_decap_8 FILLER_54_668 ();
 sg13g2_fill_1 FILLER_54_675 ();
 sg13g2_decap_4 FILLER_54_695 ();
 sg13g2_fill_1 FILLER_54_719 ();
 sg13g2_fill_1 FILLER_54_726 ();
 sg13g2_fill_2 FILLER_54_742 ();
 sg13g2_decap_4 FILLER_54_785 ();
 sg13g2_fill_1 FILLER_54_789 ();
 sg13g2_fill_1 FILLER_54_805 ();
 sg13g2_fill_2 FILLER_54_823 ();
 sg13g2_fill_1 FILLER_54_825 ();
 sg13g2_fill_2 FILLER_54_838 ();
 sg13g2_fill_1 FILLER_54_840 ();
 sg13g2_decap_8 FILLER_54_853 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_11 ();
 sg13g2_fill_2 FILLER_55_48 ();
 sg13g2_fill_2 FILLER_55_97 ();
 sg13g2_fill_1 FILLER_55_99 ();
 sg13g2_fill_1 FILLER_55_114 ();
 sg13g2_decap_4 FILLER_55_138 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_fill_1 FILLER_55_149 ();
 sg13g2_decap_8 FILLER_55_163 ();
 sg13g2_fill_1 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_183 ();
 sg13g2_fill_2 FILLER_55_204 ();
 sg13g2_fill_2 FILLER_55_212 ();
 sg13g2_fill_1 FILLER_55_214 ();
 sg13g2_fill_1 FILLER_55_265 ();
 sg13g2_fill_1 FILLER_55_274 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_fill_2 FILLER_55_287 ();
 sg13g2_fill_1 FILLER_55_306 ();
 sg13g2_decap_4 FILLER_55_388 ();
 sg13g2_fill_1 FILLER_55_430 ();
 sg13g2_fill_1 FILLER_55_470 ();
 sg13g2_fill_2 FILLER_55_486 ();
 sg13g2_fill_1 FILLER_55_501 ();
 sg13g2_decap_4 FILLER_55_514 ();
 sg13g2_fill_1 FILLER_55_518 ();
 sg13g2_fill_2 FILLER_55_523 ();
 sg13g2_fill_1 FILLER_55_525 ();
 sg13g2_decap_4 FILLER_55_534 ();
 sg13g2_fill_1 FILLER_55_538 ();
 sg13g2_fill_1 FILLER_55_551 ();
 sg13g2_decap_8 FILLER_55_556 ();
 sg13g2_decap_4 FILLER_55_563 ();
 sg13g2_decap_8 FILLER_55_572 ();
 sg13g2_decap_8 FILLER_55_602 ();
 sg13g2_fill_1 FILLER_55_621 ();
 sg13g2_fill_1 FILLER_55_684 ();
 sg13g2_fill_2 FILLER_55_690 ();
 sg13g2_fill_1 FILLER_55_692 ();
 sg13g2_fill_2 FILLER_55_697 ();
 sg13g2_fill_2 FILLER_55_724 ();
 sg13g2_decap_8 FILLER_55_737 ();
 sg13g2_decap_8 FILLER_55_753 ();
 sg13g2_fill_1 FILLER_55_760 ();
 sg13g2_fill_1 FILLER_55_778 ();
 sg13g2_fill_2 FILLER_55_785 ();
 sg13g2_fill_1 FILLER_55_787 ();
 sg13g2_decap_4 FILLER_55_810 ();
 sg13g2_fill_1 FILLER_55_814 ();
 sg13g2_decap_8 FILLER_55_835 ();
 sg13g2_decap_4 FILLER_55_842 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_11 ();
 sg13g2_fill_1 FILLER_56_39 ();
 sg13g2_fill_1 FILLER_56_54 ();
 sg13g2_fill_1 FILLER_56_73 ();
 sg13g2_fill_2 FILLER_56_103 ();
 sg13g2_fill_2 FILLER_56_118 ();
 sg13g2_fill_1 FILLER_56_120 ();
 sg13g2_decap_8 FILLER_56_139 ();
 sg13g2_fill_1 FILLER_56_146 ();
 sg13g2_decap_4 FILLER_56_152 ();
 sg13g2_fill_2 FILLER_56_156 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_fill_2 FILLER_56_212 ();
 sg13g2_fill_2 FILLER_56_217 ();
 sg13g2_fill_1 FILLER_56_219 ();
 sg13g2_fill_2 FILLER_56_276 ();
 sg13g2_fill_1 FILLER_56_278 ();
 sg13g2_fill_2 FILLER_56_308 ();
 sg13g2_decap_8 FILLER_56_315 ();
 sg13g2_fill_1 FILLER_56_322 ();
 sg13g2_decap_8 FILLER_56_328 ();
 sg13g2_fill_2 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_337 ();
 sg13g2_fill_2 FILLER_56_346 ();
 sg13g2_fill_1 FILLER_56_371 ();
 sg13g2_decap_8 FILLER_56_386 ();
 sg13g2_fill_2 FILLER_56_393 ();
 sg13g2_fill_2 FILLER_56_404 ();
 sg13g2_decap_4 FILLER_56_411 ();
 sg13g2_fill_2 FILLER_56_447 ();
 sg13g2_fill_2 FILLER_56_459 ();
 sg13g2_fill_1 FILLER_56_496 ();
 sg13g2_fill_1 FILLER_56_529 ();
 sg13g2_fill_1 FILLER_56_542 ();
 sg13g2_fill_2 FILLER_56_547 ();
 sg13g2_decap_8 FILLER_56_604 ();
 sg13g2_fill_1 FILLER_56_617 ();
 sg13g2_fill_1 FILLER_56_651 ();
 sg13g2_fill_2 FILLER_56_706 ();
 sg13g2_fill_1 FILLER_56_708 ();
 sg13g2_decap_8 FILLER_56_725 ();
 sg13g2_fill_1 FILLER_56_732 ();
 sg13g2_fill_2 FILLER_56_763 ();
 sg13g2_fill_1 FILLER_56_779 ();
 sg13g2_fill_1 FILLER_56_786 ();
 sg13g2_fill_1 FILLER_56_808 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_1 FILLER_57_44 ();
 sg13g2_fill_1 FILLER_57_50 ();
 sg13g2_fill_2 FILLER_57_96 ();
 sg13g2_fill_2 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_112 ();
 sg13g2_fill_1 FILLER_57_127 ();
 sg13g2_fill_1 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_fill_2 FILLER_57_161 ();
 sg13g2_fill_1 FILLER_57_163 ();
 sg13g2_fill_2 FILLER_57_203 ();
 sg13g2_fill_1 FILLER_57_205 ();
 sg13g2_fill_2 FILLER_57_221 ();
 sg13g2_fill_1 FILLER_57_231 ();
 sg13g2_fill_1 FILLER_57_240 ();
 sg13g2_fill_2 FILLER_57_249 ();
 sg13g2_fill_2 FILLER_57_259 ();
 sg13g2_fill_2 FILLER_57_309 ();
 sg13g2_decap_4 FILLER_57_337 ();
 sg13g2_fill_2 FILLER_57_349 ();
 sg13g2_fill_2 FILLER_57_381 ();
 sg13g2_fill_1 FILLER_57_383 ();
 sg13g2_fill_2 FILLER_57_410 ();
 sg13g2_fill_1 FILLER_57_412 ();
 sg13g2_fill_1 FILLER_57_439 ();
 sg13g2_decap_4 FILLER_57_462 ();
 sg13g2_fill_1 FILLER_57_466 ();
 sg13g2_decap_8 FILLER_57_471 ();
 sg13g2_decap_4 FILLER_57_478 ();
 sg13g2_decap_4 FILLER_57_514 ();
 sg13g2_fill_2 FILLER_57_530 ();
 sg13g2_fill_2 FILLER_57_538 ();
 sg13g2_fill_1 FILLER_57_549 ();
 sg13g2_decap_4 FILLER_57_563 ();
 sg13g2_fill_2 FILLER_57_567 ();
 sg13g2_fill_2 FILLER_57_579 ();
 sg13g2_decap_4 FILLER_57_616 ();
 sg13g2_fill_2 FILLER_57_626 ();
 sg13g2_fill_1 FILLER_57_628 ();
 sg13g2_fill_2 FILLER_57_638 ();
 sg13g2_fill_2 FILLER_57_646 ();
 sg13g2_fill_1 FILLER_57_652 ();
 sg13g2_decap_8 FILLER_57_658 ();
 sg13g2_decap_4 FILLER_57_665 ();
 sg13g2_fill_1 FILLER_57_669 ();
 sg13g2_fill_2 FILLER_57_683 ();
 sg13g2_decap_8 FILLER_57_697 ();
 sg13g2_fill_2 FILLER_57_704 ();
 sg13g2_fill_1 FILLER_57_706 ();
 sg13g2_fill_2 FILLER_57_718 ();
 sg13g2_fill_1 FILLER_57_720 ();
 sg13g2_decap_4 FILLER_57_739 ();
 sg13g2_fill_2 FILLER_57_743 ();
 sg13g2_decap_8 FILLER_57_750 ();
 sg13g2_fill_1 FILLER_57_767 ();
 sg13g2_decap_4 FILLER_57_786 ();
 sg13g2_fill_1 FILLER_57_808 ();
 sg13g2_decap_4 FILLER_57_838 ();
 sg13g2_fill_1 FILLER_57_842 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_4 FILLER_58_14 ();
 sg13g2_fill_2 FILLER_58_70 ();
 sg13g2_fill_2 FILLER_58_88 ();
 sg13g2_fill_1 FILLER_58_90 ();
 sg13g2_fill_2 FILLER_58_124 ();
 sg13g2_fill_1 FILLER_58_126 ();
 sg13g2_fill_1 FILLER_58_147 ();
 sg13g2_fill_2 FILLER_58_185 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_fill_2 FILLER_58_241 ();
 sg13g2_fill_1 FILLER_58_243 ();
 sg13g2_fill_1 FILLER_58_264 ();
 sg13g2_decap_4 FILLER_58_338 ();
 sg13g2_fill_1 FILLER_58_342 ();
 sg13g2_fill_1 FILLER_58_360 ();
 sg13g2_fill_1 FILLER_58_415 ();
 sg13g2_fill_1 FILLER_58_453 ();
 sg13g2_fill_2 FILLER_58_486 ();
 sg13g2_fill_1 FILLER_58_515 ();
 sg13g2_fill_2 FILLER_58_539 ();
 sg13g2_fill_2 FILLER_58_555 ();
 sg13g2_fill_2 FILLER_58_577 ();
 sg13g2_fill_1 FILLER_58_579 ();
 sg13g2_fill_2 FILLER_58_585 ();
 sg13g2_fill_1 FILLER_58_587 ();
 sg13g2_fill_2 FILLER_58_598 ();
 sg13g2_fill_1 FILLER_58_600 ();
 sg13g2_decap_8 FILLER_58_607 ();
 sg13g2_decap_4 FILLER_58_614 ();
 sg13g2_fill_1 FILLER_58_618 ();
 sg13g2_decap_4 FILLER_58_653 ();
 sg13g2_fill_2 FILLER_58_663 ();
 sg13g2_fill_1 FILLER_58_665 ();
 sg13g2_fill_2 FILLER_58_671 ();
 sg13g2_decap_4 FILLER_58_687 ();
 sg13g2_fill_2 FILLER_58_691 ();
 sg13g2_decap_8 FILLER_58_720 ();
 sg13g2_fill_2 FILLER_58_727 ();
 sg13g2_decap_8 FILLER_58_780 ();
 sg13g2_fill_2 FILLER_58_787 ();
 sg13g2_fill_1 FILLER_58_789 ();
 sg13g2_fill_2 FILLER_58_812 ();
 sg13g2_decap_8 FILLER_58_832 ();
 sg13g2_fill_2 FILLER_58_839 ();
 sg13g2_fill_1 FILLER_58_841 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_7 ();
 sg13g2_fill_2 FILLER_59_40 ();
 sg13g2_fill_2 FILLER_59_60 ();
 sg13g2_fill_1 FILLER_59_104 ();
 sg13g2_fill_1 FILLER_59_113 ();
 sg13g2_fill_2 FILLER_59_119 ();
 sg13g2_fill_1 FILLER_59_121 ();
 sg13g2_fill_1 FILLER_59_127 ();
 sg13g2_decap_4 FILLER_59_137 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_2 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_158 ();
 sg13g2_fill_1 FILLER_59_180 ();
 sg13g2_fill_1 FILLER_59_199 ();
 sg13g2_fill_1 FILLER_59_282 ();
 sg13g2_fill_2 FILLER_59_314 ();
 sg13g2_decap_8 FILLER_59_344 ();
 sg13g2_fill_2 FILLER_59_351 ();
 sg13g2_fill_1 FILLER_59_353 ();
 sg13g2_fill_2 FILLER_59_370 ();
 sg13g2_decap_4 FILLER_59_378 ();
 sg13g2_fill_1 FILLER_59_382 ();
 sg13g2_fill_2 FILLER_59_387 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_411 ();
 sg13g2_fill_2 FILLER_59_417 ();
 sg13g2_fill_1 FILLER_59_475 ();
 sg13g2_decap_4 FILLER_59_480 ();
 sg13g2_fill_1 FILLER_59_484 ();
 sg13g2_fill_2 FILLER_59_503 ();
 sg13g2_fill_2 FILLER_59_525 ();
 sg13g2_fill_1 FILLER_59_527 ();
 sg13g2_fill_1 FILLER_59_541 ();
 sg13g2_decap_8 FILLER_59_552 ();
 sg13g2_fill_2 FILLER_59_559 ();
 sg13g2_fill_1 FILLER_59_595 ();
 sg13g2_fill_2 FILLER_59_601 ();
 sg13g2_fill_2 FILLER_59_623 ();
 sg13g2_fill_2 FILLER_59_636 ();
 sg13g2_fill_1 FILLER_59_638 ();
 sg13g2_fill_1 FILLER_59_668 ();
 sg13g2_fill_1 FILLER_59_680 ();
 sg13g2_fill_1 FILLER_59_686 ();
 sg13g2_fill_2 FILLER_59_693 ();
 sg13g2_decap_4 FILLER_59_712 ();
 sg13g2_fill_1 FILLER_59_716 ();
 sg13g2_decap_8 FILLER_59_751 ();
 sg13g2_fill_1 FILLER_59_758 ();
 sg13g2_fill_1 FILLER_59_763 ();
 sg13g2_decap_8 FILLER_59_788 ();
 sg13g2_fill_1 FILLER_59_795 ();
 sg13g2_fill_2 FILLER_59_821 ();
 sg13g2_fill_1 FILLER_59_823 ();
 sg13g2_fill_1 FILLER_59_840 ();
 sg13g2_decap_8 FILLER_59_850 ();
 sg13g2_decap_4 FILLER_59_857 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_fill_1 FILLER_60_74 ();
 sg13g2_fill_1 FILLER_60_125 ();
 sg13g2_fill_2 FILLER_60_152 ();
 sg13g2_fill_2 FILLER_60_172 ();
 sg13g2_fill_2 FILLER_60_205 ();
 sg13g2_fill_1 FILLER_60_207 ();
 sg13g2_decap_4 FILLER_60_230 ();
 sg13g2_fill_1 FILLER_60_244 ();
 sg13g2_fill_1 FILLER_60_282 ();
 sg13g2_fill_1 FILLER_60_315 ();
 sg13g2_fill_2 FILLER_60_350 ();
 sg13g2_fill_2 FILLER_60_364 ();
 sg13g2_fill_1 FILLER_60_366 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_383 ();
 sg13g2_fill_2 FILLER_60_394 ();
 sg13g2_fill_1 FILLER_60_396 ();
 sg13g2_fill_2 FILLER_60_471 ();
 sg13g2_fill_1 FILLER_60_473 ();
 sg13g2_decap_4 FILLER_60_499 ();
 sg13g2_decap_8 FILLER_60_511 ();
 sg13g2_decap_8 FILLER_60_518 ();
 sg13g2_fill_1 FILLER_60_525 ();
 sg13g2_decap_8 FILLER_60_538 ();
 sg13g2_decap_4 FILLER_60_550 ();
 sg13g2_fill_2 FILLER_60_554 ();
 sg13g2_decap_8 FILLER_60_576 ();
 sg13g2_decap_4 FILLER_60_583 ();
 sg13g2_fill_2 FILLER_60_593 ();
 sg13g2_fill_1 FILLER_60_600 ();
 sg13g2_decap_8 FILLER_60_606 ();
 sg13g2_fill_1 FILLER_60_613 ();
 sg13g2_fill_2 FILLER_60_627 ();
 sg13g2_fill_2 FILLER_60_662 ();
 sg13g2_fill_1 FILLER_60_664 ();
 sg13g2_decap_4 FILLER_60_680 ();
 sg13g2_fill_1 FILLER_60_684 ();
 sg13g2_decap_4 FILLER_60_697 ();
 sg13g2_decap_4 FILLER_60_713 ();
 sg13g2_fill_1 FILLER_60_717 ();
 sg13g2_decap_4 FILLER_60_723 ();
 sg13g2_fill_1 FILLER_60_742 ();
 sg13g2_decap_8 FILLER_60_749 ();
 sg13g2_decap_8 FILLER_60_756 ();
 sg13g2_decap_4 FILLER_60_763 ();
 sg13g2_fill_2 FILLER_60_767 ();
 sg13g2_decap_4 FILLER_60_787 ();
 sg13g2_decap_4 FILLER_60_800 ();
 sg13g2_fill_1 FILLER_60_804 ();
 sg13g2_fill_1 FILLER_60_813 ();
 sg13g2_decap_4 FILLER_60_837 ();
 sg13g2_fill_1 FILLER_60_841 ();
 sg13g2_decap_8 FILLER_60_855 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_decap_4 FILLER_61_15 ();
 sg13g2_fill_2 FILLER_61_28 ();
 sg13g2_fill_1 FILLER_61_30 ();
 sg13g2_fill_2 FILLER_61_64 ();
 sg13g2_fill_2 FILLER_61_76 ();
 sg13g2_fill_2 FILLER_61_87 ();
 sg13g2_fill_2 FILLER_61_129 ();
 sg13g2_fill_1 FILLER_61_157 ();
 sg13g2_fill_2 FILLER_61_184 ();
 sg13g2_fill_1 FILLER_61_192 ();
 sg13g2_fill_1 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_273 ();
 sg13g2_fill_1 FILLER_61_341 ();
 sg13g2_fill_2 FILLER_61_360 ();
 sg13g2_fill_1 FILLER_61_367 ();
 sg13g2_fill_1 FILLER_61_378 ();
 sg13g2_fill_1 FILLER_61_414 ();
 sg13g2_fill_1 FILLER_61_423 ();
 sg13g2_fill_2 FILLER_61_452 ();
 sg13g2_fill_1 FILLER_61_470 ();
 sg13g2_fill_1 FILLER_61_504 ();
 sg13g2_fill_2 FILLER_61_525 ();
 sg13g2_fill_1 FILLER_61_527 ();
 sg13g2_decap_8 FILLER_61_538 ();
 sg13g2_decap_8 FILLER_61_568 ();
 sg13g2_decap_4 FILLER_61_575 ();
 sg13g2_fill_2 FILLER_61_590 ();
 sg13g2_fill_1 FILLER_61_608 ();
 sg13g2_decap_4 FILLER_61_632 ();
 sg13g2_fill_2 FILLER_61_636 ();
 sg13g2_fill_2 FILLER_61_652 ();
 sg13g2_fill_1 FILLER_61_659 ();
 sg13g2_fill_1 FILLER_61_678 ();
 sg13g2_decap_8 FILLER_61_691 ();
 sg13g2_decap_8 FILLER_61_698 ();
 sg13g2_fill_2 FILLER_61_721 ();
 sg13g2_decap_8 FILLER_61_777 ();
 sg13g2_fill_1 FILLER_61_784 ();
 sg13g2_fill_1 FILLER_61_821 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_8 FILLER_61_851 ();
 sg13g2_decap_4 FILLER_61_858 ();
 sg13g2_fill_2 FILLER_62_31 ();
 sg13g2_fill_1 FILLER_62_33 ();
 sg13g2_fill_1 FILLER_62_38 ();
 sg13g2_fill_1 FILLER_62_75 ();
 sg13g2_fill_2 FILLER_62_89 ();
 sg13g2_fill_2 FILLER_62_96 ();
 sg13g2_fill_1 FILLER_62_129 ();
 sg13g2_fill_1 FILLER_62_136 ();
 sg13g2_fill_2 FILLER_62_146 ();
 sg13g2_fill_2 FILLER_62_157 ();
 sg13g2_fill_1 FILLER_62_159 ();
 sg13g2_fill_2 FILLER_62_169 ();
 sg13g2_fill_1 FILLER_62_171 ();
 sg13g2_fill_2 FILLER_62_211 ();
 sg13g2_fill_1 FILLER_62_257 ();
 sg13g2_fill_1 FILLER_62_297 ();
 sg13g2_fill_2 FILLER_62_402 ();
 sg13g2_fill_1 FILLER_62_430 ();
 sg13g2_fill_1 FILLER_62_436 ();
 sg13g2_fill_2 FILLER_62_442 ();
 sg13g2_fill_1 FILLER_62_444 ();
 sg13g2_decap_8 FILLER_62_461 ();
 sg13g2_fill_1 FILLER_62_482 ();
 sg13g2_fill_2 FILLER_62_497 ();
 sg13g2_fill_1 FILLER_62_499 ();
 sg13g2_fill_1 FILLER_62_509 ();
 sg13g2_decap_4 FILLER_62_519 ();
 sg13g2_fill_1 FILLER_62_523 ();
 sg13g2_fill_1 FILLER_62_570 ();
 sg13g2_fill_2 FILLER_62_576 ();
 sg13g2_fill_1 FILLER_62_578 ();
 sg13g2_fill_1 FILLER_62_591 ();
 sg13g2_fill_2 FILLER_62_607 ();
 sg13g2_fill_1 FILLER_62_609 ();
 sg13g2_decap_4 FILLER_62_627 ();
 sg13g2_fill_1 FILLER_62_635 ();
 sg13g2_fill_2 FILLER_62_641 ();
 sg13g2_decap_4 FILLER_62_647 ();
 sg13g2_fill_2 FILLER_62_682 ();
 sg13g2_fill_1 FILLER_62_684 ();
 sg13g2_fill_2 FILLER_62_695 ();
 sg13g2_decap_4 FILLER_62_726 ();
 sg13g2_fill_2 FILLER_62_736 ();
 sg13g2_decap_8 FILLER_62_748 ();
 sg13g2_fill_2 FILLER_62_762 ();
 sg13g2_fill_2 FILLER_62_784 ();
 sg13g2_fill_1 FILLER_62_786 ();
 sg13g2_fill_2 FILLER_62_807 ();
 sg13g2_fill_1 FILLER_62_809 ();
 sg13g2_fill_2 FILLER_62_836 ();
 sg13g2_fill_1 FILLER_62_838 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_4 FILLER_63_17 ();
 sg13g2_fill_2 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_65 ();
 sg13g2_fill_1 FILLER_63_67 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_fill_2 FILLER_63_117 ();
 sg13g2_fill_2 FILLER_63_157 ();
 sg13g2_fill_1 FILLER_63_159 ();
 sg13g2_fill_1 FILLER_63_164 ();
 sg13g2_fill_2 FILLER_63_186 ();
 sg13g2_fill_2 FILLER_63_196 ();
 sg13g2_fill_2 FILLER_63_206 ();
 sg13g2_fill_1 FILLER_63_208 ();
 sg13g2_fill_2 FILLER_63_235 ();
 sg13g2_fill_2 FILLER_63_241 ();
 sg13g2_fill_1 FILLER_63_243 ();
 sg13g2_fill_1 FILLER_63_263 ();
 sg13g2_fill_1 FILLER_63_278 ();
 sg13g2_fill_1 FILLER_63_329 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_fill_2 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_63_423 ();
 sg13g2_fill_2 FILLER_63_436 ();
 sg13g2_fill_2 FILLER_63_471 ();
 sg13g2_decap_4 FILLER_63_487 ();
 sg13g2_fill_1 FILLER_63_491 ();
 sg13g2_fill_2 FILLER_63_501 ();
 sg13g2_fill_2 FILLER_63_521 ();
 sg13g2_fill_2 FILLER_63_529 ();
 sg13g2_fill_1 FILLER_63_531 ();
 sg13g2_decap_8 FILLER_63_541 ();
 sg13g2_fill_1 FILLER_63_548 ();
 sg13g2_fill_2 FILLER_63_559 ();
 sg13g2_fill_1 FILLER_63_561 ();
 sg13g2_fill_1 FILLER_63_571 ();
 sg13g2_decap_4 FILLER_63_592 ();
 sg13g2_fill_1 FILLER_63_612 ();
 sg13g2_decap_4 FILLER_63_623 ();
 sg13g2_decap_8 FILLER_63_642 ();
 sg13g2_fill_1 FILLER_63_649 ();
 sg13g2_decap_4 FILLER_63_657 ();
 sg13g2_fill_2 FILLER_63_670 ();
 sg13g2_decap_8 FILLER_63_690 ();
 sg13g2_fill_2 FILLER_63_697 ();
 sg13g2_fill_1 FILLER_63_699 ();
 sg13g2_fill_2 FILLER_63_711 ();
 sg13g2_fill_1 FILLER_63_713 ();
 sg13g2_fill_2 FILLER_63_730 ();
 sg13g2_decap_8 FILLER_63_756 ();
 sg13g2_fill_1 FILLER_63_763 ();
 sg13g2_fill_1 FILLER_63_768 ();
 sg13g2_fill_2 FILLER_63_784 ();
 sg13g2_fill_1 FILLER_63_786 ();
 sg13g2_fill_2 FILLER_63_791 ();
 sg13g2_fill_1 FILLER_63_793 ();
 sg13g2_fill_2 FILLER_63_806 ();
 sg13g2_fill_1 FILLER_63_808 ();
 sg13g2_decap_8 FILLER_63_842 ();
 sg13g2_decap_8 FILLER_63_849 ();
 sg13g2_decap_4 FILLER_63_856 ();
 sg13g2_fill_2 FILLER_63_860 ();
 sg13g2_fill_1 FILLER_64_31 ();
 sg13g2_fill_1 FILLER_64_77 ();
 sg13g2_fill_2 FILLER_64_133 ();
 sg13g2_fill_1 FILLER_64_135 ();
 sg13g2_fill_1 FILLER_64_157 ();
 sg13g2_fill_2 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_175 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_decap_4 FILLER_64_232 ();
 sg13g2_fill_2 FILLER_64_236 ();
 sg13g2_decap_4 FILLER_64_242 ();
 sg13g2_fill_2 FILLER_64_317 ();
 sg13g2_fill_1 FILLER_64_383 ();
 sg13g2_fill_1 FILLER_64_393 ();
 sg13g2_fill_2 FILLER_64_417 ();
 sg13g2_fill_2 FILLER_64_447 ();
 sg13g2_fill_1 FILLER_64_458 ();
 sg13g2_fill_2 FILLER_64_466 ();
 sg13g2_fill_1 FILLER_64_468 ();
 sg13g2_fill_2 FILLER_64_490 ();
 sg13g2_fill_2 FILLER_64_527 ();
 sg13g2_fill_1 FILLER_64_529 ();
 sg13g2_fill_2 FILLER_64_548 ();
 sg13g2_decap_8 FILLER_64_560 ();
 sg13g2_fill_2 FILLER_64_567 ();
 sg13g2_fill_2 FILLER_64_574 ();
 sg13g2_fill_2 FILLER_64_586 ();
 sg13g2_fill_2 FILLER_64_593 ();
 sg13g2_fill_2 FILLER_64_605 ();
 sg13g2_decap_4 FILLER_64_621 ();
 sg13g2_fill_2 FILLER_64_625 ();
 sg13g2_fill_1 FILLER_64_641 ();
 sg13g2_fill_2 FILLER_64_664 ();
 sg13g2_decap_4 FILLER_64_718 ();
 sg13g2_fill_2 FILLER_64_735 ();
 sg13g2_fill_1 FILLER_64_737 ();
 sg13g2_fill_2 FILLER_64_790 ();
 sg13g2_decap_8 FILLER_64_833 ();
 sg13g2_decap_8 FILLER_64_840 ();
 sg13g2_decap_8 FILLER_64_847 ();
 sg13g2_decap_8 FILLER_64_854 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_15 ();
 sg13g2_fill_1 FILLER_65_24 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_fill_1 FILLER_65_92 ();
 sg13g2_decap_4 FILLER_65_107 ();
 sg13g2_decap_8 FILLER_65_114 ();
 sg13g2_fill_2 FILLER_65_121 ();
 sg13g2_fill_1 FILLER_65_123 ();
 sg13g2_fill_1 FILLER_65_137 ();
 sg13g2_fill_2 FILLER_65_143 ();
 sg13g2_fill_1 FILLER_65_145 ();
 sg13g2_fill_1 FILLER_65_150 ();
 sg13g2_fill_1 FILLER_65_159 ();
 sg13g2_fill_1 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_4 FILLER_65_208 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_fill_2 FILLER_65_250 ();
 sg13g2_fill_1 FILLER_65_252 ();
 sg13g2_fill_1 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_277 ();
 sg13g2_fill_1 FILLER_65_300 ();
 sg13g2_fill_1 FILLER_65_357 ();
 sg13g2_fill_1 FILLER_65_428 ();
 sg13g2_fill_2 FILLER_65_450 ();
 sg13g2_fill_1 FILLER_65_452 ();
 sg13g2_fill_2 FILLER_65_462 ();
 sg13g2_fill_1 FILLER_65_469 ();
 sg13g2_decap_4 FILLER_65_483 ();
 sg13g2_decap_8 FILLER_65_492 ();
 sg13g2_fill_2 FILLER_65_499 ();
 sg13g2_fill_1 FILLER_65_501 ();
 sg13g2_fill_2 FILLER_65_511 ();
 sg13g2_fill_1 FILLER_65_513 ();
 sg13g2_decap_4 FILLER_65_522 ();
 sg13g2_fill_2 FILLER_65_570 ();
 sg13g2_fill_1 FILLER_65_572 ();
 sg13g2_decap_8 FILLER_65_601 ();
 sg13g2_fill_1 FILLER_65_608 ();
 sg13g2_decap_8 FILLER_65_627 ();
 sg13g2_fill_1 FILLER_65_634 ();
 sg13g2_decap_8 FILLER_65_651 ();
 sg13g2_decap_4 FILLER_65_662 ();
 sg13g2_fill_2 FILLER_65_666 ();
 sg13g2_fill_2 FILLER_65_676 ();
 sg13g2_decap_8 FILLER_65_687 ();
 sg13g2_fill_1 FILLER_65_694 ();
 sg13g2_fill_1 FILLER_65_706 ();
 sg13g2_decap_4 FILLER_65_713 ();
 sg13g2_fill_1 FILLER_65_717 ();
 sg13g2_decap_4 FILLER_65_724 ();
 sg13g2_fill_1 FILLER_65_728 ();
 sg13g2_fill_2 FILLER_65_734 ();
 sg13g2_decap_4 FILLER_65_740 ();
 sg13g2_fill_2 FILLER_65_744 ();
 sg13g2_fill_2 FILLER_65_759 ();
 sg13g2_fill_2 FILLER_65_776 ();
 sg13g2_decap_4 FILLER_65_789 ();
 sg13g2_fill_2 FILLER_65_793 ();
 sg13g2_decap_8 FILLER_65_812 ();
 sg13g2_fill_2 FILLER_65_819 ();
 sg13g2_fill_1 FILLER_65_821 ();
 sg13g2_decap_8 FILLER_65_834 ();
 sg13g2_decap_8 FILLER_65_841 ();
 sg13g2_decap_8 FILLER_65_848 ();
 sg13g2_decap_8 FILLER_65_855 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_17 ();
 sg13g2_decap_8 FILLER_66_40 ();
 sg13g2_fill_1 FILLER_66_47 ();
 sg13g2_decap_8 FILLER_66_58 ();
 sg13g2_fill_2 FILLER_66_65 ();
 sg13g2_fill_1 FILLER_66_67 ();
 sg13g2_fill_2 FILLER_66_90 ();
 sg13g2_fill_1 FILLER_66_92 ();
 sg13g2_decap_4 FILLER_66_131 ();
 sg13g2_fill_1 FILLER_66_135 ();
 sg13g2_decap_8 FILLER_66_163 ();
 sg13g2_fill_2 FILLER_66_170 ();
 sg13g2_fill_1 FILLER_66_196 ();
 sg13g2_fill_2 FILLER_66_207 ();
 sg13g2_decap_8 FILLER_66_229 ();
 sg13g2_fill_2 FILLER_66_236 ();
 sg13g2_fill_1 FILLER_66_238 ();
 sg13g2_fill_2 FILLER_66_244 ();
 sg13g2_fill_2 FILLER_66_270 ();
 sg13g2_fill_2 FILLER_66_294 ();
 sg13g2_fill_2 FILLER_66_301 ();
 sg13g2_fill_2 FILLER_66_342 ();
 sg13g2_fill_1 FILLER_66_344 ();
 sg13g2_decap_4 FILLER_66_353 ();
 sg13g2_fill_2 FILLER_66_357 ();
 sg13g2_fill_2 FILLER_66_429 ();
 sg13g2_fill_1 FILLER_66_431 ();
 sg13g2_fill_2 FILLER_66_436 ();
 sg13g2_fill_2 FILLER_66_490 ();
 sg13g2_fill_1 FILLER_66_492 ();
 sg13g2_decap_8 FILLER_66_523 ();
 sg13g2_fill_2 FILLER_66_530 ();
 sg13g2_fill_1 FILLER_66_532 ();
 sg13g2_decap_8 FILLER_66_547 ();
 sg13g2_fill_2 FILLER_66_564 ();
 sg13g2_fill_2 FILLER_66_576 ();
 sg13g2_fill_2 FILLER_66_599 ();
 sg13g2_fill_2 FILLER_66_623 ();
 sg13g2_fill_2 FILLER_66_636 ();
 sg13g2_decap_4 FILLER_66_654 ();
 sg13g2_fill_1 FILLER_66_658 ();
 sg13g2_fill_2 FILLER_66_675 ();
 sg13g2_fill_1 FILLER_66_677 ();
 sg13g2_fill_2 FILLER_66_688 ();
 sg13g2_fill_1 FILLER_66_690 ();
 sg13g2_decap_4 FILLER_66_716 ();
 sg13g2_fill_2 FILLER_66_720 ();
 sg13g2_decap_4 FILLER_66_728 ();
 sg13g2_fill_2 FILLER_66_736 ();
 sg13g2_fill_1 FILLER_66_738 ();
 sg13g2_decap_4 FILLER_66_753 ();
 sg13g2_fill_2 FILLER_66_757 ();
 sg13g2_fill_2 FILLER_66_791 ();
 sg13g2_fill_1 FILLER_66_793 ();
 sg13g2_fill_2 FILLER_66_817 ();
 sg13g2_fill_1 FILLER_66_819 ();
 sg13g2_decap_8 FILLER_66_834 ();
 sg13g2_decap_8 FILLER_66_841 ();
 sg13g2_decap_8 FILLER_66_848 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_19 ();
 sg13g2_decap_8 FILLER_67_46 ();
 sg13g2_fill_2 FILLER_67_53 ();
 sg13g2_fill_1 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_88 ();
 sg13g2_fill_1 FILLER_67_90 ();
 sg13g2_decap_8 FILLER_67_96 ();
 sg13g2_fill_1 FILLER_67_103 ();
 sg13g2_decap_4 FILLER_67_121 ();
 sg13g2_fill_1 FILLER_67_125 ();
 sg13g2_decap_4 FILLER_67_141 ();
 sg13g2_fill_2 FILLER_67_145 ();
 sg13g2_fill_2 FILLER_67_167 ();
 sg13g2_fill_1 FILLER_67_169 ();
 sg13g2_decap_4 FILLER_67_184 ();
 sg13g2_decap_4 FILLER_67_192 ();
 sg13g2_fill_2 FILLER_67_196 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_decap_4 FILLER_67_234 ();
 sg13g2_fill_1 FILLER_67_271 ();
 sg13g2_fill_2 FILLER_67_291 ();
 sg13g2_fill_2 FILLER_67_337 ();
 sg13g2_fill_1 FILLER_67_339 ();
 sg13g2_fill_1 FILLER_67_366 ();
 sg13g2_fill_2 FILLER_67_376 ();
 sg13g2_fill_1 FILLER_67_378 ();
 sg13g2_fill_1 FILLER_67_413 ();
 sg13g2_fill_2 FILLER_67_420 ();
 sg13g2_fill_1 FILLER_67_422 ();
 sg13g2_decap_8 FILLER_67_437 ();
 sg13g2_decap_4 FILLER_67_444 ();
 sg13g2_fill_1 FILLER_67_448 ();
 sg13g2_decap_8 FILLER_67_455 ();
 sg13g2_fill_2 FILLER_67_462 ();
 sg13g2_fill_1 FILLER_67_464 ();
 sg13g2_decap_8 FILLER_67_471 ();
 sg13g2_decap_8 FILLER_67_495 ();
 sg13g2_fill_2 FILLER_67_525 ();
 sg13g2_fill_1 FILLER_67_527 ();
 sg13g2_fill_1 FILLER_67_536 ();
 sg13g2_fill_1 FILLER_67_547 ();
 sg13g2_decap_8 FILLER_67_575 ();
 sg13g2_fill_1 FILLER_67_582 ();
 sg13g2_decap_4 FILLER_67_587 ();
 sg13g2_fill_1 FILLER_67_591 ();
 sg13g2_fill_2 FILLER_67_597 ();
 sg13g2_fill_1 FILLER_67_599 ();
 sg13g2_decap_8 FILLER_67_636 ();
 sg13g2_decap_4 FILLER_67_643 ();
 sg13g2_fill_2 FILLER_67_647 ();
 sg13g2_decap_8 FILLER_67_679 ();
 sg13g2_decap_4 FILLER_67_686 ();
 sg13g2_fill_1 FILLER_67_716 ();
 sg13g2_decap_8 FILLER_67_745 ();
 sg13g2_fill_2 FILLER_67_773 ();
 sg13g2_decap_8 FILLER_67_794 ();
 sg13g2_fill_1 FILLER_67_821 ();
 sg13g2_decap_8 FILLER_67_830 ();
 sg13g2_decap_8 FILLER_67_837 ();
 sg13g2_decap_8 FILLER_67_844 ();
 sg13g2_decap_8 FILLER_67_851 ();
 sg13g2_decap_4 FILLER_67_858 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_9 ();
 sg13g2_decap_4 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_fill_2 FILLER_68_45 ();
 sg13g2_decap_4 FILLER_68_75 ();
 sg13g2_fill_1 FILLER_68_79 ();
 sg13g2_fill_2 FILLER_68_93 ();
 sg13g2_fill_1 FILLER_68_95 ();
 sg13g2_decap_8 FILLER_68_101 ();
 sg13g2_fill_2 FILLER_68_118 ();
 sg13g2_fill_2 FILLER_68_146 ();
 sg13g2_fill_1 FILLER_68_154 ();
 sg13g2_fill_1 FILLER_68_171 ();
 sg13g2_decap_8 FILLER_68_176 ();
 sg13g2_fill_1 FILLER_68_193 ();
 sg13g2_fill_1 FILLER_68_199 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_216 ();
 sg13g2_decap_4 FILLER_68_223 ();
 sg13g2_fill_2 FILLER_68_227 ();
 sg13g2_fill_2 FILLER_68_343 ();
 sg13g2_fill_1 FILLER_68_345 ();
 sg13g2_fill_2 FILLER_68_352 ();
 sg13g2_fill_1 FILLER_68_354 ();
 sg13g2_fill_2 FILLER_68_364 ();
 sg13g2_fill_1 FILLER_68_389 ();
 sg13g2_fill_2 FILLER_68_417 ();
 sg13g2_fill_1 FILLER_68_419 ();
 sg13g2_fill_2 FILLER_68_446 ();
 sg13g2_fill_1 FILLER_68_448 ();
 sg13g2_fill_1 FILLER_68_474 ();
 sg13g2_fill_2 FILLER_68_497 ();
 sg13g2_decap_4 FILLER_68_519 ();
 sg13g2_fill_1 FILLER_68_529 ();
 sg13g2_decap_8 FILLER_68_536 ();
 sg13g2_fill_1 FILLER_68_543 ();
 sg13g2_fill_2 FILLER_68_591 ();
 sg13g2_fill_1 FILLER_68_605 ();
 sg13g2_fill_1 FILLER_68_612 ();
 sg13g2_fill_2 FILLER_68_617 ();
 sg13g2_fill_1 FILLER_68_619 ();
 sg13g2_decap_8 FILLER_68_639 ();
 sg13g2_fill_2 FILLER_68_646 ();
 sg13g2_decap_4 FILLER_68_662 ();
 sg13g2_fill_1 FILLER_68_666 ();
 sg13g2_decap_4 FILLER_68_713 ();
 sg13g2_fill_2 FILLER_68_722 ();
 sg13g2_fill_2 FILLER_68_730 ();
 sg13g2_fill_2 FILLER_68_759 ();
 sg13g2_fill_2 FILLER_68_767 ();
 sg13g2_fill_1 FILLER_68_769 ();
 sg13g2_fill_1 FILLER_68_782 ();
 sg13g2_decap_4 FILLER_68_791 ();
 sg13g2_fill_1 FILLER_68_795 ();
 sg13g2_decap_8 FILLER_68_808 ();
 sg13g2_decap_8 FILLER_68_815 ();
 sg13g2_decap_8 FILLER_68_822 ();
 sg13g2_decap_8 FILLER_68_829 ();
 sg13g2_decap_8 FILLER_68_836 ();
 sg13g2_decap_8 FILLER_68_843 ();
 sg13g2_decap_8 FILLER_68_850 ();
 sg13g2_decap_4 FILLER_68_857 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_fill_1 FILLER_69_30 ();
 sg13g2_decap_4 FILLER_69_44 ();
 sg13g2_fill_1 FILLER_69_48 ();
 sg13g2_decap_8 FILLER_69_62 ();
 sg13g2_fill_2 FILLER_69_69 ();
 sg13g2_fill_1 FILLER_69_71 ();
 sg13g2_decap_4 FILLER_69_96 ();
 sg13g2_fill_2 FILLER_69_119 ();
 sg13g2_fill_1 FILLER_69_121 ();
 sg13g2_fill_2 FILLER_69_128 ();
 sg13g2_fill_1 FILLER_69_141 ();
 sg13g2_decap_8 FILLER_69_162 ();
 sg13g2_decap_8 FILLER_69_169 ();
 sg13g2_fill_1 FILLER_69_176 ();
 sg13g2_decap_4 FILLER_69_195 ();
 sg13g2_fill_2 FILLER_69_199 ();
 sg13g2_fill_1 FILLER_69_218 ();
 sg13g2_fill_2 FILLER_69_245 ();
 sg13g2_fill_1 FILLER_69_273 ();
 sg13g2_fill_2 FILLER_69_335 ();
 sg13g2_fill_2 FILLER_69_354 ();
 sg13g2_fill_2 FILLER_69_376 ();
 sg13g2_fill_2 FILLER_69_393 ();
 sg13g2_fill_2 FILLER_69_413 ();
 sg13g2_fill_1 FILLER_69_415 ();
 sg13g2_decap_4 FILLER_69_427 ();
 sg13g2_fill_2 FILLER_69_431 ();
 sg13g2_decap_4 FILLER_69_439 ();
 sg13g2_fill_1 FILLER_69_443 ();
 sg13g2_decap_4 FILLER_69_472 ();
 sg13g2_fill_1 FILLER_69_476 ();
 sg13g2_fill_2 FILLER_69_493 ();
 sg13g2_fill_1 FILLER_69_495 ();
 sg13g2_fill_1 FILLER_69_510 ();
 sg13g2_fill_1 FILLER_69_524 ();
 sg13g2_decap_4 FILLER_69_544 ();
 sg13g2_fill_2 FILLER_69_548 ();
 sg13g2_fill_2 FILLER_69_560 ();
 sg13g2_fill_1 FILLER_69_562 ();
 sg13g2_decap_4 FILLER_69_584 ();
 sg13g2_fill_2 FILLER_69_588 ();
 sg13g2_fill_1 FILLER_69_600 ();
 sg13g2_fill_2 FILLER_69_607 ();
 sg13g2_fill_1 FILLER_69_619 ();
 sg13g2_decap_4 FILLER_69_631 ();
 sg13g2_fill_2 FILLER_69_635 ();
 sg13g2_fill_2 FILLER_69_643 ();
 sg13g2_fill_2 FILLER_69_649 ();
 sg13g2_decap_8 FILLER_69_666 ();
 sg13g2_fill_2 FILLER_69_673 ();
 sg13g2_fill_1 FILLER_69_675 ();
 sg13g2_decap_8 FILLER_69_681 ();
 sg13g2_fill_2 FILLER_69_688 ();
 sg13g2_decap_8 FILLER_69_706 ();
 sg13g2_fill_1 FILLER_69_713 ();
 sg13g2_fill_2 FILLER_69_746 ();
 sg13g2_fill_1 FILLER_69_748 ();
 sg13g2_fill_2 FILLER_69_766 ();
 sg13g2_decap_8 FILLER_69_781 ();
 sg13g2_decap_8 FILLER_69_788 ();
 sg13g2_decap_8 FILLER_69_795 ();
 sg13g2_decap_8 FILLER_69_810 ();
 sg13g2_decap_8 FILLER_69_817 ();
 sg13g2_decap_8 FILLER_69_824 ();
 sg13g2_decap_8 FILLER_69_831 ();
 sg13g2_decap_8 FILLER_69_838 ();
 sg13g2_decap_8 FILLER_69_845 ();
 sg13g2_decap_8 FILLER_69_852 ();
 sg13g2_fill_2 FILLER_69_859 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_25 ();
 sg13g2_fill_2 FILLER_70_32 ();
 sg13g2_fill_2 FILLER_70_60 ();
 sg13g2_fill_1 FILLER_70_62 ();
 sg13g2_decap_8 FILLER_70_92 ();
 sg13g2_fill_2 FILLER_70_118 ();
 sg13g2_fill_1 FILLER_70_120 ();
 sg13g2_decap_4 FILLER_70_142 ();
 sg13g2_fill_2 FILLER_70_146 ();
 sg13g2_fill_2 FILLER_70_162 ();
 sg13g2_fill_1 FILLER_70_164 ();
 sg13g2_fill_2 FILLER_70_175 ();
 sg13g2_fill_1 FILLER_70_177 ();
 sg13g2_fill_2 FILLER_70_183 ();
 sg13g2_fill_2 FILLER_70_190 ();
 sg13g2_fill_2 FILLER_70_198 ();
 sg13g2_fill_1 FILLER_70_200 ();
 sg13g2_fill_2 FILLER_70_212 ();
 sg13g2_fill_2 FILLER_70_291 ();
 sg13g2_fill_2 FILLER_70_304 ();
 sg13g2_fill_2 FILLER_70_323 ();
 sg13g2_fill_2 FILLER_70_348 ();
 sg13g2_fill_2 FILLER_70_369 ();
 sg13g2_fill_2 FILLER_70_444 ();
 sg13g2_fill_2 FILLER_70_472 ();
 sg13g2_decap_8 FILLER_70_482 ();
 sg13g2_fill_2 FILLER_70_489 ();
 sg13g2_fill_2 FILLER_70_502 ();
 sg13g2_fill_2 FILLER_70_515 ();
 sg13g2_fill_1 FILLER_70_548 ();
 sg13g2_fill_1 FILLER_70_558 ();
 sg13g2_fill_2 FILLER_70_575 ();
 sg13g2_fill_1 FILLER_70_577 ();
 sg13g2_decap_8 FILLER_70_602 ();
 sg13g2_fill_2 FILLER_70_633 ();
 sg13g2_fill_2 FILLER_70_640 ();
 sg13g2_fill_1 FILLER_70_662 ();
 sg13g2_fill_1 FILLER_70_672 ();
 sg13g2_decap_8 FILLER_70_679 ();
 sg13g2_decap_4 FILLER_70_686 ();
 sg13g2_fill_1 FILLER_70_690 ();
 sg13g2_fill_1 FILLER_70_698 ();
 sg13g2_decap_4 FILLER_70_709 ();
 sg13g2_fill_2 FILLER_70_713 ();
 sg13g2_decap_4 FILLER_70_727 ();
 sg13g2_fill_1 FILLER_70_731 ();
 sg13g2_fill_2 FILLER_70_740 ();
 sg13g2_decap_8 FILLER_70_747 ();
 sg13g2_decap_8 FILLER_70_754 ();
 sg13g2_decap_8 FILLER_70_761 ();
 sg13g2_decap_8 FILLER_70_768 ();
 sg13g2_decap_8 FILLER_70_775 ();
 sg13g2_decap_8 FILLER_70_782 ();
 sg13g2_decap_8 FILLER_70_789 ();
 sg13g2_decap_8 FILLER_70_796 ();
 sg13g2_decap_8 FILLER_70_803 ();
 sg13g2_decap_8 FILLER_70_810 ();
 sg13g2_decap_8 FILLER_70_817 ();
 sg13g2_decap_8 FILLER_70_824 ();
 sg13g2_decap_8 FILLER_70_831 ();
 sg13g2_decap_8 FILLER_70_838 ();
 sg13g2_decap_8 FILLER_70_845 ();
 sg13g2_decap_8 FILLER_70_852 ();
 sg13g2_fill_2 FILLER_70_859 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_18 ();
 sg13g2_fill_2 FILLER_71_28 ();
 sg13g2_fill_1 FILLER_71_46 ();
 sg13g2_fill_2 FILLER_71_67 ();
 sg13g2_fill_1 FILLER_71_69 ();
 sg13g2_decap_8 FILLER_71_74 ();
 sg13g2_fill_1 FILLER_71_81 ();
 sg13g2_decap_4 FILLER_71_90 ();
 sg13g2_fill_2 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_fill_1 FILLER_71_128 ();
 sg13g2_fill_2 FILLER_71_150 ();
 sg13g2_fill_1 FILLER_71_152 ();
 sg13g2_fill_2 FILLER_71_159 ();
 sg13g2_fill_1 FILLER_71_161 ();
 sg13g2_fill_2 FILLER_71_167 ();
 sg13g2_fill_1 FILLER_71_169 ();
 sg13g2_fill_1 FILLER_71_185 ();
 sg13g2_decap_4 FILLER_71_195 ();
 sg13g2_fill_1 FILLER_71_199 ();
 sg13g2_decap_4 FILLER_71_209 ();
 sg13g2_fill_2 FILLER_71_213 ();
 sg13g2_fill_1 FILLER_71_264 ();
 sg13g2_fill_1 FILLER_71_277 ();
 sg13g2_fill_1 FILLER_71_354 ();
 sg13g2_fill_2 FILLER_71_395 ();
 sg13g2_fill_1 FILLER_71_411 ();
 sg13g2_decap_8 FILLER_71_433 ();
 sg13g2_fill_2 FILLER_71_440 ();
 sg13g2_fill_2 FILLER_71_499 ();
 sg13g2_fill_2 FILLER_71_506 ();
 sg13g2_fill_1 FILLER_71_528 ();
 sg13g2_fill_2 FILLER_71_534 ();
 sg13g2_fill_2 FILLER_71_545 ();
 sg13g2_fill_1 FILLER_71_547 ();
 sg13g2_fill_1 FILLER_71_574 ();
 sg13g2_decap_8 FILLER_71_596 ();
 sg13g2_fill_2 FILLER_71_603 ();
 sg13g2_fill_2 FILLER_71_639 ();
 sg13g2_fill_2 FILLER_71_713 ();
 sg13g2_fill_1 FILLER_71_715 ();
 sg13g2_decap_8 FILLER_71_732 ();
 sg13g2_decap_8 FILLER_71_739 ();
 sg13g2_decap_8 FILLER_71_746 ();
 sg13g2_decap_8 FILLER_71_753 ();
 sg13g2_decap_8 FILLER_71_760 ();
 sg13g2_decap_8 FILLER_71_767 ();
 sg13g2_decap_8 FILLER_71_774 ();
 sg13g2_decap_8 FILLER_71_781 ();
 sg13g2_decap_8 FILLER_71_788 ();
 sg13g2_decap_8 FILLER_71_795 ();
 sg13g2_decap_8 FILLER_71_802 ();
 sg13g2_decap_8 FILLER_71_809 ();
 sg13g2_decap_8 FILLER_71_816 ();
 sg13g2_decap_8 FILLER_71_823 ();
 sg13g2_decap_8 FILLER_71_830 ();
 sg13g2_decap_8 FILLER_71_837 ();
 sg13g2_decap_8 FILLER_71_844 ();
 sg13g2_decap_8 FILLER_71_851 ();
 sg13g2_decap_4 FILLER_71_858 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_18 ();
 sg13g2_decap_8 FILLER_72_27 ();
 sg13g2_decap_4 FILLER_72_34 ();
 sg13g2_fill_2 FILLER_72_38 ();
 sg13g2_fill_1 FILLER_72_53 ();
 sg13g2_decap_8 FILLER_72_62 ();
 sg13g2_fill_2 FILLER_72_69 ();
 sg13g2_fill_1 FILLER_72_71 ();
 sg13g2_fill_1 FILLER_72_80 ();
 sg13g2_fill_1 FILLER_72_95 ();
 sg13g2_fill_2 FILLER_72_104 ();
 sg13g2_fill_1 FILLER_72_106 ();
 sg13g2_decap_4 FILLER_72_125 ();
 sg13g2_fill_2 FILLER_72_129 ();
 sg13g2_fill_2 FILLER_72_157 ();
 sg13g2_decap_4 FILLER_72_168 ();
 sg13g2_fill_1 FILLER_72_180 ();
 sg13g2_fill_1 FILLER_72_185 ();
 sg13g2_fill_2 FILLER_72_212 ();
 sg13g2_fill_1 FILLER_72_240 ();
 sg13g2_fill_1 FILLER_72_344 ();
 sg13g2_decap_4 FILLER_72_428 ();
 sg13g2_fill_1 FILLER_72_465 ();
 sg13g2_decap_8 FILLER_72_491 ();
 sg13g2_fill_2 FILLER_72_498 ();
 sg13g2_fill_2 FILLER_72_512 ();
 sg13g2_fill_1 FILLER_72_514 ();
 sg13g2_fill_2 FILLER_72_535 ();
 sg13g2_fill_1 FILLER_72_537 ();
 sg13g2_fill_2 FILLER_72_542 ();
 sg13g2_decap_4 FILLER_72_563 ();
 sg13g2_fill_1 FILLER_72_574 ();
 sg13g2_fill_1 FILLER_72_581 ();
 sg13g2_fill_2 FILLER_72_596 ();
 sg13g2_fill_2 FILLER_72_607 ();
 sg13g2_fill_1 FILLER_72_609 ();
 sg13g2_fill_1 FILLER_72_628 ();
 sg13g2_decap_4 FILLER_72_634 ();
 sg13g2_fill_1 FILLER_72_638 ();
 sg13g2_fill_2 FILLER_72_650 ();
 sg13g2_fill_1 FILLER_72_652 ();
 sg13g2_decap_4 FILLER_72_686 ();
 sg13g2_fill_2 FILLER_72_698 ();
 sg13g2_fill_1 FILLER_72_700 ();
 sg13g2_decap_8 FILLER_72_727 ();
 sg13g2_decap_8 FILLER_72_734 ();
 sg13g2_decap_8 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_748 ();
 sg13g2_decap_8 FILLER_72_755 ();
 sg13g2_decap_8 FILLER_72_762 ();
 sg13g2_decap_8 FILLER_72_769 ();
 sg13g2_decap_8 FILLER_72_776 ();
 sg13g2_decap_8 FILLER_72_783 ();
 sg13g2_decap_8 FILLER_72_790 ();
 sg13g2_decap_8 FILLER_72_797 ();
 sg13g2_decap_8 FILLER_72_804 ();
 sg13g2_decap_8 FILLER_72_811 ();
 sg13g2_decap_8 FILLER_72_818 ();
 sg13g2_decap_8 FILLER_72_825 ();
 sg13g2_decap_8 FILLER_72_832 ();
 sg13g2_decap_8 FILLER_72_839 ();
 sg13g2_decap_8 FILLER_72_846 ();
 sg13g2_decap_8 FILLER_72_853 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_7 ();
 sg13g2_decap_4 FILLER_73_32 ();
 sg13g2_fill_2 FILLER_73_36 ();
 sg13g2_fill_1 FILLER_73_46 ();
 sg13g2_decap_8 FILLER_73_57 ();
 sg13g2_decap_4 FILLER_73_64 ();
 sg13g2_fill_2 FILLER_73_68 ();
 sg13g2_decap_4 FILLER_73_104 ();
 sg13g2_fill_1 FILLER_73_108 ();
 sg13g2_fill_2 FILLER_73_119 ();
 sg13g2_fill_1 FILLER_73_121 ();
 sg13g2_decap_8 FILLER_73_144 ();
 sg13g2_decap_4 FILLER_73_151 ();
 sg13g2_fill_2 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_170 ();
 sg13g2_fill_2 FILLER_73_187 ();
 sg13g2_fill_2 FILLER_73_209 ();
 sg13g2_fill_1 FILLER_73_211 ();
 sg13g2_fill_2 FILLER_73_221 ();
 sg13g2_fill_1 FILLER_73_223 ();
 sg13g2_fill_1 FILLER_73_305 ();
 sg13g2_fill_2 FILLER_73_335 ();
 sg13g2_fill_1 FILLER_73_381 ();
 sg13g2_fill_2 FILLER_73_400 ();
 sg13g2_fill_1 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_73_414 ();
 sg13g2_decap_4 FILLER_73_425 ();
 sg13g2_fill_2 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_73_447 ();
 sg13g2_decap_4 FILLER_73_454 ();
 sg13g2_fill_1 FILLER_73_458 ();
 sg13g2_fill_2 FILLER_73_469 ();
 sg13g2_fill_2 FILLER_73_507 ();
 sg13g2_fill_1 FILLER_73_509 ();
 sg13g2_decap_8 FILLER_73_519 ();
 sg13g2_fill_1 FILLER_73_526 ();
 sg13g2_fill_2 FILLER_73_551 ();
 sg13g2_fill_1 FILLER_73_553 ();
 sg13g2_fill_1 FILLER_73_561 ();
 sg13g2_decap_8 FILLER_73_567 ();
 sg13g2_decap_4 FILLER_73_574 ();
 sg13g2_fill_1 FILLER_73_578 ();
 sg13g2_decap_4 FILLER_73_587 ();
 sg13g2_fill_1 FILLER_73_591 ();
 sg13g2_decap_4 FILLER_73_633 ();
 sg13g2_fill_2 FILLER_73_650 ();
 sg13g2_fill_1 FILLER_73_652 ();
 sg13g2_decap_4 FILLER_73_661 ();
 sg13g2_fill_2 FILLER_73_665 ();
 sg13g2_fill_1 FILLER_73_693 ();
 sg13g2_fill_2 FILLER_73_703 ();
 sg13g2_fill_1 FILLER_73_705 ();
 sg13g2_decap_8 FILLER_73_711 ();
 sg13g2_decap_8 FILLER_73_718 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_decap_8 FILLER_73_732 ();
 sg13g2_decap_8 FILLER_73_739 ();
 sg13g2_decap_8 FILLER_73_746 ();
 sg13g2_decap_8 FILLER_73_753 ();
 sg13g2_decap_8 FILLER_73_760 ();
 sg13g2_decap_8 FILLER_73_767 ();
 sg13g2_decap_8 FILLER_73_774 ();
 sg13g2_decap_8 FILLER_73_781 ();
 sg13g2_decap_8 FILLER_73_788 ();
 sg13g2_decap_8 FILLER_73_795 ();
 sg13g2_decap_8 FILLER_73_802 ();
 sg13g2_decap_8 FILLER_73_809 ();
 sg13g2_decap_8 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_830 ();
 sg13g2_decap_8 FILLER_73_837 ();
 sg13g2_decap_8 FILLER_73_844 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_decap_4 FILLER_73_858 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_36 ();
 sg13g2_fill_2 FILLER_74_40 ();
 sg13g2_decap_4 FILLER_74_71 ();
 sg13g2_decap_8 FILLER_74_92 ();
 sg13g2_decap_8 FILLER_74_99 ();
 sg13g2_decap_4 FILLER_74_106 ();
 sg13g2_fill_2 FILLER_74_127 ();
 sg13g2_fill_2 FILLER_74_133 ();
 sg13g2_fill_2 FILLER_74_140 ();
 sg13g2_fill_2 FILLER_74_179 ();
 sg13g2_fill_1 FILLER_74_181 ();
 sg13g2_fill_2 FILLER_74_245 ();
 sg13g2_fill_1 FILLER_74_247 ();
 sg13g2_fill_1 FILLER_74_295 ();
 sg13g2_fill_1 FILLER_74_306 ();
 sg13g2_fill_2 FILLER_74_337 ();
 sg13g2_fill_2 FILLER_74_368 ();
 sg13g2_fill_1 FILLER_74_375 ();
 sg13g2_fill_1 FILLER_74_424 ();
 sg13g2_decap_4 FILLER_74_438 ();
 sg13g2_fill_1 FILLER_74_446 ();
 sg13g2_fill_1 FILLER_74_464 ();
 sg13g2_fill_1 FILLER_74_541 ();
 sg13g2_fill_1 FILLER_74_553 ();
 sg13g2_decap_8 FILLER_74_560 ();
 sg13g2_decap_4 FILLER_74_567 ();
 sg13g2_fill_1 FILLER_74_587 ();
 sg13g2_decap_8 FILLER_74_612 ();
 sg13g2_fill_2 FILLER_74_619 ();
 sg13g2_decap_8 FILLER_74_626 ();
 sg13g2_decap_4 FILLER_74_633 ();
 sg13g2_fill_1 FILLER_74_637 ();
 sg13g2_decap_8 FILLER_74_651 ();
 sg13g2_decap_8 FILLER_74_658 ();
 sg13g2_decap_8 FILLER_74_665 ();
 sg13g2_fill_1 FILLER_74_672 ();
 sg13g2_decap_8 FILLER_74_678 ();
 sg13g2_decap_8 FILLER_74_685 ();
 sg13g2_decap_8 FILLER_74_692 ();
 sg13g2_decap_8 FILLER_74_699 ();
 sg13g2_decap_8 FILLER_74_706 ();
 sg13g2_decap_8 FILLER_74_713 ();
 sg13g2_decap_8 FILLER_74_720 ();
 sg13g2_decap_8 FILLER_74_727 ();
 sg13g2_decap_8 FILLER_74_734 ();
 sg13g2_decap_8 FILLER_74_741 ();
 sg13g2_decap_8 FILLER_74_748 ();
 sg13g2_decap_8 FILLER_74_755 ();
 sg13g2_decap_8 FILLER_74_762 ();
 sg13g2_decap_8 FILLER_74_769 ();
 sg13g2_decap_8 FILLER_74_776 ();
 sg13g2_decap_8 FILLER_74_783 ();
 sg13g2_decap_8 FILLER_74_790 ();
 sg13g2_decap_8 FILLER_74_797 ();
 sg13g2_decap_8 FILLER_74_804 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_decap_8 FILLER_74_818 ();
 sg13g2_decap_8 FILLER_74_825 ();
 sg13g2_decap_8 FILLER_74_832 ();
 sg13g2_decap_8 FILLER_74_839 ();
 sg13g2_decap_8 FILLER_74_846 ();
 sg13g2_decap_8 FILLER_74_853 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_51 ();
 sg13g2_fill_1 FILLER_75_53 ();
 sg13g2_fill_1 FILLER_75_58 ();
 sg13g2_decap_8 FILLER_75_73 ();
 sg13g2_fill_1 FILLER_75_106 ();
 sg13g2_fill_2 FILLER_75_118 ();
 sg13g2_fill_1 FILLER_75_120 ();
 sg13g2_fill_1 FILLER_75_129 ();
 sg13g2_fill_2 FILLER_75_156 ();
 sg13g2_decap_8 FILLER_75_162 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_decap_4 FILLER_75_177 ();
 sg13g2_fill_1 FILLER_75_191 ();
 sg13g2_fill_2 FILLER_75_239 ();
 sg13g2_fill_1 FILLER_75_246 ();
 sg13g2_decap_4 FILLER_75_424 ();
 sg13g2_fill_1 FILLER_75_442 ();
 sg13g2_fill_1 FILLER_75_460 ();
 sg13g2_fill_2 FILLER_75_477 ();
 sg13g2_fill_2 FILLER_75_483 ();
 sg13g2_decap_8 FILLER_75_532 ();
 sg13g2_fill_1 FILLER_75_539 ();
 sg13g2_fill_2 FILLER_75_588 ();
 sg13g2_fill_1 FILLER_75_590 ();
 sg13g2_fill_2 FILLER_75_599 ();
 sg13g2_decap_8 FILLER_75_627 ();
 sg13g2_decap_8 FILLER_75_634 ();
 sg13g2_decap_8 FILLER_75_641 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_decap_8 FILLER_75_655 ();
 sg13g2_decap_8 FILLER_75_662 ();
 sg13g2_decap_8 FILLER_75_669 ();
 sg13g2_decap_8 FILLER_75_676 ();
 sg13g2_decap_8 FILLER_75_683 ();
 sg13g2_decap_8 FILLER_75_690 ();
 sg13g2_decap_8 FILLER_75_697 ();
 sg13g2_decap_8 FILLER_75_704 ();
 sg13g2_decap_8 FILLER_75_711 ();
 sg13g2_decap_8 FILLER_75_718 ();
 sg13g2_decap_8 FILLER_75_725 ();
 sg13g2_decap_8 FILLER_75_732 ();
 sg13g2_decap_8 FILLER_75_739 ();
 sg13g2_decap_8 FILLER_75_746 ();
 sg13g2_decap_8 FILLER_75_753 ();
 sg13g2_decap_8 FILLER_75_760 ();
 sg13g2_decap_8 FILLER_75_767 ();
 sg13g2_decap_8 FILLER_75_774 ();
 sg13g2_decap_8 FILLER_75_781 ();
 sg13g2_decap_8 FILLER_75_788 ();
 sg13g2_decap_8 FILLER_75_795 ();
 sg13g2_decap_8 FILLER_75_802 ();
 sg13g2_decap_8 FILLER_75_809 ();
 sg13g2_decap_8 FILLER_75_816 ();
 sg13g2_decap_8 FILLER_75_823 ();
 sg13g2_decap_8 FILLER_75_830 ();
 sg13g2_decap_8 FILLER_75_837 ();
 sg13g2_decap_8 FILLER_75_844 ();
 sg13g2_decap_8 FILLER_75_851 ();
 sg13g2_decap_4 FILLER_75_858 ();
 sg13g2_decap_4 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_4 ();
 sg13g2_fill_2 FILLER_76_50 ();
 sg13g2_fill_1 FILLER_76_52 ();
 sg13g2_fill_2 FILLER_76_73 ();
 sg13g2_fill_1 FILLER_76_91 ();
 sg13g2_fill_2 FILLER_76_105 ();
 sg13g2_fill_2 FILLER_76_116 ();
 sg13g2_fill_1 FILLER_76_118 ();
 sg13g2_fill_1 FILLER_76_132 ();
 sg13g2_decap_4 FILLER_76_149 ();
 sg13g2_fill_2 FILLER_76_158 ();
 sg13g2_fill_1 FILLER_76_170 ();
 sg13g2_fill_2 FILLER_76_188 ();
 sg13g2_fill_2 FILLER_76_205 ();
 sg13g2_fill_2 FILLER_76_217 ();
 sg13g2_fill_2 FILLER_76_260 ();
 sg13g2_fill_1 FILLER_76_262 ();
 sg13g2_fill_2 FILLER_76_308 ();
 sg13g2_fill_1 FILLER_76_379 ();
 sg13g2_fill_1 FILLER_76_393 ();
 sg13g2_fill_2 FILLER_76_403 ();
 sg13g2_fill_2 FILLER_76_422 ();
 sg13g2_fill_2 FILLER_76_476 ();
 sg13g2_fill_1 FILLER_76_503 ();
 sg13g2_fill_2 FILLER_76_509 ();
 sg13g2_fill_2 FILLER_76_521 ();
 sg13g2_fill_1 FILLER_76_523 ();
 sg13g2_fill_2 FILLER_76_532 ();
 sg13g2_fill_2 FILLER_76_552 ();
 sg13g2_fill_2 FILLER_76_585 ();
 sg13g2_decap_8 FILLER_76_608 ();
 sg13g2_decap_8 FILLER_76_615 ();
 sg13g2_decap_8 FILLER_76_622 ();
 sg13g2_decap_8 FILLER_76_629 ();
 sg13g2_decap_8 FILLER_76_636 ();
 sg13g2_decap_8 FILLER_76_643 ();
 sg13g2_decap_8 FILLER_76_650 ();
 sg13g2_decap_8 FILLER_76_657 ();
 sg13g2_decap_8 FILLER_76_664 ();
 sg13g2_decap_8 FILLER_76_671 ();
 sg13g2_decap_8 FILLER_76_678 ();
 sg13g2_decap_8 FILLER_76_685 ();
 sg13g2_decap_8 FILLER_76_692 ();
 sg13g2_decap_8 FILLER_76_699 ();
 sg13g2_decap_8 FILLER_76_706 ();
 sg13g2_decap_8 FILLER_76_713 ();
 sg13g2_decap_8 FILLER_76_720 ();
 sg13g2_decap_8 FILLER_76_727 ();
 sg13g2_decap_8 FILLER_76_734 ();
 sg13g2_decap_8 FILLER_76_741 ();
 sg13g2_decap_8 FILLER_76_748 ();
 sg13g2_decap_8 FILLER_76_755 ();
 sg13g2_decap_8 FILLER_76_762 ();
 sg13g2_decap_8 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_776 ();
 sg13g2_decap_8 FILLER_76_783 ();
 sg13g2_decap_8 FILLER_76_790 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_804 ();
 sg13g2_decap_8 FILLER_76_811 ();
 sg13g2_decap_8 FILLER_76_818 ();
 sg13g2_decap_8 FILLER_76_825 ();
 sg13g2_decap_8 FILLER_76_832 ();
 sg13g2_decap_8 FILLER_76_839 ();
 sg13g2_decap_8 FILLER_76_846 ();
 sg13g2_decap_8 FILLER_76_853 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_7 ();
 sg13g2_fill_1 FILLER_77_9 ();
 sg13g2_decap_8 FILLER_77_18 ();
 sg13g2_decap_8 FILLER_77_25 ();
 sg13g2_decap_4 FILLER_77_32 ();
 sg13g2_fill_1 FILLER_77_61 ();
 sg13g2_fill_1 FILLER_77_66 ();
 sg13g2_decap_8 FILLER_77_74 ();
 sg13g2_fill_2 FILLER_77_81 ();
 sg13g2_decap_8 FILLER_77_106 ();
 sg13g2_fill_2 FILLER_77_136 ();
 sg13g2_fill_1 FILLER_77_138 ();
 sg13g2_fill_2 FILLER_77_144 ();
 sg13g2_fill_2 FILLER_77_161 ();
 sg13g2_decap_4 FILLER_77_173 ();
 sg13g2_fill_2 FILLER_77_248 ();
 sg13g2_fill_2 FILLER_77_306 ();
 sg13g2_fill_2 FILLER_77_339 ();
 sg13g2_decap_4 FILLER_77_401 ();
 sg13g2_fill_1 FILLER_77_405 ();
 sg13g2_fill_2 FILLER_77_432 ();
 sg13g2_fill_1 FILLER_77_455 ();
 sg13g2_fill_2 FILLER_77_466 ();
 sg13g2_fill_2 FILLER_77_474 ();
 sg13g2_decap_8 FILLER_77_558 ();
 sg13g2_decap_8 FILLER_77_565 ();
 sg13g2_decap_8 FILLER_77_572 ();
 sg13g2_fill_1 FILLER_77_579 ();
 sg13g2_decap_8 FILLER_77_589 ();
 sg13g2_decap_8 FILLER_77_596 ();
 sg13g2_decap_8 FILLER_77_603 ();
 sg13g2_decap_8 FILLER_77_610 ();
 sg13g2_decap_8 FILLER_77_617 ();
 sg13g2_decap_8 FILLER_77_624 ();
 sg13g2_decap_8 FILLER_77_631 ();
 sg13g2_decap_8 FILLER_77_638 ();
 sg13g2_decap_8 FILLER_77_645 ();
 sg13g2_decap_8 FILLER_77_652 ();
 sg13g2_decap_8 FILLER_77_659 ();
 sg13g2_decap_8 FILLER_77_666 ();
 sg13g2_decap_8 FILLER_77_673 ();
 sg13g2_decap_8 FILLER_77_680 ();
 sg13g2_decap_8 FILLER_77_687 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_decap_8 FILLER_77_701 ();
 sg13g2_decap_8 FILLER_77_708 ();
 sg13g2_decap_8 FILLER_77_715 ();
 sg13g2_decap_8 FILLER_77_722 ();
 sg13g2_decap_8 FILLER_77_729 ();
 sg13g2_decap_8 FILLER_77_736 ();
 sg13g2_decap_8 FILLER_77_743 ();
 sg13g2_decap_8 FILLER_77_750 ();
 sg13g2_decap_8 FILLER_77_757 ();
 sg13g2_decap_8 FILLER_77_764 ();
 sg13g2_decap_8 FILLER_77_771 ();
 sg13g2_decap_8 FILLER_77_778 ();
 sg13g2_decap_8 FILLER_77_785 ();
 sg13g2_decap_8 FILLER_77_792 ();
 sg13g2_decap_8 FILLER_77_799 ();
 sg13g2_decap_8 FILLER_77_806 ();
 sg13g2_decap_8 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_820 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_decap_8 FILLER_77_834 ();
 sg13g2_decap_8 FILLER_77_841 ();
 sg13g2_decap_8 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_855 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_26 ();
 sg13g2_fill_1 FILLER_78_28 ();
 sg13g2_decap_4 FILLER_78_46 ();
 sg13g2_decap_4 FILLER_78_64 ();
 sg13g2_fill_1 FILLER_78_77 ();
 sg13g2_decap_4 FILLER_78_98 ();
 sg13g2_fill_2 FILLER_78_102 ();
 sg13g2_fill_2 FILLER_78_111 ();
 sg13g2_fill_2 FILLER_78_132 ();
 sg13g2_fill_1 FILLER_78_237 ();
 sg13g2_fill_1 FILLER_78_264 ();
 sg13g2_fill_2 FILLER_78_306 ();
 sg13g2_fill_2 FILLER_78_329 ();
 sg13g2_fill_1 FILLER_78_392 ();
 sg13g2_fill_1 FILLER_78_545 ();
 sg13g2_decap_4 FILLER_78_555 ();
 sg13g2_fill_1 FILLER_78_559 ();
 sg13g2_decap_8 FILLER_78_568 ();
 sg13g2_decap_8 FILLER_78_575 ();
 sg13g2_decap_8 FILLER_78_582 ();
 sg13g2_decap_8 FILLER_78_589 ();
 sg13g2_decap_8 FILLER_78_596 ();
 sg13g2_decap_8 FILLER_78_603 ();
 sg13g2_decap_8 FILLER_78_610 ();
 sg13g2_decap_8 FILLER_78_617 ();
 sg13g2_decap_8 FILLER_78_624 ();
 sg13g2_decap_8 FILLER_78_631 ();
 sg13g2_decap_8 FILLER_78_638 ();
 sg13g2_decap_8 FILLER_78_645 ();
 sg13g2_decap_8 FILLER_78_652 ();
 sg13g2_decap_8 FILLER_78_659 ();
 sg13g2_decap_8 FILLER_78_666 ();
 sg13g2_decap_8 FILLER_78_673 ();
 sg13g2_decap_8 FILLER_78_680 ();
 sg13g2_decap_8 FILLER_78_687 ();
 sg13g2_decap_8 FILLER_78_694 ();
 sg13g2_decap_8 FILLER_78_701 ();
 sg13g2_decap_8 FILLER_78_708 ();
 sg13g2_decap_8 FILLER_78_715 ();
 sg13g2_decap_8 FILLER_78_722 ();
 sg13g2_decap_8 FILLER_78_729 ();
 sg13g2_decap_8 FILLER_78_736 ();
 sg13g2_decap_8 FILLER_78_743 ();
 sg13g2_decap_8 FILLER_78_750 ();
 sg13g2_decap_8 FILLER_78_757 ();
 sg13g2_decap_8 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_771 ();
 sg13g2_decap_8 FILLER_78_778 ();
 sg13g2_decap_8 FILLER_78_785 ();
 sg13g2_decap_8 FILLER_78_792 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_806 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_8 FILLER_78_820 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_9 ();
 sg13g2_decap_8 FILLER_79_18 ();
 sg13g2_fill_2 FILLER_79_25 ();
 sg13g2_fill_2 FILLER_79_53 ();
 sg13g2_decap_8 FILLER_79_89 ();
 sg13g2_fill_1 FILLER_79_126 ();
 sg13g2_fill_1 FILLER_79_191 ();
 sg13g2_fill_1 FILLER_79_201 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_fill_2 FILLER_79_335 ();
 sg13g2_fill_2 FILLER_79_372 ();
 sg13g2_fill_2 FILLER_79_506 ();
 sg13g2_decap_8 FILLER_79_547 ();
 sg13g2_decap_8 FILLER_79_554 ();
 sg13g2_decap_8 FILLER_79_561 ();
 sg13g2_decap_8 FILLER_79_568 ();
 sg13g2_decap_8 FILLER_79_575 ();
 sg13g2_decap_8 FILLER_79_582 ();
 sg13g2_decap_8 FILLER_79_589 ();
 sg13g2_decap_8 FILLER_79_596 ();
 sg13g2_decap_8 FILLER_79_603 ();
 sg13g2_decap_8 FILLER_79_610 ();
 sg13g2_decap_8 FILLER_79_617 ();
 sg13g2_decap_8 FILLER_79_624 ();
 sg13g2_decap_8 FILLER_79_631 ();
 sg13g2_decap_8 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_645 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_8 FILLER_79_659 ();
 sg13g2_decap_8 FILLER_79_666 ();
 sg13g2_decap_8 FILLER_79_673 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_687 ();
 sg13g2_decap_8 FILLER_79_694 ();
 sg13g2_decap_8 FILLER_79_701 ();
 sg13g2_decap_8 FILLER_79_708 ();
 sg13g2_decap_8 FILLER_79_715 ();
 sg13g2_decap_8 FILLER_79_722 ();
 sg13g2_decap_8 FILLER_79_729 ();
 sg13g2_decap_8 FILLER_79_736 ();
 sg13g2_decap_8 FILLER_79_743 ();
 sg13g2_decap_8 FILLER_79_750 ();
 sg13g2_decap_8 FILLER_79_757 ();
 sg13g2_decap_8 FILLER_79_764 ();
 sg13g2_decap_8 FILLER_79_771 ();
 sg13g2_decap_8 FILLER_79_778 ();
 sg13g2_decap_8 FILLER_79_785 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_827 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_fill_2 FILLER_80_35 ();
 sg13g2_fill_1 FILLER_80_37 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_fill_2 FILLER_80_49 ();
 sg13g2_fill_1 FILLER_80_51 ();
 sg13g2_fill_2 FILLER_80_78 ();
 sg13g2_fill_2 FILLER_80_111 ();
 sg13g2_fill_2 FILLER_80_175 ();
 sg13g2_fill_2 FILLER_80_260 ();
 sg13g2_fill_1 FILLER_80_309 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_fill_1 FILLER_80_426 ();
 sg13g2_decap_8 FILLER_80_435 ();
 sg13g2_decap_4 FILLER_80_442 ();
 sg13g2_fill_1 FILLER_80_446 ();
 sg13g2_fill_2 FILLER_80_454 ();
 sg13g2_fill_1 FILLER_80_491 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_decap_8 FILLER_80_547 ();
 sg13g2_decap_8 FILLER_80_554 ();
 sg13g2_decap_8 FILLER_80_561 ();
 sg13g2_decap_8 FILLER_80_568 ();
 sg13g2_decap_8 FILLER_80_575 ();
 sg13g2_decap_8 FILLER_80_582 ();
 sg13g2_decap_8 FILLER_80_589 ();
 sg13g2_decap_8 FILLER_80_596 ();
 sg13g2_decap_8 FILLER_80_603 ();
 sg13g2_decap_8 FILLER_80_610 ();
 sg13g2_decap_8 FILLER_80_617 ();
 sg13g2_decap_8 FILLER_80_624 ();
 sg13g2_decap_8 FILLER_80_631 ();
 sg13g2_decap_8 FILLER_80_638 ();
 sg13g2_decap_8 FILLER_80_645 ();
 sg13g2_decap_8 FILLER_80_652 ();
 sg13g2_decap_8 FILLER_80_659 ();
 sg13g2_decap_8 FILLER_80_666 ();
 sg13g2_decap_8 FILLER_80_673 ();
 sg13g2_decap_8 FILLER_80_680 ();
 sg13g2_decap_8 FILLER_80_687 ();
 sg13g2_decap_8 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_701 ();
 sg13g2_decap_8 FILLER_80_708 ();
 sg13g2_decap_8 FILLER_80_715 ();
 sg13g2_decap_8 FILLER_80_722 ();
 sg13g2_decap_8 FILLER_80_729 ();
 sg13g2_decap_8 FILLER_80_736 ();
 sg13g2_decap_8 FILLER_80_743 ();
 sg13g2_decap_8 FILLER_80_750 ();
 sg13g2_decap_8 FILLER_80_757 ();
 sg13g2_decap_8 FILLER_80_764 ();
 sg13g2_decap_8 FILLER_80_771 ();
 sg13g2_decap_8 FILLER_80_778 ();
 sg13g2_decap_8 FILLER_80_785 ();
 sg13g2_decap_8 FILLER_80_792 ();
 sg13g2_decap_8 FILLER_80_799 ();
 sg13g2_decap_8 FILLER_80_806 ();
 sg13g2_decap_8 FILLER_80_813 ();
 sg13g2_decap_8 FILLER_80_820 ();
 sg13g2_decap_8 FILLER_80_827 ();
 sg13g2_decap_8 FILLER_80_834 ();
 sg13g2_decap_8 FILLER_80_841 ();
 sg13g2_decap_8 FILLER_80_848 ();
 sg13g2_decap_8 FILLER_80_855 ();
endmodule

module tt_um_brandonramos_VGA_Pong_with_NES_Controllers (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \Pong.b ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[0] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[10] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[11] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[12] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[13] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[14] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[15] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[16] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[17] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[18] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[1] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[2] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[3] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[4] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[5] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[6] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[7] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[8] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[9] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[0] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[10] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[11] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[12] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[13] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[14] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[15] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[16] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[17] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[18] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[1] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[2] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[3] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[4] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[5] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[6] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[7] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[8] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[9] ;
 wire \Pong.control_unit.state_ballMovement[0] ;
 wire \Pong.control_unit.state_ballMovement[1] ;
 wire \Pong.control_unit.state_ballMovement[2] ;
 wire \Pong.control_unit.state_ballMovement[3] ;
 wire \Pong.control_unit.state_ballMovement[4] ;
 wire \Pong.datapath.Ball_Clock.Q[0] ;
 wire \Pong.datapath.Ball_Clock.Q[10] ;
 wire \Pong.datapath.Ball_Clock.Q[11] ;
 wire \Pong.datapath.Ball_Clock.Q[12] ;
 wire \Pong.datapath.Ball_Clock.Q[13] ;
 wire \Pong.datapath.Ball_Clock.Q[14] ;
 wire \Pong.datapath.Ball_Clock.Q[15] ;
 wire \Pong.datapath.Ball_Clock.Q[16] ;
 wire \Pong.datapath.Ball_Clock.Q[1] ;
 wire \Pong.datapath.Ball_Clock.Q[2] ;
 wire \Pong.datapath.Ball_Clock.Q[3] ;
 wire \Pong.datapath.Ball_Clock.Q[4] ;
 wire \Pong.datapath.Ball_Clock.Q[5] ;
 wire \Pong.datapath.Ball_Clock.Q[6] ;
 wire \Pong.datapath.Ball_Clock.Q[7] ;
 wire \Pong.datapath.Ball_Clock.Q[8] ;
 wire \Pong.datapath.Ball_Clock.Q[9] ;
 wire \Pong.datapath.Ball_Clock.roll ;
 wire \Pong.datapath.NES_activity_Left[2] ;
 wire \Pong.datapath.NES_activity_Left[3] ;
 wire \Pong.datapath.NES_activity_Left[4] ;
 wire \Pong.datapath.NES_activity_Left[5] ;
 wire \Pong.datapath.NES_activity_Right[2] ;
 wire \Pong.datapath.NES_activity_Right[3] ;
 wire \Pong.datapath.NES_activity_Right[4] ;
 wire \Pong.datapath.NES_activity_Right[5] ;
 wire \Pong.datapath.NES_counter_left.Q[0] ;
 wire \Pong.datapath.NES_counter_left.Q[1] ;
 wire \Pong.datapath.NES_counter_left.Q[2] ;
 wire \Pong.datapath.NES_counter_left.Q[3] ;
 wire \Pong.datapath.NES_counter_left.Q[4] ;
 wire \Pong.datapath.NES_counter_left.Q[5] ;
 wire \Pong.datapath.NES_counter_left.Q[6] ;
 wire \Pong.datapath.NES_counter_left.Q[7] ;
 wire \Pong.datapath.NES_counter_right.Q[0] ;
 wire \Pong.datapath.NES_counter_right.Q[1] ;
 wire \Pong.datapath.NES_counter_right.Q[2] ;
 wire \Pong.datapath.NES_counter_right.Q[3] ;
 wire \Pong.datapath.NES_counter_right.Q[4] ;
 wire \Pong.datapath.NES_counter_right.Q[5] ;
 wire \Pong.datapath.NES_counter_right.Q[6] ;
 wire \Pong.datapath.NES_counter_right.Q[7] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[0] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[10] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[11] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[12] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[13] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[14] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[15] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[16] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[17] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[18] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[1] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[2] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[3] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[4] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[5] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[6] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[7] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[8] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[9] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[0] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[10] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[11] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[12] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[13] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[14] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[15] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[16] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[17] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[18] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[1] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[2] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[3] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[4] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[5] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[6] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[7] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[8] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[9] ;
 wire \Pong.datapath.NES_wire_Left[2] ;
 wire \Pong.datapath.NES_wire_Left[3] ;
 wire \Pong.datapath.NES_wire_Left[4] ;
 wire \Pong.datapath.NES_wire_Left[5] ;
 wire \Pong.datapath.NES_wire_Right[2] ;
 wire \Pong.datapath.NES_wire_Right[3] ;
 wire \Pong.datapath.NES_wire_Right[4] ;
 wire \Pong.datapath.NES_wire_Right[5] ;
 wire \Pong.datapath.ballFunction.ball_center_x[0] ;
 wire \Pong.datapath.ballFunction.ball_center_x[1] ;
 wire \Pong.datapath.ballFunction.ball_center_x[2] ;
 wire \Pong.datapath.ballFunction.ball_center_x[3] ;
 wire \Pong.datapath.ballFunction.ball_center_x[4] ;
 wire \Pong.datapath.ballFunction.ball_center_x[5] ;
 wire \Pong.datapath.ballFunction.ball_center_x[6] ;
 wire \Pong.datapath.ballFunction.ball_center_x[7] ;
 wire \Pong.datapath.ballFunction.ball_center_x[8] ;
 wire \Pong.datapath.ballFunction.ball_center_x[9] ;
 wire \Pong.datapath.ballFunction.ball_center_y[0] ;
 wire \Pong.datapath.ballFunction.ball_center_y[1] ;
 wire \Pong.datapath.ballFunction.ball_center_y[2] ;
 wire \Pong.datapath.ballFunction.ball_center_y[3] ;
 wire \Pong.datapath.ballFunction.ball_center_y[4] ;
 wire \Pong.datapath.ballFunction.ball_center_y[5] ;
 wire \Pong.datapath.ballFunction.ball_center_y[6] ;
 wire \Pong.datapath.ballFunction.ball_center_y[7] ;
 wire \Pong.datapath.ballFunction.ball_center_y[8] ;
 wire \Pong.datapath.ballFunction.ball_center_y[9] ;
 wire \Pong.datapath.ballFunction.reset_n ;
 wire \Pong.datapath.h_sync ;
 wire \Pong.datapath.leftPaddle[0] ;
 wire \Pong.datapath.leftPaddle[1] ;
 wire \Pong.datapath.leftPaddle[2] ;
 wire \Pong.datapath.leftPaddle[3] ;
 wire \Pong.datapath.leftPaddle[4] ;
 wire \Pong.datapath.leftPaddle[5] ;
 wire \Pong.datapath.leftPaddle[6] ;
 wire \Pong.datapath.leftPaddle[7] ;
 wire \Pong.datapath.leftPaddle[8] ;
 wire \Pong.datapath.leftPaddle[9] ;
 wire \Pong.datapath.old_NES_Left[2] ;
 wire \Pong.datapath.old_NES_Left[3] ;
 wire \Pong.datapath.old_NES_Left[4] ;
 wire \Pong.datapath.old_NES_Left[5] ;
 wire \Pong.datapath.old_NES_Right[2] ;
 wire \Pong.datapath.old_NES_Right[3] ;
 wire \Pong.datapath.old_NES_Right[4] ;
 wire \Pong.datapath.old_NES_Right[5] ;
 wire \Pong.datapath.rightPaddle[0] ;
 wire \Pong.datapath.rightPaddle[1] ;
 wire \Pong.datapath.rightPaddle[2] ;
 wire \Pong.datapath.rightPaddle[3] ;
 wire \Pong.datapath.rightPaddle[4] ;
 wire \Pong.datapath.rightPaddle[5] ;
 wire \Pong.datapath.rightPaddle[6] ;
 wire \Pong.datapath.rightPaddle[7] ;
 wire \Pong.datapath.rightPaddle[8] ;
 wire \Pong.datapath.rightPaddle[9] ;
 wire \Pong.datapath.scoreLeft[0] ;
 wire \Pong.datapath.scoreLeft[1] ;
 wire \Pong.datapath.scoreLeft[2] ;
 wire \Pong.datapath.scoreLeft[3] ;
 wire \Pong.datapath.scoreRight[0] ;
 wire \Pong.datapath.scoreRight[1] ;
 wire \Pong.datapath.scoreRight[2] ;
 wire \Pong.datapath.scoreRight[3] ;
 wire \Pong.datapath.score_flag ;
 wire \Pong.datapath.sw_ballMovement_reg[0] ;
 wire \Pong.datapath.sw_ballMovement_reg[2] ;
 wire \Pong.datapath.sw_ballMovement_reg[3] ;
 wire \Pong.datapath.sw_ballMovement_reg[4] ;
 wire \Pong.datapath.sw_ballMovement_reg[5] ;
 wire \Pong.datapath.v_sync ;
 wire \Pong.datapath.vga.Column_Counter.Q[0] ;
 wire \Pong.datapath.vga.Column_Counter.Q[1] ;
 wire \Pong.datapath.vga.Column_Counter.Q[2] ;
 wire \Pong.datapath.vga.Column_Counter.Q[3] ;
 wire \Pong.datapath.vga.Column_Counter.Q[4] ;
 wire \Pong.datapath.vga.Column_Counter.Q[5] ;
 wire \Pong.datapath.vga.Column_Counter.Q[6] ;
 wire \Pong.datapath.vga.Column_Counter.Q[7] ;
 wire \Pong.datapath.vga.Column_Counter.Q[8] ;
 wire \Pong.datapath.vga.Column_Counter.Q[9] ;
 wire \Pong.datapath.vga.Row_Counter.Q[0] ;
 wire \Pong.datapath.vga.Row_Counter.Q[1] ;
 wire \Pong.datapath.vga.Row_Counter.Q[2] ;
 wire \Pong.datapath.vga.Row_Counter.Q[3] ;
 wire \Pong.datapath.vga.Row_Counter.Q[4] ;
 wire \Pong.datapath.vga.Row_Counter.Q[5] ;
 wire \Pong.datapath.vga.Row_Counter.Q[6] ;
 wire \Pong.datapath.vga.Row_Counter.Q[7] ;
 wire \Pong.datapath.vga.Row_Counter.Q[8] ;
 wire \Pong.datapath.vga.Row_Counter.Q[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net5;
 wire net226;
 wire net227;
 wire net6;
 wire net228;
 wire clknet_0_clk;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;

 sg13g2_inv_1 _2543_ (.Y(_1774_),
    .A(net608));
 sg13g2_inv_2 _2544_ (.Y(_1775_),
    .A(net618));
 sg13g2_inv_2 _2545_ (.Y(_1776_),
    .A(net620));
 sg13g2_inv_2 _2546_ (.Y(_1777_),
    .A(\Pong.datapath.ballFunction.ball_center_y[3] ));
 sg13g2_inv_1 _2547_ (.Y(_1778_),
    .A(\Pong.datapath.Ball_Clock.Q[5] ));
 sg13g2_inv_1 _2548_ (.Y(_1779_),
    .A(\Pong.datapath.Ball_Clock.Q[0] ));
 sg13g2_inv_1 _2549_ (.Y(_1780_),
    .A(net328));
 sg13g2_inv_1 _2550_ (.Y(_1781_),
    .A(net349));
 sg13g2_inv_1 _2551_ (.Y(_1782_),
    .A(net459));
 sg13g2_inv_1 _2552_ (.Y(_1783_),
    .A(net506));
 sg13g2_inv_1 _2553_ (.Y(_1784_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[8] ));
 sg13g2_inv_1 _2554_ (.Y(_1785_),
    .A(net482));
 sg13g2_inv_1 _2555_ (.Y(_1786_),
    .A(net473));
 sg13g2_inv_1 _2556_ (.Y(_1787_),
    .A(net668));
 sg13g2_inv_2 _2557_ (.Y(_1788_),
    .A(net677));
 sg13g2_inv_1 _2558_ (.Y(_1789_),
    .A(net681));
 sg13g2_inv_1 _2559_ (.Y(_1790_),
    .A(net683));
 sg13g2_inv_2 _2560_ (.Y(_1791_),
    .A(net686));
 sg13g2_inv_1 _2561_ (.Y(_1792_),
    .A(net690));
 sg13g2_inv_2 _2562_ (.Y(_1793_),
    .A(net693));
 sg13g2_inv_4 _2563_ (.A(net697),
    .Y(_1794_));
 sg13g2_inv_2 _2564_ (.Y(_1795_),
    .A(net698));
 sg13g2_inv_1 _2565_ (.Y(_1796_),
    .A(net743));
 sg13g2_inv_1 _2566_ (.Y(_1797_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[11] ));
 sg13g2_inv_1 _2567_ (.Y(_1798_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[13] ));
 sg13g2_inv_1 _2568_ (.Y(_1799_),
    .A(\Pong.control_unit.state_ballMovement[3] ));
 sg13g2_inv_1 _2569_ (.Y(_1800_),
    .A(\Pong.control_unit.state_ballMovement[0] ));
 sg13g2_inv_2 _2570_ (.Y(_1801_),
    .A(net433));
 sg13g2_inv_1 _2571_ (.Y(_1802_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ));
 sg13g2_inv_1 _2572_ (.Y(_1803_),
    .A(net337));
 sg13g2_inv_1 _2573_ (.Y(_1804_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[11] ));
 sg13g2_inv_1 _2574_ (.Y(_1805_),
    .A(_0113_));
 sg13g2_inv_1 _2575_ (.Y(_1806_),
    .A(net257));
 sg13g2_inv_1 _2576_ (.Y(_1807_),
    .A(net526));
 sg13g2_inv_2 _2577_ (.Y(_1808_),
    .A(\Pong.datapath.NES_activity_Left[5] ));
 sg13g2_inv_1 _2578_ (.Y(_1809_),
    .A(\Pong.datapath.rightPaddle[8] ));
 sg13g2_inv_2 _2579_ (.Y(_1810_),
    .A(\Pong.datapath.rightPaddle[6] ));
 sg13g2_inv_2 _2580_ (.Y(_1811_),
    .A(\Pong.datapath.rightPaddle[5] ));
 sg13g2_inv_4 _2581_ (.A(\Pong.datapath.rightPaddle[3] ),
    .Y(_1812_));
 sg13g2_inv_2 _2582_ (.Y(_1813_),
    .A(\Pong.datapath.rightPaddle[4] ));
 sg13g2_inv_1 _2583_ (.Y(_1814_),
    .A(_0059_));
 sg13g2_inv_1 _2584_ (.Y(_1815_),
    .A(_0066_));
 sg13g2_inv_1 _2585_ (.Y(_1816_),
    .A(net622));
 sg13g2_inv_2 _2586_ (.Y(_1817_),
    .A(\Pong.datapath.leftPaddle[7] ));
 sg13g2_inv_2 _2587_ (.Y(_1818_),
    .A(net707));
 sg13g2_inv_1 _2588_ (.Y(_1819_),
    .A(net710));
 sg13g2_inv_1 _2589_ (.Y(_1820_),
    .A(\Pong.datapath.leftPaddle[9] ));
 sg13g2_inv_2 _2590_ (.Y(_1821_),
    .A(net718));
 sg13g2_inv_1 _2591_ (.Y(_1822_),
    .A(net721));
 sg13g2_inv_1 _2592_ (.Y(_1823_),
    .A(\Pong.datapath.scoreRight[3] ));
 sg13g2_inv_1 _2593_ (.Y(_1824_),
    .A(net373));
 sg13g2_inv_1 _2594_ (.Y(_1825_),
    .A(net523));
 sg13g2_inv_1 _2595_ (.Y(_1826_),
    .A(\Pong.datapath.NES_activity_Right[2] ));
 sg13g2_inv_2 _2596_ (.Y(_1827_),
    .A(net723));
 sg13g2_inv_1 _2597_ (.Y(_1828_),
    .A(\Pong.datapath.NES_activity_Left[2] ));
 sg13g2_inv_2 _2598_ (.Y(_1829_),
    .A(net705));
 sg13g2_inv_1 _2599_ (.Y(_1830_),
    .A(_0083_));
 sg13g2_inv_1 _2600_ (.Y(_1831_),
    .A(net685));
 sg13g2_inv_1 _2601_ (.Y(_1832_),
    .A(_0092_));
 sg13g2_inv_1 _2602_ (.Y(_1833_),
    .A(_0097_));
 sg13g2_inv_1 _2603_ (.Y(_1834_),
    .A(_0106_));
 sg13g2_nand2b_1 _2604_ (.Y(_1835_),
    .B(\Pong.datapath.NES_counter_left.Q[3] ),
    .A_N(\Pong.datapath.NES_counter_left.Q[2] ));
 sg13g2_nor2_1 _2605_ (.A(\Pong.datapath.NES_counter_left.Q[6] ),
    .B(\Pong.datapath.NES_counter_left.Q[5] ),
    .Y(_1836_));
 sg13g2_nand3_1 _2606_ (.B(\Pong.datapath.NES_counter_left.Q[4] ),
    .C(_1836_),
    .A(\Pong.datapath.NES_counter_left.Q[7] ),
    .Y(_1837_));
 sg13g2_nor4_2 _2607_ (.A(net424),
    .B(\Pong.datapath.NES_counter_left.Q[0] ),
    .C(_1835_),
    .Y(_1838_),
    .D(_1837_));
 sg13g2_nor2_1 _2608_ (.A(net741),
    .B(_1838_),
    .Y(_1839_));
 sg13g2_and2_1 _2609_ (.A(net748),
    .B(_1838_),
    .X(_1840_));
 sg13g2_a22oi_1 _2610_ (.Y(_1841_),
    .B1(net645),
    .B2(net270),
    .A2(net648),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[11] ));
 sg13g2_inv_1 _2611_ (.Y(_0002_),
    .A(net271));
 sg13g2_a22oi_1 _2612_ (.Y(_1842_),
    .B1(net645),
    .B2(net342),
    .A2(net648),
    .A1(net311));
 sg13g2_inv_1 _2613_ (.Y(_0013_),
    .A(_1842_));
 sg13g2_a22oi_1 _2614_ (.Y(_1843_),
    .B1(net647),
    .B2(net261),
    .A2(net650),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[5] ));
 sg13g2_inv_1 _2615_ (.Y(_0014_),
    .A(net262));
 sg13g2_a22oi_1 _2616_ (.Y(_1844_),
    .B1(net646),
    .B2(net384),
    .A2(net649),
    .A1(net381));
 sg13g2_inv_1 _2617_ (.Y(_0017_),
    .A(_1844_));
 sg13g2_a22oi_1 _2618_ (.Y(_1845_),
    .B1(net646),
    .B2(net380),
    .A2(net649),
    .A1(net309));
 sg13g2_inv_1 _2619_ (.Y(_0016_),
    .A(_1845_));
 sg13g2_a22oi_1 _2620_ (.Y(_1846_),
    .B1(net647),
    .B2(net345),
    .A2(net650),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ));
 sg13g2_inv_1 _2621_ (.Y(_0012_),
    .A(net346));
 sg13g2_a22oi_1 _2622_ (.Y(_1847_),
    .B1(net645),
    .B2(net293),
    .A2(net648),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[6] ));
 sg13g2_inv_1 _2623_ (.Y(_0015_),
    .A(net294));
 sg13g2_nand2_2 _2624_ (.Y(_1848_),
    .A(net459),
    .B(\Pong.datapath.NES_delay_counter_left.Q[13] ));
 sg13g2_nand2_2 _2625_ (.Y(_1849_),
    .A(net298),
    .B(\Pong.datapath.NES_delay_counter_left.Q[9] ));
 sg13g2_or2_1 _2626_ (.X(_1850_),
    .B(\Pong.datapath.NES_delay_counter_left.Q[11] ),
    .A(\Pong.datapath.NES_delay_counter_left.Q[12] ));
 sg13g2_nor4_2 _2627_ (.A(\Pong.datapath.NES_delay_counter_left.Q[15] ),
    .B(_1848_),
    .C(_1849_),
    .Y(_1851_),
    .D(_1850_));
 sg13g2_nand2_1 _2628_ (.Y(_1852_),
    .A(net259),
    .B(\Pong.datapath.NES_delay_counter_left.Q[17] ));
 sg13g2_nand4_1 _2629_ (.B(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .C(net539),
    .A(net306),
    .Y(_1853_),
    .D(\Pong.datapath.NES_delay_counter_left.Q[0] ));
 sg13g2_and2_1 _2630_ (.A(\Pong.datapath.NES_delay_counter_left.Q[2] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[1] ),
    .X(_1854_));
 sg13g2_nand3_1 _2631_ (.B(net326),
    .C(_1854_),
    .A(net279),
    .Y(_1855_));
 sg13g2_and4_1 _2632_ (.A(\Pong.datapath.NES_delay_counter_left.Q[6] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[5] ),
    .C(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .D(\Pong.datapath.NES_delay_counter_left.Q[3] ),
    .X(_1856_));
 sg13g2_nand4_1 _2633_ (.B(\Pong.datapath.NES_delay_counter_left.Q[0] ),
    .C(_1854_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[7] ),
    .Y(_1857_),
    .D(_1856_));
 sg13g2_nor4_2 _2634_ (.A(net537),
    .B(net409),
    .C(_1852_),
    .Y(_1858_),
    .D(_1857_));
 sg13g2_nand3_1 _2635_ (.B(_1851_),
    .C(_1858_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[0] ),
    .Y(_1859_));
 sg13g2_inv_2 _2636_ (.Y(_1860_),
    .A(net338));
 sg13g2_a22oi_1 _2637_ (.Y(_1861_),
    .B1(_1860_),
    .B2(net748),
    .A2(net650),
    .A1(net261));
 sg13g2_inv_1 _2638_ (.Y(_0001_),
    .A(_1861_));
 sg13g2_a21oi_1 _2639_ (.A1(_1851_),
    .A2(_1858_),
    .Y(_1862_),
    .B1(_1803_));
 sg13g2_a21oi_2 _2640_ (.B1(net741),
    .Y(_1863_),
    .A2(_1838_),
    .A1(net451));
 sg13g2_nand2b_1 _2641_ (.Y(_0000_),
    .B(net452),
    .A_N(net538));
 sg13g2_a22oi_1 _2642_ (.Y(_1864_),
    .B1(net645),
    .B2(net295),
    .A2(net648),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ));
 sg13g2_inv_1 _2643_ (.Y(_0018_),
    .A(net296));
 sg13g2_a22oi_1 _2644_ (.Y(_1865_),
    .B1(net645),
    .B2(net314),
    .A2(net648),
    .A1(net270));
 sg13g2_inv_1 _2645_ (.Y(_0010_),
    .A(_1865_));
 sg13g2_a22oi_1 _2646_ (.Y(_1866_),
    .B1(net647),
    .B2(net339),
    .A2(net650),
    .A1(net322));
 sg13g2_inv_1 _2647_ (.Y(_0011_),
    .A(_1866_));
 sg13g2_nand2b_1 _2648_ (.Y(_1867_),
    .B(net405),
    .A_N(\Pong.datapath.NES_counter_right.Q[2] ));
 sg13g2_nor2_1 _2649_ (.A(\Pong.datapath.NES_counter_right.Q[6] ),
    .B(\Pong.datapath.NES_counter_right.Q[5] ),
    .Y(_1868_));
 sg13g2_nand3_1 _2650_ (.B(\Pong.datapath.NES_counter_right.Q[4] ),
    .C(_1868_),
    .A(net365),
    .Y(_1869_));
 sg13g2_nor4_2 _2651_ (.A(\Pong.datapath.NES_counter_right.Q[1] ),
    .B(\Pong.datapath.NES_counter_right.Q[0] ),
    .C(_1867_),
    .Y(_1870_),
    .D(_1869_));
 sg13g2_and2_1 _2652_ (.A(net747),
    .B(_1870_),
    .X(_1871_));
 sg13g2_nor2_2 _2653_ (.A(net741),
    .B(_1870_),
    .Y(_1872_));
 sg13g2_a22oi_1 _2654_ (.Y(_1873_),
    .B1(net642),
    .B2(net297),
    .A2(net644),
    .A1(net289));
 sg13g2_inv_1 _2655_ (.Y(_0033_),
    .A(_1873_));
 sg13g2_a22oi_1 _2656_ (.Y(_1874_),
    .B1(net641),
    .B2(net341),
    .A2(net643),
    .A1(net265));
 sg13g2_inv_1 _2657_ (.Y(_0034_),
    .A(_1874_));
 sg13g2_a22oi_1 _2658_ (.Y(_1875_),
    .B1(net642),
    .B2(net263),
    .A2(net644),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[12] ));
 sg13g2_inv_1 _2659_ (.Y(_0035_),
    .A(net264));
 sg13g2_a22oi_1 _2660_ (.Y(_1876_),
    .B1(net641),
    .B2(net394),
    .A2(_1871_),
    .A1(net360));
 sg13g2_inv_1 _2661_ (.Y(_0036_),
    .A(_1876_));
 sg13g2_a22oi_1 _2662_ (.Y(_1877_),
    .B1(_1872_),
    .B2(net278),
    .A2(net643),
    .A1(net272));
 sg13g2_inv_1 _2663_ (.Y(_0037_),
    .A(_1877_));
 sg13g2_nand2_1 _2664_ (.Y(_1878_),
    .A(net255),
    .B(net328));
 sg13g2_nor2_1 _2665_ (.A(\Pong.datapath.NES_delay_counter_right.Q[16] ),
    .B(_1878_),
    .Y(_1879_));
 sg13g2_and2_1 _2666_ (.A(net457),
    .B(net408),
    .X(_1880_));
 sg13g2_nand4_1 _2667_ (.B(\Pong.datapath.NES_delay_counter_right.Q[2] ),
    .C(\Pong.datapath.NES_delay_counter_right.Q[1] ),
    .A(net267),
    .Y(_1881_),
    .D(\Pong.datapath.NES_delay_counter_right.Q[0] ));
 sg13g2_nand4_1 _2668_ (.B(\Pong.datapath.NES_delay_counter_right.Q[6] ),
    .C(\Pong.datapath.NES_delay_counter_right.Q[5] ),
    .A(\Pong.datapath.NES_delay_counter_right.Q[7] ),
    .Y(_1882_),
    .D(\Pong.datapath.NES_delay_counter_right.Q[4] ));
 sg13g2_or2_1 _2669_ (.X(_1883_),
    .B(_1882_),
    .A(_1881_));
 sg13g2_nor2_1 _2670_ (.A(\Pong.datapath.NES_delay_counter_right.Q[12] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[11] ),
    .Y(_1884_));
 sg13g2_and2_1 _2671_ (.A(\Pong.datapath.NES_delay_counter_right.Q[14] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[13] ),
    .X(_1885_));
 sg13g2_nand2_1 _2672_ (.Y(_1886_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[10] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[9] ));
 sg13g2_nor4_1 _2673_ (.A(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[8] ),
    .C(_1883_),
    .D(_1886_),
    .Y(_1887_));
 sg13g2_nand3_1 _2674_ (.B(_1885_),
    .C(_1887_),
    .A(_1884_),
    .Y(_1888_));
 sg13g2_nor3_1 _2675_ (.A(\Pong.datapath.NES_delay_counter_right.Q[16] ),
    .B(_1878_),
    .C(_1888_),
    .Y(_1889_));
 sg13g2_nand2_1 _2676_ (.Y(_1890_),
    .A(net289),
    .B(net642));
 sg13g2_nor2b_1 _2677_ (.A(\Pong.datapath.NES_delay_counter_right.Q[11] ),
    .B_N(\Pong.datapath.NES_delay_counter_right.Q[10] ),
    .Y(_1891_));
 sg13g2_nor2_1 _2678_ (.A(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[12] ),
    .Y(_1892_));
 sg13g2_nand4_1 _2679_ (.B(_1885_),
    .C(_1891_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[9] ),
    .Y(_1893_),
    .D(_1892_));
 sg13g2_nor3_1 _2680_ (.A(\Pong.datapath.NES_delay_counter_right.Q[8] ),
    .B(_1883_),
    .C(_1893_),
    .Y(_1894_));
 sg13g2_nand3_1 _2681_ (.B(_1879_),
    .C(_1894_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[0] ),
    .Y(_1895_));
 sg13g2_o21ai_1 _2682_ (.B1(_1890_),
    .Y(_0020_),
    .A1(net741),
    .A2(_1895_));
 sg13g2_a22oi_1 _2683_ (.Y(_1896_),
    .B1(_1872_),
    .B2(net265),
    .A2(net643),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ));
 sg13g2_inv_1 _2684_ (.Y(_0021_),
    .A(net266));
 sg13g2_a22oi_1 _2685_ (.Y(_1897_),
    .B1(net642),
    .B2(net276),
    .A2(net644),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[2] ));
 sg13g2_inv_1 _2686_ (.Y(_0022_),
    .A(net277));
 sg13g2_a22oi_1 _2687_ (.Y(_1898_),
    .B1(net641),
    .B2(net360),
    .A2(_1871_),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ));
 sg13g2_inv_1 _2688_ (.Y(_0023_),
    .A(net361));
 sg13g2_a22oi_1 _2689_ (.Y(_1899_),
    .B1(net641),
    .B2(net272),
    .A2(net643),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[4] ));
 sg13g2_inv_1 _2690_ (.Y(_0024_),
    .A(net273));
 sg13g2_a22oi_1 _2691_ (.Y(_1900_),
    .B1(net642),
    .B2(net333),
    .A2(net644),
    .A1(net297));
 sg13g2_inv_1 _2692_ (.Y(_0025_),
    .A(_1900_));
 sg13g2_a22oi_1 _2693_ (.Y(_1901_),
    .B1(net642),
    .B2(net340),
    .A2(net644),
    .A1(net263));
 sg13g2_inv_1 _2694_ (.Y(_0026_),
    .A(_1901_));
 sg13g2_nand2_2 _2695_ (.Y(_1902_),
    .A(net623),
    .B(net624));
 sg13g2_nand4_1 _2696_ (.B(\Pong.datapath.ballFunction.ball_center_y[4] ),
    .C(net624),
    .A(_1774_),
    .Y(_1903_),
    .D(net632));
 sg13g2_nor4_1 _2697_ (.A(net613),
    .B(net615),
    .C(net618),
    .D(\Pong.datapath.ballFunction.ball_center_y[5] ),
    .Y(_1904_));
 sg13g2_nor2_2 _2698_ (.A(net626),
    .B(net628),
    .Y(_1905_));
 sg13g2_o21ai_1 _2699_ (.B1(_1904_),
    .Y(_1906_),
    .A1(_1902_),
    .A2(_1905_));
 sg13g2_a21oi_2 _2700_ (.B1(_1906_),
    .Y(_0043_),
    .A2(_1903_),
    .A1(_1805_));
 sg13g2_nand2_1 _2701_ (.Y(_1907_),
    .A(net745),
    .B(\Pong.control_unit.state_ballMovement[0] ));
 sg13g2_nor2_1 _2702_ (.A(\Pong.datapath.sw_ballMovement_reg[3] ),
    .B(_1907_),
    .Y(_1908_));
 sg13g2_nor2b_1 _2703_ (.A(\Pong.datapath.sw_ballMovement_reg[3] ),
    .B_N(\Pong.control_unit.state_ballMovement[2] ),
    .Y(_1909_));
 sg13g2_nor2_1 _2704_ (.A(net738),
    .B(\Pong.datapath.sw_ballMovement_reg[2] ),
    .Y(_1910_));
 sg13g2_and2_1 _2705_ (.A(_1909_),
    .B(_1910_),
    .X(_1911_));
 sg13g2_nand3_1 _2706_ (.B(\Pong.datapath.sw_ballMovement_reg[4] ),
    .C(net418),
    .A(net745),
    .Y(_1912_));
 sg13g2_a22oi_1 _2707_ (.Y(_1913_),
    .B1(_1911_),
    .B2(_1806_),
    .A2(_1908_),
    .A1(net439));
 sg13g2_nand2_1 _2708_ (.Y(_0040_),
    .A(_1912_),
    .B(net440));
 sg13g2_nor3_1 _2709_ (.A(\Pong.datapath.sw_ballMovement_reg[3] ),
    .B(\Pong.datapath.sw_ballMovement_reg[0] ),
    .C(_1907_),
    .Y(_1914_));
 sg13g2_nand2b_1 _2710_ (.Y(_1915_),
    .B(_1914_),
    .A_N(net257));
 sg13g2_a21oi_1 _2711_ (.A1(\Pong.datapath.sw_ballMovement_reg[2] ),
    .A2(_1909_),
    .Y(_1916_),
    .B1(net738));
 sg13g2_a21oi_1 _2712_ (.A1(\Pong.control_unit.state_ballMovement[3] ),
    .A2(\Pong.datapath.sw_ballMovement_reg[4] ),
    .Y(_1917_),
    .B1(net402));
 sg13g2_nand3_1 _2713_ (.B(_1916_),
    .C(net403),
    .A(_1915_),
    .Y(_0038_));
 sg13g2_nor3_1 _2714_ (.A(net738),
    .B(_1799_),
    .C(net439),
    .Y(_1918_));
 sg13g2_nor2_1 _2715_ (.A(net257),
    .B(\Pong.datapath.sw_ballMovement_reg[4] ),
    .Y(_1919_));
 sg13g2_nand2_1 _2716_ (.Y(_1920_),
    .A(_1918_),
    .B(_1919_));
 sg13g2_nor2_1 _2717_ (.A(net738),
    .B(\Pong.datapath.sw_ballMovement_reg[4] ),
    .Y(_1921_));
 sg13g2_nand3_1 _2718_ (.B(net418),
    .C(_1921_),
    .A(net447),
    .Y(_1922_));
 sg13g2_nand3_1 _2719_ (.B(\Pong.control_unit.state_ballMovement[0] ),
    .C(\Pong.datapath.sw_ballMovement_reg[3] ),
    .A(net745),
    .Y(_1923_));
 sg13g2_nand3_1 _2720_ (.B(_1922_),
    .C(_1923_),
    .A(_1920_),
    .Y(_0041_));
 sg13g2_a21oi_1 _2721_ (.A1(\Pong.control_unit.state_ballMovement[4] ),
    .A2(_1910_),
    .Y(_1924_),
    .B1(_1918_));
 sg13g2_nor2_1 _2722_ (.A(_1911_),
    .B(_1914_),
    .Y(_1925_));
 sg13g2_o21ai_1 _2723_ (.B1(_1925_),
    .Y(_1926_),
    .A1(\Pong.datapath.sw_ballMovement_reg[4] ),
    .A2(_1924_));
 sg13g2_and2_1 _2724_ (.A(net257),
    .B(_1926_),
    .X(_0039_));
 sg13g2_nand3_1 _2725_ (.B(_1910_),
    .C(_1919_),
    .A(net418),
    .Y(_1927_));
 sg13g2_nand3_1 _2726_ (.B(\Pong.datapath.sw_ballMovement_reg[0] ),
    .C(_1921_),
    .A(\Pong.control_unit.state_ballMovement[3] ),
    .Y(_1928_));
 sg13g2_nand3_1 _2727_ (.B(\Pong.control_unit.state_ballMovement[2] ),
    .C(\Pong.datapath.sw_ballMovement_reg[3] ),
    .A(net745),
    .Y(_1929_));
 sg13g2_nand3_1 _2728_ (.B(_1928_),
    .C(_1929_),
    .A(net419),
    .Y(_0042_));
 sg13g2_nand2_1 _2729_ (.Y(_1930_),
    .A(\Pong.datapath.Ball_Clock.Q[10] ),
    .B(\Pong.datapath.Ball_Clock.Q[9] ));
 sg13g2_nand3_1 _2730_ (.B(\Pong.datapath.Ball_Clock.Q[15] ),
    .C(\Pong.datapath.Ball_Clock.Q[7] ),
    .A(\Pong.datapath.Ball_Clock.Q[16] ),
    .Y(_1931_));
 sg13g2_nor3_1 _2731_ (.A(\Pong.datapath.Ball_Clock.Q[8] ),
    .B(_1930_),
    .C(_1931_),
    .Y(_1932_));
 sg13g2_nor4_2 _2732_ (.A(\Pong.datapath.Ball_Clock.Q[14] ),
    .B(\Pong.datapath.Ball_Clock.Q[13] ),
    .C(\Pong.datapath.Ball_Clock.Q[12] ),
    .Y(_1933_),
    .D(\Pong.datapath.Ball_Clock.Q[11] ));
 sg13g2_nor3_1 _2733_ (.A(\Pong.datapath.Ball_Clock.Q[2] ),
    .B(\Pong.datapath.Ball_Clock.Q[1] ),
    .C(\Pong.datapath.Ball_Clock.Q[0] ),
    .Y(_1934_));
 sg13g2_nor4_1 _2734_ (.A(\Pong.datapath.Ball_Clock.Q[6] ),
    .B(_1778_),
    .C(\Pong.datapath.Ball_Clock.Q[4] ),
    .D(\Pong.datapath.Ball_Clock.Q[3] ),
    .Y(_1935_));
 sg13g2_and4_1 _2735_ (.A(_1932_),
    .B(_1933_),
    .C(_1934_),
    .D(_1935_),
    .X(\Pong.datapath.Ball_Clock.roll ));
 sg13g2_a22oi_1 _2736_ (.Y(_1936_),
    .B1(_1872_),
    .B2(net303),
    .A2(net643),
    .A1(net278));
 sg13g2_inv_1 _2737_ (.Y(_0028_),
    .A(_1936_));
 sg13g2_a22oi_1 _2738_ (.Y(_1937_),
    .B1(net641),
    .B2(net320),
    .A2(net643),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[8] ));
 sg13g2_inv_1 _2739_ (.Y(_0027_),
    .A(net321));
 sg13g2_a22oi_1 _2740_ (.Y(_1938_),
    .B1(net642),
    .B2(net312),
    .A2(net644),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[16] ));
 sg13g2_inv_1 _2741_ (.Y(_0032_),
    .A(net313));
 sg13g2_a22oi_1 _2742_ (.Y(_1939_),
    .B1(net641),
    .B2(net395),
    .A2(net643),
    .A1(net333));
 sg13g2_inv_1 _2743_ (.Y(_0031_),
    .A(_1939_));
 sg13g2_a22oi_1 _2744_ (.Y(_1940_),
    .B1(net641),
    .B2(net304),
    .A2(net644),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ));
 sg13g2_inv_1 _2745_ (.Y(_0030_),
    .A(net305));
 sg13g2_a22oi_1 _2746_ (.Y(_1941_),
    .B1(net641),
    .B2(net291),
    .A2(net643),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ));
 sg13g2_inv_1 _2747_ (.Y(_0029_),
    .A(net292));
 sg13g2_a21oi_1 _2748_ (.A1(net341),
    .A2(_1870_),
    .Y(_1942_),
    .B1(net741));
 sg13g2_o21ai_1 _2749_ (.B1(_1942_),
    .Y(_0019_),
    .A1(_1801_),
    .A2(_1889_));
 sg13g2_a22oi_1 _2750_ (.Y(_1943_),
    .B1(net645),
    .B2(net301),
    .A2(net648),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[18] ));
 sg13g2_inv_1 _2751_ (.Y(_0009_),
    .A(net302));
 sg13g2_a22oi_1 _2752_ (.Y(_1944_),
    .B1(net646),
    .B2(net381),
    .A2(net649),
    .A1(net339));
 sg13g2_inv_1 _2753_ (.Y(_0008_),
    .A(_1944_));
 sg13g2_a22oi_1 _2754_ (.Y(_1945_),
    .B1(net646),
    .B2(net309),
    .A2(net649),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ));
 sg13g2_inv_1 _2755_ (.Y(_0007_),
    .A(net310));
 sg13g2_a22oi_1 _2756_ (.Y(_1946_),
    .B1(net647),
    .B2(net281),
    .A2(net650),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ));
 sg13g2_inv_1 _2757_ (.Y(_0006_),
    .A(net282));
 sg13g2_a22oi_1 _2758_ (.Y(_1947_),
    .B1(net645),
    .B2(net311),
    .A2(net648),
    .A1(net295));
 sg13g2_inv_1 _2759_ (.Y(_0005_),
    .A(_1947_));
 sg13g2_a22oi_1 _2760_ (.Y(_1948_),
    .B1(net645),
    .B2(net399),
    .A2(net648),
    .A1(net384));
 sg13g2_inv_1 _2761_ (.Y(_0004_),
    .A(_1948_));
 sg13g2_a22oi_1 _2762_ (.Y(_1949_),
    .B1(net647),
    .B2(net322),
    .A2(net650),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ));
 sg13g2_inv_1 _2763_ (.Y(_0003_),
    .A(net323));
 sg13g2_nor2_2 _2764_ (.A(net628),
    .B(net631),
    .Y(_1950_));
 sg13g2_or2_1 _2765_ (.X(_1951_),
    .B(net631),
    .A(net628));
 sg13g2_nor2_1 _2766_ (.A(net624),
    .B(net626),
    .Y(_1952_));
 sg13g2_or2_2 _2767_ (.X(_1953_),
    .B(net626),
    .A(net624));
 sg13g2_nor2_1 _2768_ (.A(net629),
    .B(_1953_),
    .Y(_1954_));
 sg13g2_nor2_1 _2769_ (.A(net625),
    .B(net593),
    .Y(_1955_));
 sg13g2_nor2_2 _2770_ (.A(_1951_),
    .B(_1953_),
    .Y(_1956_));
 sg13g2_nor3_1 _2771_ (.A(\Pong.datapath.ballFunction.ball_center_y[4] ),
    .B(net629),
    .C(_1953_),
    .Y(_1957_));
 sg13g2_nand2b_2 _2772_ (.Y(_1958_),
    .B(_1956_),
    .A_N(net623));
 sg13g2_nand2_1 _2773_ (.Y(_1959_),
    .A(net613),
    .B(net615));
 sg13g2_nand3_1 _2774_ (.B(_1775_),
    .C(net620),
    .A(_1774_),
    .Y(_1960_));
 sg13g2_nor3_2 _2775_ (.A(_1958_),
    .B(_1959_),
    .C(_1960_),
    .Y(_0044_));
 sg13g2_or2_1 _2776_ (.X(_1961_),
    .B(_0044_),
    .A(_0043_));
 sg13g2_nand2_1 _2777_ (.Y(_1962_),
    .A(net728),
    .B(net727));
 sg13g2_nand4_1 _2778_ (.B(\Pong.datapath.rightPaddle[4] ),
    .C(net728),
    .A(\Pong.datapath.rightPaddle[3] ),
    .Y(_1963_),
    .D(net727));
 sg13g2_nand3_1 _2779_ (.B(_1811_),
    .C(_1963_),
    .A(_1810_),
    .Y(_1964_));
 sg13g2_nor2_1 _2780_ (.A(net724),
    .B(_1964_),
    .Y(_1965_));
 sg13g2_nor3_2 _2781_ (.A(\Pong.datapath.rightPaddle[8] ),
    .B(net724),
    .C(_1964_),
    .Y(_1966_));
 sg13g2_xnor2_1 _2782_ (.Y(_1967_),
    .A(_0056_),
    .B(_1966_));
 sg13g2_inv_1 _2783_ (.Y(_1968_),
    .A(_1967_));
 sg13g2_xnor2_1 _2784_ (.Y(_1969_),
    .A(_0058_),
    .B(_1965_));
 sg13g2_xnor2_1 _2785_ (.Y(_1970_),
    .A(_0113_),
    .B(_1967_));
 sg13g2_a21oi_1 _2786_ (.A1(net611),
    .A2(_1969_),
    .Y(_1971_),
    .B1(_1970_));
 sg13g2_xnor2_1 _2787_ (.Y(_1972_),
    .A(_0059_),
    .B(_1964_));
 sg13g2_nand2_1 _2788_ (.Y(_1973_),
    .A(net615),
    .B(_1972_));
 sg13g2_o21ai_1 _2789_ (.B1(_1973_),
    .Y(_1974_),
    .A1(net611),
    .A2(_1969_));
 sg13g2_inv_1 _2790_ (.Y(_1975_),
    .A(_1974_));
 sg13g2_nor2_1 _2791_ (.A(net614),
    .B(_1972_),
    .Y(_1976_));
 sg13g2_nand2_1 _2792_ (.Y(_1977_),
    .A(_0061_),
    .B(_1963_));
 sg13g2_xor2_1 _2793_ (.B(_1977_),
    .A(_0060_),
    .X(_1978_));
 sg13g2_inv_1 _2794_ (.Y(_1979_),
    .A(_1978_));
 sg13g2_xnor2_1 _2795_ (.Y(_1980_),
    .A(_1811_),
    .B(_1963_));
 sg13g2_nor2_1 _2796_ (.A(_0066_),
    .B(_1962_),
    .Y(_1981_));
 sg13g2_xor2_1 _2797_ (.B(_1981_),
    .A(_0065_),
    .X(_1982_));
 sg13g2_nor2_1 _2798_ (.A(_1816_),
    .B(_1982_),
    .Y(_1983_));
 sg13g2_xnor2_1 _2799_ (.Y(_1984_),
    .A(_0063_),
    .B(_1980_));
 sg13g2_nor2_1 _2800_ (.A(_1983_),
    .B(_1984_),
    .Y(_1985_));
 sg13g2_and2_1 _2801_ (.A(net630),
    .B(net728),
    .X(_1986_));
 sg13g2_nand2b_1 _2802_ (.Y(_1987_),
    .B(net730),
    .A_N(net632));
 sg13g2_xor2_1 _2803_ (.B(net728),
    .A(net630),
    .X(_1988_));
 sg13g2_a21oi_1 _2804_ (.A1(_1987_),
    .A2(_1988_),
    .Y(_1989_),
    .B1(_1986_));
 sg13g2_xnor2_1 _2805_ (.Y(_1990_),
    .A(_1815_),
    .B(_1962_));
 sg13g2_nand2_1 _2806_ (.Y(_1991_),
    .A(_1777_),
    .B(_1990_));
 sg13g2_nor2_1 _2807_ (.A(net728),
    .B(net727),
    .Y(_1992_));
 sg13g2_xnor2_1 _2808_ (.Y(_1993_),
    .A(net728),
    .B(net727));
 sg13g2_or2_1 _2809_ (.X(_1994_),
    .B(_1993_),
    .A(_0067_));
 sg13g2_and2_1 _2810_ (.A(_0067_),
    .B(_1993_),
    .X(_1995_));
 sg13g2_nand2_1 _2811_ (.Y(_1996_),
    .A(_0067_),
    .B(_1993_));
 sg13g2_nand2b_1 _2812_ (.Y(_1997_),
    .B(\Pong.datapath.ballFunction.ball_center_y[3] ),
    .A_N(_1990_));
 sg13g2_a22oi_1 _2813_ (.Y(_1998_),
    .B1(_1994_),
    .B2(_1996_),
    .A2(_1990_),
    .A1(_1777_));
 sg13g2_nand2_1 _2814_ (.Y(_1999_),
    .A(_1997_),
    .B(_1998_));
 sg13g2_nor2_1 _2815_ (.A(_1989_),
    .B(_1999_),
    .Y(_2000_));
 sg13g2_nand3_1 _2816_ (.B(_1991_),
    .C(_1993_),
    .A(net627),
    .Y(_2001_));
 sg13g2_nand2_1 _2817_ (.Y(_2002_),
    .A(_1816_),
    .B(_1982_));
 sg13g2_nand3_1 _2818_ (.B(_2001_),
    .C(_2002_),
    .A(_1997_),
    .Y(_2003_));
 sg13g2_o21ai_1 _2819_ (.B1(_1985_),
    .Y(_2004_),
    .A1(_2000_),
    .A2(_2003_));
 sg13g2_o21ai_1 _2820_ (.B1(_2004_),
    .Y(_2005_),
    .A1(_1776_),
    .A2(_1980_));
 sg13g2_xor2_1 _2821_ (.B(_1978_),
    .A(net617),
    .X(_2006_));
 sg13g2_a22oi_1 _2822_ (.Y(_2007_),
    .B1(_2005_),
    .B2(_2006_),
    .A2(_1979_),
    .A1(\Pong.datapath.ballFunction.ball_center_y[6] ));
 sg13g2_o21ai_1 _2823_ (.B1(_1975_),
    .Y(_2008_),
    .A1(_1976_),
    .A2(_2007_));
 sg13g2_a22oi_1 _2824_ (.Y(_2009_),
    .B1(_1971_),
    .B2(_2008_),
    .A2(_1968_),
    .A1(net609));
 sg13g2_nand2_1 _2825_ (.Y(_2010_),
    .A(_1812_),
    .B(_1992_));
 sg13g2_nor4_2 _2826_ (.A(\Pong.datapath.rightPaddle[3] ),
    .B(\Pong.datapath.rightPaddle[4] ),
    .C(net729),
    .Y(_2011_),
    .D(net727));
 sg13g2_nor2_2 _2827_ (.A(_1811_),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_xnor2_1 _2828_ (.Y(_2013_),
    .A(\Pong.datapath.rightPaddle[5] ),
    .B(_2011_));
 sg13g2_nor2_1 _2829_ (.A(_1776_),
    .B(_2013_),
    .Y(_2014_));
 sg13g2_xnor2_1 _2830_ (.Y(_2015_),
    .A(_1815_),
    .B(_1992_));
 sg13g2_xnor2_1 _2831_ (.Y(_2016_),
    .A(_0068_),
    .B(_2015_));
 sg13g2_a21oi_1 _2832_ (.A1(_1989_),
    .A2(_1994_),
    .Y(_2017_),
    .B1(_1995_));
 sg13g2_xor2_1 _2833_ (.B(_2010_),
    .A(_0065_),
    .X(_2018_));
 sg13g2_nor2_1 _2834_ (.A(net622),
    .B(_2018_),
    .Y(_2019_));
 sg13g2_xor2_1 _2835_ (.B(_2013_),
    .A(net619),
    .X(_2020_));
 sg13g2_a22oi_1 _2836_ (.Y(_2021_),
    .B1(_2016_),
    .B2(_2017_),
    .A2(_2015_),
    .A1(\Pong.datapath.ballFunction.ball_center_y[3] ));
 sg13g2_a21oi_1 _2837_ (.A1(net622),
    .A2(_2018_),
    .Y(_2022_),
    .B1(_2021_));
 sg13g2_o21ai_1 _2838_ (.B1(_2020_),
    .Y(_2023_),
    .A1(_2019_),
    .A2(_2022_));
 sg13g2_nor2b_1 _2839_ (.A(_2014_),
    .B_N(_2023_),
    .Y(_2024_));
 sg13g2_xnor2_1 _2840_ (.Y(_2025_),
    .A(_0060_),
    .B(_2012_));
 sg13g2_xnor2_1 _2841_ (.Y(_2026_),
    .A(net617),
    .B(_2025_));
 sg13g2_nor2_1 _2842_ (.A(_1775_),
    .B(_2025_),
    .Y(_2027_));
 sg13g2_nand2_1 _2843_ (.Y(_2028_),
    .A(net726),
    .B(_2012_));
 sg13g2_nor2_1 _2844_ (.A(_0059_),
    .B(_2028_),
    .Y(_2029_));
 sg13g2_xnor2_1 _2845_ (.Y(_2030_),
    .A(_0059_),
    .B(_2028_));
 sg13g2_a21oi_1 _2846_ (.A1(net614),
    .A2(_2030_),
    .Y(_2031_),
    .B1(_2027_));
 sg13g2_o21ai_1 _2847_ (.B1(_2031_),
    .Y(_2032_),
    .A1(_2024_),
    .A2(_2026_));
 sg13g2_xor2_1 _2848_ (.B(_2029_),
    .A(_0058_),
    .X(_2033_));
 sg13g2_xnor2_1 _2849_ (.Y(_2034_),
    .A(net611),
    .B(_2033_));
 sg13g2_o21ai_1 _2850_ (.B1(_2034_),
    .Y(_2035_),
    .A1(net614),
    .A2(_2030_));
 sg13g2_nand2b_1 _2851_ (.Y(_2036_),
    .B(_2032_),
    .A_N(_2035_));
 sg13g2_nand4_1 _2852_ (.B(net724),
    .C(net726),
    .A(\Pong.datapath.rightPaddle[8] ),
    .Y(_2037_),
    .D(_2012_));
 sg13g2_xnor2_1 _2853_ (.Y(_2038_),
    .A(_0056_),
    .B(_2037_));
 sg13g2_a22oi_1 _2854_ (.Y(_2039_),
    .B1(_2038_),
    .B2(net609),
    .A2(_2033_),
    .A1(net613));
 sg13g2_nor2_1 _2855_ (.A(net609),
    .B(_2038_),
    .Y(_2040_));
 sg13g2_nand4_1 _2856_ (.B(net724),
    .C(net726),
    .A(\Pong.datapath.rightPaddle[8] ),
    .Y(_2041_),
    .D(\Pong.datapath.rightPaddle[9] ));
 sg13g2_inv_1 _2857_ (.Y(_2042_),
    .A(_2041_));
 sg13g2_a221oi_1 _2858_ (.B2(_2012_),
    .C1(_2040_),
    .B1(_2042_),
    .A1(_2036_),
    .Y(_2043_),
    .A2(_2039_));
 sg13g2_nand2b_1 _2859_ (.Y(_2044_),
    .B(net632),
    .A_N(net730));
 sg13g2_and4_1 _2860_ (.A(_1987_),
    .B(_1988_),
    .C(_2002_),
    .D(_2044_),
    .X(_2045_));
 sg13g2_nand2b_1 _2861_ (.Y(_2046_),
    .B(_2045_),
    .A_N(_1976_));
 sg13g2_nand2_1 _2862_ (.Y(_2047_),
    .A(_1985_),
    .B(_2006_));
 sg13g2_nor4_1 _2863_ (.A(_1974_),
    .B(_1999_),
    .C(_2046_),
    .D(_2047_),
    .Y(_2048_));
 sg13g2_nor2_1 _2864_ (.A(net604),
    .B(net605),
    .Y(_2049_));
 sg13g2_nor2_2 _2865_ (.A(net601),
    .B(net603),
    .Y(_2050_));
 sg13g2_nor2_1 _2866_ (.A(\Pong.datapath.ballFunction.ball_center_x[8] ),
    .B(net595),
    .Y(_2051_));
 sg13g2_nand3_1 _2867_ (.B(net597),
    .C(_2051_),
    .A(\Pong.datapath.ballFunction.ball_center_x[9] ),
    .Y(_2052_));
 sg13g2_nor2b_1 _2868_ (.A(net598),
    .B_N(net600),
    .Y(_2053_));
 sg13g2_nor4_1 _2869_ (.A(net601),
    .B(net603),
    .C(net607),
    .D(_2052_),
    .Y(_2054_));
 sg13g2_nor2b_1 _2870_ (.A(\Pong.datapath.rightPaddle[9] ),
    .B_N(_1966_),
    .Y(_2055_));
 sg13g2_a21oi_2 _2871_ (.B1(_2055_),
    .Y(_2056_),
    .A2(_2048_),
    .A1(_1971_));
 sg13g2_nand4_1 _2872_ (.B(_2053_),
    .C(_2054_),
    .A(\Pong.datapath.ballFunction.ball_center_x[0] ),
    .Y(_2057_),
    .D(_2056_));
 sg13g2_nor3_2 _2873_ (.A(_2009_),
    .B(_2043_),
    .C(_2057_),
    .Y(_2058_));
 sg13g2_nor2_2 _2874_ (.A(net716),
    .B(net713),
    .Y(_2059_));
 sg13g2_nor3_2 _2875_ (.A(net711),
    .B(net715),
    .C(net713),
    .Y(_2060_));
 sg13g2_and2_1 _2876_ (.A(_1819_),
    .B(_2060_),
    .X(_2061_));
 sg13g2_nand2b_1 _2877_ (.Y(_2062_),
    .B(net708),
    .A_N(_2061_));
 sg13g2_xor2_1 _2878_ (.B(_2061_),
    .A(net708),
    .X(_2063_));
 sg13g2_xor2_1 _2879_ (.B(_2063_),
    .A(net619),
    .X(_2064_));
 sg13g2_xnor2_1 _2880_ (.Y(_2065_),
    .A(_0074_),
    .B(_2060_));
 sg13g2_or2_1 _2881_ (.X(_2066_),
    .B(_2065_),
    .A(net622));
 sg13g2_xnor2_1 _2882_ (.Y(_2067_),
    .A(_0075_),
    .B(_2059_));
 sg13g2_xor2_1 _2883_ (.B(_2067_),
    .A(_0068_),
    .X(_2068_));
 sg13g2_nand2_1 _2884_ (.Y(_2069_),
    .A(net630),
    .B(net715));
 sg13g2_nor2b_1 _2885_ (.A(net632),
    .B_N(net717),
    .Y(_2070_));
 sg13g2_nor2_1 _2886_ (.A(net630),
    .B(net715),
    .Y(_2071_));
 sg13g2_a21oi_1 _2887_ (.A1(net630),
    .A2(net715),
    .Y(_2072_),
    .B1(_2070_));
 sg13g2_nand2b_1 _2888_ (.Y(_2073_),
    .B(_2072_),
    .A_N(_2071_));
 sg13g2_o21ai_1 _2889_ (.B1(_2069_),
    .Y(_2074_),
    .A1(_2070_),
    .A2(_2071_));
 sg13g2_nand2_1 _2890_ (.Y(_2075_),
    .A(net715),
    .B(net713));
 sg13g2_xnor2_1 _2891_ (.Y(_2076_),
    .A(net715),
    .B(net713));
 sg13g2_nor2_1 _2892_ (.A(_0067_),
    .B(_2076_),
    .Y(_2077_));
 sg13g2_nor2_1 _2893_ (.A(_2074_),
    .B(_2077_),
    .Y(_2078_));
 sg13g2_a21oi_1 _2894_ (.A1(_0067_),
    .A2(_2076_),
    .Y(_2079_),
    .B1(_2078_));
 sg13g2_o21ai_1 _2895_ (.B1(_2066_),
    .Y(_2080_),
    .A1(_1777_),
    .A2(_2067_));
 sg13g2_a21o_1 _2896_ (.A2(_2079_),
    .A1(_2068_),
    .B1(_2080_),
    .X(_2081_));
 sg13g2_a21oi_1 _2897_ (.A1(net622),
    .A2(_2065_),
    .Y(_2082_),
    .B1(_2064_));
 sg13g2_a22oi_1 _2898_ (.Y(_2083_),
    .B1(_2081_),
    .B2(_2082_),
    .A2(_2063_),
    .A1(net620));
 sg13g2_xor2_1 _2899_ (.B(_2062_),
    .A(_0072_),
    .X(_2084_));
 sg13g2_xnor2_1 _2900_ (.Y(_2085_),
    .A(net617),
    .B(_2084_));
 sg13g2_nor2_1 _2901_ (.A(_1775_),
    .B(_2084_),
    .Y(_2086_));
 sg13g2_or2_1 _2902_ (.X(_2087_),
    .B(_2062_),
    .A(_1818_));
 sg13g2_nor2_1 _2903_ (.A(_0071_),
    .B(_2087_),
    .Y(_2088_));
 sg13g2_xnor2_1 _2904_ (.Y(_2089_),
    .A(_0071_),
    .B(_2087_));
 sg13g2_a21oi_1 _2905_ (.A1(net614),
    .A2(_2089_),
    .Y(_2090_),
    .B1(_2086_));
 sg13g2_o21ai_1 _2906_ (.B1(_2090_),
    .Y(_2091_),
    .A1(_2083_),
    .A2(_2085_));
 sg13g2_xor2_1 _2907_ (.B(_2088_),
    .A(_0070_),
    .X(_2092_));
 sg13g2_xor2_1 _2908_ (.B(_2092_),
    .A(net611),
    .X(_2093_));
 sg13g2_o21ai_1 _2909_ (.B1(_2091_),
    .Y(_2094_),
    .A1(net614),
    .A2(_2089_));
 sg13g2_nand3_1 _2910_ (.B(\Pong.datapath.leftPaddle[7] ),
    .C(\Pong.datapath.leftPaddle[6] ),
    .A(\Pong.datapath.leftPaddle[8] ),
    .Y(_2095_));
 sg13g2_or2_1 _2911_ (.X(_2096_),
    .B(_2095_),
    .A(_2062_));
 sg13g2_inv_1 _2912_ (.Y(_2097_),
    .A(_2096_));
 sg13g2_xnor2_1 _2913_ (.Y(_2098_),
    .A(net706),
    .B(_2096_));
 sg13g2_a22oi_1 _2914_ (.Y(_2099_),
    .B1(_2098_),
    .B2(net609),
    .A2(_2092_),
    .A1(net613));
 sg13g2_o21ai_1 _2915_ (.B1(_2099_),
    .Y(_2100_),
    .A1(_2093_),
    .A2(_2094_));
 sg13g2_o21ai_1 _2916_ (.B1(_2100_),
    .Y(_2101_),
    .A1(net608),
    .A2(_2098_));
 sg13g2_a21oi_2 _2917_ (.B1(_2101_),
    .Y(_2102_),
    .A2(_2097_),
    .A1(net529));
 sg13g2_and2_2 _2918_ (.A(net711),
    .B(net710),
    .X(_2103_));
 sg13g2_nand2b_2 _2919_ (.Y(_2104_),
    .B(_2103_),
    .A_N(_2075_));
 sg13g2_nor2_1 _2920_ (.A(net707),
    .B(net708),
    .Y(_2105_));
 sg13g2_nand2_1 _2921_ (.Y(_2106_),
    .A(_2104_),
    .B(_2105_));
 sg13g2_nand3_1 _2922_ (.B(_2104_),
    .C(_2105_),
    .A(_1817_),
    .Y(_2107_));
 sg13g2_nor2_1 _2923_ (.A(\Pong.datapath.leftPaddle[8] ),
    .B(_2107_),
    .Y(_2108_));
 sg13g2_xnor2_1 _2924_ (.Y(_2109_),
    .A(net706),
    .B(_2108_));
 sg13g2_nand2b_1 _2925_ (.Y(_2110_),
    .B(net608),
    .A_N(_2109_));
 sg13g2_xor2_1 _2926_ (.B(_2106_),
    .A(_0071_),
    .X(_2111_));
 sg13g2_nand2b_1 _2927_ (.Y(_2112_),
    .B(_2111_),
    .A_N(net614));
 sg13g2_nand2_1 _2928_ (.Y(_2113_),
    .A(_0073_),
    .B(_2104_));
 sg13g2_xnor2_1 _2929_ (.Y(_2114_),
    .A(_0072_),
    .B(_2113_));
 sg13g2_nand2_1 _2930_ (.Y(_2115_),
    .A(net618),
    .B(_2114_));
 sg13g2_xnor2_1 _2931_ (.Y(_2116_),
    .A(net617),
    .B(_2114_));
 sg13g2_xor2_1 _2932_ (.B(_2104_),
    .A(net708),
    .X(_2117_));
 sg13g2_nor2_1 _2933_ (.A(_1776_),
    .B(_2117_),
    .Y(_2118_));
 sg13g2_nor2_1 _2934_ (.A(_0075_),
    .B(_2075_),
    .Y(_2119_));
 sg13g2_xor2_1 _2935_ (.B(_2119_),
    .A(_0074_),
    .X(_2120_));
 sg13g2_nand2b_1 _2936_ (.Y(_2121_),
    .B(net622),
    .A_N(_2120_));
 sg13g2_xor2_1 _2937_ (.B(_2117_),
    .A(net619),
    .X(_2122_));
 sg13g2_nand2_1 _2938_ (.Y(_2123_),
    .A(_2121_),
    .B(_2122_));
 sg13g2_xor2_1 _2939_ (.B(_2075_),
    .A(_0075_),
    .X(_2124_));
 sg13g2_nand2_1 _2940_ (.Y(_2125_),
    .A(_1777_),
    .B(_2124_));
 sg13g2_nor2_1 _2941_ (.A(_1777_),
    .B(_2124_),
    .Y(_2126_));
 sg13g2_xor2_1 _2942_ (.B(_2076_),
    .A(_0067_),
    .X(_2127_));
 sg13g2_a21oi_1 _2943_ (.A1(_1777_),
    .A2(_2124_),
    .Y(_2128_),
    .B1(_2127_));
 sg13g2_nor2b_1 _2944_ (.A(_2126_),
    .B_N(_2128_),
    .Y(_2129_));
 sg13g2_nand2_1 _2945_ (.Y(_2130_),
    .A(_2074_),
    .B(_2129_));
 sg13g2_and2_1 _2946_ (.A(net627),
    .B(_2076_),
    .X(_2131_));
 sg13g2_a221oi_1 _2947_ (.B2(_2131_),
    .C1(_2126_),
    .B1(_2125_),
    .A1(_1816_),
    .Y(_2132_),
    .A2(_2120_));
 sg13g2_a21oi_1 _2948_ (.A1(_2130_),
    .A2(_2132_),
    .Y(_2133_),
    .B1(_2123_));
 sg13g2_o21ai_1 _2949_ (.B1(_2116_),
    .Y(_2134_),
    .A1(_2118_),
    .A2(_2133_));
 sg13g2_nand2_1 _2950_ (.Y(_2135_),
    .A(_2115_),
    .B(_2134_));
 sg13g2_nand2b_1 _2951_ (.Y(_2136_),
    .B(net614),
    .A_N(_2111_));
 sg13g2_xor2_1 _2952_ (.B(_2107_),
    .A(_0070_),
    .X(_2137_));
 sg13g2_o21ai_1 _2953_ (.B1(_2136_),
    .Y(_2138_),
    .A1(net611),
    .A2(_2137_));
 sg13g2_a21oi_1 _2954_ (.A1(_2112_),
    .A2(_2135_),
    .Y(_2139_),
    .B1(_2138_));
 sg13g2_xnor2_1 _2955_ (.Y(_2140_),
    .A(_0113_),
    .B(_2109_));
 sg13g2_a21o_1 _2956_ (.A2(_2137_),
    .A1(net611),
    .B1(_2140_),
    .X(_2141_));
 sg13g2_o21ai_1 _2957_ (.B1(_2110_),
    .Y(_2142_),
    .A1(_2139_),
    .A2(_2141_));
 sg13g2_a221oi_1 _2958_ (.B2(_1816_),
    .C1(_2073_),
    .B1(_2120_),
    .A1(net632),
    .Y(_2143_),
    .A2(_1821_));
 sg13g2_nand3_1 _2959_ (.B(_2129_),
    .C(_2143_),
    .A(_2112_),
    .Y(_2144_));
 sg13g2_nand3_1 _2960_ (.B(_2121_),
    .C(_2122_),
    .A(_2116_),
    .Y(_2145_));
 sg13g2_nor4_1 _2961_ (.A(_2138_),
    .B(_2141_),
    .C(_2144_),
    .D(_2145_),
    .Y(_2146_));
 sg13g2_nor3_1 _2962_ (.A(\Pong.datapath.leftPaddle[8] ),
    .B(\Pong.datapath.leftPaddle[9] ),
    .C(_2107_),
    .Y(_2147_));
 sg13g2_or2_1 _2963_ (.X(_2148_),
    .B(net594),
    .A(\Pong.datapath.ballFunction.ball_center_x[9] ));
 sg13g2_nor3_2 _2964_ (.A(\Pong.datapath.ballFunction.ball_center_x[7] ),
    .B(net597),
    .C(_2148_),
    .Y(_2149_));
 sg13g2_nand2_1 _2965_ (.Y(_2150_),
    .A(net606),
    .B(\Pong.datapath.ballFunction.ball_center_x[0] ));
 sg13g2_and2_2 _2966_ (.A(net601),
    .B(net603),
    .X(_2151_));
 sg13g2_nand2b_2 _2967_ (.Y(_2152_),
    .B(_2151_),
    .A_N(net592));
 sg13g2_nand2b_2 _2968_ (.Y(_2153_),
    .B(net598),
    .A_N(net600));
 sg13g2_nor2_1 _2969_ (.A(_2152_),
    .B(_2153_),
    .Y(_2154_));
 sg13g2_nand2_2 _2970_ (.Y(_2155_),
    .A(_2149_),
    .B(_2154_));
 sg13g2_nor3_1 _2971_ (.A(_2146_),
    .B(_2147_),
    .C(_2155_),
    .Y(_2156_));
 sg13g2_nand2_2 _2972_ (.Y(_2157_),
    .A(_2142_),
    .B(_2156_));
 sg13g2_nor4_2 _2973_ (.A(_1961_),
    .B(_2058_),
    .C(_2102_),
    .Y(_0045_),
    .D(_2157_));
 sg13g2_nor2b_1 _2974_ (.A(_1961_),
    .B_N(_2058_),
    .Y(_0046_));
 sg13g2_nor2_1 _2975_ (.A(\Pong.datapath.ballFunction.ball_center_x[4] ),
    .B(net602),
    .Y(_2158_));
 sg13g2_nand2_1 _2976_ (.Y(_2159_),
    .A(net597),
    .B(\Pong.datapath.ballFunction.ball_center_x[5] ));
 sg13g2_o21ai_1 _2977_ (.B1(_2051_),
    .Y(_2160_),
    .A1(_2158_),
    .A2(_2159_));
 sg13g2_nor2_2 _2978_ (.A(net606),
    .B(\Pong.datapath.ballFunction.ball_center_x[0] ),
    .Y(_2161_));
 sg13g2_or2_1 _2979_ (.X(_2162_),
    .B(\Pong.datapath.ballFunction.ball_center_x[0] ),
    .A(net606));
 sg13g2_nor2_2 _2980_ (.A(net604),
    .B(net590),
    .Y(_2163_));
 sg13g2_nand3b_1 _2981_ (.B(net602),
    .C(\Pong.datapath.ballFunction.ball_center_x[4] ),
    .Y(_2164_),
    .A_N(_2163_));
 sg13g2_nor2b_1 _2982_ (.A(net598),
    .B_N(_2149_),
    .Y(_2165_));
 sg13g2_a22oi_1 _2983_ (.Y(_2166_),
    .B1(_2164_),
    .B2(_2165_),
    .A2(_2160_),
    .A1(\Pong.datapath.ballFunction.ball_center_x[9] ));
 sg13g2_nor3_1 _2984_ (.A(_1961_),
    .B(_2058_),
    .C(_2166_),
    .Y(_0047_));
 sg13g2_nor2_1 _2985_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[5] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[10] ),
    .Y(_2167_));
 sg13g2_nand2_1 _2986_ (.Y(_2168_),
    .A(_0115_),
    .B(_2167_));
 sg13g2_or2_1 _2987_ (.X(_2169_),
    .B(_2168_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ));
 sg13g2_nand2b_1 _2988_ (.Y(_2170_),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[18] ),
    .A_N(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ));
 sg13g2_nand2_1 _2989_ (.Y(_2171_),
    .A(_0121_),
    .B(_2170_));
 sg13g2_or2_1 _2990_ (.X(_2172_),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[1] ));
 sg13g2_a21oi_1 _2991_ (.A1(_1797_),
    .A2(\Pong.control_unit.NES_Controller_Left.state_NESController[6] ),
    .Y(_2173_),
    .B1(_2172_));
 sg13g2_o21ai_1 _2992_ (.B1(_0120_),
    .Y(_2174_),
    .A1(_2171_),
    .A2(_2173_));
 sg13g2_nand2_1 _2993_ (.Y(_2175_),
    .A(_0119_),
    .B(_2174_));
 sg13g2_nand2_1 _2994_ (.Y(_2176_),
    .A(_0123_),
    .B(_2175_));
 sg13g2_nand2_1 _2995_ (.Y(_2177_),
    .A(_0122_),
    .B(_2176_));
 sg13g2_a21oi_1 _2996_ (.A1(_0118_),
    .A2(_2177_),
    .Y(_2178_),
    .B1(\Pong.control_unit.NES_Controller_Left.state_NESController[17] ));
 sg13g2_o21ai_1 _2997_ (.B1(_1798_),
    .Y(_2179_),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[8] ),
    .A2(_2178_));
 sg13g2_a21oi_2 _2998_ (.B1(_2169_),
    .Y(uio_out[1]),
    .A2(_2179_),
    .A1(_1802_));
 sg13g2_nor2b_2 _2999_ (.A(_2167_),
    .B_N(_0115_),
    .Y(uio_out[2]));
 sg13g2_nor2_1 _3000_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[5] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[10] ),
    .Y(_2180_));
 sg13g2_nand2_1 _3001_ (.Y(_2181_),
    .A(_0116_),
    .B(_2180_));
 sg13g2_or2_1 _3002_ (.X(_2182_),
    .B(_2181_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ));
 sg13g2_nand2b_1 _3003_ (.Y(_2183_),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ),
    .A_N(\Pong.control_unit.NES_Controller_Right.state_NESController[9] ));
 sg13g2_nand2_1 _3004_ (.Y(_2184_),
    .A(_0128_),
    .B(_2183_));
 sg13g2_or2_1 _3005_ (.X(_2185_),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[9] ));
 sg13g2_a21oi_1 _3006_ (.A1(\Pong.control_unit.NES_Controller_Right.state_NESController[6] ),
    .A2(_1804_),
    .Y(_2186_),
    .B1(_2185_));
 sg13g2_o21ai_1 _3007_ (.B1(_0127_),
    .Y(_2187_),
    .A1(_2184_),
    .A2(_2186_));
 sg13g2_nand2_1 _3008_ (.Y(_2188_),
    .A(_0126_),
    .B(_2187_));
 sg13g2_nand2_1 _3009_ (.Y(_2189_),
    .A(_0130_),
    .B(_2188_));
 sg13g2_nand2_1 _3010_ (.Y(_2190_),
    .A(_0129_),
    .B(_2189_));
 sg13g2_a21oi_1 _3011_ (.A1(_0125_),
    .A2(_2190_),
    .Y(_2191_),
    .B1(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ));
 sg13g2_nor2b_1 _3012_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ),
    .B_N(\Pong.control_unit.NES_Controller_Right.state_NESController[13] ),
    .Y(_2192_));
 sg13g2_nor3_1 _3013_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[8] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ),
    .C(_2191_),
    .Y(_2193_));
 sg13g2_nor3_2 _3014_ (.A(_2182_),
    .B(_2192_),
    .C(_2193_),
    .Y(uio_out[4]));
 sg13g2_nor2b_2 _3015_ (.A(_2180_),
    .B_N(_0116_),
    .Y(uio_out[5]));
 sg13g2_nand2_1 _3016_ (.Y(_2194_),
    .A(net716),
    .B(net717));
 sg13g2_nand3_1 _3017_ (.B(net713),
    .C(net717),
    .A(net716),
    .Y(_2195_));
 sg13g2_o21ai_1 _3018_ (.B1(_0075_),
    .Y(_2196_),
    .A1(net711),
    .A2(_2195_));
 sg13g2_o21ai_1 _3019_ (.B1(net708),
    .Y(_2197_),
    .A1(net710),
    .A2(_2196_));
 sg13g2_nor2_1 _3020_ (.A(_1818_),
    .B(_2197_),
    .Y(_2198_));
 sg13g2_nor3_1 _3021_ (.A(_1817_),
    .B(_1818_),
    .C(_2197_),
    .Y(_2199_));
 sg13g2_nor2_1 _3022_ (.A(_2095_),
    .B(_2197_),
    .Y(_0296_));
 sg13g2_xnor2_1 _3023_ (.Y(_0297_),
    .A(\Pong.datapath.leftPaddle[8] ),
    .B(_2199_));
 sg13g2_xor2_1 _3024_ (.B(_2198_),
    .A(_0071_),
    .X(_0298_));
 sg13g2_xnor2_1 _3025_ (.Y(_0299_),
    .A(_1818_),
    .B(_2197_));
 sg13g2_xor2_1 _3026_ (.B(_0299_),
    .A(_0085_),
    .X(_0300_));
 sg13g2_xor2_1 _3027_ (.B(_0297_),
    .A(_0087_),
    .X(_0301_));
 sg13g2_xnor2_1 _3028_ (.Y(_0302_),
    .A(net681),
    .B(_0298_));
 sg13g2_nor3_1 _3029_ (.A(_0300_),
    .B(_0301_),
    .C(_0302_),
    .Y(_0303_));
 sg13g2_or3_1 _3030_ (.A(net708),
    .B(net710),
    .C(_2196_),
    .X(_0304_));
 sg13g2_nand2_1 _3031_ (.Y(_0305_),
    .A(_2197_),
    .B(_0304_));
 sg13g2_xnor2_1 _3032_ (.Y(_0306_),
    .A(_0084_),
    .B(_0305_));
 sg13g2_xor2_1 _3033_ (.B(_2196_),
    .A(_0074_),
    .X(_0307_));
 sg13g2_nor2_1 _3034_ (.A(_0083_),
    .B(_0307_),
    .Y(_0308_));
 sg13g2_xnor2_1 _3035_ (.Y(_0309_),
    .A(_1830_),
    .B(_0307_));
 sg13g2_nand2_1 _3036_ (.Y(_0310_),
    .A(_0306_),
    .B(_0309_));
 sg13g2_nor2_1 _3037_ (.A(_0079_),
    .B(_2194_),
    .Y(_0311_));
 sg13g2_xor2_1 _3038_ (.B(_0311_),
    .A(net711),
    .X(_0312_));
 sg13g2_nand2b_1 _3039_ (.Y(_0313_),
    .B(_1793_),
    .A_N(_0312_));
 sg13g2_and2_1 _3040_ (.A(net693),
    .B(_0312_),
    .X(_0314_));
 sg13g2_nand2_1 _3041_ (.Y(_0315_),
    .A(_0079_),
    .B(_2194_));
 sg13g2_xor2_1 _3042_ (.B(_2194_),
    .A(_0079_),
    .X(_0316_));
 sg13g2_xor2_1 _3043_ (.B(_0316_),
    .A(_0081_),
    .X(_0317_));
 sg13g2_o21ai_1 _3044_ (.B1(_0317_),
    .Y(_0318_),
    .A1(net693),
    .A2(_0312_));
 sg13g2_nor2_1 _3045_ (.A(_0314_),
    .B(_0318_),
    .Y(_0319_));
 sg13g2_nor2_1 _3046_ (.A(net699),
    .B(net717),
    .Y(_0320_));
 sg13g2_nor2_1 _3047_ (.A(net716),
    .B(net718),
    .Y(_0321_));
 sg13g2_or2_1 _3048_ (.X(_0322_),
    .B(net717),
    .A(net716));
 sg13g2_xnor2_1 _3049_ (.Y(_0323_),
    .A(net716),
    .B(net718));
 sg13g2_xnor2_1 _3050_ (.Y(_0324_),
    .A(_0096_),
    .B(_0323_));
 sg13g2_nand2b_1 _3051_ (.Y(_0325_),
    .B(_0324_),
    .A_N(_0320_));
 sg13g2_nand2_1 _3052_ (.Y(_0326_),
    .A(\Pong.datapath.vga.Row_Counter.Q[1] ),
    .B(_0323_));
 sg13g2_nand2_1 _3053_ (.Y(_0327_),
    .A(_0325_),
    .B(_0326_));
 sg13g2_nor2b_1 _3054_ (.A(_0316_),
    .B_N(net696),
    .Y(_0328_));
 sg13g2_a221oi_1 _3055_ (.B2(_0313_),
    .C1(_0314_),
    .B1(_0328_),
    .A1(_0319_),
    .Y(_0329_),
    .A2(_0327_));
 sg13g2_a22oi_1 _3056_ (.Y(_0330_),
    .B1(_0306_),
    .B2(_0308_),
    .A2(_0305_),
    .A1(\Pong.datapath.vga.Row_Counter.Q[5] ));
 sg13g2_o21ai_1 _3057_ (.B1(_0330_),
    .Y(_0331_),
    .A1(_0310_),
    .A2(_0329_));
 sg13g2_a22oi_1 _3058_ (.Y(_0332_),
    .B1(_0299_),
    .B2(net684),
    .A2(_0298_),
    .A1(net681));
 sg13g2_nor2_1 _3059_ (.A(_0301_),
    .B(_0332_),
    .Y(_0333_));
 sg13g2_o21ai_1 _3060_ (.B1(_0333_),
    .Y(_0334_),
    .A1(net681),
    .A2(_0298_));
 sg13g2_a22oi_1 _3061_ (.Y(_0335_),
    .B1(_0303_),
    .B2(_0331_),
    .A2(_0297_),
    .A1(net679));
 sg13g2_o21ai_1 _3062_ (.B1(_0319_),
    .Y(_0336_),
    .A1(_1795_),
    .A2(_1821_));
 sg13g2_nor3_1 _3063_ (.A(_0310_),
    .B(_0325_),
    .C(_0336_),
    .Y(_0337_));
 sg13g2_a22oi_1 _3064_ (.Y(_0338_),
    .B1(_0337_),
    .B2(_0303_),
    .A2(_0335_),
    .A1(_0334_));
 sg13g2_xnor2_1 _3065_ (.Y(_0339_),
    .A(net706),
    .B(_0296_));
 sg13g2_nor2_1 _3066_ (.A(_1788_),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_a22oi_1 _3067_ (.Y(_0341_),
    .B1(_0339_),
    .B2(_1788_),
    .A2(_0296_),
    .A1(\Pong.datapath.leftPaddle[9] ));
 sg13g2_o21ai_1 _3068_ (.B1(_0341_),
    .Y(_0342_),
    .A1(_0338_),
    .A2(_0340_));
 sg13g2_nor3_1 _3069_ (.A(net715),
    .B(net713),
    .C(net717),
    .Y(_0343_));
 sg13g2_nor2b_1 _3070_ (.A(_0343_),
    .B_N(net711),
    .Y(_0344_));
 sg13g2_nand2b_2 _3071_ (.Y(_0345_),
    .B(_2103_),
    .A_N(_0343_));
 sg13g2_nand2_1 _3072_ (.Y(_0346_),
    .A(_2108_),
    .B(_0345_));
 sg13g2_xor2_1 _3073_ (.B(_0346_),
    .A(net706),
    .X(_0347_));
 sg13g2_nor2b_1 _3074_ (.A(_2107_),
    .B_N(_0345_),
    .Y(_0348_));
 sg13g2_xnor2_1 _3075_ (.Y(_0349_),
    .A(_0070_),
    .B(_0348_));
 sg13g2_or2_1 _3076_ (.X(_0350_),
    .B(_0349_),
    .A(_0087_));
 sg13g2_o21ai_1 _3077_ (.B1(_0073_),
    .Y(_0351_),
    .A1(net708),
    .A2(_0345_));
 sg13g2_nor2_1 _3078_ (.A(net707),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_xnor2_1 _3079_ (.Y(_0353_),
    .A(_0071_),
    .B(_0352_));
 sg13g2_nand2_1 _3080_ (.Y(_0354_),
    .A(_1789_),
    .B(_0353_));
 sg13g2_xor2_1 _3081_ (.B(_0345_),
    .A(net709),
    .X(_0355_));
 sg13g2_nand2b_1 _3082_ (.Y(_0356_),
    .B(\Pong.datapath.vga.Row_Counter.Q[5] ),
    .A_N(_0355_));
 sg13g2_xnor2_1 _3083_ (.Y(_0357_),
    .A(_0079_),
    .B(_0322_));
 sg13g2_or2_1 _3084_ (.X(_0358_),
    .B(_0323_),
    .A(_1794_));
 sg13g2_o21ai_1 _3085_ (.B1(_0358_),
    .Y(_0359_),
    .A1(_0320_),
    .A2(_0324_));
 sg13g2_xnor2_1 _3086_ (.Y(_0360_),
    .A(_0081_),
    .B(_0357_));
 sg13g2_a22oi_1 _3087_ (.Y(_0361_),
    .B1(_0359_),
    .B2(_0360_),
    .A2(_0357_),
    .A1(net696));
 sg13g2_and2_1 _3088_ (.A(_1821_),
    .B(_2060_),
    .X(_0362_));
 sg13g2_nor2_1 _3089_ (.A(_0344_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_a21oi_1 _3090_ (.A1(_1793_),
    .A2(_0363_),
    .Y(_0364_),
    .B1(_0361_));
 sg13g2_xnor2_1 _3091_ (.Y(_0365_),
    .A(_1819_),
    .B(_0344_));
 sg13g2_o21ai_1 _3092_ (.B1(net693),
    .Y(_0366_),
    .A1(_0344_),
    .A2(_0362_));
 sg13g2_o21ai_1 _3093_ (.B1(_0366_),
    .Y(_0367_),
    .A1(net688),
    .A2(_0365_));
 sg13g2_xnor2_1 _3094_ (.Y(_0368_),
    .A(_0084_),
    .B(_0355_));
 sg13g2_a21oi_1 _3095_ (.A1(net688),
    .A2(_0365_),
    .Y(_0369_),
    .B1(_0368_));
 sg13g2_o21ai_1 _3096_ (.B1(_0369_),
    .Y(_0370_),
    .A1(_0364_),
    .A2(_0367_));
 sg13g2_xor2_1 _3097_ (.B(_0351_),
    .A(_0072_),
    .X(_0371_));
 sg13g2_xnor2_1 _3098_ (.Y(_0372_),
    .A(_0085_),
    .B(_0371_));
 sg13g2_a21oi_1 _3099_ (.A1(_0356_),
    .A2(_0370_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_nand2b_1 _3100_ (.Y(_0374_),
    .B(net684),
    .A_N(_0371_));
 sg13g2_o21ai_1 _3101_ (.B1(_0374_),
    .Y(_0375_),
    .A1(_1789_),
    .A2(_0353_));
 sg13g2_o21ai_1 _3102_ (.B1(_0354_),
    .Y(_0376_),
    .A1(_0373_),
    .A2(_0375_));
 sg13g2_xnor2_1 _3103_ (.Y(_0377_),
    .A(net675),
    .B(_0347_));
 sg13g2_a21o_1 _3104_ (.A2(_0349_),
    .A1(_0087_),
    .B1(_0377_),
    .X(_0378_));
 sg13g2_a21o_1 _3105_ (.A2(_0376_),
    .A1(_0350_),
    .B1(_0378_),
    .X(_0379_));
 sg13g2_o21ai_1 _3106_ (.B1(_0379_),
    .Y(_0380_),
    .A1(_1788_),
    .A2(_0347_));
 sg13g2_o21ai_1 _3107_ (.B1(_2147_),
    .Y(_0381_),
    .A1(net708),
    .A2(_0345_));
 sg13g2_nor2_1 _3108_ (.A(\Pong.datapath.vga.Column_Counter.Q[1] ),
    .B(net674),
    .Y(_0382_));
 sg13g2_or2_1 _3109_ (.X(_0383_),
    .B(net674),
    .A(\Pong.datapath.vga.Column_Counter.Q[1] ));
 sg13g2_nand3b_1 _3110_ (.B(_0382_),
    .C(net669),
    .Y(_0384_),
    .A_N(net672));
 sg13g2_nand2_2 _3111_ (.Y(_0385_),
    .A(\Pong.datapath.vga.Column_Counter.Q[5] ),
    .B(_1787_));
 sg13g2_o21ai_1 _3112_ (.B1(_1832_),
    .Y(_0386_),
    .A1(net670),
    .A2(_0385_));
 sg13g2_o21ai_1 _3113_ (.B1(_0386_),
    .Y(_0387_),
    .A1(_0384_),
    .A2(_0385_));
 sg13g2_nor2_2 _3114_ (.A(net659),
    .B(net660),
    .Y(_0388_));
 sg13g2_nor2_1 _3115_ (.A(net662),
    .B(net664),
    .Y(_0389_));
 sg13g2_nand2_1 _3116_ (.Y(_0390_),
    .A(net666),
    .B(net668));
 sg13g2_and2_1 _3117_ (.A(net669),
    .B(net671),
    .X(_0391_));
 sg13g2_o21ai_1 _3118_ (.B1(net666),
    .Y(_0392_),
    .A1(net667),
    .A2(_0391_));
 sg13g2_and4_2 _3119_ (.A(_0387_),
    .B(_0388_),
    .C(_0389_),
    .D(_0392_),
    .X(_0393_));
 sg13g2_nand4_1 _3120_ (.B(_0380_),
    .C(_0381_),
    .A(_0342_),
    .Y(_0394_),
    .D(_0393_));
 sg13g2_nand2_1 _3121_ (.Y(_0395_),
    .A(net729),
    .B(net731));
 sg13g2_and3_1 _3122_ (.X(_0396_),
    .A(net728),
    .B(net727),
    .C(net730));
 sg13g2_a21oi_2 _3123_ (.B1(_1815_),
    .Y(_0397_),
    .A2(_0396_),
    .A1(_1812_));
 sg13g2_a21oi_2 _3124_ (.B1(_1811_),
    .Y(_0398_),
    .A2(_0397_),
    .A1(_1813_));
 sg13g2_a21o_1 _3125_ (.A2(_0397_),
    .A1(_1813_),
    .B1(_1811_),
    .X(_0399_));
 sg13g2_a21oi_1 _3126_ (.A1(net726),
    .A2(_0398_),
    .Y(_0400_),
    .B1(_1814_));
 sg13g2_nor3_1 _3127_ (.A(_1810_),
    .B(_0059_),
    .C(_0399_),
    .Y(_0401_));
 sg13g2_nor3_1 _3128_ (.A(net681),
    .B(_0400_),
    .C(_0401_),
    .Y(_0402_));
 sg13g2_o21ai_1 _3129_ (.B1(net681),
    .Y(_0403_),
    .A1(_0400_),
    .A2(_0401_));
 sg13g2_xnor2_1 _3130_ (.Y(_0404_),
    .A(net726),
    .B(_0398_));
 sg13g2_xnor2_1 _3131_ (.Y(_0405_),
    .A(net682),
    .B(_0404_));
 sg13g2_nand3b_1 _3132_ (.B(_0403_),
    .C(_0405_),
    .Y(_0406_),
    .A_N(_0402_));
 sg13g2_nand3_1 _3133_ (.B(_1813_),
    .C(_0397_),
    .A(_1811_),
    .Y(_0407_));
 sg13g2_a21oi_1 _3134_ (.A1(_0399_),
    .A2(_0407_),
    .Y(_0408_),
    .B1(net685));
 sg13g2_and3_1 _3135_ (.X(_0409_),
    .A(net685),
    .B(_0399_),
    .C(_0407_));
 sg13g2_nor2_1 _3136_ (.A(_0408_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_xnor2_1 _3137_ (.Y(_0411_),
    .A(_0065_),
    .B(_0397_));
 sg13g2_and2_1 _3138_ (.A(net688),
    .B(_0411_),
    .X(_0412_));
 sg13g2_nor2_1 _3139_ (.A(net688),
    .B(_0411_),
    .Y(_0413_));
 sg13g2_nor4_1 _3140_ (.A(_0408_),
    .B(_0409_),
    .C(_0412_),
    .D(_0413_),
    .Y(_0414_));
 sg13g2_nand3b_1 _3141_ (.B(net731),
    .C(net729),
    .Y(_0415_),
    .A_N(_0077_));
 sg13g2_xnor2_1 _3142_ (.Y(_0416_),
    .A(\Pong.datapath.rightPaddle[3] ),
    .B(_0415_));
 sg13g2_and2_1 _3143_ (.A(net693),
    .B(_0416_),
    .X(_0417_));
 sg13g2_nand2b_1 _3144_ (.Y(_0418_),
    .B(_1793_),
    .A_N(_0416_));
 sg13g2_nand2_1 _3145_ (.Y(_0419_),
    .A(_0077_),
    .B(_0395_));
 sg13g2_xor2_1 _3146_ (.B(_0395_),
    .A(_0077_),
    .X(_0420_));
 sg13g2_xor2_1 _3147_ (.B(_0420_),
    .A(_0081_),
    .X(_0421_));
 sg13g2_nand3b_1 _3148_ (.B(_0418_),
    .C(_0421_),
    .Y(_0422_),
    .A_N(_0417_));
 sg13g2_nor2_1 _3149_ (.A(net699),
    .B(net730),
    .Y(_0423_));
 sg13g2_or2_1 _3150_ (.X(_0424_),
    .B(net730),
    .A(net699));
 sg13g2_or2_1 _3151_ (.X(_0425_),
    .B(net731),
    .A(net729));
 sg13g2_xnor2_1 _3152_ (.Y(_0426_),
    .A(net729),
    .B(net731));
 sg13g2_xnor2_1 _3153_ (.Y(_0427_),
    .A(_0096_),
    .B(_0426_));
 sg13g2_a22oi_1 _3154_ (.Y(_0428_),
    .B1(_0427_),
    .B2(_0424_),
    .A2(_0426_),
    .A1(\Pong.datapath.vga.Row_Counter.Q[1] ));
 sg13g2_nor2b_1 _3155_ (.A(_0420_),
    .B_N(net696),
    .Y(_0429_));
 sg13g2_o21ai_1 _3156_ (.B1(_0418_),
    .Y(_0430_),
    .A1(_0417_),
    .A2(_0429_));
 sg13g2_o21ai_1 _3157_ (.B1(_0430_),
    .Y(_0431_),
    .A1(_0422_),
    .A2(_0428_));
 sg13g2_a21oi_1 _3158_ (.A1(_0399_),
    .A2(_0407_),
    .Y(_0432_),
    .B1(_1791_));
 sg13g2_a221oi_1 _3159_ (.B2(_0431_),
    .C1(_0432_),
    .B1(_0414_),
    .A1(_0410_),
    .Y(_0433_),
    .A2(_0413_));
 sg13g2_nand2_1 _3160_ (.Y(_0434_),
    .A(net684),
    .B(_0404_));
 sg13g2_a21o_1 _3161_ (.A2(_0434_),
    .A1(_0403_),
    .B1(_0402_),
    .X(_0435_));
 sg13g2_o21ai_1 _3162_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0406_),
    .A2(_0433_));
 sg13g2_nand3_1 _3163_ (.B(net726),
    .C(_0398_),
    .A(net724),
    .Y(_0437_));
 sg13g2_nor2_1 _3164_ (.A(_1809_),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_xnor2_1 _3165_ (.Y(_0439_),
    .A(_1809_),
    .B(_0437_));
 sg13g2_xnor2_1 _3166_ (.Y(_0440_),
    .A(net678),
    .B(_0439_));
 sg13g2_a22oi_1 _3167_ (.Y(_0441_),
    .B1(_0440_),
    .B2(_0436_),
    .A2(_0439_),
    .A1(\Pong.datapath.vga.Row_Counter.Q[8] ));
 sg13g2_xor2_1 _3168_ (.B(_0438_),
    .A(_0056_),
    .X(_0442_));
 sg13g2_nand2_1 _3169_ (.Y(_0443_),
    .A(net699),
    .B(net730));
 sg13g2_nand3_1 _3170_ (.B(_0427_),
    .C(_0443_),
    .A(_0424_),
    .Y(_0444_));
 sg13g2_nor2_1 _3171_ (.A(_0422_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_and2_1 _3172_ (.A(_0414_),
    .B(_0445_),
    .X(_0446_));
 sg13g2_nand3b_1 _3173_ (.B(_0440_),
    .C(_0446_),
    .Y(_0447_),
    .A_N(_0406_));
 sg13g2_o21ai_1 _3174_ (.B1(_0447_),
    .Y(_0448_),
    .A1(net677),
    .A2(_0442_));
 sg13g2_nand2_1 _3175_ (.Y(_0449_),
    .A(net677),
    .B(_0442_));
 sg13g2_o21ai_1 _3176_ (.B1(_0449_),
    .Y(_0450_),
    .A1(_0441_),
    .A2(_0448_));
 sg13g2_nand2_1 _3177_ (.Y(_0451_),
    .A(\Pong.datapath.rightPaddle[9] ),
    .B(_0438_));
 sg13g2_or3_1 _3178_ (.A(net728),
    .B(net727),
    .C(net730),
    .X(_0452_));
 sg13g2_nand2_1 _3179_ (.Y(_0453_),
    .A(\Pong.datapath.rightPaddle[3] ),
    .B(_0452_));
 sg13g2_nand3_1 _3180_ (.B(\Pong.datapath.rightPaddle[4] ),
    .C(_0452_),
    .A(\Pong.datapath.rightPaddle[3] ),
    .Y(_0454_));
 sg13g2_xnor2_1 _3181_ (.Y(_0455_),
    .A(_1811_),
    .B(_0454_));
 sg13g2_nor2_1 _3182_ (.A(_1791_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_xnor2_1 _3183_ (.Y(_0457_),
    .A(_0077_),
    .B(_0425_));
 sg13g2_or2_1 _3184_ (.X(_0458_),
    .B(_0426_),
    .A(_1794_));
 sg13g2_o21ai_1 _3185_ (.B1(_0458_),
    .Y(_0459_),
    .A1(_0423_),
    .A2(_0427_));
 sg13g2_xnor2_1 _3186_ (.Y(_0460_),
    .A(net694),
    .B(_0457_));
 sg13g2_a22oi_1 _3187_ (.Y(_0461_),
    .B1(_0459_),
    .B2(_0460_),
    .A2(_0457_),
    .A1(net696));
 sg13g2_o21ai_1 _3188_ (.B1(_0453_),
    .Y(_0462_),
    .A1(net730),
    .A2(_2010_));
 sg13g2_nor2_1 _3189_ (.A(net693),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_xnor2_1 _3190_ (.Y(_0464_),
    .A(_1813_),
    .B(_0453_));
 sg13g2_a22oi_1 _3191_ (.Y(_0465_),
    .B1(_0464_),
    .B2(_1830_),
    .A2(_0462_),
    .A1(net693));
 sg13g2_o21ai_1 _3192_ (.B1(_0465_),
    .Y(_0466_),
    .A1(_0461_),
    .A2(_0463_));
 sg13g2_nor2_1 _3193_ (.A(_1830_),
    .B(_0464_),
    .Y(_0467_));
 sg13g2_xnor2_1 _3194_ (.Y(_0468_),
    .A(net685),
    .B(_0455_));
 sg13g2_nor2_1 _3195_ (.A(_0467_),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_a21o_1 _3196_ (.A2(_0469_),
    .A1(_0466_),
    .B1(_0456_),
    .X(_0470_));
 sg13g2_o21ai_1 _3197_ (.B1(_0061_),
    .Y(_0471_),
    .A1(\Pong.datapath.rightPaddle[5] ),
    .A2(_0454_));
 sg13g2_xnor2_1 _3198_ (.Y(_0472_),
    .A(_0060_),
    .B(_0471_));
 sg13g2_xnor2_1 _3199_ (.Y(_0473_),
    .A(net682),
    .B(_0472_));
 sg13g2_nor2_1 _3200_ (.A(net726),
    .B(_0471_),
    .Y(_0474_));
 sg13g2_xnor2_1 _3201_ (.Y(_0475_),
    .A(_0059_),
    .B(_0474_));
 sg13g2_nor2_1 _3202_ (.A(_1789_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_a221oi_1 _3203_ (.B2(_0470_),
    .C1(_0476_),
    .B1(_0473_),
    .A1(net684),
    .Y(_0477_),
    .A2(_0472_));
 sg13g2_a21oi_1 _3204_ (.A1(_1789_),
    .A2(_0475_),
    .Y(_0478_),
    .B1(_0477_));
 sg13g2_nand2_1 _3205_ (.Y(_0479_),
    .A(_1965_),
    .B(_0454_));
 sg13g2_xor2_1 _3206_ (.B(_0479_),
    .A(_0058_),
    .X(_0480_));
 sg13g2_nor2_1 _3207_ (.A(net678),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_nand2_1 _3208_ (.Y(_0482_),
    .A(_1966_),
    .B(_0454_));
 sg13g2_xor2_1 _3209_ (.B(_0482_),
    .A(_0056_),
    .X(_0483_));
 sg13g2_xnor2_1 _3210_ (.Y(_0484_),
    .A(net675),
    .B(_0483_));
 sg13g2_a21oi_1 _3211_ (.A1(net678),
    .A2(_0480_),
    .Y(_0485_),
    .B1(_0484_));
 sg13g2_o21ai_1 _3212_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_0478_),
    .A2(_0481_));
 sg13g2_nand2b_1 _3213_ (.Y(_0487_),
    .B(net677),
    .A_N(_0483_));
 sg13g2_nand2b_2 _3214_ (.Y(_0488_),
    .B(net665),
    .A_N(net663));
 sg13g2_nand2b_1 _3215_ (.Y(_0489_),
    .B(net671),
    .A_N(net669));
 sg13g2_o21ai_1 _3216_ (.B1(_0090_),
    .Y(_0490_),
    .A1(_0382_),
    .A2(_0489_));
 sg13g2_nand3b_1 _3217_ (.B(net667),
    .C(_0490_),
    .Y(_0491_),
    .A_N(net666));
 sg13g2_a21o_1 _3218_ (.A2(_0491_),
    .A1(_0092_),
    .B1(_0488_),
    .X(_0492_));
 sg13g2_nor2b_1 _3219_ (.A(net660),
    .B_N(_0094_),
    .Y(_0493_));
 sg13g2_o21ai_1 _3220_ (.B1(_2055_),
    .Y(_0494_),
    .A1(\Pong.datapath.rightPaddle[5] ),
    .A2(_0454_));
 sg13g2_nand2_1 _3221_ (.Y(_0495_),
    .A(net658),
    .B(_0095_));
 sg13g2_nand2_1 _3222_ (.Y(_0496_),
    .A(net667),
    .B(net669));
 sg13g2_nand4_1 _3223_ (.B(net667),
    .C(net669),
    .A(net664),
    .Y(_0497_),
    .D(_0384_));
 sg13g2_nor2b_1 _3224_ (.A(net660),
    .B_N(net658),
    .Y(_0498_));
 sg13g2_a21oi_1 _3225_ (.A1(net664),
    .A2(net666),
    .Y(_0499_),
    .B1(net663));
 sg13g2_nand3_1 _3226_ (.B(_0498_),
    .C(_0499_),
    .A(_0497_),
    .Y(_0500_));
 sg13g2_a22oi_1 _3227_ (.Y(_0501_),
    .B1(_0495_),
    .B2(_0500_),
    .A2(_0493_),
    .A1(_0492_));
 sg13g2_nand2_1 _3228_ (.Y(_0502_),
    .A(_0494_),
    .B(_0501_));
 sg13g2_a221oi_1 _3229_ (.B2(_0487_),
    .C1(_0502_),
    .B1(_0486_),
    .A1(_0450_),
    .Y(_0503_),
    .A2(_0451_));
 sg13g2_nor2_1 _3230_ (.A(net676),
    .B(_1795_),
    .Y(_0504_));
 sg13g2_a21oi_1 _3231_ (.A1(net695),
    .A2(_0504_),
    .Y(_0505_),
    .B1(_0088_));
 sg13g2_or2_1 _3232_ (.X(_0506_),
    .B(net695),
    .A(net692));
 sg13g2_nor2_1 _3233_ (.A(net686),
    .B(_0506_),
    .Y(_0507_));
 sg13g2_nand2_1 _3234_ (.Y(_0508_),
    .A(net680),
    .B(net683));
 sg13g2_and3_2 _3235_ (.X(_0509_),
    .A(net679),
    .B(net680),
    .C(net683));
 sg13g2_nand3_1 _3236_ (.B(net680),
    .C(net683),
    .A(net679),
    .Y(_0510_));
 sg13g2_a21oi_1 _3237_ (.A1(_1791_),
    .A2(_1792_),
    .Y(_0511_),
    .B1(_0510_));
 sg13g2_o21ai_1 _3238_ (.B1(_0509_),
    .Y(_0512_),
    .A1(net686),
    .A2(net689));
 sg13g2_o21ai_1 _3239_ (.B1(_0088_),
    .Y(_0513_),
    .A1(_0507_),
    .A2(_0512_));
 sg13g2_nand2_1 _3240_ (.Y(_0514_),
    .A(net689),
    .B(_1794_));
 sg13g2_nor4_1 _3241_ (.A(net686),
    .B(net692),
    .C(_0510_),
    .D(_0514_),
    .Y(_0515_));
 sg13g2_nand2b_1 _3242_ (.Y(_0516_),
    .B(_0515_),
    .A_N(_0505_));
 sg13g2_nor2_1 _3243_ (.A(net676),
    .B(_0509_),
    .Y(_0517_));
 sg13g2_nor2_1 _3244_ (.A(net676),
    .B(net689),
    .Y(_0518_));
 sg13g2_and2_1 _3245_ (.A(_0507_),
    .B(_0509_),
    .X(_0519_));
 sg13g2_and2_1 _3246_ (.A(_1794_),
    .B(_0519_),
    .X(_0520_));
 sg13g2_a221oi_1 _3247_ (.B2(_0520_),
    .C1(_0517_),
    .B1(_0518_),
    .A1(_0513_),
    .Y(_0521_),
    .A2(_0516_));
 sg13g2_nor2_1 _3248_ (.A(\Pong.datapath.scoreLeft[2] ),
    .B(\Pong.datapath.scoreLeft[1] ),
    .Y(_0522_));
 sg13g2_nor2_1 _3249_ (.A(_1824_),
    .B(_0522_),
    .Y(_0523_));
 sg13g2_nor2b_1 _3250_ (.A(\Pong.datapath.scoreLeft[1] ),
    .B_N(\Pong.datapath.scoreLeft[2] ),
    .Y(_0524_));
 sg13g2_nor3_1 _3251_ (.A(\Pong.datapath.scoreLeft[0] ),
    .B(_0523_),
    .C(_0524_),
    .Y(_0525_));
 sg13g2_and3_1 _3252_ (.X(_0526_),
    .A(net679),
    .B(net680),
    .C(net687));
 sg13g2_nand3_1 _3253_ (.B(net680),
    .C(net686),
    .A(net679),
    .Y(_0527_));
 sg13g2_nand2_1 _3254_ (.Y(_0528_),
    .A(_0517_),
    .B(_0527_));
 sg13g2_nor4_2 _3255_ (.A(net676),
    .B(net683),
    .C(net690),
    .Y(_0529_),
    .D(_0527_));
 sg13g2_nand2_2 _3256_ (.Y(_0530_),
    .A(net697),
    .B(net698));
 sg13g2_nand3_1 _3257_ (.B(net697),
    .C(net698),
    .A(net691),
    .Y(_0531_));
 sg13g2_nand4_1 _3258_ (.B(net695),
    .C(net697),
    .A(net691),
    .Y(_0532_),
    .D(net698));
 sg13g2_a22oi_1 _3259_ (.Y(_0533_),
    .B1(_0529_),
    .B2(_0532_),
    .A2(_0527_),
    .A1(_0517_));
 sg13g2_and4_1 _3260_ (.A(net691),
    .B(net696),
    .C(net697),
    .D(_1795_),
    .X(_0534_));
 sg13g2_a21oi_2 _3261_ (.B1(_0533_),
    .Y(_0535_),
    .A2(_0534_),
    .A1(_0529_));
 sg13g2_and2_1 _3262_ (.A(net675),
    .B(_0510_),
    .X(_0536_));
 sg13g2_nor2_1 _3263_ (.A(net675),
    .B(_0504_),
    .Y(_0537_));
 sg13g2_a21oi_1 _3264_ (.A1(_1792_),
    .A2(_0520_),
    .Y(_0538_),
    .B1(_0536_));
 sg13g2_nor3_2 _3265_ (.A(_0535_),
    .B(_0537_),
    .C(_0538_),
    .Y(_0539_));
 sg13g2_a21oi_1 _3266_ (.A1(\Pong.datapath.scoreLeft[2] ),
    .A2(_1824_),
    .Y(_0540_),
    .B1(_0522_));
 sg13g2_nand2_1 _3267_ (.Y(_0541_),
    .A(_1824_),
    .B(\Pong.datapath.scoreLeft[0] ));
 sg13g2_nor2_1 _3268_ (.A(_0524_),
    .B(_0541_),
    .Y(_0542_));
 sg13g2_nor2_1 _3269_ (.A(_0540_),
    .B(_0542_),
    .Y(_0543_));
 sg13g2_a22oi_1 _3270_ (.Y(_0544_),
    .B1(_0539_),
    .B2(_0543_),
    .A2(_0525_),
    .A1(_0521_));
 sg13g2_nand2_1 _3271_ (.Y(_0545_),
    .A(net671),
    .B(_0383_));
 sg13g2_a21oi_1 _3272_ (.A1(net671),
    .A2(_0383_),
    .Y(_0546_),
    .B1(net669));
 sg13g2_nor2_1 _3273_ (.A(_0388_),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_nor3_2 _3274_ (.A(net662),
    .B(net664),
    .C(net666),
    .Y(_0548_));
 sg13g2_nand2b_1 _3275_ (.Y(_0549_),
    .B(net660),
    .A_N(net659));
 sg13g2_nor2_1 _3276_ (.A(net667),
    .B(_0549_),
    .Y(_0550_));
 sg13g2_nor3_1 _3277_ (.A(net664),
    .B(net666),
    .C(net668),
    .Y(_0551_));
 sg13g2_nand2_1 _3278_ (.Y(_0552_),
    .A(_0548_),
    .B(_0550_));
 sg13g2_a21oi_1 _3279_ (.A1(_0548_),
    .A2(_0550_),
    .Y(_0553_),
    .B1(_0388_));
 sg13g2_or2_1 _3280_ (.X(_0554_),
    .B(_0489_),
    .A(_0383_));
 sg13g2_nor2_1 _3281_ (.A(_0552_),
    .B(_0554_),
    .Y(_0555_));
 sg13g2_nor3_1 _3282_ (.A(_0547_),
    .B(_0553_),
    .C(_0555_),
    .Y(_0556_));
 sg13g2_nand2b_1 _3283_ (.Y(_0557_),
    .B(_0095_),
    .A_N(net661));
 sg13g2_nand2_1 _3284_ (.Y(_0558_),
    .A(net661),
    .B(_0548_));
 sg13g2_or2_1 _3285_ (.X(_0559_),
    .B(_0558_),
    .A(net670));
 sg13g2_nor2b_1 _3286_ (.A(net659),
    .B_N(net674),
    .Y(_0560_));
 sg13g2_and3_1 _3287_ (.X(_0561_),
    .A(net671),
    .B(net673),
    .C(_0560_));
 sg13g2_o21ai_1 _3288_ (.B1(_0557_),
    .Y(_0562_),
    .A1(net667),
    .A2(_0559_));
 sg13g2_o21ai_1 _3289_ (.B1(_0562_),
    .Y(_0563_),
    .A1(net657),
    .A2(_0561_));
 sg13g2_nor3_1 _3290_ (.A(_0544_),
    .B(_0556_),
    .C(_0563_),
    .Y(_0564_));
 sg13g2_nor2b_1 _3291_ (.A(\Pong.datapath.scoreRight[3] ),
    .B_N(\Pong.datapath.scoreRight[0] ),
    .Y(_0565_));
 sg13g2_nand2_1 _3292_ (.Y(_0566_),
    .A(_1823_),
    .B(\Pong.datapath.scoreRight[0] ));
 sg13g2_nor2_2 _3293_ (.A(\Pong.datapath.scoreRight[2] ),
    .B(\Pong.datapath.scoreRight[1] ),
    .Y(_0567_));
 sg13g2_or2_1 _3294_ (.X(_0568_),
    .B(\Pong.datapath.scoreRight[1] ),
    .A(\Pong.datapath.scoreRight[2] ));
 sg13g2_a21oi_1 _3295_ (.A1(\Pong.datapath.scoreRight[2] ),
    .A2(_1823_),
    .Y(_0569_),
    .B1(_0567_));
 sg13g2_nand2_1 _3296_ (.Y(_0570_),
    .A(_0566_),
    .B(_0569_));
 sg13g2_and2_1 _3297_ (.A(\Pong.datapath.scoreRight[2] ),
    .B(\Pong.datapath.scoreRight[1] ),
    .X(_0571_));
 sg13g2_nand2_1 _3298_ (.Y(_0572_),
    .A(_0565_),
    .B(_0571_));
 sg13g2_nand3_1 _3299_ (.B(\Pong.datapath.scoreRight[0] ),
    .C(_0567_),
    .A(\Pong.datapath.scoreRight[3] ),
    .Y(_0573_));
 sg13g2_nand2_1 _3300_ (.Y(_0574_),
    .A(_0572_),
    .B(_0573_));
 sg13g2_o21ai_1 _3301_ (.B1(\Pong.datapath.scoreRight[3] ),
    .Y(_0575_),
    .A1(\Pong.datapath.scoreRight[0] ),
    .A2(_0568_));
 sg13g2_o21ai_1 _3302_ (.B1(\Pong.datapath.scoreRight[2] ),
    .Y(_0576_),
    .A1(\Pong.datapath.scoreRight[1] ),
    .A2(\Pong.datapath.scoreRight[0] ));
 sg13g2_a21o_1 _3303_ (.A2(_0576_),
    .A1(_0575_),
    .B1(_0574_),
    .X(_0577_));
 sg13g2_a22oi_1 _3304_ (.Y(_0578_),
    .B1(_0577_),
    .B2(_0539_),
    .A2(_0570_),
    .A1(_0521_));
 sg13g2_nand4_1 _3305_ (.B(net666),
    .C(net668),
    .A(net664),
    .Y(_0579_),
    .D(net669));
 sg13g2_nor2_1 _3306_ (.A(net659),
    .B(net662),
    .Y(_0580_));
 sg13g2_o21ai_1 _3307_ (.B1(_0580_),
    .Y(_0581_),
    .A1(_0545_),
    .A2(_0579_));
 sg13g2_nand2b_1 _3308_ (.Y(_0582_),
    .B(_0581_),
    .A_N(_0388_));
 sg13g2_nor2b_1 _3309_ (.A(net662),
    .B_N(net657),
    .Y(_0583_));
 sg13g2_nor3_1 _3310_ (.A(net671),
    .B(net673),
    .C(_0560_),
    .Y(_0584_));
 sg13g2_o21ai_1 _3311_ (.B1(_0583_),
    .Y(_0585_),
    .A1(_0579_),
    .A2(_0584_));
 sg13g2_nand3_1 _3312_ (.B(_0582_),
    .C(_0585_),
    .A(_0557_),
    .Y(_0586_));
 sg13g2_nor2_1 _3313_ (.A(_0578_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_nand2_2 _3314_ (.Y(_0588_),
    .A(net667),
    .B(_0548_));
 sg13g2_o21ai_1 _3315_ (.B1(_0388_),
    .Y(_0589_),
    .A1(_0554_),
    .A2(_0588_));
 sg13g2_o21ai_1 _3316_ (.B1(_0548_),
    .Y(_0590_),
    .A1(_1787_),
    .A2(_0546_));
 sg13g2_o21ai_1 _3317_ (.B1(_0493_),
    .Y(_0591_),
    .A1(_0392_),
    .A2(_0488_));
 sg13g2_nor2_1 _3318_ (.A(_0385_),
    .B(_0488_),
    .Y(_0592_));
 sg13g2_nand4_1 _3319_ (.B(_0391_),
    .C(_0498_),
    .A(_0382_),
    .Y(_0593_),
    .D(_0592_));
 sg13g2_nand3_1 _3320_ (.B(_0591_),
    .C(_0593_),
    .A(net658),
    .Y(_0594_));
 sg13g2_o21ai_1 _3321_ (.B1(_0594_),
    .Y(_0595_),
    .A1(_0589_),
    .A2(_0590_));
 sg13g2_nand2_2 _3322_ (.Y(_0596_),
    .A(_1794_),
    .B(_1795_));
 sg13g2_nand2_2 _3323_ (.Y(_0597_),
    .A(_1793_),
    .B(net696));
 sg13g2_nor4_2 _3324_ (.A(net679),
    .B(net680),
    .C(net683),
    .Y(_0598_),
    .D(net686));
 sg13g2_and2_1 _3325_ (.A(_1788_),
    .B(_0598_),
    .X(_0599_));
 sg13g2_a21oi_1 _3326_ (.A1(net689),
    .A2(_0599_),
    .Y(_0600_),
    .B1(_0529_));
 sg13g2_nor4_1 _3327_ (.A(_0595_),
    .B(_0596_),
    .C(_0597_),
    .D(_0600_),
    .Y(_0601_));
 sg13g2_a21oi_1 _3328_ (.A1(net695),
    .A2(_0596_),
    .Y(_0602_),
    .B1(net691));
 sg13g2_nand2_1 _3329_ (.Y(_0603_),
    .A(_0529_),
    .B(_0602_));
 sg13g2_nand2_1 _3330_ (.Y(_0604_),
    .A(net689),
    .B(_0506_));
 sg13g2_and2_1 _3331_ (.A(_0599_),
    .B(_0604_),
    .X(_0605_));
 sg13g2_or4_1 _3332_ (.A(net658),
    .B(net660),
    .C(_0554_),
    .D(_0588_),
    .X(_0606_));
 sg13g2_a221oi_1 _3333_ (.B2(_0593_),
    .C1(_0605_),
    .B1(_0606_),
    .A1(_0528_),
    .Y(_0607_),
    .A2(_0603_));
 sg13g2_nor4_1 _3334_ (.A(_0564_),
    .B(_0587_),
    .C(_0601_),
    .D(_0607_),
    .Y(_0608_));
 sg13g2_xnor2_1 _3335_ (.Y(_0609_),
    .A(net619),
    .B(net685));
 sg13g2_xnor2_1 _3336_ (.Y(_0610_),
    .A(_1958_),
    .B(net589));
 sg13g2_xnor2_1 _3337_ (.Y(_0611_),
    .A(_0086_),
    .B(_0097_));
 sg13g2_nor3_1 _3338_ (.A(net620),
    .B(net623),
    .C(_1953_),
    .Y(_0612_));
 sg13g2_or3_2 _3339_ (.A(net620),
    .B(net623),
    .C(_1953_),
    .X(_0613_));
 sg13g2_nor2_1 _3340_ (.A(net593),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_nor3_2 _3341_ (.A(net618),
    .B(net593),
    .C(_0613_),
    .Y(_0615_));
 sg13g2_xor2_1 _3342_ (.B(net678),
    .A(net610),
    .X(_0616_));
 sg13g2_xnor2_1 _3343_ (.Y(_0617_),
    .A(net610),
    .B(net678));
 sg13g2_or3_2 _3344_ (.A(net615),
    .B(net618),
    .C(_0613_),
    .X(_0618_));
 sg13g2_nor2_1 _3345_ (.A(net629),
    .B(_0618_),
    .Y(_0619_));
 sg13g2_or2_1 _3346_ (.X(_0620_),
    .B(_0618_),
    .A(net593));
 sg13g2_nand2_1 _3347_ (.Y(_0621_),
    .A(_0616_),
    .B(_0620_));
 sg13g2_nor2b_2 _3348_ (.A(net617),
    .B_N(net682),
    .Y(_0622_));
 sg13g2_nor2b_2 _3349_ (.A(net682),
    .B_N(net616),
    .Y(_0623_));
 sg13g2_nor2_2 _3350_ (.A(_0622_),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_or2_2 _3351_ (.X(_0625_),
    .B(_0623_),
    .A(_0622_));
 sg13g2_nor2_1 _3352_ (.A(net629),
    .B(_0613_),
    .Y(_0626_));
 sg13g2_xnor2_1 _3353_ (.Y(_0627_),
    .A(_0068_),
    .B(_0082_));
 sg13g2_a22oi_1 _3354_ (.Y(_0628_),
    .B1(_0627_),
    .B2(_1905_),
    .A2(_0626_),
    .A1(_0624_));
 sg13g2_xor2_1 _3355_ (.B(net698),
    .A(net631),
    .X(_0629_));
 sg13g2_and2_1 _3356_ (.A(net628),
    .B(net631),
    .X(_0630_));
 sg13g2_nand2_2 _3357_ (.Y(_0631_),
    .A(net628),
    .B(net631));
 sg13g2_nor2_2 _3358_ (.A(_1950_),
    .B(net585),
    .Y(_0632_));
 sg13g2_xnor2_1 _3359_ (.Y(_0633_),
    .A(_0096_),
    .B(_0632_));
 sg13g2_and2_1 _3360_ (.A(_0629_),
    .B(_0633_),
    .X(_0634_));
 sg13g2_xor2_1 _3361_ (.B(net688),
    .A(net621),
    .X(_0635_));
 sg13g2_nand2b_1 _3362_ (.Y(_0636_),
    .B(_0625_),
    .A_N(_0614_));
 sg13g2_xor2_1 _3363_ (.B(net694),
    .A(_0067_),
    .X(_0637_));
 sg13g2_o21ai_1 _3364_ (.B1(_0616_),
    .Y(_0638_),
    .A1(net608),
    .A2(net612));
 sg13g2_inv_1 _3365_ (.Y(_0639_),
    .A(_0638_));
 sg13g2_o21ai_1 _3366_ (.B1(_0637_),
    .Y(_0640_),
    .A1(_0618_),
    .A2(_0639_));
 sg13g2_xnor2_1 _3367_ (.Y(_0641_),
    .A(_1950_),
    .B(_0637_));
 sg13g2_nand2b_1 _3368_ (.Y(_0642_),
    .B(_0113_),
    .A_N(net675));
 sg13g2_xnor2_1 _3369_ (.Y(_0643_),
    .A(_0113_),
    .B(net675));
 sg13g2_nor3_1 _3370_ (.A(net612),
    .B(net628),
    .C(_0618_),
    .Y(_0644_));
 sg13g2_nor2_1 _3371_ (.A(net612),
    .B(_0620_),
    .Y(_0645_));
 sg13g2_inv_1 _3372_ (.Y(_0646_),
    .A(_0645_));
 sg13g2_xnor2_1 _3373_ (.Y(_0647_),
    .A(net582),
    .B(_0645_));
 sg13g2_xnor2_1 _3374_ (.Y(_0648_),
    .A(net627),
    .B(net696));
 sg13g2_xnor2_1 _3375_ (.Y(_0649_),
    .A(net613),
    .B(net679));
 sg13g2_xnor2_1 _3376_ (.Y(_0650_),
    .A(net608),
    .B(net676));
 sg13g2_xnor2_1 _3377_ (.Y(_0651_),
    .A(net623),
    .B(\Pong.datapath.vga.Row_Counter.Q[4] ));
 sg13g2_xor2_1 _3378_ (.B(net697),
    .A(net630),
    .X(_0652_));
 sg13g2_xnor2_1 _3379_ (.Y(_0653_),
    .A(\Pong.datapath.ballFunction.ball_center_y[1] ),
    .B(net697));
 sg13g2_xnor2_1 _3380_ (.Y(_0654_),
    .A(net614),
    .B(net680));
 sg13g2_xnor2_1 _3381_ (.Y(_0655_),
    .A(\Pong.datapath.ballFunction.ball_center_y[6] ),
    .B(net683));
 sg13g2_xnor2_1 _3382_ (.Y(_0656_),
    .A(net624),
    .B(net692));
 sg13g2_xnor2_1 _3383_ (.Y(_0657_),
    .A(net620),
    .B(net687));
 sg13g2_nand4_1 _3384_ (.B(_0654_),
    .C(_0655_),
    .A(_0649_),
    .Y(_0658_),
    .D(_0657_));
 sg13g2_nand4_1 _3385_ (.B(_0650_),
    .C(_0651_),
    .A(_0648_),
    .Y(_0659_),
    .D(_0656_));
 sg13g2_nor4_1 _3386_ (.A(_0629_),
    .B(_0652_),
    .C(_0658_),
    .D(_0659_),
    .Y(_0660_));
 sg13g2_nand2_2 _3387_ (.Y(_0661_),
    .A(net624),
    .B(net626));
 sg13g2_nor2_1 _3388_ (.A(net621),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_nand2_2 _3389_ (.Y(_0663_),
    .A(net627),
    .B(net628));
 sg13g2_nand2_1 _3390_ (.Y(_0664_),
    .A(net625),
    .B(net585));
 sg13g2_or2_1 _3391_ (.X(_0665_),
    .B(_0661_),
    .A(_0631_));
 sg13g2_nor2_1 _3392_ (.A(net621),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_xnor2_1 _3393_ (.Y(_0667_),
    .A(net619),
    .B(_0666_));
 sg13g2_nor2_1 _3394_ (.A(net685),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_nor2_1 _3395_ (.A(net625),
    .B(net585),
    .Y(_0669_));
 sg13g2_xnor2_1 _3396_ (.Y(_0670_),
    .A(net625),
    .B(net585));
 sg13g2_xor2_1 _3397_ (.B(_0664_),
    .A(net586),
    .X(_0671_));
 sg13g2_and2_1 _3398_ (.A(net685),
    .B(_0667_),
    .X(_0672_));
 sg13g2_nand2_1 _3399_ (.Y(_0673_),
    .A(net615),
    .B(net618));
 sg13g2_nand4_1 _3400_ (.B(net623),
    .C(net624),
    .A(net620),
    .Y(_0674_),
    .D(net625));
 sg13g2_nor2_1 _3401_ (.A(_0631_),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_or2_2 _3402_ (.X(_0676_),
    .B(_0674_),
    .A(_0673_));
 sg13g2_nor2_1 _3403_ (.A(_0631_),
    .B(_0676_),
    .Y(_0677_));
 sg13g2_nor2_1 _3404_ (.A(net610),
    .B(_0676_),
    .Y(_0678_));
 sg13g2_nor3_2 _3405_ (.A(net610),
    .B(_0631_),
    .C(_0676_),
    .Y(_0679_));
 sg13g2_xnor2_1 _3406_ (.Y(_0680_),
    .A(net584),
    .B(_0665_));
 sg13g2_nand2b_1 _3407_ (.Y(_0681_),
    .B(_0629_),
    .A_N(_0633_));
 sg13g2_a21oi_1 _3408_ (.A1(net608),
    .A2(net612),
    .Y(_0682_),
    .B1(_0617_));
 sg13g2_nor2_1 _3409_ (.A(_0676_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_nor3_2 _3410_ (.A(net616),
    .B(_0631_),
    .C(_0674_),
    .Y(_0684_));
 sg13g2_xnor2_1 _3411_ (.Y(_0685_),
    .A(_0625_),
    .B(_0675_));
 sg13g2_nor2_1 _3412_ (.A(net616),
    .B(_0674_),
    .Y(_0686_));
 sg13g2_nor2_1 _3413_ (.A(_0617_),
    .B(_0677_),
    .Y(_0687_));
 sg13g2_xnor2_1 _3414_ (.Y(_0688_),
    .A(net587),
    .B(_0684_));
 sg13g2_or4_1 _3415_ (.A(_0668_),
    .B(_0671_),
    .C(_0680_),
    .D(_0681_),
    .X(_0689_));
 sg13g2_a21oi_1 _3416_ (.A1(_0630_),
    .A2(_0683_),
    .Y(_0690_),
    .B1(_0687_));
 sg13g2_xor2_1 _3417_ (.B(_0679_),
    .A(net582),
    .X(_0691_));
 sg13g2_xnor2_1 _3418_ (.Y(_0692_),
    .A(net694),
    .B(_0670_));
 sg13g2_nand4_1 _3419_ (.B(_0690_),
    .C(_0691_),
    .A(_0685_),
    .Y(_0693_),
    .D(_0692_));
 sg13g2_nor4_1 _3420_ (.A(_0672_),
    .B(_0688_),
    .C(_0689_),
    .D(_0693_),
    .Y(_0694_));
 sg13g2_xor2_1 _3421_ (.B(_0615_),
    .A(net587),
    .X(_0695_));
 sg13g2_o21ai_1 _3422_ (.B1(_0695_),
    .Y(_0696_),
    .A1(net631),
    .A2(_0628_));
 sg13g2_nand4_1 _3423_ (.B(_0634_),
    .C(_0636_),
    .A(_0610_),
    .Y(_0697_),
    .D(_0641_));
 sg13g2_or2_1 _3424_ (.X(_0698_),
    .B(_0697_),
    .A(_0696_));
 sg13g2_nor2_1 _3425_ (.A(_1955_),
    .B(net586),
    .Y(_0699_));
 sg13g2_nor3_1 _3426_ (.A(_1956_),
    .B(net584),
    .C(_0699_),
    .Y(_0700_));
 sg13g2_a21oi_1 _3427_ (.A1(_1956_),
    .A2(net584),
    .Y(_0701_),
    .B1(_0700_));
 sg13g2_o21ai_1 _3428_ (.B1(_0621_),
    .Y(_0702_),
    .A1(_0620_),
    .A2(_0639_));
 sg13g2_nor4_1 _3429_ (.A(_0647_),
    .B(_0698_),
    .C(_0701_),
    .D(_0702_),
    .Y(_0703_));
 sg13g2_or3_1 _3430_ (.A(_0660_),
    .B(_0694_),
    .C(_0703_),
    .X(_0704_));
 sg13g2_nor2_1 _3431_ (.A(net657),
    .B(_1834_),
    .Y(_0705_));
 sg13g2_xnor2_1 _3432_ (.Y(_0706_),
    .A(net657),
    .B(_0106_));
 sg13g2_xor2_1 _3433_ (.B(_0106_),
    .A(net657),
    .X(_0707_));
 sg13g2_nand2b_2 _3434_ (.Y(_0708_),
    .B(_2050_),
    .A_N(net600));
 sg13g2_nor4_2 _3435_ (.A(net598),
    .B(net600),
    .C(net601),
    .Y(_0709_),
    .D(net603));
 sg13g2_nand2b_2 _3436_ (.Y(_0710_),
    .B(_0709_),
    .A_N(net596));
 sg13g2_or2_2 _3437_ (.X(_0711_),
    .B(_0710_),
    .A(net595));
 sg13g2_or2_1 _3438_ (.X(_0712_),
    .B(_0711_),
    .A(net594));
 sg13g2_xor2_1 _3439_ (.B(_0103_),
    .A(_0093_),
    .X(_0713_));
 sg13g2_xnor2_1 _3440_ (.Y(_0714_),
    .A(_0093_),
    .B(_0103_));
 sg13g2_nor2_1 _3441_ (.A(_0709_),
    .B(_0714_),
    .Y(_0715_));
 sg13g2_nand2b_1 _3442_ (.Y(_0716_),
    .B(_0109_),
    .A_N(_0105_));
 sg13g2_nor2b_1 _3443_ (.A(_0109_),
    .B_N(_0105_),
    .Y(_0717_));
 sg13g2_xnor2_1 _3444_ (.Y(_0718_),
    .A(_0109_),
    .B(_0105_));
 sg13g2_xor2_1 _3445_ (.B(_0105_),
    .A(_0109_),
    .X(_0719_));
 sg13g2_a221oi_1 _3446_ (.B2(_0711_),
    .C1(_0715_),
    .B1(net581),
    .A1(_0707_),
    .Y(_0720_),
    .A2(_0712_));
 sg13g2_nor2b_1 _3447_ (.A(_0104_),
    .B_N(_0094_),
    .Y(_0721_));
 sg13g2_xor2_1 _3448_ (.B(_0104_),
    .A(_0094_),
    .X(_0722_));
 sg13g2_xnor2_1 _3449_ (.Y(_0723_),
    .A(_0091_),
    .B(net599));
 sg13g2_xor2_1 _3450_ (.B(net599),
    .A(_0091_),
    .X(_0724_));
 sg13g2_xor2_1 _3451_ (.B(_0102_),
    .A(_0092_),
    .X(_0725_));
 sg13g2_nor2_1 _3452_ (.A(_0724_),
    .B(net579),
    .Y(_0726_));
 sg13g2_nor2_1 _3453_ (.A(_2050_),
    .B(_0723_),
    .Y(_0727_));
 sg13g2_a221oi_1 _3454_ (.B2(_0708_),
    .C1(_0727_),
    .B1(_0725_),
    .A1(_0710_),
    .Y(_0728_),
    .A2(net580));
 sg13g2_nor2_1 _3455_ (.A(_0708_),
    .B(net579),
    .Y(_0729_));
 sg13g2_a21oi_1 _3456_ (.A1(_2050_),
    .A2(_0723_),
    .Y(_0730_),
    .B1(_0729_));
 sg13g2_o21ai_1 _3457_ (.B1(_0713_),
    .Y(_0731_),
    .A1(net596),
    .A2(net580));
 sg13g2_nand2_1 _3458_ (.Y(_0732_),
    .A(_0709_),
    .B(_0731_));
 sg13g2_nand2_1 _3459_ (.Y(_0733_),
    .A(_0730_),
    .B(_0732_));
 sg13g2_xnor2_1 _3460_ (.Y(_0734_),
    .A(\Pong.datapath.ballFunction.ball_center_x[0] ),
    .B(net674));
 sg13g2_xnor2_1 _3461_ (.Y(_0735_),
    .A(net605),
    .B(net673));
 sg13g2_nand2_2 _3462_ (.Y(_0736_),
    .A(_0734_),
    .B(_0735_));
 sg13g2_xnor2_1 _3463_ (.Y(_0737_),
    .A(net603),
    .B(net672));
 sg13g2_nor2_1 _3464_ (.A(_0736_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_nor2_1 _3465_ (.A(_2050_),
    .B(_2151_),
    .Y(_0739_));
 sg13g2_xor2_1 _3466_ (.B(_0739_),
    .A(_0090_),
    .X(_0740_));
 sg13g2_nor4_1 _3467_ (.A(_0733_),
    .B(_0736_),
    .C(_0737_),
    .D(_0740_),
    .Y(_0741_));
 sg13g2_nor3_2 _3468_ (.A(net594),
    .B(_0707_),
    .C(_0711_),
    .Y(_0742_));
 sg13g2_a21oi_1 _3469_ (.A1(_2148_),
    .A2(net581),
    .Y(_0743_),
    .B1(_0711_));
 sg13g2_nor2_1 _3470_ (.A(_0742_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nand4_1 _3471_ (.B(_0728_),
    .C(_0741_),
    .A(_0720_),
    .Y(_0745_),
    .D(_0744_));
 sg13g2_and3_2 _3472_ (.X(_0746_),
    .A(net600),
    .B(net602),
    .C(net603));
 sg13g2_and2_1 _3473_ (.A(net598),
    .B(_0746_),
    .X(_0747_));
 sg13g2_nand3_1 _3474_ (.B(net596),
    .C(net576),
    .A(net595),
    .Y(_0748_));
 sg13g2_nor2_1 _3475_ (.A(net581),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_or2_1 _3476_ (.X(_0750_),
    .B(_0748_),
    .A(net581));
 sg13g2_nand2b_1 _3477_ (.Y(_0751_),
    .B(net576),
    .A_N(_0103_));
 sg13g2_a22oi_1 _3478_ (.Y(_0752_),
    .B1(_0751_),
    .B2(_0722_),
    .A2(_0748_),
    .A1(net581));
 sg13g2_nand4_1 _3479_ (.B(_0740_),
    .C(_0750_),
    .A(_0738_),
    .Y(_0753_),
    .D(_0752_));
 sg13g2_nand4_1 _3480_ (.B(net594),
    .C(net595),
    .A(\Pong.datapath.ballFunction.ball_center_x[9] ),
    .Y(_0754_),
    .D(net596));
 sg13g2_o21ai_1 _3481_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0103_),
    .A2(net580));
 sg13g2_o21ai_1 _3482_ (.B1(net576),
    .Y(_0756_),
    .A1(_0714_),
    .A2(_0755_));
 sg13g2_inv_1 _3483_ (.Y(_0757_),
    .A(_0756_));
 sg13g2_xor2_1 _3484_ (.B(_2151_),
    .A(net600),
    .X(_0758_));
 sg13g2_xnor2_1 _3485_ (.Y(_0759_),
    .A(_0091_),
    .B(_0758_));
 sg13g2_xnor2_1 _3486_ (.Y(_0760_),
    .A(net579),
    .B(_0746_));
 sg13g2_o21ai_1 _3487_ (.B1(_0760_),
    .Y(_0761_),
    .A1(_0714_),
    .A2(net576));
 sg13g2_nor2_1 _3488_ (.A(_0105_),
    .B(_0748_),
    .Y(_0762_));
 sg13g2_xnor2_1 _3489_ (.Y(_0763_),
    .A(_0706_),
    .B(_0762_));
 sg13g2_or4_1 _3490_ (.A(_0757_),
    .B(_0759_),
    .C(_0761_),
    .D(_0763_),
    .X(_0764_));
 sg13g2_o21ai_1 _3491_ (.B1(_0745_),
    .Y(_0765_),
    .A1(_0753_),
    .A2(_0764_));
 sg13g2_nor2_1 _3492_ (.A(_0613_),
    .B(net585),
    .Y(_0766_));
 sg13g2_nor3_1 _3493_ (.A(net612),
    .B(_0618_),
    .C(net585),
    .Y(_0767_));
 sg13g2_xnor2_1 _3494_ (.Y(_0768_),
    .A(net582),
    .B(_0767_));
 sg13g2_xor2_1 _3495_ (.B(net688),
    .A(net623),
    .X(_0769_));
 sg13g2_a21oi_1 _3496_ (.A1(net621),
    .A2(net589),
    .Y(_0770_),
    .B1(_0769_));
 sg13g2_nor2_1 _3497_ (.A(_1953_),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_nor2_1 _3498_ (.A(_0631_),
    .B(_0637_),
    .Y(_0772_));
 sg13g2_nand3_1 _3499_ (.B(_0769_),
    .C(_0772_),
    .A(net589),
    .Y(_0773_));
 sg13g2_o21ai_1 _3500_ (.B1(_0773_),
    .Y(_0774_),
    .A1(net585),
    .A2(_0771_));
 sg13g2_xnor2_1 _3501_ (.Y(_0775_),
    .A(net618),
    .B(net682));
 sg13g2_xnor2_1 _3502_ (.Y(_0776_),
    .A(_0766_),
    .B(_0775_));
 sg13g2_a21oi_2 _3503_ (.B1(net589),
    .Y(_0777_),
    .A2(_1952_),
    .A1(net621));
 sg13g2_xnor2_1 _3504_ (.Y(_0778_),
    .A(net586),
    .B(_0669_));
 sg13g2_nor3_1 _3505_ (.A(_0681_),
    .B(_0777_),
    .C(_0778_),
    .Y(_0779_));
 sg13g2_nand3_1 _3506_ (.B(_0776_),
    .C(_0779_),
    .A(_0774_),
    .Y(_0780_));
 sg13g2_nor2_1 _3507_ (.A(_1952_),
    .B(_0769_),
    .Y(_0781_));
 sg13g2_o21ai_1 _3508_ (.B1(_0631_),
    .Y(_0782_),
    .A1(_0640_),
    .A2(_0781_));
 sg13g2_nand3_1 _3509_ (.B(net587),
    .C(_0766_),
    .A(net616),
    .Y(_0783_));
 sg13g2_a21o_1 _3510_ (.A2(_0766_),
    .A1(net616),
    .B1(net587),
    .X(_0784_));
 sg13g2_o21ai_1 _3511_ (.B1(_0616_),
    .Y(_0785_),
    .A1(_0618_),
    .A2(net585));
 sg13g2_nand4_1 _3512_ (.B(_0783_),
    .C(_0784_),
    .A(_0782_),
    .Y(_0786_),
    .D(_0785_));
 sg13g2_nor3_2 _3513_ (.A(_0768_),
    .B(_0780_),
    .C(_0786_),
    .Y(_0787_));
 sg13g2_nor3_1 _3514_ (.A(net593),
    .B(_0616_),
    .C(net584),
    .Y(_0788_));
 sg13g2_nand2_1 _3515_ (.Y(_0789_),
    .A(net589),
    .B(_0788_));
 sg13g2_nand2_1 _3516_ (.Y(_0790_),
    .A(_0624_),
    .B(net582));
 sg13g2_a21oi_1 _3517_ (.A1(net582),
    .A2(_0678_),
    .Y(_0791_),
    .B1(_0683_));
 sg13g2_nor2_1 _3518_ (.A(_0623_),
    .B(_0674_),
    .Y(_0792_));
 sg13g2_nand2_1 _3519_ (.Y(_0793_),
    .A(net587),
    .B(_0792_));
 sg13g2_nand2_1 _3520_ (.Y(_0794_),
    .A(net589),
    .B(_0662_));
 sg13g2_nand4_1 _3521_ (.B(_0791_),
    .C(_0793_),
    .A(net593),
    .Y(_0795_),
    .D(_0794_));
 sg13g2_o21ai_1 _3522_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0789_),
    .A2(_0790_));
 sg13g2_a22oi_1 _3523_ (.Y(_0797_),
    .B1(net586),
    .B2(net694),
    .A2(net593),
    .A1(net625));
 sg13g2_o21ai_1 _3524_ (.B1(net586),
    .Y(_0798_),
    .A1(net625),
    .A2(net593));
 sg13g2_nor2_1 _3525_ (.A(net582),
    .B(_0678_),
    .Y(_0799_));
 sg13g2_a21oi_1 _3526_ (.A1(_0797_),
    .A2(_0798_),
    .Y(_0800_),
    .B1(_0799_));
 sg13g2_a21oi_1 _3527_ (.A1(net694),
    .A2(_0798_),
    .Y(_0801_),
    .B1(_0797_));
 sg13g2_xnor2_1 _3528_ (.Y(_0802_),
    .A(net584),
    .B(_0661_));
 sg13g2_a21oi_1 _3529_ (.A1(_0789_),
    .A2(_0802_),
    .Y(_0803_),
    .B1(_0801_));
 sg13g2_and2_1 _3530_ (.A(_0625_),
    .B(_0674_),
    .X(_0804_));
 sg13g2_o21ai_1 _3531_ (.B1(_0676_),
    .Y(_0805_),
    .A1(_0616_),
    .A2(_0804_));
 sg13g2_o21ai_1 _3532_ (.B1(_0805_),
    .Y(_0806_),
    .A1(net589),
    .A2(_0662_));
 sg13g2_o21ai_1 _3533_ (.B1(_0634_),
    .Y(_0807_),
    .A1(net587),
    .A2(_0622_));
 sg13g2_nor2_1 _3534_ (.A(_0806_),
    .B(_0807_),
    .Y(_0808_));
 sg13g2_nand4_1 _3535_ (.B(_0800_),
    .C(_0803_),
    .A(_0796_),
    .Y(_0809_),
    .D(_0808_));
 sg13g2_nor2b_1 _3536_ (.A(_0787_),
    .B_N(_0809_),
    .Y(_0810_));
 sg13g2_nand2b_1 _3537_ (.Y(_0811_),
    .B(_0809_),
    .A_N(_0787_));
 sg13g2_nor2_2 _3538_ (.A(net606),
    .B(_0710_),
    .Y(_0812_));
 sg13g2_a21oi_1 _3539_ (.A1(_0104_),
    .A2(_0812_),
    .Y(_0813_),
    .B1(_0718_));
 sg13g2_nand2b_1 _3540_ (.Y(_0814_),
    .B(_0734_),
    .A_N(_0735_));
 sg13g2_xnor2_1 _3541_ (.Y(_0815_),
    .A(net604),
    .B(_0089_));
 sg13g2_xnor2_1 _3542_ (.Y(_0816_),
    .A(net605),
    .B(_0815_));
 sg13g2_xor2_1 _3543_ (.B(_2049_),
    .A(net602),
    .X(_0817_));
 sg13g2_xnor2_1 _3544_ (.Y(_0818_),
    .A(_0090_),
    .B(_0817_));
 sg13g2_or3_1 _3545_ (.A(_0814_),
    .B(_0816_),
    .C(_0818_),
    .X(_0819_));
 sg13g2_nor2_1 _3546_ (.A(net607),
    .B(_0708_),
    .Y(_0820_));
 sg13g2_nand2_1 _3547_ (.Y(_0821_),
    .A(_0102_),
    .B(_0820_));
 sg13g2_xnor2_1 _3548_ (.Y(_0822_),
    .A(_0713_),
    .B(_0821_));
 sg13g2_nand3_1 _3549_ (.B(_0718_),
    .C(_0812_),
    .A(_0104_),
    .Y(_0823_));
 sg13g2_nor3_1 _3550_ (.A(net594),
    .B(net606),
    .C(_0711_),
    .Y(_0824_));
 sg13g2_o21ai_1 _3551_ (.B1(_0823_),
    .Y(_0825_),
    .A1(_0706_),
    .A2(_0824_));
 sg13g2_nor4_1 _3552_ (.A(_0813_),
    .B(_0819_),
    .C(_0822_),
    .D(_0825_),
    .Y(_0826_));
 sg13g2_a21oi_1 _3553_ (.A1(_2149_),
    .A2(_0709_),
    .Y(_0827_),
    .B1(_0742_));
 sg13g2_nor2_1 _3554_ (.A(net605),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_xor2_1 _3555_ (.B(_0094_),
    .A(net595),
    .X(_0829_));
 sg13g2_and2_1 _3556_ (.A(_0812_),
    .B(_0829_),
    .X(_0830_));
 sg13g2_xor2_1 _3557_ (.B(_0092_),
    .A(net598),
    .X(_0831_));
 sg13g2_nand2_1 _3558_ (.Y(_0832_),
    .A(_0100_),
    .B(_2049_));
 sg13g2_xnor2_1 _3559_ (.Y(_0833_),
    .A(_0723_),
    .B(_0832_));
 sg13g2_o21ai_1 _3560_ (.B1(_0833_),
    .Y(_0834_),
    .A1(_0820_),
    .A2(_0831_));
 sg13g2_a21oi_1 _3561_ (.A1(_0820_),
    .A2(_0831_),
    .Y(_0835_),
    .B1(_0834_));
 sg13g2_o21ai_1 _3562_ (.B1(_0835_),
    .Y(_0836_),
    .A1(_0812_),
    .A2(_0829_));
 sg13g2_nor3_1 _3563_ (.A(_0828_),
    .B(_0830_),
    .C(_0836_),
    .Y(_0837_));
 sg13g2_nand3_1 _3564_ (.B(net596),
    .C(_0713_),
    .A(net595),
    .Y(_0838_));
 sg13g2_nand4_1 _3565_ (.B(\Pong.datapath.ballFunction.ball_center_x[7] ),
    .C(net596),
    .A(net594),
    .Y(_0839_),
    .D(_0713_));
 sg13g2_xnor2_1 _3566_ (.Y(_0840_),
    .A(_0705_),
    .B(_0839_));
 sg13g2_a21oi_1 _3567_ (.A1(net605),
    .A2(_0746_),
    .Y(_0841_),
    .B1(_0831_));
 sg13g2_a221oi_1 _3568_ (.B2(_0100_),
    .C1(_0841_),
    .B1(_0724_),
    .A1(_0718_),
    .Y(_0842_),
    .A2(_0721_));
 sg13g2_a21oi_1 _3569_ (.A1(net657),
    .A2(_1834_),
    .Y(_0843_),
    .B1(_0814_));
 sg13g2_nand3_1 _3570_ (.B(_0746_),
    .C(_0831_),
    .A(net607),
    .Y(_0844_));
 sg13g2_or2_1 _3571_ (.X(_0845_),
    .B(_0721_),
    .A(_0718_));
 sg13g2_nand4_1 _3572_ (.B(_0843_),
    .C(_0844_),
    .A(_0842_),
    .Y(_0846_),
    .D(_0845_));
 sg13g2_nand3_1 _3573_ (.B(net606),
    .C(net576),
    .A(net596),
    .Y(_0847_));
 sg13g2_nand3_1 _3574_ (.B(_0714_),
    .C(_0747_),
    .A(net606),
    .Y(_0848_));
 sg13g2_o21ai_1 _3575_ (.B1(_0848_),
    .Y(_0849_),
    .A1(_0722_),
    .A2(_0847_));
 sg13g2_a21oi_1 _3576_ (.A1(net580),
    .A2(_0847_),
    .Y(_0850_),
    .B1(_0849_));
 sg13g2_nand2b_1 _3577_ (.Y(_0851_),
    .B(_0100_),
    .A_N(_0090_));
 sg13g2_xnor2_1 _3578_ (.Y(_0852_),
    .A(_0090_),
    .B(_0100_));
 sg13g2_a22oi_1 _3579_ (.Y(_0853_),
    .B1(_0723_),
    .B2(_0852_),
    .A2(net605),
    .A1(net603));
 sg13g2_nor2b_1 _3580_ (.A(_0853_),
    .B_N(_0816_),
    .Y(_0854_));
 sg13g2_a21o_1 _3581_ (.A2(net576),
    .A1(net605),
    .B1(_0714_),
    .X(_0855_));
 sg13g2_nand3b_1 _3582_ (.B(_0724_),
    .C(_0090_),
    .Y(_0856_),
    .A_N(_0100_));
 sg13g2_nand4_1 _3583_ (.B(net605),
    .C(_0851_),
    .A(net603),
    .Y(_0857_),
    .D(_0856_));
 sg13g2_nand4_1 _3584_ (.B(_0854_),
    .C(_0855_),
    .A(_0850_),
    .Y(_0858_),
    .D(_0857_));
 sg13g2_nor3_1 _3585_ (.A(_0840_),
    .B(_0846_),
    .C(_0858_),
    .Y(_0859_));
 sg13g2_a21oi_1 _3586_ (.A1(_0826_),
    .A2(_0837_),
    .Y(_0860_),
    .B1(_0859_));
 sg13g2_a21o_1 _3587_ (.A2(_0837_),
    .A1(_0826_),
    .B1(_0859_),
    .X(_0861_));
 sg13g2_a22oi_1 _3588_ (.Y(_0862_),
    .B1(_0811_),
    .B2(_0861_),
    .A2(_0765_),
    .A1(_0704_));
 sg13g2_a21oi_1 _3589_ (.A1(_0732_),
    .A2(_0744_),
    .Y(_0863_),
    .B1(net590));
 sg13g2_nand2_1 _3590_ (.Y(_0864_),
    .A(_2050_),
    .B(_2161_));
 sg13g2_nor2_1 _3591_ (.A(_2162_),
    .B(_0708_),
    .Y(_0865_));
 sg13g2_nand2_1 _3592_ (.Y(_0866_),
    .A(_2161_),
    .B(_0709_));
 sg13g2_nor2_1 _3593_ (.A(net590),
    .B(_0711_),
    .Y(_0867_));
 sg13g2_or2_1 _3594_ (.X(_0868_),
    .B(_0710_),
    .A(_2162_));
 sg13g2_nor3_2 _3595_ (.A(net594),
    .B(net595),
    .C(_0868_),
    .Y(_0869_));
 sg13g2_nor2_1 _3596_ (.A(_0706_),
    .B(_0869_),
    .Y(_0870_));
 sg13g2_xnor2_1 _3597_ (.Y(_0871_),
    .A(net579),
    .B(_0865_));
 sg13g2_and2_1 _3598_ (.A(net591),
    .B(net590),
    .X(_0872_));
 sg13g2_xnor2_1 _3599_ (.Y(_0873_),
    .A(_0098_),
    .B(_0872_));
 sg13g2_nand2b_1 _3600_ (.Y(_0874_),
    .B(_0873_),
    .A_N(_0734_));
 sg13g2_xor2_1 _3601_ (.B(_0852_),
    .A(_2163_),
    .X(_0875_));
 sg13g2_xnor2_1 _3602_ (.Y(_0876_),
    .A(_0099_),
    .B(_2161_));
 sg13g2_xnor2_1 _3603_ (.Y(_0877_),
    .A(net598),
    .B(\Pong.datapath.vga.Column_Counter.Q[5] ));
 sg13g2_xnor2_1 _3604_ (.Y(_0878_),
    .A(\Pong.datapath.ballFunction.ball_center_x[9] ),
    .B(\Pong.datapath.vga.Column_Counter.Q[9] ));
 sg13g2_xnor2_1 _3605_ (.Y(_0879_),
    .A(\Pong.datapath.ballFunction.ball_center_x[8] ),
    .B(net660));
 sg13g2_xnor2_1 _3606_ (.Y(_0880_),
    .A(net601),
    .B(net670));
 sg13g2_nand4_1 _3607_ (.B(_0878_),
    .C(_0879_),
    .A(_0877_),
    .Y(_0881_),
    .D(_0880_));
 sg13g2_xnor2_1 _3608_ (.Y(_0882_),
    .A(\Pong.datapath.ballFunction.ball_center_x[7] ),
    .B(net663));
 sg13g2_xnor2_1 _3609_ (.Y(_0883_),
    .A(net600),
    .B(net668));
 sg13g2_xnor2_1 _3610_ (.Y(_0884_),
    .A(net597),
    .B(net665));
 sg13g2_nand4_1 _3611_ (.B(_0882_),
    .C(_0883_),
    .A(_0737_),
    .Y(_0885_),
    .D(_0884_));
 sg13g2_nor3_2 _3612_ (.A(_0736_),
    .B(_0881_),
    .C(_0885_),
    .Y(_0886_));
 sg13g2_o21ai_1 _3613_ (.B1(_0724_),
    .Y(_0887_),
    .A1(net599),
    .A2(net579));
 sg13g2_a21oi_1 _3614_ (.A1(_2151_),
    .A2(_0887_),
    .Y(_0888_),
    .B1(_0757_));
 sg13g2_a21oi_1 _3615_ (.A1(_0706_),
    .A2(_0762_),
    .Y(_0889_),
    .B1(_0749_));
 sg13g2_a21oi_1 _3616_ (.A1(_0888_),
    .A2(_0889_),
    .Y(_0890_),
    .B1(net592));
 sg13g2_nand2b_2 _3617_ (.Y(_0891_),
    .B(net576),
    .A_N(net591));
 sg13g2_nor2_1 _3618_ (.A(_0103_),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_o21ai_1 _3619_ (.B1(net580),
    .Y(_0893_),
    .A1(_0103_),
    .A2(_0891_));
 sg13g2_o21ai_1 _3620_ (.B1(net581),
    .Y(_0894_),
    .A1(net591),
    .A2(_0748_));
 sg13g2_o21ai_1 _3621_ (.B1(_2152_),
    .Y(_0895_),
    .A1(_0724_),
    .A2(net579));
 sg13g2_nor2_2 _3622_ (.A(_0099_),
    .B(net591),
    .Y(_0896_));
 sg13g2_nand2_1 _3623_ (.Y(_0897_),
    .A(_0099_),
    .B(net591));
 sg13g2_nor2b_1 _3624_ (.A(_0896_),
    .B_N(_0897_),
    .Y(_0898_));
 sg13g2_nor3_2 _3625_ (.A(_0105_),
    .B(net591),
    .C(_0748_),
    .Y(_0899_));
 sg13g2_nor2_1 _3626_ (.A(_0734_),
    .B(_0873_),
    .Y(_0900_));
 sg13g2_xor2_1 _3627_ (.B(_0898_),
    .A(_0089_),
    .X(_0901_));
 sg13g2_xor2_1 _3628_ (.B(_0896_),
    .A(_0852_),
    .X(_0902_));
 sg13g2_nand4_1 _3629_ (.B(_0894_),
    .C(_0901_),
    .A(_0893_),
    .Y(_0903_),
    .D(_0902_));
 sg13g2_a22oi_1 _3630_ (.Y(_0904_),
    .B1(_0891_),
    .B2(_0713_),
    .A2(net579),
    .A1(net599));
 sg13g2_nand2_1 _3631_ (.Y(_0905_),
    .A(_0900_),
    .B(_0904_));
 sg13g2_o21ai_1 _3632_ (.B1(_0895_),
    .Y(_0906_),
    .A1(_0706_),
    .A2(_0899_));
 sg13g2_nor4_1 _3633_ (.A(_0890_),
    .B(_0903_),
    .C(_0905_),
    .D(_0906_),
    .Y(_0907_));
 sg13g2_a21oi_1 _3634_ (.A1(_0713_),
    .A2(_0866_),
    .Y(_0908_),
    .B1(_0874_));
 sg13g2_nand2_1 _3635_ (.Y(_0909_),
    .A(_0871_),
    .B(_0908_));
 sg13g2_o21ai_1 _3636_ (.B1(net581),
    .Y(_0910_),
    .A1(net590),
    .A2(_0711_));
 sg13g2_xnor2_1 _3637_ (.Y(_0911_),
    .A(_0723_),
    .B(_0864_));
 sg13g2_xnor2_1 _3638_ (.Y(_0912_),
    .A(_0089_),
    .B(_0876_));
 sg13g2_a21oi_1 _3639_ (.A1(net580),
    .A2(_0868_),
    .Y(_0913_),
    .B1(_0912_));
 sg13g2_nand4_1 _3640_ (.B(_0910_),
    .C(_0911_),
    .A(_0875_),
    .Y(_0914_),
    .D(_0913_));
 sg13g2_nor4_1 _3641_ (.A(_0863_),
    .B(_0870_),
    .C(_0909_),
    .D(_0914_),
    .Y(_0915_));
 sg13g2_nor2_1 _3642_ (.A(_0101_),
    .B(_2152_),
    .Y(_0916_));
 sg13g2_nor3_2 _3643_ (.A(_0886_),
    .B(_0907_),
    .C(_0915_),
    .Y(_0917_));
 sg13g2_o21ai_1 _3644_ (.B1(_0794_),
    .Y(_0918_),
    .A1(_0625_),
    .A2(_0674_));
 sg13g2_nor3_1 _3645_ (.A(_0629_),
    .B(_0648_),
    .C(_0652_),
    .Y(_0919_));
 sg13g2_nand2_1 _3646_ (.Y(_0920_),
    .A(_1953_),
    .B(_0661_));
 sg13g2_xnor2_1 _3647_ (.Y(_0921_),
    .A(_0082_),
    .B(_0920_));
 sg13g2_nor4_2 _3648_ (.A(_0799_),
    .B(_0802_),
    .C(_0806_),
    .Y(_0922_),
    .D(_0918_));
 sg13g2_xor2_1 _3649_ (.B(_0686_),
    .A(net587),
    .X(_0923_));
 sg13g2_and4_1 _3650_ (.A(_0791_),
    .B(_0919_),
    .C(_0921_),
    .D(_0923_),
    .X(_0924_));
 sg13g2_a21oi_1 _3651_ (.A1(net588),
    .A2(_0624_),
    .Y(_0925_),
    .B1(_0612_));
 sg13g2_nand2b_1 _3652_ (.Y(_0926_),
    .B(_0623_),
    .A_N(net588));
 sg13g2_nand3b_1 _3653_ (.B(_0926_),
    .C(_0612_),
    .Y(_0927_),
    .A_N(_0622_));
 sg13g2_xnor2_1 _3654_ (.Y(_0928_),
    .A(net612),
    .B(net678));
 sg13g2_nand2_1 _3655_ (.Y(_0929_),
    .A(net610),
    .B(net583));
 sg13g2_or2_1 _3656_ (.X(_0930_),
    .B(net588),
    .A(net617));
 sg13g2_o21ai_1 _3657_ (.B1(_0930_),
    .Y(_0931_),
    .A1(net611),
    .A2(net583));
 sg13g2_a21o_1 _3658_ (.A2(net583),
    .A1(_0618_),
    .B1(_0928_),
    .X(_0932_));
 sg13g2_or4_1 _3659_ (.A(_0777_),
    .B(_0781_),
    .C(_0921_),
    .D(_0931_),
    .X(_0933_));
 sg13g2_o21ai_1 _3660_ (.B1(_0929_),
    .Y(_0934_),
    .A1(net608),
    .A2(net612));
 sg13g2_o21ai_1 _3661_ (.B1(_0928_),
    .Y(_0935_),
    .A1(_0618_),
    .A2(_0934_));
 sg13g2_nand3_1 _3662_ (.B(_0927_),
    .C(_0935_),
    .A(_0919_),
    .Y(_0936_));
 sg13g2_nor4_1 _3663_ (.A(_0771_),
    .B(_0925_),
    .C(_0933_),
    .D(_0936_),
    .Y(_0937_));
 sg13g2_a22oi_1 _3664_ (.Y(_0938_),
    .B1(_0932_),
    .B2(_0937_),
    .A2(_0924_),
    .A1(_0922_));
 sg13g2_a21o_1 _3665_ (.A2(_0938_),
    .A1(_0810_),
    .B1(_0917_),
    .X(_0939_));
 sg13g2_nand3_1 _3666_ (.B(_0862_),
    .C(_0939_),
    .A(_0608_),
    .Y(_0940_));
 sg13g2_nor3_1 _3667_ (.A(_0707_),
    .B(_0717_),
    .C(_0748_),
    .Y(_0941_));
 sg13g2_nand2_1 _3668_ (.Y(_0942_),
    .A(_0815_),
    .B(_0888_));
 sg13g2_o21ai_1 _3669_ (.B1(net590),
    .Y(_0943_),
    .A1(_0941_),
    .A2(_0942_));
 sg13g2_nand2_1 _3670_ (.Y(_0944_),
    .A(net604),
    .B(net590));
 sg13g2_xnor2_1 _3671_ (.Y(_0945_),
    .A(_0852_),
    .B(_0944_));
 sg13g2_a21oi_1 _3672_ (.A1(_2151_),
    .A2(net590),
    .Y(_0946_),
    .B1(_0726_));
 sg13g2_a21oi_1 _3673_ (.A1(_0719_),
    .A2(_0838_),
    .Y(_0947_),
    .B1(_0946_));
 sg13g2_or3_1 _3674_ (.A(_0713_),
    .B(net580),
    .C(_0815_),
    .X(_0948_));
 sg13g2_a21oi_1 _3675_ (.A1(_2161_),
    .A2(_0948_),
    .Y(_0949_),
    .B1(_0874_));
 sg13g2_a22oi_1 _3676_ (.Y(_0950_),
    .B1(net579),
    .B2(net599),
    .A2(_0716_),
    .A1(_0707_));
 sg13g2_o21ai_1 _3677_ (.B1(_0950_),
    .Y(_0951_),
    .A1(_0714_),
    .A2(net576));
 sg13g2_a21oi_1 _3678_ (.A1(net580),
    .A2(_0751_),
    .Y(_0952_),
    .B1(_0951_));
 sg13g2_and2_1 _3679_ (.A(_0949_),
    .B(_0952_),
    .X(_0953_));
 sg13g2_nand4_1 _3680_ (.B(_0945_),
    .C(_0947_),
    .A(_0943_),
    .Y(_0954_),
    .D(_0953_));
 sg13g2_nor2_1 _3681_ (.A(net592),
    .B(net581),
    .Y(_0955_));
 sg13g2_or2_1 _3682_ (.X(_0956_),
    .B(_0955_),
    .A(_0815_));
 sg13g2_xnor2_1 _3683_ (.Y(_0957_),
    .A(_0852_),
    .B(_0897_));
 sg13g2_and4_1 _3684_ (.A(_0728_),
    .B(_0900_),
    .C(_0956_),
    .D(_0957_),
    .X(_0958_));
 sg13g2_nor2_1 _3685_ (.A(_0707_),
    .B(_0948_),
    .Y(_0959_));
 sg13g2_a21oi_1 _3686_ (.A1(_0726_),
    .A2(_0959_),
    .Y(_0960_),
    .B1(net592));
 sg13g2_a21oi_1 _3687_ (.A1(_0743_),
    .A2(_0815_),
    .Y(_0961_),
    .B1(_0960_));
 sg13g2_o21ai_1 _3688_ (.B1(net591),
    .Y(_0962_),
    .A1(_0733_),
    .A2(_0742_));
 sg13g2_nand4_1 _3689_ (.B(_0958_),
    .C(_0961_),
    .A(_0720_),
    .Y(_0963_),
    .D(_0962_));
 sg13g2_nand4_1 _3690_ (.B(_0917_),
    .C(_0954_),
    .A(_0860_),
    .Y(_0964_),
    .D(_0963_));
 sg13g2_xnor2_1 _3691_ (.Y(_0965_),
    .A(_1957_),
    .B(_0609_));
 sg13g2_xnor2_1 _3692_ (.Y(_0966_),
    .A(_1775_),
    .B(net588));
 sg13g2_and2_1 _3693_ (.A(_0626_),
    .B(_0966_),
    .X(_0967_));
 sg13g2_a21oi_1 _3694_ (.A1(net587),
    .A2(_0624_),
    .Y(_0968_),
    .B1(_0626_));
 sg13g2_xnor2_1 _3695_ (.Y(_0969_),
    .A(_1954_),
    .B(_0635_));
 sg13g2_nor2b_1 _3696_ (.A(_1905_),
    .B_N(_0663_),
    .Y(_0970_));
 sg13g2_xnor2_1 _3697_ (.Y(_0971_),
    .A(net694),
    .B(_0970_));
 sg13g2_nor2_1 _3698_ (.A(_1905_),
    .B(net586),
    .Y(_0972_));
 sg13g2_nor3_1 _3699_ (.A(_0629_),
    .B(_0653_),
    .C(_0972_),
    .Y(_0973_));
 sg13g2_nand4_1 _3700_ (.B(_0969_),
    .C(_0971_),
    .A(_0628_),
    .Y(_0974_),
    .D(_0973_));
 sg13g2_nor4_1 _3701_ (.A(_0965_),
    .B(_0967_),
    .C(_0968_),
    .D(_0974_),
    .Y(_0975_));
 sg13g2_xnor2_1 _3702_ (.Y(_0976_),
    .A(_0616_),
    .B(_0619_));
 sg13g2_o21ai_1 _3703_ (.B1(_0644_),
    .Y(_0977_),
    .A1(_1774_),
    .A2(net582));
 sg13g2_or2_1 _3704_ (.X(_0978_),
    .B(_0644_),
    .A(net582));
 sg13g2_nand4_1 _3705_ (.B(_0976_),
    .C(_0977_),
    .A(_0975_),
    .Y(_0979_),
    .D(_0978_));
 sg13g2_nor2_1 _3706_ (.A(_1902_),
    .B(_0663_),
    .Y(_0980_));
 sg13g2_nor4_2 _3707_ (.A(_1775_),
    .B(_1776_),
    .C(_1902_),
    .Y(_0981_),
    .D(_0663_));
 sg13g2_nand2b_1 _3708_ (.Y(_0982_),
    .B(_0981_),
    .A_N(_1959_));
 sg13g2_nand2b_1 _3709_ (.Y(_0983_),
    .B(_0982_),
    .A_N(net583));
 sg13g2_o21ai_1 _3710_ (.B1(_0981_),
    .Y(_0984_),
    .A1(_0097_),
    .A2(_0616_));
 sg13g2_nand2b_1 _3711_ (.Y(_0985_),
    .B(_0984_),
    .A_N(net588));
 sg13g2_nand2_1 _3712_ (.Y(_0986_),
    .A(net586),
    .B(_0663_));
 sg13g2_nor2_1 _3713_ (.A(net586),
    .B(_0663_),
    .Y(_0987_));
 sg13g2_o21ai_1 _3714_ (.B1(_0987_),
    .Y(_0988_),
    .A1(_0068_),
    .A2(net584));
 sg13g2_o21ai_1 _3715_ (.B1(_0988_),
    .Y(_0989_),
    .A1(net584),
    .A2(_0986_));
 sg13g2_nand3_1 _3716_ (.B(_0985_),
    .C(_0989_),
    .A(_0983_),
    .Y(_0990_));
 sg13g2_a21oi_1 _3717_ (.A1(net619),
    .A2(_1831_),
    .Y(_0991_),
    .B1(_0625_));
 sg13g2_a22oi_1 _3718_ (.Y(_0992_),
    .B1(_0991_),
    .B2(_0980_),
    .A2(_0981_),
    .A1(net588));
 sg13g2_a21oi_1 _3719_ (.A1(_0086_),
    .A2(_1833_),
    .Y(_0993_),
    .B1(_0617_));
 sg13g2_nor4_1 _3720_ (.A(_0629_),
    .B(_0653_),
    .C(_0971_),
    .D(_0993_),
    .Y(_0994_));
 sg13g2_nand2b_1 _3721_ (.Y(_0995_),
    .B(_0642_),
    .A_N(_0982_));
 sg13g2_o21ai_1 _3722_ (.B1(_0625_),
    .Y(_0996_),
    .A1(net619),
    .A2(_1831_));
 sg13g2_o21ai_1 _3723_ (.B1(_0996_),
    .Y(_0997_),
    .A1(net589),
    .A2(_0980_));
 sg13g2_a21oi_1 _3724_ (.A1(_0068_),
    .A2(net584),
    .Y(_0998_),
    .B1(_0997_));
 sg13g2_nand4_1 _3725_ (.B(_0994_),
    .C(_0995_),
    .A(_0992_),
    .Y(_0999_),
    .D(_0998_));
 sg13g2_o21ai_1 _3726_ (.B1(_0979_),
    .Y(_1000_),
    .A1(_0990_),
    .A2(_0999_));
 sg13g2_or2_1 _3727_ (.X(_1001_),
    .B(_1000_),
    .A(_0704_));
 sg13g2_and2_1 _3728_ (.A(_0964_),
    .B(_1001_),
    .X(_1002_));
 sg13g2_nor4_1 _3729_ (.A(_0384_),
    .B(_0385_),
    .C(_0488_),
    .D(_0549_),
    .Y(_1003_));
 sg13g2_nand2_1 _3730_ (.Y(_1004_),
    .A(net669),
    .B(_0384_));
 sg13g2_nand2_1 _3731_ (.Y(_1005_),
    .A(_0592_),
    .B(_1004_));
 sg13g2_nor2_1 _3732_ (.A(_0388_),
    .B(_0499_),
    .Y(_1006_));
 sg13g2_a21oi_1 _3733_ (.A1(_1005_),
    .A2(_1006_),
    .Y(_1007_),
    .B1(_1003_));
 sg13g2_nand2_1 _3734_ (.Y(_1008_),
    .A(_1823_),
    .B(\Pong.datapath.scoreRight[1] ));
 sg13g2_nand2b_1 _3735_ (.Y(_1009_),
    .B(\Pong.datapath.scoreRight[2] ),
    .A_N(\Pong.datapath.scoreRight[1] ));
 sg13g2_a21oi_1 _3736_ (.A1(_0568_),
    .A2(_1008_),
    .Y(_1010_),
    .B1(\Pong.datapath.scoreRight[0] ));
 sg13g2_a21oi_1 _3737_ (.A1(_0565_),
    .A2(_1009_),
    .Y(_1011_),
    .B1(_0569_));
 sg13g2_a22oi_1 _3738_ (.Y(_1012_),
    .B1(_1011_),
    .B2(_0539_),
    .A2(_1010_),
    .A1(_0521_));
 sg13g2_nor3_1 _3739_ (.A(_0488_),
    .B(_0549_),
    .C(_1012_),
    .Y(_1013_));
 sg13g2_nand2_1 _3740_ (.Y(_1014_),
    .A(net689),
    .B(_0526_));
 sg13g2_nor2_1 _3741_ (.A(_0506_),
    .B(_0514_),
    .Y(_1015_));
 sg13g2_o21ai_1 _3742_ (.B1(_0536_),
    .Y(_1016_),
    .A1(_1014_),
    .A2(_1015_));
 sg13g2_nand4_1 _3743_ (.B(_0504_),
    .C(_0526_),
    .A(_1790_),
    .Y(_1017_),
    .D(_1015_));
 sg13g2_a21oi_1 _3744_ (.A1(_1016_),
    .A2(_1017_),
    .Y(_1018_),
    .B1(_0535_));
 sg13g2_nand4_1 _3745_ (.B(net697),
    .C(_1795_),
    .A(net689),
    .Y(_1019_),
    .D(_0519_));
 sg13g2_nand3_1 _3746_ (.B(_0507_),
    .C(_0530_),
    .A(net689),
    .Y(_1020_));
 sg13g2_a21oi_1 _3747_ (.A1(_0511_),
    .A2(_1020_),
    .Y(_1021_),
    .B1(net676));
 sg13g2_a22oi_1 _3748_ (.Y(_1022_),
    .B1(_1019_),
    .B2(_1021_),
    .A2(_0516_),
    .A1(_0513_));
 sg13g2_or2_1 _3749_ (.X(_1023_),
    .B(_1022_),
    .A(_1018_));
 sg13g2_nor3_1 _3750_ (.A(_0566_),
    .B(_0567_),
    .C(_0571_),
    .Y(_1024_));
 sg13g2_o21ai_1 _3751_ (.B1(_1023_),
    .Y(_1025_),
    .A1(_1010_),
    .A2(_1024_));
 sg13g2_nand2_1 _3752_ (.Y(_1026_),
    .A(_0574_),
    .B(_1018_));
 sg13g2_nand2_1 _3753_ (.Y(_1027_),
    .A(_0518_),
    .B(_0519_));
 sg13g2_xnor2_1 _3754_ (.Y(_1028_),
    .A(\Pong.datapath.scoreRight[3] ),
    .B(_0567_));
 sg13g2_nand4_1 _3755_ (.B(_0519_),
    .C(_0572_),
    .A(_0518_),
    .Y(_1029_),
    .D(_1028_));
 sg13g2_nand3_1 _3756_ (.B(_1026_),
    .C(_1029_),
    .A(_1025_),
    .Y(_1030_));
 sg13g2_a22oi_1 _3757_ (.Y(_1031_),
    .B1(_1030_),
    .B2(_0582_),
    .A2(_1013_),
    .A1(_0392_));
 sg13g2_nand2b_1 _3758_ (.Y(_1032_),
    .B(_1004_),
    .A_N(net658));
 sg13g2_o21ai_1 _3759_ (.B1(_0553_),
    .Y(_1033_),
    .A1(_0588_),
    .A2(_1032_));
 sg13g2_nand2_1 _3760_ (.Y(_1034_),
    .A(_0540_),
    .B(_0541_));
 sg13g2_nand3_1 _3761_ (.B(\Pong.datapath.scoreLeft[0] ),
    .C(_0522_),
    .A(\Pong.datapath.scoreLeft[3] ),
    .Y(_1035_));
 sg13g2_and2_1 _3762_ (.A(\Pong.datapath.scoreLeft[2] ),
    .B(\Pong.datapath.scoreLeft[1] ),
    .X(_1036_));
 sg13g2_nand3_1 _3763_ (.B(\Pong.datapath.scoreLeft[0] ),
    .C(_1036_),
    .A(_1824_),
    .Y(_1037_));
 sg13g2_nand2_1 _3764_ (.Y(_1038_),
    .A(_1035_),
    .B(_1037_));
 sg13g2_a21oi_2 _3765_ (.B1(_0523_),
    .Y(_1039_),
    .A2(\Pong.datapath.scoreLeft[0] ),
    .A1(\Pong.datapath.scoreLeft[3] ));
 sg13g2_o21ai_1 _3766_ (.B1(\Pong.datapath.scoreLeft[2] ),
    .Y(_1040_),
    .A1(\Pong.datapath.scoreLeft[0] ),
    .A2(\Pong.datapath.scoreLeft[1] ));
 sg13g2_a21o_1 _3767_ (.A2(_1040_),
    .A1(_1039_),
    .B1(_1038_),
    .X(_1041_));
 sg13g2_a22oi_1 _3768_ (.Y(_1042_),
    .B1(_1041_),
    .B2(_0539_),
    .A2(_1034_),
    .A1(_0521_));
 sg13g2_nand3_1 _3769_ (.B(_0496_),
    .C(_0548_),
    .A(net657),
    .Y(_1043_));
 sg13g2_nand3_1 _3770_ (.B(net671),
    .C(net673),
    .A(net661),
    .Y(_1044_));
 sg13g2_nand3b_1 _3771_ (.B(_0560_),
    .C(net671),
    .Y(_1045_),
    .A_N(net673));
 sg13g2_o21ai_1 _3772_ (.B1(_1044_),
    .Y(_1046_),
    .A1(_0559_),
    .A2(_1045_));
 sg13g2_a22oi_1 _3773_ (.Y(_1047_),
    .B1(_1046_),
    .B2(net667),
    .A2(_1043_),
    .A1(_0557_));
 sg13g2_nor2_1 _3774_ (.A(_1042_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_nor3_1 _3775_ (.A(_0522_),
    .B(_0541_),
    .C(_1036_),
    .Y(_1049_));
 sg13g2_o21ai_1 _3776_ (.B1(_1023_),
    .Y(_1050_),
    .A1(_0525_),
    .A2(_1049_));
 sg13g2_nor3_1 _3777_ (.A(\Pong.datapath.scoreLeft[2] ),
    .B(\Pong.datapath.scoreLeft[3] ),
    .C(\Pong.datapath.scoreLeft[1] ),
    .Y(_1051_));
 sg13g2_nor3_1 _3778_ (.A(_0523_),
    .B(_1027_),
    .C(_1051_),
    .Y(_1052_));
 sg13g2_a22oi_1 _3779_ (.Y(_1053_),
    .B1(_1052_),
    .B2(_1037_),
    .A2(_1038_),
    .A1(_1018_));
 sg13g2_a21oi_1 _3780_ (.A1(_1050_),
    .A2(_1053_),
    .Y(_1054_),
    .B1(_0556_));
 sg13g2_o21ai_1 _3781_ (.B1(_1033_),
    .Y(_1055_),
    .A1(_1048_),
    .A2(_1054_));
 sg13g2_o21ai_1 _3782_ (.B1(_1055_),
    .Y(_1056_),
    .A1(_1007_),
    .A2(_1031_));
 sg13g2_nor4_1 _3783_ (.A(_0503_),
    .B(_0940_),
    .C(_1002_),
    .D(_1056_),
    .Y(_1057_));
 sg13g2_nand2_1 _3784_ (.Y(_1058_),
    .A(net686),
    .B(_0509_));
 sg13g2_nand2_1 _3785_ (.Y(_1059_),
    .A(net658),
    .B(net660));
 sg13g2_o21ai_1 _3786_ (.B1(net658),
    .Y(_1060_),
    .A1(net660),
    .A2(net662));
 sg13g2_nand3_1 _3787_ (.B(net695),
    .C(_0596_),
    .A(net691),
    .Y(_1061_));
 sg13g2_o21ai_1 _3788_ (.B1(_0512_),
    .Y(_1062_),
    .A1(_0510_),
    .A2(_1061_));
 sg13g2_o21ai_1 _3789_ (.B1(_0595_),
    .Y(_1063_),
    .A1(_0605_),
    .A2(_1062_));
 sg13g2_nand4_1 _3790_ (.B(_1058_),
    .C(_1060_),
    .A(_1788_),
    .Y(_1064_),
    .D(_1063_));
 sg13g2_a21oi_2 _3791_ (.B1(_1064_),
    .Y(\Pong.b ),
    .A2(_1057_),
    .A1(_0394_));
 sg13g2_nand4_1 _3792_ (.B(net692),
    .C(_0509_),
    .A(net686),
    .Y(_1065_),
    .D(_0596_));
 sg13g2_a21oi_1 _3793_ (.A1(net691),
    .A2(net695),
    .Y(_1066_),
    .B1(net690));
 sg13g2_a21oi_1 _3794_ (.A1(_0531_),
    .A2(_1066_),
    .Y(_1067_),
    .B1(_1058_));
 sg13g2_a21oi_1 _3795_ (.A1(net675),
    .A2(_1065_),
    .Y(_1068_),
    .B1(_1067_));
 sg13g2_nand2_1 _3796_ (.Y(\Pong.datapath.v_sync ),
    .A(_1788_),
    .B(_1068_));
 sg13g2_nand2_1 _3797_ (.Y(_1069_),
    .A(net673),
    .B(net674));
 sg13g2_nand3_1 _3798_ (.B(net674),
    .C(_0391_),
    .A(net673),
    .Y(_1070_));
 sg13g2_nand2_1 _3799_ (.Y(_1071_),
    .A(_0551_),
    .B(_1070_));
 sg13g2_nand2_1 _3800_ (.Y(_1072_),
    .A(net662),
    .B(_1071_));
 sg13g2_or2_1 _3801_ (.X(_1073_),
    .B(_0385_),
    .A(net661));
 sg13g2_o21ai_1 _3802_ (.B1(_0390_),
    .Y(_1074_),
    .A1(_1070_),
    .A2(_1073_));
 sg13g2_nand4_1 _3803_ (.B(net662),
    .C(net664),
    .A(net658),
    .Y(_1075_),
    .D(_1074_));
 sg13g2_nand2_1 _3804_ (.Y(_1076_),
    .A(\Pong.datapath.vga.Column_Counter.Q[9] ),
    .B(_0551_));
 sg13g2_a22oi_1 _3805_ (.Y(_1077_),
    .B1(_1076_),
    .B2(net657),
    .A2(_1072_),
    .A1(_0498_));
 sg13g2_nand3_1 _3806_ (.B(_1075_),
    .C(_1077_),
    .A(_1059_),
    .Y(\Pong.datapath.h_sync ));
 sg13g2_a221oi_1 _3807_ (.B2(_1807_),
    .C1(\Pong.datapath.score_flag ),
    .B1(net721),
    .A1(net656),
    .Y(_1078_),
    .A2(net471));
 sg13g2_and2_1 _3808_ (.A(_0573_),
    .B(_1035_),
    .X(_1079_));
 sg13g2_nand2_2 _3809_ (.Y(_1080_),
    .A(net601),
    .B(_2163_));
 sg13g2_nand2_1 _3810_ (.Y(_1081_),
    .A(_2053_),
    .B(_2149_));
 sg13g2_or2_1 _3811_ (.X(_1082_),
    .B(_2153_),
    .A(_2052_));
 sg13g2_a21oi_2 _3812_ (.B1(_1080_),
    .Y(_1083_),
    .A2(_1082_),
    .A1(_1081_));
 sg13g2_nand3b_1 _3813_ (.B(_1083_),
    .C(\Pong.datapath.score_flag ),
    .Y(_1084_),
    .A_N(_1079_));
 sg13g2_nor3_2 _3814_ (.A(_2052_),
    .B(_2153_),
    .C(_1080_),
    .Y(_1085_));
 sg13g2_and2_1 _3815_ (.A(\Pong.datapath.score_flag ),
    .B(_1085_),
    .X(_1086_));
 sg13g2_nand2_1 _3816_ (.Y(_1087_),
    .A(\Pong.datapath.score_flag ),
    .B(_1085_));
 sg13g2_and4_2 _3817_ (.A(net601),
    .B(_2053_),
    .C(_2149_),
    .D(_2163_),
    .X(_1088_));
 sg13g2_nor2_1 _3818_ (.A(_1085_),
    .B(_1088_),
    .Y(_1089_));
 sg13g2_nor2_1 _3819_ (.A(_1079_),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_or2_1 _3820_ (.X(_1091_),
    .B(_1089_),
    .A(_1079_));
 sg13g2_and3_1 _3821_ (.X(_1092_),
    .A(\Pong.datapath.score_flag ),
    .B(_0575_),
    .C(_1088_));
 sg13g2_a221oi_1 _3822_ (.B2(\Pong.datapath.score_flag ),
    .C1(_1092_),
    .B1(_1090_),
    .A1(_1039_),
    .Y(_1093_),
    .A2(_1086_));
 sg13g2_inv_1 _3823_ (.Y(_1094_),
    .A(_1093_));
 sg13g2_nor3_2 _3824_ (.A(_2052_),
    .B(_2153_),
    .C(_1080_),
    .Y(_1095_));
 sg13g2_nand3_1 _3825_ (.B(_1039_),
    .C(_1095_),
    .A(\Pong.datapath.score_flag ),
    .Y(_1096_));
 sg13g2_o21ai_1 _3826_ (.B1(net749),
    .Y(_0131_),
    .A1(net527),
    .A2(_1094_));
 sg13g2_nor3_1 _3827_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[8] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[13] ),
    .C(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ),
    .Y(_1097_));
 sg13g2_nor2_1 _3828_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[7] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[12] ),
    .Y(_1098_));
 sg13g2_nand2_1 _3829_ (.Y(_1099_),
    .A(_0128_),
    .B(_0127_));
 sg13g2_o21ai_1 _3830_ (.B1(_0126_),
    .Y(_1100_),
    .A1(_2183_),
    .A2(_1099_));
 sg13g2_nand3_1 _3831_ (.B(_1098_),
    .C(_1100_),
    .A(_0125_),
    .Y(_1101_));
 sg13g2_nand2_1 _3832_ (.Y(_1102_),
    .A(_0124_),
    .B(_1101_));
 sg13g2_a21oi_1 _3833_ (.A1(_1097_),
    .A2(_1102_),
    .Y(_1103_),
    .B1(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ));
 sg13g2_nor2_1 _3834_ (.A(_2181_),
    .B(_1103_),
    .Y(_1104_));
 sg13g2_nor2_1 _3835_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[4] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[16] ),
    .Y(_1105_));
 sg13g2_a21oi_1 _3836_ (.A1(_0128_),
    .A2(_2183_),
    .Y(_1106_),
    .B1(\Pong.control_unit.NES_Controller_Right.state_NESController[4] ));
 sg13g2_nand4_1 _3837_ (.B(_2184_),
    .C(_1098_),
    .A(_0125_),
    .Y(_1107_),
    .D(_1105_));
 sg13g2_a21oi_1 _3838_ (.A1(_0124_),
    .A2(_1107_),
    .Y(_1108_),
    .B1(\Pong.control_unit.NES_Controller_Right.state_NESController[8] ));
 sg13g2_nor2_1 _3839_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ),
    .B(_2182_),
    .Y(_1109_));
 sg13g2_o21ai_1 _3840_ (.B1(_1109_),
    .Y(_1110_),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[13] ),
    .A2(_1108_));
 sg13g2_nand2b_2 _3841_ (.Y(_1111_),
    .B(_1110_),
    .A_N(_1104_));
 sg13g2_nor2_1 _3842_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[2] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ),
    .Y(_1112_));
 sg13g2_nand2_1 _3843_ (.Y(_1113_),
    .A(_1097_),
    .B(_1112_));
 sg13g2_nor2_1 _3844_ (.A(_2182_),
    .B(_1113_),
    .Y(_1114_));
 sg13g2_o21ai_1 _3845_ (.B1(_0130_),
    .Y(_1115_),
    .A1(\Pong.control_unit.NES_Controller_Right.state_NESController[16] ),
    .A2(_1106_));
 sg13g2_nand2_1 _3846_ (.Y(_1116_),
    .A(_0129_),
    .B(_1115_));
 sg13g2_and2_1 _3847_ (.A(_1114_),
    .B(_1116_),
    .X(_1117_));
 sg13g2_inv_1 _3848_ (.Y(_1118_),
    .A(_1117_));
 sg13g2_nor3_1 _3849_ (.A(_1804_),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[14] ),
    .C(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ),
    .Y(_1119_));
 sg13g2_nor2b_1 _3850_ (.A(_2185_),
    .B_N(_1098_),
    .Y(_1120_));
 sg13g2_nand4_1 _3851_ (.B(_1114_),
    .C(_1119_),
    .A(_1105_),
    .Y(_1121_),
    .D(_1120_));
 sg13g2_inv_1 _3852_ (.Y(_1122_),
    .A(_1121_));
 sg13g2_nand3_1 _3853_ (.B(_1118_),
    .C(_1121_),
    .A(_1111_),
    .Y(_1123_));
 sg13g2_nand2_1 _3854_ (.Y(_1124_),
    .A(_1118_),
    .B(_1122_));
 sg13g2_nor2_1 _3855_ (.A(_1111_),
    .B(_1124_),
    .Y(_1125_));
 sg13g2_o21ai_1 _3856_ (.B1(_1123_),
    .Y(_1126_),
    .A1(_1111_),
    .A2(_1124_));
 sg13g2_or2_1 _3857_ (.X(_1127_),
    .B(_1110_),
    .A(_1104_));
 sg13g2_nor2_1 _3858_ (.A(_1118_),
    .B(_1122_),
    .Y(_1128_));
 sg13g2_nand2_1 _3859_ (.Y(_1129_),
    .A(_1117_),
    .B(_1121_));
 sg13g2_a21oi_1 _3860_ (.A1(_1127_),
    .A2(_1128_),
    .Y(_1130_),
    .B1(_1126_));
 sg13g2_nor3_1 _3861_ (.A(net3),
    .B(_1127_),
    .C(_1129_),
    .Y(_1131_));
 sg13g2_o21ai_1 _3862_ (.B1(net747),
    .Y(_1132_),
    .A1(net387),
    .A2(_1130_));
 sg13g2_nor2_1 _3863_ (.A(_1131_),
    .B(_1132_),
    .Y(_0132_));
 sg13g2_nor3_2 _3864_ (.A(net322),
    .B(net339),
    .C(_2169_),
    .Y(_1133_));
 sg13g2_nor2_1 _3865_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[13] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ),
    .Y(_1134_));
 sg13g2_nor3_1 _3866_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[13] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[8] ),
    .C(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ),
    .Y(_1135_));
 sg13g2_a21oi_1 _3867_ (.A1(_0121_),
    .A2(_2170_),
    .Y(_1136_),
    .B1(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ));
 sg13g2_o21ai_1 _3868_ (.B1(_0123_),
    .Y(_1137_),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ),
    .A2(_1136_));
 sg13g2_nand2_1 _3869_ (.Y(_1138_),
    .A(_0122_),
    .B(_1137_));
 sg13g2_and2_1 _3870_ (.A(_1135_),
    .B(_1138_),
    .X(_1139_));
 sg13g2_nor4_1 _3871_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[8] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ),
    .C(\Pong.control_unit.NES_Controller_Left.state_NESController[14] ),
    .D(\Pong.control_unit.NES_Controller_Left.state_NESController[18] ),
    .Y(_1140_));
 sg13g2_nor2_1 _3872_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ),
    .Y(_1141_));
 sg13g2_nor3_1 _3873_ (.A(_1797_),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ),
    .C(_2172_),
    .Y(_1142_));
 sg13g2_and4_1 _3874_ (.A(_1134_),
    .B(_1140_),
    .C(_1141_),
    .D(_1142_),
    .X(_1143_));
 sg13g2_nand3b_1 _3875_ (.B(_1139_),
    .C(_1133_),
    .Y(_1144_),
    .A_N(_1143_));
 sg13g2_nand2_1 _3876_ (.Y(_1145_),
    .A(_0121_),
    .B(_0120_));
 sg13g2_o21ai_1 _3877_ (.B1(_0119_),
    .Y(_1146_),
    .A1(_2170_),
    .A2(_1145_));
 sg13g2_nor2b_1 _3878_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ),
    .B_N(_0118_),
    .Y(_1147_));
 sg13g2_nand3b_1 _3879_ (.B(_1146_),
    .C(_1147_),
    .Y(_1148_),
    .A_N(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ));
 sg13g2_nand2_1 _3880_ (.Y(_1149_),
    .A(_0117_),
    .B(_1148_));
 sg13g2_a21oi_1 _3881_ (.A1(_1135_),
    .A2(_1149_),
    .Y(_1150_),
    .B1(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ));
 sg13g2_nor2_1 _3882_ (.A(_2168_),
    .B(_1150_),
    .Y(_1151_));
 sg13g2_inv_1 _3883_ (.Y(_1152_),
    .A(_1151_));
 sg13g2_nand3_1 _3884_ (.B(_1141_),
    .C(_1147_),
    .A(_1136_),
    .Y(_1153_));
 sg13g2_a21oi_1 _3885_ (.A1(_0117_),
    .A2(_1153_),
    .Y(_1154_),
    .B1(\Pong.control_unit.NES_Controller_Left.state_NESController[8] ));
 sg13g2_nor2_1 _3886_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ),
    .B(_2169_),
    .Y(_1155_));
 sg13g2_o21ai_1 _3887_ (.B1(_1155_),
    .Y(_1156_),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[13] ),
    .A2(_1154_));
 sg13g2_nand3b_1 _3888_ (.B(_1143_),
    .C(_1133_),
    .Y(_1157_),
    .A_N(_1139_));
 sg13g2_and3_1 _3889_ (.X(_1158_),
    .A(_1152_),
    .B(_1156_),
    .C(_1157_));
 sg13g2_o21ai_1 _3890_ (.B1(_1133_),
    .Y(_1159_),
    .A1(_1139_),
    .A2(_1143_));
 sg13g2_a21oi_1 _3891_ (.A1(_1152_),
    .A2(_1156_),
    .Y(_1160_),
    .B1(_1159_));
 sg13g2_o21ai_1 _3892_ (.B1(_1144_),
    .Y(_1161_),
    .A1(_1158_),
    .A2(_1160_));
 sg13g2_nor2_1 _3893_ (.A(_1152_),
    .B(_1156_),
    .Y(_1162_));
 sg13g2_a21oi_1 _3894_ (.A1(_1144_),
    .A2(_1162_),
    .Y(_1163_),
    .B1(net398));
 sg13g2_nor3_1 _3895_ (.A(net2),
    .B(_1152_),
    .C(_1156_),
    .Y(_1164_));
 sg13g2_a221oi_1 _3896_ (.B2(_1159_),
    .C1(net742),
    .B1(_1164_),
    .A1(_1161_),
    .Y(_0133_),
    .A2(_1163_));
 sg13g2_mux2_1 _3897_ (.A0(net497),
    .A1(net2),
    .S(_1158_),
    .X(_1165_));
 sg13g2_nor2b_1 _3898_ (.A(_1165_),
    .B_N(_1161_),
    .Y(_1166_));
 sg13g2_nor2_1 _3899_ (.A(net742),
    .B(_1166_),
    .Y(_0134_));
 sg13g2_nand3b_1 _3900_ (.B(_1151_),
    .C(_1156_),
    .Y(_1167_),
    .A_N(_1159_));
 sg13g2_mux2_1 _3901_ (.A0(net2),
    .A1(net501),
    .S(_1167_),
    .X(_1168_));
 sg13g2_nor2b_1 _3902_ (.A(_1168_),
    .B_N(_1161_),
    .Y(_1169_));
 sg13g2_nor2_1 _3903_ (.A(net742),
    .B(_1169_),
    .Y(_0135_));
 sg13g2_nor3_1 _3904_ (.A(_1151_),
    .B(_1156_),
    .C(_1159_),
    .Y(_1170_));
 sg13g2_mux2_1 _3905_ (.A0(net500),
    .A1(net2),
    .S(_1170_),
    .X(_1171_));
 sg13g2_nor2b_1 _3906_ (.A(_1171_),
    .B_N(_1161_),
    .Y(_1172_));
 sg13g2_nor2_1 _3907_ (.A(net742),
    .B(_1172_),
    .Y(_0136_));
 sg13g2_nand2_1 _3908_ (.Y(_1173_),
    .A(_1104_),
    .B(_1110_));
 sg13g2_a21oi_1 _3909_ (.A1(_1128_),
    .A2(_1173_),
    .Y(_1174_),
    .B1(_1126_));
 sg13g2_nor3_1 _3910_ (.A(net3),
    .B(_1129_),
    .C(_1173_),
    .Y(_1175_));
 sg13g2_o21ai_1 _3911_ (.B1(net747),
    .Y(_1176_),
    .A1(net400),
    .A2(_1174_));
 sg13g2_nor2_1 _3912_ (.A(_1175_),
    .B(_1176_),
    .Y(_0137_));
 sg13g2_a21oi_1 _3913_ (.A1(_1111_),
    .A2(_1128_),
    .Y(_1177_),
    .B1(_1126_));
 sg13g2_nor3_1 _3914_ (.A(net3),
    .B(_1111_),
    .C(_1129_),
    .Y(_1178_));
 sg13g2_o21ai_1 _3915_ (.B1(net747),
    .Y(_1179_),
    .A1(net389),
    .A2(_1177_));
 sg13g2_nor2_1 _3916_ (.A(_1178_),
    .B(_1179_),
    .Y(_0138_));
 sg13g2_or3_1 _3917_ (.A(_2181_),
    .B(_1103_),
    .C(_1110_),
    .X(_1180_));
 sg13g2_nor2b_1 _3918_ (.A(_1123_),
    .B_N(_1180_),
    .Y(_1181_));
 sg13g2_nor3_1 _3919_ (.A(_1125_),
    .B(_1128_),
    .C(_1181_),
    .Y(_1182_));
 sg13g2_nor4_1 _3920_ (.A(net3),
    .B(_1117_),
    .C(_1122_),
    .D(_1180_),
    .Y(_1183_));
 sg13g2_o21ai_1 _3921_ (.B1(net747),
    .Y(_1184_),
    .A1(net415),
    .A2(_1182_));
 sg13g2_nor2_1 _3922_ (.A(_1183_),
    .B(_1184_),
    .Y(_0139_));
 sg13g2_nand2_1 _3923_ (.Y(_1185_),
    .A(net749),
    .B(_1084_));
 sg13g2_nor2b_1 _3924_ (.A(\Pong.datapath.NES_activity_Left[5] ),
    .B_N(net455),
    .Y(_1186_));
 sg13g2_nand2_1 _3925_ (.Y(_1187_),
    .A(net656),
    .B(net455));
 sg13g2_nand2b_1 _3926_ (.Y(_1188_),
    .B(_1187_),
    .A_N(_1092_));
 sg13g2_a21oi_1 _3927_ (.A1(net487),
    .A2(_1186_),
    .Y(_1189_),
    .B1(_1092_));
 sg13g2_and2_1 _3928_ (.A(\Pong.datapath.scoreRight[0] ),
    .B(_1092_),
    .X(_1190_));
 sg13g2_nor3_1 _3929_ (.A(_1185_),
    .B(_1189_),
    .C(_1190_),
    .Y(_0140_));
 sg13g2_a21oi_1 _3930_ (.A1(net481),
    .A2(_1188_),
    .Y(_1191_),
    .B1(_1190_));
 sg13g2_and2_1 _3931_ (.A(net481),
    .B(_1190_),
    .X(_1192_));
 sg13g2_nor3_1 _3932_ (.A(_1185_),
    .B(_1191_),
    .C(_1192_),
    .Y(_0141_));
 sg13g2_a22oi_1 _3933_ (.Y(_1193_),
    .B1(_1190_),
    .B2(_0571_),
    .A2(_1090_),
    .A1(\Pong.datapath.score_flag ));
 sg13g2_nand2_1 _3934_ (.Y(_1194_),
    .A(_1188_),
    .B(_1193_));
 sg13g2_nor2_1 _3935_ (.A(net469),
    .B(_1192_),
    .Y(_1195_));
 sg13g2_nor3_1 _3936_ (.A(net742),
    .B(_1194_),
    .C(net470),
    .Y(_0142_));
 sg13g2_nand3_1 _3937_ (.B(_1091_),
    .C(_1190_),
    .A(_0571_),
    .Y(_1196_));
 sg13g2_a21o_1 _3938_ (.A2(_1196_),
    .A1(_1823_),
    .B1(net742),
    .X(_1197_));
 sg13g2_a21oi_1 _3939_ (.A1(net426),
    .A2(_1194_),
    .Y(_0143_),
    .B1(_1197_));
 sg13g2_nand2_1 _3940_ (.Y(_1198_),
    .A(_1096_),
    .B(_1187_));
 sg13g2_nand2b_1 _3941_ (.Y(_1199_),
    .B(_1198_),
    .A_N(_1185_));
 sg13g2_and2_1 _3942_ (.A(_1825_),
    .B(_1096_),
    .X(_1200_));
 sg13g2_nor2_1 _3943_ (.A(_1825_),
    .B(_1096_),
    .Y(_1201_));
 sg13g2_nor2_1 _3944_ (.A(_0541_),
    .B(_1087_),
    .Y(_1202_));
 sg13g2_nor3_1 _3945_ (.A(_1199_),
    .B(_1200_),
    .C(_1201_),
    .Y(_0144_));
 sg13g2_xnor2_1 _3946_ (.Y(_1203_),
    .A(net485),
    .B(_1201_));
 sg13g2_nor2_1 _3947_ (.A(_1199_),
    .B(net486),
    .Y(_0145_));
 sg13g2_a21oi_1 _3948_ (.A1(\Pong.datapath.scoreLeft[1] ),
    .A2(_1202_),
    .Y(_1204_),
    .B1(net421));
 sg13g2_nor2_1 _3949_ (.A(_1037_),
    .B(_1087_),
    .Y(_1205_));
 sg13g2_nor3_1 _3950_ (.A(_1199_),
    .B(net422),
    .C(_1205_),
    .Y(_0146_));
 sg13g2_a21oi_1 _3951_ (.A1(_1084_),
    .A2(_1198_),
    .Y(_1206_),
    .B1(_1824_));
 sg13g2_a21oi_1 _3952_ (.A1(_1091_),
    .A2(_1205_),
    .Y(_1207_),
    .B1(net373));
 sg13g2_nor3_1 _3953_ (.A(net742),
    .B(_1206_),
    .C(_1207_),
    .Y(_0147_));
 sg13g2_nand2_2 _3954_ (.Y(_1208_),
    .A(net749),
    .B(_1093_));
 sg13g2_nand3_1 _3955_ (.B(net455),
    .C(_1093_),
    .A(net749),
    .Y(_1209_));
 sg13g2_o21ai_1 _3956_ (.B1(net656),
    .Y(_1210_),
    .A1(net471),
    .A2(\Pong.datapath.ballFunction.reset_n ));
 sg13g2_a21oi_1 _3957_ (.A1(_1822_),
    .A2(net472),
    .Y(_0148_),
    .B1(_1209_));
 sg13g2_a21oi_2 _3958_ (.B1(\Pong.datapath.rightPaddle[2] ),
    .Y(_1211_),
    .A2(net731),
    .A1(net729));
 sg13g2_nor2_1 _3959_ (.A(_1812_),
    .B(_1211_),
    .Y(_1212_));
 sg13g2_nor3_2 _3960_ (.A(_1812_),
    .B(_1813_),
    .C(_1211_),
    .Y(_1213_));
 sg13g2_nand2_1 _3961_ (.Y(_1214_),
    .A(\Pong.datapath.rightPaddle[5] ),
    .B(_1213_));
 sg13g2_nor2_1 _3962_ (.A(_2041_),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_nand4_1 _3963_ (.B(\Pong.datapath.rightPaddle[6] ),
    .C(\Pong.datapath.rightPaddle[5] ),
    .A(net724),
    .Y(_1216_),
    .D(_1213_));
 sg13g2_nor2_1 _3964_ (.A(_0058_),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_xnor2_1 _3965_ (.Y(_1218_),
    .A(_0056_),
    .B(_1217_));
 sg13g2_nor2_2 _3966_ (.A(_1215_),
    .B(_1218_),
    .Y(_1219_));
 sg13g2_nor2_1 _3967_ (.A(_0060_),
    .B(_1214_),
    .Y(_1220_));
 sg13g2_xnor2_1 _3968_ (.Y(_1221_),
    .A(_1814_),
    .B(_1220_));
 sg13g2_xor2_1 _3969_ (.B(_1216_),
    .A(_0058_),
    .X(_1222_));
 sg13g2_xnor2_1 _3970_ (.Y(_1223_),
    .A(_1810_),
    .B(_1214_));
 sg13g2_xor2_1 _3971_ (.B(_1212_),
    .A(_0065_),
    .X(_1224_));
 sg13g2_xor2_1 _3972_ (.B(_1213_),
    .A(_0061_),
    .X(_1225_));
 sg13g2_or2_1 _3973_ (.X(_1226_),
    .B(_1211_),
    .A(_0396_));
 sg13g2_xnor2_1 _3974_ (.Y(_1227_),
    .A(_1812_),
    .B(_0419_));
 sg13g2_nand2_1 _3975_ (.Y(_1228_),
    .A(_1226_),
    .B(_1227_));
 sg13g2_nand4_1 _3976_ (.B(_1224_),
    .C(_1225_),
    .A(_1223_),
    .Y(_1229_),
    .D(_1228_));
 sg13g2_nand3b_1 _3977_ (.B(_1222_),
    .C(_1229_),
    .Y(_1230_),
    .A_N(_1221_));
 sg13g2_nand2_2 _3978_ (.Y(_1231_),
    .A(_1219_),
    .B(_1230_));
 sg13g2_nor2_2 _3979_ (.A(net655),
    .B(_1231_),
    .Y(_1232_));
 sg13g2_nand2_1 _3980_ (.Y(_1233_),
    .A(net731),
    .B(_1232_));
 sg13g2_nand2_1 _3981_ (.Y(_1234_),
    .A(_1808_),
    .B(net731));
 sg13g2_o21ai_1 _3982_ (.B1(_1234_),
    .Y(_1235_),
    .A1(_1826_),
    .A2(_1231_));
 sg13g2_nand3_1 _3983_ (.B(_1233_),
    .C(_1235_),
    .A(_1827_),
    .Y(_1236_));
 sg13g2_nand2_2 _3984_ (.Y(_1237_),
    .A(\Pong.datapath.rightPaddle[2] ),
    .B(_0425_));
 sg13g2_nand2_2 _3985_ (.Y(_1238_),
    .A(_1812_),
    .B(_1237_));
 sg13g2_nand3_1 _3986_ (.B(_0065_),
    .C(_1237_),
    .A(_1812_),
    .Y(_1239_));
 sg13g2_xnor2_1 _3987_ (.Y(_1240_),
    .A(_0065_),
    .B(_1238_));
 sg13g2_o21ai_1 _3988_ (.B1(_1240_),
    .Y(_1241_),
    .A1(_0065_),
    .A2(_1992_));
 sg13g2_xor2_1 _3989_ (.B(_1239_),
    .A(_0061_),
    .X(_1242_));
 sg13g2_nor3_2 _3990_ (.A(\Pong.datapath.rightPaddle[5] ),
    .B(\Pong.datapath.rightPaddle[4] ),
    .C(_1238_),
    .Y(_1243_));
 sg13g2_nand2_2 _3991_ (.Y(_1244_),
    .A(_1810_),
    .B(_1243_));
 sg13g2_xnor2_1 _3992_ (.Y(_1245_),
    .A(net726),
    .B(_1243_));
 sg13g2_a21oi_1 _3993_ (.A1(_1241_),
    .A2(_1242_),
    .Y(_1246_),
    .B1(net725));
 sg13g2_and3_1 _3994_ (.X(_1247_),
    .A(_0056_),
    .B(_1245_),
    .C(_1246_));
 sg13g2_nor2_1 _3995_ (.A(net725),
    .B(_1244_),
    .Y(_1248_));
 sg13g2_xnor2_1 _3996_ (.Y(_1249_),
    .A(_0058_),
    .B(_1248_));
 sg13g2_nor2b_1 _3997_ (.A(_1249_),
    .B_N(_1247_),
    .Y(_1250_));
 sg13g2_nand2b_1 _3998_ (.Y(_1251_),
    .B(net731),
    .A_N(net573));
 sg13g2_a21oi_1 _3999_ (.A1(_1234_),
    .A2(net572),
    .Y(_1252_),
    .B1(_1827_));
 sg13g2_a21oi_1 _4000_ (.A1(_1251_),
    .A2(_1252_),
    .Y(_1253_),
    .B1(net719));
 sg13g2_a221oi_1 _4001_ (.B2(_1253_),
    .C1(_1209_),
    .B1(_1236_),
    .A1(net719),
    .Y(_0149_),
    .A2(_1234_));
 sg13g2_nand2_1 _4002_ (.Y(_1254_),
    .A(_1808_),
    .B(net729));
 sg13g2_o21ai_1 _4003_ (.B1(_1254_),
    .Y(_1255_),
    .A1(net655),
    .A2(_1231_));
 sg13g2_a21oi_1 _4004_ (.A1(_0426_),
    .A2(_1232_),
    .Y(_1256_),
    .B1(net723));
 sg13g2_nand2_1 _4005_ (.Y(_1257_),
    .A(_1255_),
    .B(_1256_));
 sg13g2_nor2_1 _4006_ (.A(_0426_),
    .B(net572),
    .Y(_1258_));
 sg13g2_a21oi_1 _4007_ (.A1(net572),
    .A2(_1254_),
    .Y(_1259_),
    .B1(_1258_));
 sg13g2_a21oi_1 _4008_ (.A1(net723),
    .A2(_1259_),
    .Y(_1260_),
    .B1(net720));
 sg13g2_a221oi_1 _4009_ (.B2(_1260_),
    .C1(_1209_),
    .B1(_1257_),
    .A1(net720),
    .Y(_0150_),
    .A2(_1254_));
 sg13g2_or2_1 _4010_ (.X(_1261_),
    .B(net727),
    .A(\Pong.datapath.NES_activity_Left[5] ));
 sg13g2_mux2_1 _4011_ (.A0(_1226_),
    .A1(_1261_),
    .S(_1231_),
    .X(_1262_));
 sg13g2_a21o_1 _4012_ (.A2(_1261_),
    .A1(_1826_),
    .B1(net723),
    .X(_1263_));
 sg13g2_a21oi_1 _4013_ (.A1(\Pong.datapath.NES_activity_Right[2] ),
    .A2(_1262_),
    .Y(_1264_),
    .B1(_1263_));
 sg13g2_nand2_1 _4014_ (.Y(_1265_),
    .A(_0452_),
    .B(_1237_));
 sg13g2_o21ai_1 _4015_ (.B1(net723),
    .Y(_1266_),
    .A1(net572),
    .A2(_1265_));
 sg13g2_a21oi_1 _4016_ (.A1(net572),
    .A2(_1261_),
    .Y(_1267_),
    .B1(_1266_));
 sg13g2_or3_1 _4017_ (.A(net719),
    .B(_1264_),
    .C(_1267_),
    .X(_1268_));
 sg13g2_nand2_1 _4018_ (.Y(_1269_),
    .A(net719),
    .B(_1261_));
 sg13g2_nand2_2 _4019_ (.Y(_1270_),
    .A(net749),
    .B(_1807_));
 sg13g2_nor2_2 _4020_ (.A(net463),
    .B(_1208_),
    .Y(_1271_));
 sg13g2_nand3_1 _4021_ (.B(_1269_),
    .C(_1271_),
    .A(_1268_),
    .Y(_0151_));
 sg13g2_nand2_2 _4022_ (.Y(_1272_),
    .A(net656),
    .B(_1812_));
 sg13g2_mux2_1 _4023_ (.A0(_1227_),
    .A1(_1272_),
    .S(_1231_),
    .X(_1273_));
 sg13g2_nand2_1 _4024_ (.Y(_1274_),
    .A(net508),
    .B(_1273_));
 sg13g2_a21oi_1 _4025_ (.A1(net655),
    .A2(_1272_),
    .Y(_1275_),
    .B1(net723));
 sg13g2_nand2_1 _4026_ (.Y(_1276_),
    .A(net572),
    .B(_1272_));
 sg13g2_nand3_1 _4027_ (.B(\Pong.datapath.rightPaddle[2] ),
    .C(_0425_),
    .A(\Pong.datapath.rightPaddle[3] ),
    .Y(_1277_));
 sg13g2_a21oi_1 _4028_ (.A1(_1238_),
    .A2(_1277_),
    .Y(_1278_),
    .B1(net572));
 sg13g2_nor2_1 _4029_ (.A(_1827_),
    .B(_1278_),
    .Y(_1279_));
 sg13g2_a221oi_1 _4030_ (.B2(_1279_),
    .C1(net719),
    .B1(_1276_),
    .A1(_1274_),
    .Y(_1280_),
    .A2(_1275_));
 sg13g2_nand2_1 _4031_ (.Y(_1281_),
    .A(net719),
    .B(_1272_));
 sg13g2_nand3b_1 _4032_ (.B(_1281_),
    .C(_1271_),
    .Y(_0152_),
    .A_N(_1280_));
 sg13g2_nand2_1 _4033_ (.Y(_1282_),
    .A(net656),
    .B(_1813_));
 sg13g2_a21oi_1 _4034_ (.A1(_1219_),
    .A2(_1230_),
    .Y(_1283_),
    .B1(_1282_));
 sg13g2_nand3_1 _4035_ (.B(_1224_),
    .C(_1230_),
    .A(_1219_),
    .Y(_1284_));
 sg13g2_nor2_1 _4036_ (.A(net655),
    .B(_1283_),
    .Y(_1285_));
 sg13g2_a221oi_1 _4037_ (.B2(_1285_),
    .C1(net722),
    .B1(_1284_),
    .A1(net655),
    .Y(_1286_),
    .A2(_1282_));
 sg13g2_o21ai_1 _4038_ (.B1(net722),
    .Y(_1287_),
    .A1(_1240_),
    .A2(net573));
 sg13g2_a21oi_1 _4039_ (.A1(net572),
    .A2(_1282_),
    .Y(_1288_),
    .B1(_1287_));
 sg13g2_or3_1 _4040_ (.A(net719),
    .B(_1286_),
    .C(_1288_),
    .X(_1289_));
 sg13g2_nand2_1 _4041_ (.Y(_1290_),
    .A(net719),
    .B(_1282_));
 sg13g2_nand3_1 _4042_ (.B(_1289_),
    .C(_1290_),
    .A(_1271_),
    .Y(_0153_));
 sg13g2_nand2_1 _4043_ (.Y(_1291_),
    .A(net656),
    .B(\Pong.datapath.rightPaddle[5] ));
 sg13g2_o21ai_1 _4044_ (.B1(_1291_),
    .Y(_1292_),
    .A1(net655),
    .A2(_1231_));
 sg13g2_a21oi_1 _4045_ (.A1(_1225_),
    .A2(_1232_),
    .Y(_1293_),
    .B1(net722));
 sg13g2_nor2_1 _4046_ (.A(_1242_),
    .B(net573),
    .Y(_1294_));
 sg13g2_a21oi_1 _4047_ (.A1(net573),
    .A2(_1291_),
    .Y(_1295_),
    .B1(_1294_));
 sg13g2_a221oi_1 _4048_ (.B2(net722),
    .C1(net720),
    .B1(_1295_),
    .A1(_1292_),
    .Y(_1296_),
    .A2(_1293_));
 sg13g2_a21oi_1 _4049_ (.A1(net720),
    .A2(_1291_),
    .Y(_1297_),
    .B1(_1209_));
 sg13g2_nor2b_1 _4050_ (.A(_1296_),
    .B_N(_1297_),
    .Y(_0154_));
 sg13g2_nand2_1 _4051_ (.Y(_1298_),
    .A(net656),
    .B(_1810_));
 sg13g2_a21oi_1 _4052_ (.A1(_1219_),
    .A2(_1230_),
    .Y(_1299_),
    .B1(_1298_));
 sg13g2_nand3_1 _4053_ (.B(_1223_),
    .C(_1230_),
    .A(_1219_),
    .Y(_1300_));
 sg13g2_nor2_1 _4054_ (.A(net655),
    .B(_1299_),
    .Y(_1301_));
 sg13g2_a221oi_1 _4055_ (.B2(_1301_),
    .C1(net722),
    .B1(_1300_),
    .A1(net655),
    .Y(_1302_),
    .A2(_1298_));
 sg13g2_a21oi_1 _4056_ (.A1(net573),
    .A2(_1298_),
    .Y(_1303_),
    .B1(_1827_));
 sg13g2_a21oi_1 _4057_ (.A1(_1245_),
    .A2(_1303_),
    .Y(_1304_),
    .B1(net720));
 sg13g2_nand2b_1 _4058_ (.Y(_1305_),
    .B(_1304_),
    .A_N(_1302_));
 sg13g2_nand2_1 _4059_ (.Y(_1306_),
    .A(net720),
    .B(_1298_));
 sg13g2_nand3_1 _4060_ (.B(_1305_),
    .C(_1306_),
    .A(_1271_),
    .Y(_0155_));
 sg13g2_nor2_2 _4061_ (.A(\Pong.datapath.NES_activity_Left[5] ),
    .B(net725),
    .Y(_1307_));
 sg13g2_a22oi_1 _4062_ (.Y(_1308_),
    .B1(_1231_),
    .B2(_1307_),
    .A2(_1221_),
    .A1(_1219_));
 sg13g2_o21ai_1 _4063_ (.B1(_1827_),
    .Y(_1309_),
    .A1(\Pong.datapath.NES_activity_Right[2] ),
    .A2(_1307_));
 sg13g2_a21oi_1 _4064_ (.A1(\Pong.datapath.NES_activity_Right[2] ),
    .A2(_1308_),
    .Y(_1310_),
    .B1(_1309_));
 sg13g2_o21ai_1 _4065_ (.B1(net722),
    .Y(_1311_),
    .A1(net725),
    .A2(_1244_));
 sg13g2_a21oi_1 _4066_ (.A1(net724),
    .A2(_1244_),
    .Y(_1312_),
    .B1(net573));
 sg13g2_nor2_1 _4067_ (.A(_1307_),
    .B(_1312_),
    .Y(_1313_));
 sg13g2_o21ai_1 _4068_ (.B1(_1822_),
    .Y(_1314_),
    .A1(_1311_),
    .A2(_1313_));
 sg13g2_nor2_1 _4069_ (.A(_1822_),
    .B(_1307_),
    .Y(_1315_));
 sg13g2_nor3_1 _4070_ (.A(net463),
    .B(_1208_),
    .C(_1315_),
    .Y(_1316_));
 sg13g2_o21ai_1 _4071_ (.B1(_1316_),
    .Y(_0156_),
    .A1(_1310_),
    .A2(_1314_));
 sg13g2_nor2_1 _4072_ (.A(net477),
    .B(_1809_),
    .Y(_1317_));
 sg13g2_mux2_1 _4073_ (.A0(_1317_),
    .A1(_1222_),
    .S(_1232_),
    .X(_1318_));
 sg13g2_a21oi_1 _4074_ (.A1(_1247_),
    .A2(_1317_),
    .Y(_1319_),
    .B1(_1249_));
 sg13g2_o21ai_1 _4075_ (.B1(_1822_),
    .Y(_1320_),
    .A1(_1827_),
    .A2(_1319_));
 sg13g2_a21oi_1 _4076_ (.A1(_1827_),
    .A2(_1318_),
    .Y(_1321_),
    .B1(_1320_));
 sg13g2_nor2_1 _4077_ (.A(_1822_),
    .B(_1317_),
    .Y(_1322_));
 sg13g2_nor3_1 _4078_ (.A(_1209_),
    .B(_1321_),
    .C(_1322_),
    .Y(_0157_));
 sg13g2_nand2_1 _4079_ (.Y(_1323_),
    .A(net656),
    .B(\Pong.datapath.rightPaddle[9] ));
 sg13g2_or3_1 _4080_ (.A(net722),
    .B(_1232_),
    .C(_1323_),
    .X(_1324_));
 sg13g2_nor3_1 _4081_ (.A(\Pong.datapath.rightPaddle[8] ),
    .B(net724),
    .C(_1244_),
    .Y(_1325_));
 sg13g2_xnor2_1 _4082_ (.Y(_1326_),
    .A(_0056_),
    .B(_1325_));
 sg13g2_o21ai_1 _4083_ (.B1(net722),
    .Y(_1327_),
    .A1(net573),
    .A2(_1326_));
 sg13g2_a21oi_1 _4084_ (.A1(net573),
    .A2(_1323_),
    .Y(_1328_),
    .B1(_1327_));
 sg13g2_nor2_1 _4085_ (.A(net721),
    .B(_1328_),
    .Y(_1329_));
 sg13g2_a221oi_1 _4086_ (.B2(_1329_),
    .C1(_1209_),
    .B1(_1324_),
    .A1(net721),
    .Y(_0158_),
    .A2(_1323_));
 sg13g2_and2_1 _4087_ (.A(net747),
    .B(net229),
    .X(_0159_));
 sg13g2_and2_1 _4088_ (.A(net746),
    .B(net232),
    .X(_0160_));
 sg13g2_and2_1 _4089_ (.A(net746),
    .B(net230),
    .X(_0161_));
 sg13g2_and2_1 _4090_ (.A(net746),
    .B(net244),
    .X(_0162_));
 sg13g2_nor3_1 _4091_ (.A(\Pong.datapath.NES_wire_Right[2] ),
    .B(net240),
    .C(_1270_),
    .Y(_0163_));
 sg13g2_nor3_1 _4092_ (.A(\Pong.datapath.NES_wire_Right[3] ),
    .B(net249),
    .C(_1270_),
    .Y(_0164_));
 sg13g2_nor3_1 _4093_ (.A(\Pong.datapath.NES_wire_Right[4] ),
    .B(net236),
    .C(_1270_),
    .Y(_0165_));
 sg13g2_nor3_1 _4094_ (.A(\Pong.datapath.NES_wire_Right[5] ),
    .B(net242),
    .C(_1270_),
    .Y(_0166_));
 sg13g2_a21o_1 _4095_ (.A2(net717),
    .A1(net715),
    .B1(net713),
    .X(_1330_));
 sg13g2_nand2_1 _4096_ (.Y(_1331_),
    .A(net712),
    .B(_1330_));
 sg13g2_and2_1 _4097_ (.A(_2103_),
    .B(_1330_),
    .X(_1332_));
 sg13g2_nand2_1 _4098_ (.Y(_1333_),
    .A(net709),
    .B(_1332_));
 sg13g2_xnor2_1 _4099_ (.Y(_1334_),
    .A(_1818_),
    .B(_1333_));
 sg13g2_xor2_1 _4100_ (.B(_1332_),
    .A(_0073_),
    .X(_1335_));
 sg13g2_nand2_1 _4101_ (.Y(_1336_),
    .A(_2195_),
    .B(_1330_));
 sg13g2_xor2_1 _4102_ (.B(_0315_),
    .A(net712),
    .X(_1337_));
 sg13g2_nand2_1 _4103_ (.Y(_1338_),
    .A(_1336_),
    .B(_1337_));
 sg13g2_xnor2_1 _4104_ (.Y(_1339_),
    .A(_0074_),
    .B(_1331_));
 sg13g2_nand4_1 _4105_ (.B(_1335_),
    .C(_1338_),
    .A(_1334_),
    .Y(_1340_),
    .D(_1339_));
 sg13g2_nand4_1 _4106_ (.B(net707),
    .C(net709),
    .A(\Pong.datapath.leftPaddle[7] ),
    .Y(_1341_),
    .D(_1332_));
 sg13g2_nor2_1 _4107_ (.A(_0070_),
    .B(_1341_),
    .Y(_1342_));
 sg13g2_xor2_1 _4108_ (.B(_1341_),
    .A(_0070_),
    .X(_1343_));
 sg13g2_nor2_1 _4109_ (.A(_0072_),
    .B(_1333_),
    .Y(_1344_));
 sg13g2_xnor2_1 _4110_ (.Y(_1345_),
    .A(_0071_),
    .B(_1344_));
 sg13g2_nand3_1 _4111_ (.B(_1343_),
    .C(_1345_),
    .A(_1340_),
    .Y(_1346_));
 sg13g2_or3_1 _4112_ (.A(_1820_),
    .B(_2095_),
    .C(_1333_),
    .X(_1347_));
 sg13g2_xor2_1 _4113_ (.B(_1342_),
    .A(_0069_),
    .X(_1348_));
 sg13g2_nand3_1 _4114_ (.B(_1347_),
    .C(_1348_),
    .A(_1346_),
    .Y(_1349_));
 sg13g2_xnor2_1 _4115_ (.Y(_1350_),
    .A(net718),
    .B(_1349_));
 sg13g2_o21ai_1 _4116_ (.B1(_1829_),
    .Y(_1351_),
    .A1(net352),
    .A2(\Pong.datapath.NES_activity_Left[2] ));
 sg13g2_a21oi_1 _4117_ (.A1(\Pong.datapath.NES_activity_Left[2] ),
    .A2(_1350_),
    .Y(_1352_),
    .B1(_1351_));
 sg13g2_o21ai_1 _4118_ (.B1(net714),
    .Y(_1353_),
    .A1(net716),
    .A2(net717));
 sg13g2_nand2b_1 _4119_ (.Y(_1354_),
    .B(_1353_),
    .A_N(net712));
 sg13g2_nor3_1 _4120_ (.A(net709),
    .B(\Pong.datapath.leftPaddle[4] ),
    .C(_1354_),
    .Y(_1355_));
 sg13g2_or4_2 _4121_ (.A(\Pong.datapath.leftPaddle[6] ),
    .B(net709),
    .C(\Pong.datapath.leftPaddle[4] ),
    .D(_1354_),
    .X(_1356_));
 sg13g2_nor2_1 _4122_ (.A(\Pong.datapath.leftPaddle[7] ),
    .B(_1356_),
    .Y(_1357_));
 sg13g2_xnor2_1 _4123_ (.Y(_1358_),
    .A(_0070_),
    .B(_1357_));
 sg13g2_xnor2_1 _4124_ (.Y(_1359_),
    .A(net707),
    .B(_1355_));
 sg13g2_nand2_1 _4125_ (.Y(_1360_),
    .A(net706),
    .B(_1359_));
 sg13g2_nand3b_1 _4126_ (.B(_0074_),
    .C(_1353_),
    .Y(_1361_),
    .A_N(net712));
 sg13g2_xnor2_1 _4127_ (.Y(_1362_),
    .A(_0074_),
    .B(_1354_));
 sg13g2_o21ai_1 _4128_ (.B1(_1362_),
    .Y(_1363_),
    .A1(_0074_),
    .A2(_2059_));
 sg13g2_xor2_1 _4129_ (.B(_1361_),
    .A(_0073_),
    .X(_1364_));
 sg13g2_and2_1 _4130_ (.A(_1363_),
    .B(_1364_),
    .X(_1365_));
 sg13g2_nor4_2 _4131_ (.A(\Pong.datapath.leftPaddle[7] ),
    .B(_1358_),
    .C(_1360_),
    .Y(_1366_),
    .D(_1365_));
 sg13g2_xnor2_1 _4132_ (.Y(_1367_),
    .A(_1821_),
    .B(_1366_));
 sg13g2_a21oi_1 _4133_ (.A1(net705),
    .A2(_1367_),
    .Y(_1368_),
    .B1(_1352_));
 sg13g2_nand3_1 _4134_ (.B(_1093_),
    .C(_1186_),
    .A(net749),
    .Y(_1369_));
 sg13g2_nand2_1 _4135_ (.Y(_1370_),
    .A(net701),
    .B(net352));
 sg13g2_o21ai_1 _4136_ (.B1(_1370_),
    .Y(_1371_),
    .A1(net701),
    .A2(_1368_));
 sg13g2_nor2_1 _4137_ (.A(_1369_),
    .B(_1371_),
    .Y(_0167_));
 sg13g2_or2_1 _4138_ (.X(_1372_),
    .B(_1349_),
    .A(_1828_));
 sg13g2_nand2b_1 _4139_ (.Y(_1373_),
    .B(_0323_),
    .A_N(net571));
 sg13g2_a21oi_1 _4140_ (.A1(net253),
    .A2(net571),
    .Y(_1374_),
    .B1(net705));
 sg13g2_nand2_1 _4141_ (.Y(_1375_),
    .A(_1373_),
    .B(_1374_));
 sg13g2_o21ai_1 _4142_ (.B1(net704),
    .Y(_1376_),
    .A1(_0323_),
    .A2(net575));
 sg13g2_a21oi_1 _4143_ (.A1(net253),
    .A2(net575),
    .Y(_1377_),
    .B1(_1376_));
 sg13g2_nor2_1 _4144_ (.A(net702),
    .B(_1377_),
    .Y(_1378_));
 sg13g2_a221oi_1 _4145_ (.B2(_1378_),
    .C1(_1369_),
    .B1(_1375_),
    .A1(net702),
    .Y(_0168_),
    .A2(net253));
 sg13g2_mux2_1 _4146_ (.A0(_1336_),
    .A1(net714),
    .S(net571),
    .X(_1379_));
 sg13g2_o21ai_1 _4147_ (.B1(net714),
    .Y(_1380_),
    .A1(_0321_),
    .A2(net575));
 sg13g2_nor3_1 _4148_ (.A(net714),
    .B(_0321_),
    .C(net575),
    .Y(_1381_));
 sg13g2_nor2_1 _4149_ (.A(_1829_),
    .B(_1381_),
    .Y(_1382_));
 sg13g2_a21oi_1 _4150_ (.A1(_1380_),
    .A2(_1382_),
    .Y(_1383_),
    .B1(net700));
 sg13g2_o21ai_1 _4151_ (.B1(_1383_),
    .Y(_1384_),
    .A1(net704),
    .A2(_1379_));
 sg13g2_nand2_1 _4152_ (.Y(_1385_),
    .A(net714),
    .B(net703));
 sg13g2_nor3_2 _4153_ (.A(net463),
    .B(net502),
    .C(_1208_),
    .Y(_1386_));
 sg13g2_nand3_1 _4154_ (.B(_1385_),
    .C(_1386_),
    .A(_1384_),
    .Y(_0169_));
 sg13g2_mux2_1 _4155_ (.A0(_1337_),
    .A1(net712),
    .S(net571),
    .X(_1387_));
 sg13g2_a21oi_1 _4156_ (.A1(net713),
    .A2(_0322_),
    .Y(_1388_),
    .B1(net575));
 sg13g2_o21ai_1 _4157_ (.B1(net704),
    .Y(_1389_),
    .A1(net711),
    .A2(_1388_));
 sg13g2_a21oi_1 _4158_ (.A1(net711),
    .A2(_1388_),
    .Y(_1390_),
    .B1(_1389_));
 sg13g2_a21oi_1 _4159_ (.A1(_1829_),
    .A2(_1387_),
    .Y(_1391_),
    .B1(_1390_));
 sg13g2_o21ai_1 _4160_ (.B1(_1386_),
    .Y(_1392_),
    .A1(net703),
    .A2(_1391_));
 sg13g2_a21o_1 _4161_ (.A2(net703),
    .A1(net711),
    .B1(_1392_),
    .X(_0170_));
 sg13g2_nor2_1 _4162_ (.A(_1339_),
    .B(_1349_),
    .Y(_1393_));
 sg13g2_and2_1 _4163_ (.A(net710),
    .B(_1349_),
    .X(_1394_));
 sg13g2_o21ai_1 _4164_ (.B1(\Pong.datapath.NES_activity_Left[2] ),
    .Y(_1395_),
    .A1(_1393_),
    .A2(_1394_));
 sg13g2_a21oi_1 _4165_ (.A1(net710),
    .A2(_1828_),
    .Y(_1396_),
    .B1(net705));
 sg13g2_nor2_1 _4166_ (.A(_1362_),
    .B(_1366_),
    .Y(_1397_));
 sg13g2_a21oi_1 _4167_ (.A1(net710),
    .A2(net575),
    .Y(_1398_),
    .B1(_1397_));
 sg13g2_a221oi_1 _4168_ (.B2(net705),
    .C1(net700),
    .B1(_1398_),
    .A1(_1395_),
    .Y(_1399_),
    .A2(_1396_));
 sg13g2_a21oi_1 _4169_ (.A1(net710),
    .A2(net700),
    .Y(_1400_),
    .B1(_1399_));
 sg13g2_nand2_1 _4170_ (.Y(_0171_),
    .A(_1386_),
    .B(_1400_));
 sg13g2_nand2b_1 _4171_ (.Y(_1401_),
    .B(_1335_),
    .A_N(_1372_));
 sg13g2_a21oi_1 _4172_ (.A1(_0073_),
    .A2(net571),
    .Y(_1402_),
    .B1(net705));
 sg13g2_nand2_1 _4173_ (.Y(_1403_),
    .A(_1401_),
    .B(_1402_));
 sg13g2_o21ai_1 _4174_ (.B1(net704),
    .Y(_1404_),
    .A1(_1364_),
    .A2(_1366_));
 sg13g2_a21oi_1 _4175_ (.A1(_0073_),
    .A2(net575),
    .Y(_1405_),
    .B1(_1404_));
 sg13g2_nor2_1 _4176_ (.A(net700),
    .B(_1405_),
    .Y(_1406_));
 sg13g2_a221oi_1 _4177_ (.B2(_1406_),
    .C1(_1369_),
    .B1(_1403_),
    .A1(net519),
    .Y(_0172_),
    .A2(net700));
 sg13g2_nand2_1 _4178_ (.Y(_1407_),
    .A(net707),
    .B(_1349_));
 sg13g2_o21ai_1 _4179_ (.B1(_1407_),
    .Y(_1408_),
    .A1(_1334_),
    .A2(_1349_));
 sg13g2_o21ai_1 _4180_ (.B1(_1829_),
    .Y(_1409_),
    .A1(_1818_),
    .A2(\Pong.datapath.NES_activity_Left[2] ));
 sg13g2_a21oi_1 _4181_ (.A1(\Pong.datapath.NES_activity_Left[2] ),
    .A2(_1408_),
    .Y(_1410_),
    .B1(_1409_));
 sg13g2_nand2_1 _4182_ (.Y(_1411_),
    .A(net704),
    .B(_1359_));
 sg13g2_a21oi_1 _4183_ (.A1(net707),
    .A2(net575),
    .Y(_1412_),
    .B1(_1411_));
 sg13g2_or3_1 _4184_ (.A(net700),
    .B(_1410_),
    .C(_1412_),
    .X(_1413_));
 sg13g2_nand2_1 _4185_ (.Y(_1414_),
    .A(net707),
    .B(net703));
 sg13g2_nand3_1 _4186_ (.B(_1413_),
    .C(_1414_),
    .A(_1386_),
    .Y(_0173_));
 sg13g2_mux2_1 _4187_ (.A0(_1345_),
    .A1(\Pong.datapath.leftPaddle[7] ),
    .S(net571),
    .X(_1415_));
 sg13g2_xnor2_1 _4188_ (.Y(_1416_),
    .A(_1817_),
    .B(_1356_));
 sg13g2_a21oi_1 _4189_ (.A1(net704),
    .A2(_1416_),
    .Y(_1417_),
    .B1(net703));
 sg13g2_o21ai_1 _4190_ (.B1(_1417_),
    .Y(_1418_),
    .A1(net704),
    .A2(_1415_));
 sg13g2_nand2_1 _4191_ (.Y(_1419_),
    .A(net512),
    .B(net703));
 sg13g2_nand3_1 _4192_ (.B(_1418_),
    .C(_1419_),
    .A(_1386_),
    .Y(_0174_));
 sg13g2_o21ai_1 _4193_ (.B1(_1829_),
    .Y(_1420_),
    .A1(_1343_),
    .A2(net571));
 sg13g2_a21o_1 _4194_ (.A2(_1372_),
    .A1(_0070_),
    .B1(_1420_),
    .X(_1421_));
 sg13g2_a21oi_1 _4195_ (.A1(net705),
    .A2(_1358_),
    .Y(_1422_),
    .B1(net701));
 sg13g2_a221oi_1 _4196_ (.B2(_1422_),
    .C1(_1369_),
    .B1(_1421_),
    .A1(_0070_),
    .Y(_0175_),
    .A2(net701));
 sg13g2_nor4_1 _4197_ (.A(\Pong.datapath.leftPaddle[8] ),
    .B(\Pong.datapath.leftPaddle[7] ),
    .C(_1829_),
    .D(_1356_),
    .Y(_1423_));
 sg13g2_nor2_1 _4198_ (.A(net706),
    .B(_1423_),
    .Y(_1424_));
 sg13g2_o21ai_1 _4199_ (.B1(_1424_),
    .Y(_1425_),
    .A1(net704),
    .A2(net571));
 sg13g2_a21oi_1 _4200_ (.A1(net706),
    .A2(_1423_),
    .Y(_1426_),
    .B1(net700));
 sg13g2_a22oi_1 _4201_ (.Y(_1427_),
    .B1(_1425_),
    .B2(_1426_),
    .A2(net700),
    .A1(net706));
 sg13g2_nor2b_1 _4202_ (.A(_1369_),
    .B_N(_1427_),
    .Y(_0176_));
 sg13g2_nand2_2 _4203_ (.Y(_1428_),
    .A(net749),
    .B(_1808_));
 sg13g2_nor3_1 _4204_ (.A(\Pong.datapath.NES_wire_Left[2] ),
    .B(net247),
    .C(_1428_),
    .Y(_0177_));
 sg13g2_nor3_1 _4205_ (.A(\Pong.datapath.NES_wire_Left[3] ),
    .B(net251),
    .C(_1428_),
    .Y(_0178_));
 sg13g2_nor3_1 _4206_ (.A(\Pong.datapath.NES_wire_Left[4] ),
    .B(net238),
    .C(_1428_),
    .Y(_0179_));
 sg13g2_nor3_1 _4207_ (.A(\Pong.datapath.NES_wire_Left[5] ),
    .B(net245),
    .C(_1428_),
    .Y(_0180_));
 sg13g2_and2_1 _4208_ (.A(net750),
    .B(net233),
    .X(_0181_));
 sg13g2_and2_1 _4209_ (.A(net750),
    .B(net234),
    .X(_0182_));
 sg13g2_and2_1 _4210_ (.A(net749),
    .B(net235),
    .X(_0183_));
 sg13g2_and2_1 _4211_ (.A(net750),
    .B(net231),
    .X(_0184_));
 sg13g2_nor3_2 _4212_ (.A(_0588_),
    .B(_1059_),
    .C(_1070_),
    .Y(_1429_));
 sg13g2_nand3_1 _4213_ (.B(net691),
    .C(net695),
    .A(net676),
    .Y(_1430_));
 sg13g2_nand2_1 _4214_ (.Y(_1431_),
    .A(_1792_),
    .B(_0598_));
 sg13g2_a21o_1 _4215_ (.A2(_1066_),
    .A1(_0598_),
    .B1(_1788_),
    .X(_1432_));
 sg13g2_nor3_1 _4216_ (.A(_0596_),
    .B(_1430_),
    .C(_1431_),
    .Y(_1433_));
 sg13g2_and2_1 _4217_ (.A(_1429_),
    .B(_1432_),
    .X(_1434_));
 sg13g2_o21ai_1 _4218_ (.B1(_1429_),
    .Y(_1435_),
    .A1(_1432_),
    .A2(_1433_));
 sg13g2_inv_1 _4219_ (.Y(_1436_),
    .A(net639));
 sg13g2_nand2_1 _4220_ (.Y(_1437_),
    .A(net698),
    .B(_1436_));
 sg13g2_o21ai_1 _4221_ (.B1(net745),
    .Y(_1438_),
    .A1(net698),
    .A2(net640));
 sg13g2_a21oi_1 _4222_ (.A1(net698),
    .A2(_1436_),
    .Y(_0185_),
    .B1(_1438_));
 sg13g2_o21ai_1 _4223_ (.B1(net745),
    .Y(_1439_),
    .A1(_0530_),
    .A2(net639));
 sg13g2_a21oi_1 _4224_ (.A1(_1794_),
    .A2(_1437_),
    .Y(_0186_),
    .B1(_1439_));
 sg13g2_nor2_1 _4225_ (.A(net694),
    .B(_0530_),
    .Y(_1440_));
 sg13g2_xor2_1 _4226_ (.B(_0530_),
    .A(net694),
    .X(_1441_));
 sg13g2_a22oi_1 _4227_ (.Y(_1442_),
    .B1(_1441_),
    .B2(net640),
    .A2(net639),
    .A1(net695));
 sg13g2_nor2_1 _4228_ (.A(net739),
    .B(_1442_),
    .Y(_0187_));
 sg13g2_xnor2_1 _4229_ (.Y(_1443_),
    .A(net516),
    .B(_1440_));
 sg13g2_a22oi_1 _4230_ (.Y(_1444_),
    .B1(_1443_),
    .B2(_1434_),
    .A2(_1435_),
    .A1(net691));
 sg13g2_nor2_1 _4231_ (.A(net739),
    .B(_1444_),
    .Y(_0188_));
 sg13g2_nor2_1 _4232_ (.A(net688),
    .B(_0532_),
    .Y(_1445_));
 sg13g2_xnor2_1 _4233_ (.Y(_1446_),
    .A(net688),
    .B(_0532_));
 sg13g2_o21ai_1 _4234_ (.B1(net1),
    .Y(_1447_),
    .A1(net690),
    .A2(_1434_));
 sg13g2_a21oi_1 _4235_ (.A1(net640),
    .A2(_1446_),
    .Y(_0189_),
    .B1(_1447_));
 sg13g2_xnor2_1 _4236_ (.Y(_1448_),
    .A(net685),
    .B(_1445_));
 sg13g2_a22oi_1 _4237_ (.Y(_1449_),
    .B1(_1448_),
    .B2(net640),
    .A2(net639),
    .A1(net687));
 sg13g2_nor2_1 _4238_ (.A(net739),
    .B(_1449_),
    .Y(_0190_));
 sg13g2_or3_2 _4239_ (.A(_1791_),
    .B(_1792_),
    .C(_0532_),
    .X(_1450_));
 sg13g2_xor2_1 _4240_ (.B(_1450_),
    .A(net682),
    .X(_1451_));
 sg13g2_a22oi_1 _4241_ (.Y(_1452_),
    .B1(_1451_),
    .B2(net640),
    .A2(net639),
    .A1(net683));
 sg13g2_nor2_1 _4242_ (.A(net738),
    .B(_1452_),
    .Y(_0191_));
 sg13g2_o21ai_1 _4243_ (.B1(net475),
    .Y(_1453_),
    .A1(net682),
    .A2(_1450_));
 sg13g2_nor3_1 _4244_ (.A(net682),
    .B(net475),
    .C(_1450_),
    .Y(_1454_));
 sg13g2_nor2b_1 _4245_ (.A(_1454_),
    .B_N(net640),
    .Y(_1455_));
 sg13g2_a22oi_1 _4246_ (.Y(_1456_),
    .B1(_1453_),
    .B2(_1455_),
    .A2(net639),
    .A1(net680));
 sg13g2_nor2_1 _4247_ (.A(net738),
    .B(net476),
    .Y(_0192_));
 sg13g2_o21ai_1 _4248_ (.B1(net678),
    .Y(_1457_),
    .A1(_0508_),
    .A2(_1450_));
 sg13g2_nor3_1 _4249_ (.A(net678),
    .B(_0508_),
    .C(_1450_),
    .Y(_1458_));
 sg13g2_nor2b_1 _4250_ (.A(_1458_),
    .B_N(net640),
    .Y(_1459_));
 sg13g2_a22oi_1 _4251_ (.Y(_1460_),
    .B1(_1457_),
    .B2(_1459_),
    .A2(net639),
    .A1(net679));
 sg13g2_nor2_1 _4252_ (.A(net738),
    .B(_1460_),
    .Y(_0193_));
 sg13g2_xnor2_1 _4253_ (.Y(_1461_),
    .A(net675),
    .B(_1458_));
 sg13g2_a22oi_1 _4254_ (.Y(_1462_),
    .B1(_1461_),
    .B2(net640),
    .A2(net639),
    .A1(net676));
 sg13g2_nor2_1 _4255_ (.A(net738),
    .B(_1462_),
    .Y(_0194_));
 sg13g2_nor2b_2 _4256_ (.A(_0109_),
    .B_N(net659),
    .Y(_1463_));
 sg13g2_and2_2 _4257_ (.A(_0558_),
    .B(_1463_),
    .X(_1464_));
 sg13g2_nand2_2 _4258_ (.Y(_1465_),
    .A(_0558_),
    .B(_1463_));
 sg13g2_o21ai_1 _4259_ (.B1(net745),
    .Y(_1466_),
    .A1(net388),
    .A2(_1465_));
 sg13g2_a21oi_1 _4260_ (.A1(net674),
    .A2(_1465_),
    .Y(_0195_),
    .B1(_1466_));
 sg13g2_a21oi_1 _4261_ (.A1(net674),
    .A2(_1465_),
    .Y(_1467_),
    .B1(net673));
 sg13g2_o21ai_1 _4262_ (.B1(net744),
    .Y(_1468_),
    .A1(_1069_),
    .A2(_1464_));
 sg13g2_nor2_1 _4263_ (.A(_1467_),
    .B(_1468_),
    .Y(_0196_));
 sg13g2_nor2_2 _4264_ (.A(_1429_),
    .B(_1464_),
    .Y(_1469_));
 sg13g2_nor2_1 _4265_ (.A(_0089_),
    .B(_1069_),
    .Y(_1470_));
 sg13g2_xor2_1 _4266_ (.B(_1069_),
    .A(_0089_),
    .X(_1471_));
 sg13g2_a22oi_1 _4267_ (.Y(_1472_),
    .B1(_1469_),
    .B2(_1471_),
    .A2(_1464_),
    .A1(net672));
 sg13g2_nor2_1 _4268_ (.A(net735),
    .B(net496),
    .Y(_0197_));
 sg13g2_xnor2_1 _4269_ (.Y(_1473_),
    .A(_0090_),
    .B(_1470_));
 sg13g2_a22oi_1 _4270_ (.Y(_1474_),
    .B1(_1469_),
    .B2(_1473_),
    .A2(_1464_),
    .A1(net670));
 sg13g2_nor2_1 _4271_ (.A(net735),
    .B(net493),
    .Y(_0198_));
 sg13g2_nor2_1 _4272_ (.A(_0091_),
    .B(_1070_),
    .Y(_1475_));
 sg13g2_xor2_1 _4273_ (.B(_1070_),
    .A(_0091_),
    .X(_1476_));
 sg13g2_a22oi_1 _4274_ (.Y(_1477_),
    .B1(_1469_),
    .B2(_1476_),
    .A2(_1464_),
    .A1(net668));
 sg13g2_nor2_1 _4275_ (.A(net735),
    .B(net504),
    .Y(_0199_));
 sg13g2_xnor2_1 _4276_ (.Y(_1478_),
    .A(_0092_),
    .B(_1475_));
 sg13g2_a22oi_1 _4277_ (.Y(_1479_),
    .B1(_1469_),
    .B2(_1478_),
    .A2(_1463_),
    .A1(net666));
 sg13g2_nor2_1 _4278_ (.A(net735),
    .B(net535),
    .Y(_0200_));
 sg13g2_nor2_1 _4279_ (.A(_0390_),
    .B(_1070_),
    .Y(_1480_));
 sg13g2_nor3_1 _4280_ (.A(_0093_),
    .B(_0390_),
    .C(_1070_),
    .Y(_1481_));
 sg13g2_xnor2_1 _4281_ (.Y(_1482_),
    .A(_0093_),
    .B(_1480_));
 sg13g2_a22oi_1 _4282_ (.Y(_1483_),
    .B1(_1469_),
    .B2(_1482_),
    .A2(_1464_),
    .A1(net665));
 sg13g2_nor2_1 _4283_ (.A(net735),
    .B(net480),
    .Y(_0201_));
 sg13g2_xnor2_1 _4284_ (.Y(_1484_),
    .A(_0094_),
    .B(_1481_));
 sg13g2_a22oi_1 _4285_ (.Y(_1485_),
    .B1(_1469_),
    .B2(_1484_),
    .A2(_1463_),
    .A1(net663));
 sg13g2_nor2_1 _4286_ (.A(net735),
    .B(net499),
    .Y(_0202_));
 sg13g2_and3_1 _4287_ (.X(_1486_),
    .A(net662),
    .B(net664),
    .C(_1480_));
 sg13g2_nor2b_1 _4288_ (.A(_0109_),
    .B_N(_1486_),
    .Y(_1487_));
 sg13g2_xnor2_1 _4289_ (.Y(_1488_),
    .A(_0109_),
    .B(_1486_));
 sg13g2_a22oi_1 _4290_ (.Y(_1489_),
    .B1(_1469_),
    .B2(_1488_),
    .A2(_1464_),
    .A1(net661));
 sg13g2_nor2_1 _4291_ (.A(net736),
    .B(_1489_),
    .Y(_0203_));
 sg13g2_xor2_1 _4292_ (.B(_1487_),
    .A(net533),
    .X(_1490_));
 sg13g2_o21ai_1 _4293_ (.B1(_1465_),
    .Y(_1491_),
    .A1(_1429_),
    .A2(_1490_));
 sg13g2_and2_1 _4294_ (.A(net743),
    .B(_1491_),
    .X(_0204_));
 sg13g2_nand3_1 _4295_ (.B(\Pong.datapath.NES_counter_left.Q[4] ),
    .C(\Pong.datapath.NES_counter_left.Q[3] ),
    .A(\Pong.datapath.NES_counter_left.Q[7] ),
    .Y(_1492_));
 sg13g2_o21ai_1 _4296_ (.B1(\Pong.datapath.NES_counter_left.Q[7] ),
    .Y(_1493_),
    .A1(\Pong.datapath.NES_counter_left.Q[6] ),
    .A2(\Pong.datapath.NES_counter_left.Q[5] ));
 sg13g2_nand3_1 _4297_ (.B(_1492_),
    .C(_1493_),
    .A(_0115_),
    .Y(_1494_));
 sg13g2_nand2_1 _4298_ (.Y(_1495_),
    .A(_0115_),
    .B(_1838_));
 sg13g2_a21oi_2 _4299_ (.B1(_1786_),
    .Y(_1496_),
    .A2(_1495_),
    .A1(_1494_));
 sg13g2_nand2_2 _4300_ (.Y(_1497_),
    .A(net748),
    .B(_1803_));
 sg13g2_a21oi_1 _4301_ (.A1(_1786_),
    .A2(_1494_),
    .Y(_1498_),
    .B1(_1497_));
 sg13g2_nor2b_1 _4302_ (.A(_1496_),
    .B_N(_1498_),
    .Y(_0205_));
 sg13g2_xnor2_1 _4303_ (.Y(_1499_),
    .A(net424),
    .B(_1496_));
 sg13g2_nor2_1 _4304_ (.A(_1497_),
    .B(net425),
    .Y(_0206_));
 sg13g2_a21oi_1 _4305_ (.A1(\Pong.datapath.NES_counter_left.Q[1] ),
    .A2(_1496_),
    .Y(_1500_),
    .B1(net317));
 sg13g2_and3_1 _4306_ (.X(_1501_),
    .A(net317),
    .B(net424),
    .C(_1496_));
 sg13g2_nor3_1 _4307_ (.A(_1497_),
    .B(net318),
    .C(_1501_),
    .Y(_0207_));
 sg13g2_nor2_1 _4308_ (.A(net430),
    .B(_1501_),
    .Y(_1502_));
 sg13g2_nand2b_1 _4309_ (.Y(_1503_),
    .B(_1495_),
    .A_N(_1497_));
 sg13g2_and2_1 _4310_ (.A(net430),
    .B(_1501_),
    .X(_1504_));
 sg13g2_nor3_1 _4311_ (.A(_1502_),
    .B(_1503_),
    .C(_1504_),
    .Y(_0208_));
 sg13g2_nor2_1 _4312_ (.A(net410),
    .B(_1504_),
    .Y(_1505_));
 sg13g2_and2_1 _4313_ (.A(net410),
    .B(_1504_),
    .X(_1506_));
 sg13g2_nor3_1 _4314_ (.A(_1503_),
    .B(net411),
    .C(_1506_),
    .Y(_0209_));
 sg13g2_nor2_1 _4315_ (.A(net392),
    .B(_1506_),
    .Y(_1507_));
 sg13g2_and2_1 _4316_ (.A(net392),
    .B(_1506_),
    .X(_1508_));
 sg13g2_nor3_1 _4317_ (.A(_1497_),
    .B(net393),
    .C(_1508_),
    .Y(_0210_));
 sg13g2_xnor2_1 _4318_ (.Y(_1509_),
    .A(net382),
    .B(_1508_));
 sg13g2_nor2_1 _4319_ (.A(_1497_),
    .B(_1509_),
    .Y(_0211_));
 sg13g2_a22oi_1 _4320_ (.Y(_1510_),
    .B1(_1508_),
    .B2(net382),
    .A2(_1495_),
    .A1(\Pong.datapath.NES_counter_left.Q[7] ));
 sg13g2_nor2_1 _4321_ (.A(_1497_),
    .B(net383),
    .Y(_0212_));
 sg13g2_nand3_1 _4322_ (.B(\Pong.datapath.NES_counter_right.Q[4] ),
    .C(\Pong.datapath.NES_counter_right.Q[3] ),
    .A(\Pong.datapath.NES_counter_right.Q[7] ),
    .Y(_1511_));
 sg13g2_o21ai_1 _4323_ (.B1(\Pong.datapath.NES_counter_right.Q[7] ),
    .Y(_1512_),
    .A1(\Pong.datapath.NES_counter_right.Q[6] ),
    .A2(\Pong.datapath.NES_counter_right.Q[5] ));
 sg13g2_nand3_1 _4324_ (.B(_1511_),
    .C(_1512_),
    .A(_0116_),
    .Y(_1513_));
 sg13g2_nand2_1 _4325_ (.Y(_1514_),
    .A(_0116_),
    .B(_1870_));
 sg13g2_a21oi_1 _4326_ (.A1(_1513_),
    .A2(_1514_),
    .Y(_1515_),
    .B1(_1785_));
 sg13g2_nand2_2 _4327_ (.Y(_1516_),
    .A(net747),
    .B(_1801_));
 sg13g2_inv_1 _4328_ (.Y(_1517_),
    .A(_1516_));
 sg13g2_a21oi_1 _4329_ (.A1(_1785_),
    .A2(_1513_),
    .Y(_1518_),
    .B1(_1516_));
 sg13g2_nor2b_1 _4330_ (.A(_1515_),
    .B_N(net483),
    .Y(_0213_));
 sg13g2_and2_1 _4331_ (.A(net449),
    .B(_1515_),
    .X(_1519_));
 sg13g2_o21ai_1 _4332_ (.B1(_1517_),
    .Y(_1520_),
    .A1(net449),
    .A2(_1515_));
 sg13g2_nor2_1 _4333_ (.A(_1519_),
    .B(net450),
    .Y(_0214_));
 sg13g2_nor2_1 _4334_ (.A(net357),
    .B(_1519_),
    .Y(_1521_));
 sg13g2_and2_1 _4335_ (.A(net357),
    .B(_1519_),
    .X(_1522_));
 sg13g2_nor3_1 _4336_ (.A(_1516_),
    .B(net358),
    .C(_1522_),
    .Y(_0215_));
 sg13g2_nor2_1 _4337_ (.A(net405),
    .B(_1522_),
    .Y(_1523_));
 sg13g2_nand2_1 _4338_ (.Y(_1524_),
    .A(_1514_),
    .B(_1517_));
 sg13g2_and2_1 _4339_ (.A(net405),
    .B(_1522_),
    .X(_1525_));
 sg13g2_nor3_1 _4340_ (.A(_1523_),
    .B(_1524_),
    .C(_1525_),
    .Y(_0216_));
 sg13g2_nor2_1 _4341_ (.A(net377),
    .B(_1525_),
    .Y(_1526_));
 sg13g2_and2_1 _4342_ (.A(net377),
    .B(_1525_),
    .X(_1527_));
 sg13g2_nor3_1 _4343_ (.A(_1524_),
    .B(net378),
    .C(_1527_),
    .Y(_0217_));
 sg13g2_and2_1 _4344_ (.A(net446),
    .B(_1527_),
    .X(_1528_));
 sg13g2_o21ai_1 _4345_ (.B1(_1517_),
    .Y(_1529_),
    .A1(net446),
    .A2(_1527_));
 sg13g2_nor2_1 _4346_ (.A(_1528_),
    .B(_1529_),
    .Y(_0218_));
 sg13g2_o21ai_1 _4347_ (.B1(_1517_),
    .Y(_1530_),
    .A1(net375),
    .A2(_1528_));
 sg13g2_a21oi_1 _4348_ (.A1(net375),
    .A2(_1528_),
    .Y(_0219_),
    .B1(_1530_));
 sg13g2_a22oi_1 _4349_ (.Y(_1531_),
    .B1(_1528_),
    .B2(\Pong.datapath.NES_counter_right.Q[6] ),
    .A2(_1514_),
    .A1(net365));
 sg13g2_nor2_1 _4350_ (.A(_1516_),
    .B(net366),
    .Y(_0220_));
 sg13g2_nand2_1 _4351_ (.Y(_1532_),
    .A(_1784_),
    .B(_1857_));
 sg13g2_nor2_1 _4352_ (.A(\Pong.datapath.NES_delay_counter_left.Q[16] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[15] ),
    .Y(_1533_));
 sg13g2_nor2b_1 _4353_ (.A(\Pong.datapath.NES_delay_counter_left.Q[12] ),
    .B_N(_0112_),
    .Y(_1534_));
 sg13g2_o21ai_1 _4354_ (.B1(_1533_),
    .Y(_1535_),
    .A1(_1848_),
    .A2(_1534_));
 sg13g2_a21oi_1 _4355_ (.A1(_1851_),
    .A2(_1532_),
    .Y(_1536_),
    .B1(_1535_));
 sg13g2_o21ai_1 _4356_ (.B1(net337),
    .Y(_1537_),
    .A1(_1852_),
    .A2(_1536_));
 sg13g2_inv_1 _4357_ (.Y(_1538_),
    .A(_1537_));
 sg13g2_nand2_2 _4358_ (.Y(_1539_),
    .A(_1859_),
    .B(_1537_));
 sg13g2_inv_1 _4359_ (.Y(_1540_),
    .A(_1539_));
 sg13g2_nor2_1 _4360_ (.A(net444),
    .B(_1539_),
    .Y(_1541_));
 sg13g2_a21oi_1 _4361_ (.A1(net444),
    .A2(_1539_),
    .Y(_1542_),
    .B1(net735));
 sg13g2_nor2b_1 _4362_ (.A(_1541_),
    .B_N(_1542_),
    .Y(_0221_));
 sg13g2_a21oi_1 _4363_ (.A1(\Pong.datapath.NES_delay_counter_left.Q[0] ),
    .A2(_1539_),
    .Y(_1543_),
    .B1(net286));
 sg13g2_and3_1 _4364_ (.X(_1544_),
    .A(net286),
    .B(\Pong.datapath.NES_delay_counter_left.Q[0] ),
    .C(_1539_));
 sg13g2_nor3_1 _4365_ (.A(net736),
    .B(net287),
    .C(_1544_),
    .Y(_0222_));
 sg13g2_and2_1 _4366_ (.A(net428),
    .B(_1544_),
    .X(_1545_));
 sg13g2_o21ai_1 _4367_ (.B1(net743),
    .Y(_1546_),
    .A1(net428),
    .A2(_1544_));
 sg13g2_nor2_1 _4368_ (.A(_1545_),
    .B(net429),
    .Y(_0223_));
 sg13g2_and2_1 _4369_ (.A(net445),
    .B(_1545_),
    .X(_1547_));
 sg13g2_o21ai_1 _4370_ (.B1(net743),
    .Y(_1548_),
    .A1(net445),
    .A2(_1545_));
 sg13g2_nor2_1 _4371_ (.A(_1547_),
    .B(_1548_),
    .Y(_0224_));
 sg13g2_xnor2_1 _4372_ (.Y(_1549_),
    .A(net435),
    .B(_1547_));
 sg13g2_nor2_1 _4373_ (.A(net736),
    .B(net436),
    .Y(_0225_));
 sg13g2_a21oi_1 _4374_ (.A1(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .A2(_1547_),
    .Y(_1550_),
    .B1(net306));
 sg13g2_and3_1 _4375_ (.X(_1551_),
    .A(net306),
    .B(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .C(_1547_));
 sg13g2_nor3_1 _4376_ (.A(net736),
    .B(net307),
    .C(_1551_),
    .Y(_0226_));
 sg13g2_o21ai_1 _4377_ (.B1(net743),
    .Y(_1552_),
    .A1(net326),
    .A2(_1551_));
 sg13g2_a21oi_1 _4378_ (.A1(net326),
    .A2(_1551_),
    .Y(_0227_),
    .B1(_1552_));
 sg13g2_a21oi_1 _4379_ (.A1(\Pong.datapath.NES_delay_counter_left.Q[6] ),
    .A2(_1551_),
    .Y(_1553_),
    .B1(net279));
 sg13g2_nor3_2 _4380_ (.A(net540),
    .B(_1855_),
    .C(_1540_),
    .Y(_1554_));
 sg13g2_nor3_1 _4381_ (.A(net736),
    .B(net280),
    .C(_1554_),
    .Y(_0228_));
 sg13g2_nor2_1 _4382_ (.A(net409),
    .B(_1554_),
    .Y(_1555_));
 sg13g2_nand2_2 _4383_ (.Y(_1556_),
    .A(net743),
    .B(_1859_));
 sg13g2_and2_1 _4384_ (.A(net409),
    .B(_1554_),
    .X(_1557_));
 sg13g2_nor3_1 _4385_ (.A(_1555_),
    .B(_1556_),
    .C(_1557_),
    .Y(_0229_));
 sg13g2_a21oi_1 _4386_ (.A1(net453),
    .A2(_1557_),
    .Y(_1558_),
    .B1(_1556_));
 sg13g2_o21ai_1 _4387_ (.B1(_1558_),
    .Y(_1559_),
    .A1(net453),
    .A2(_1557_));
 sg13g2_inv_1 _4388_ (.Y(_0230_),
    .A(_1559_));
 sg13g2_a21oi_1 _4389_ (.A1(\Pong.datapath.NES_delay_counter_left.Q[9] ),
    .A2(_1557_),
    .Y(_1560_),
    .B1(net298));
 sg13g2_nor3_1 _4390_ (.A(_1784_),
    .B(_1849_),
    .C(_1857_),
    .Y(_1561_));
 sg13g2_nor2b_1 _4391_ (.A(_1849_),
    .B_N(_1557_),
    .Y(_1562_));
 sg13g2_nor3_1 _4392_ (.A(_1556_),
    .B(net299),
    .C(_1562_),
    .Y(_0231_));
 sg13g2_nor4_2 _4393_ (.A(_1784_),
    .B(_1849_),
    .C(_1853_),
    .Y(_1563_),
    .D(_1855_));
 sg13g2_xnor2_1 _4394_ (.Y(_1564_),
    .A(net414),
    .B(_1563_));
 sg13g2_a22oi_1 _4395_ (.Y(_1565_),
    .B1(_1564_),
    .B2(_1538_),
    .A2(_1540_),
    .A1(net396));
 sg13g2_nor2_1 _4396_ (.A(net736),
    .B(_1565_),
    .Y(_0232_));
 sg13g2_nand3_1 _4397_ (.B(\Pong.datapath.NES_delay_counter_left.Q[11] ),
    .C(_1563_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[12] ),
    .Y(_1566_));
 sg13g2_a21oi_1 _4398_ (.A1(net396),
    .A2(_1562_),
    .Y(_1567_),
    .B1(\Pong.datapath.NES_delay_counter_left.Q[12] ));
 sg13g2_nand4_1 _4399_ (.B(\Pong.datapath.NES_delay_counter_left.Q[11] ),
    .C(_1538_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[12] ),
    .Y(_1568_),
    .D(_1561_));
 sg13g2_nand2_1 _4400_ (.Y(_1569_),
    .A(net743),
    .B(_1568_));
 sg13g2_nor2_1 _4401_ (.A(net397),
    .B(_1569_),
    .Y(_0233_));
 sg13g2_o21ai_1 _4402_ (.B1(_1568_),
    .Y(_1570_),
    .A1(_1783_),
    .A2(_1860_));
 sg13g2_o21ai_1 _4403_ (.B1(_1570_),
    .Y(_1571_),
    .A1(_1783_),
    .A2(_1568_));
 sg13g2_nor2_1 _4404_ (.A(net739),
    .B(net507),
    .Y(_0234_));
 sg13g2_o21ai_1 _4405_ (.B1(_1782_),
    .Y(_1572_),
    .A1(_1783_),
    .A2(_1568_));
 sg13g2_inv_1 _4406_ (.Y(_1573_),
    .A(net460));
 sg13g2_nor2_2 _4407_ (.A(_1848_),
    .B(_1568_),
    .Y(_1574_));
 sg13g2_nor3_1 _4408_ (.A(_1556_),
    .B(_1573_),
    .C(_1574_),
    .Y(_0235_));
 sg13g2_xnor2_1 _4409_ (.Y(_1575_),
    .A(net467),
    .B(_1574_));
 sg13g2_nor2_1 _4410_ (.A(net736),
    .B(net468),
    .Y(_0236_));
 sg13g2_a21o_1 _4411_ (.A2(_1574_),
    .A1(net467),
    .B1(net514),
    .X(_1576_));
 sg13g2_nand3_1 _4412_ (.B(\Pong.datapath.NES_delay_counter_left.Q[15] ),
    .C(_1574_),
    .A(net514),
    .Y(_1577_));
 sg13g2_and3_1 _4413_ (.X(_0237_),
    .A(net743),
    .B(_1576_),
    .C(_1577_));
 sg13g2_nand3_1 _4414_ (.B(\Pong.datapath.NES_delay_counter_left.Q[16] ),
    .C(\Pong.datapath.NES_delay_counter_left.Q[15] ),
    .A(\Pong.datapath.NES_delay_counter_left.Q[17] ),
    .Y(_1578_));
 sg13g2_nor3_1 _4415_ (.A(_1848_),
    .B(_1566_),
    .C(_1578_),
    .Y(_1579_));
 sg13g2_or2_1 _4416_ (.X(_1580_),
    .B(_1579_),
    .A(_1537_));
 sg13g2_a221oi_1 _4417_ (.B2(_1539_),
    .C1(net735),
    .B1(_1580_),
    .A1(_1781_),
    .Y(_0238_),
    .A2(_1577_));
 sg13g2_a21oi_1 _4418_ (.A1(\Pong.control_unit.NES_Controller_Left.state_NESController[0] ),
    .A2(_1579_),
    .Y(_1581_),
    .B1(net259));
 sg13g2_nor2_1 _4419_ (.A(_1556_),
    .B(net260),
    .Y(_0239_));
 sg13g2_nand3_1 _4420_ (.B(\Pong.datapath.NES_delay_counter_right.Q[9] ),
    .C(\Pong.datapath.NES_delay_counter_right.Q[8] ),
    .A(\Pong.datapath.NES_delay_counter_right.Q[10] ),
    .Y(_1582_));
 sg13g2_nor2b_1 _4421_ (.A(\Pong.datapath.NES_delay_counter_right.Q[12] ),
    .B_N(_0111_),
    .Y(_1583_));
 sg13g2_o21ai_1 _4422_ (.B1(_1583_),
    .Y(_1584_),
    .A1(\Pong.datapath.NES_delay_counter_right.Q[11] ),
    .A2(_1582_));
 sg13g2_and2_1 _4423_ (.A(_1885_),
    .B(_1584_),
    .X(_1585_));
 sg13g2_nor4_1 _4424_ (.A(\Pong.datapath.NES_delay_counter_right.Q[16] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .C(_1894_),
    .D(_1585_),
    .Y(_1586_));
 sg13g2_nor2_1 _4425_ (.A(_1878_),
    .B(_1586_),
    .Y(_1587_));
 sg13g2_nor2_1 _4426_ (.A(_1801_),
    .B(_1587_),
    .Y(_1588_));
 sg13g2_inv_1 _4427_ (.Y(_1589_),
    .A(_1588_));
 sg13g2_o21ai_1 _4428_ (.B1(_1895_),
    .Y(_1590_),
    .A1(_1801_),
    .A2(_1587_));
 sg13g2_inv_1 _4429_ (.Y(_1591_),
    .A(_1590_));
 sg13g2_nor2_1 _4430_ (.A(net370),
    .B(_1590_),
    .Y(_1592_));
 sg13g2_and2_1 _4431_ (.A(net370),
    .B(_1590_),
    .X(_1593_));
 sg13g2_nor3_1 _4432_ (.A(net740),
    .B(_1592_),
    .C(_1593_),
    .Y(_0240_));
 sg13g2_xnor2_1 _4433_ (.Y(_1594_),
    .A(net408),
    .B(_1593_));
 sg13g2_nor2_1 _4434_ (.A(net740),
    .B(_1594_),
    .Y(_0241_));
 sg13g2_a21oi_1 _4435_ (.A1(net408),
    .A2(_1593_),
    .Y(_1595_),
    .B1(net457));
 sg13g2_a21oi_1 _4436_ (.A1(_1880_),
    .A2(_1593_),
    .Y(_1596_),
    .B1(_1595_));
 sg13g2_and2_1 _4437_ (.A(net746),
    .B(_1596_),
    .X(_0242_));
 sg13g2_a21oi_1 _4438_ (.A1(_1880_),
    .A2(_1593_),
    .Y(_1597_),
    .B1(net267));
 sg13g2_nor2_1 _4439_ (.A(_1881_),
    .B(_1591_),
    .Y(_1598_));
 sg13g2_nor3_1 _4440_ (.A(net740),
    .B(net268),
    .C(_1598_),
    .Y(_0243_));
 sg13g2_nor2_1 _4441_ (.A(net368),
    .B(_1598_),
    .Y(_1599_));
 sg13g2_and2_1 _4442_ (.A(net368),
    .B(_1598_),
    .X(_1600_));
 sg13g2_nor3_1 _4443_ (.A(net740),
    .B(net369),
    .C(_1600_),
    .Y(_0244_));
 sg13g2_nand2_1 _4444_ (.Y(_1601_),
    .A(net407),
    .B(_1600_));
 sg13g2_xnor2_1 _4445_ (.Y(_1602_),
    .A(net407),
    .B(_1600_));
 sg13g2_nor2_1 _4446_ (.A(net740),
    .B(_1602_),
    .Y(_0245_));
 sg13g2_nand2b_1 _4447_ (.Y(_1603_),
    .B(_1601_),
    .A_N(net462));
 sg13g2_nand3_1 _4448_ (.B(net407),
    .C(_1600_),
    .A(net462),
    .Y(_1604_));
 sg13g2_and3_1 _4449_ (.X(_0246_),
    .A(net746),
    .B(_1603_),
    .C(_1604_));
 sg13g2_nor2b_1 _4450_ (.A(net324),
    .B_N(_1604_),
    .Y(_1605_));
 sg13g2_nor2_2 _4451_ (.A(_1883_),
    .B(_1591_),
    .Y(_1606_));
 sg13g2_nor3_1 _4452_ (.A(net740),
    .B(net325),
    .C(_1606_),
    .Y(_0247_));
 sg13g2_nand2_2 _4453_ (.Y(_1607_),
    .A(net747),
    .B(_1895_));
 sg13g2_xnor2_1 _4454_ (.Y(_1608_),
    .A(net466),
    .B(_1606_));
 sg13g2_nor2_1 _4455_ (.A(_1607_),
    .B(_1608_),
    .Y(_0248_));
 sg13g2_and3_1 _4456_ (.X(_1609_),
    .A(net362),
    .B(\Pong.datapath.NES_delay_counter_right.Q[8] ),
    .C(_1606_));
 sg13g2_a21oi_1 _4457_ (.A1(\Pong.datapath.NES_delay_counter_right.Q[8] ),
    .A2(_1606_),
    .Y(_1610_),
    .B1(net362));
 sg13g2_nor3_1 _4458_ (.A(_1607_),
    .B(_1609_),
    .C(net363),
    .Y(_0249_));
 sg13g2_nor2_1 _4459_ (.A(net385),
    .B(_1609_),
    .Y(_1611_));
 sg13g2_nor2_1 _4460_ (.A(_1883_),
    .B(_1582_),
    .Y(_1612_));
 sg13g2_and2_1 _4461_ (.A(_1590_),
    .B(_1612_),
    .X(_1613_));
 sg13g2_nor3_1 _4462_ (.A(_1607_),
    .B(net386),
    .C(_1613_),
    .Y(_0250_));
 sg13g2_xnor2_1 _4463_ (.Y(_1614_),
    .A(net412),
    .B(_1612_));
 sg13g2_a22oi_1 _4464_ (.Y(_1615_),
    .B1(_1614_),
    .B2(_1588_),
    .A2(_1591_),
    .A1(\Pong.datapath.NES_delay_counter_right.Q[11] ));
 sg13g2_nor2_1 _4465_ (.A(net740),
    .B(net413),
    .Y(_0251_));
 sg13g2_nand3_1 _4466_ (.B(\Pong.datapath.NES_delay_counter_right.Q[11] ),
    .C(_1612_),
    .A(net347),
    .Y(_1616_));
 sg13g2_nor2_2 _4467_ (.A(_1589_),
    .B(_1616_),
    .Y(_1617_));
 sg13g2_a21oi_1 _4468_ (.A1(\Pong.datapath.NES_delay_counter_right.Q[11] ),
    .A2(_1613_),
    .Y(_1618_),
    .B1(net347));
 sg13g2_nor3_1 _4469_ (.A(net740),
    .B(_1617_),
    .C(net348),
    .Y(_0252_));
 sg13g2_a21oi_1 _4470_ (.A1(net437),
    .A2(_1895_),
    .Y(_1619_),
    .B1(_1617_));
 sg13g2_a21oi_1 _4471_ (.A1(net437),
    .A2(_1617_),
    .Y(_1620_),
    .B1(net741));
 sg13g2_nor2b_1 _4472_ (.A(net438),
    .B_N(_1620_),
    .Y(_0253_));
 sg13g2_a21oi_1 _4473_ (.A1(\Pong.datapath.NES_delay_counter_right.Q[13] ),
    .A2(_1617_),
    .Y(_1621_),
    .B1(net283));
 sg13g2_and3_1 _4474_ (.X(_1622_),
    .A(net283),
    .B(\Pong.datapath.NES_delay_counter_right.Q[13] ),
    .C(_1617_));
 sg13g2_nor3_1 _4475_ (.A(_1607_),
    .B(net284),
    .C(_1622_),
    .Y(_0254_));
 sg13g2_or2_1 _4476_ (.X(_1623_),
    .B(_1622_),
    .A(net528));
 sg13g2_nand2_1 _4477_ (.Y(_1624_),
    .A(net528),
    .B(_1622_));
 sg13g2_and3_1 _4478_ (.X(_0255_),
    .A(net746),
    .B(_1623_),
    .C(_1624_));
 sg13g2_nand2b_1 _4479_ (.Y(_1625_),
    .B(_1624_),
    .A_N(net517));
 sg13g2_nand3_1 _4480_ (.B(net541),
    .C(_1622_),
    .A(net517),
    .Y(_1626_));
 sg13g2_and3_1 _4481_ (.X(_0256_),
    .A(net746),
    .B(net518),
    .C(_1626_));
 sg13g2_nand4_1 _4482_ (.B(\Pong.datapath.NES_delay_counter_right.Q[16] ),
    .C(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .A(\Pong.datapath.NES_delay_counter_right.Q[17] ),
    .Y(_1627_),
    .D(_1885_));
 sg13g2_nor2_1 _4483_ (.A(_1616_),
    .B(_1627_),
    .Y(_1628_));
 sg13g2_o21ai_1 _4484_ (.B1(_1590_),
    .Y(_1629_),
    .A1(_1589_),
    .A2(_1628_));
 sg13g2_nand2_1 _4485_ (.Y(_1630_),
    .A(net746),
    .B(_1629_));
 sg13g2_a21oi_1 _4486_ (.A1(_1780_),
    .A2(_1626_),
    .Y(_0257_),
    .B1(_1630_));
 sg13g2_a21oi_1 _4487_ (.A1(\Pong.control_unit.NES_Controller_Right.state_NESController[0] ),
    .A2(_1628_),
    .Y(_1631_),
    .B1(net255));
 sg13g2_nor2_1 _4488_ (.A(_1607_),
    .B(net256),
    .Y(_0258_));
 sg13g2_o21ai_1 _4489_ (.B1(_1932_),
    .Y(_1632_),
    .A1(\Pong.datapath.Ball_Clock.Q[6] ),
    .A2(\Pong.datapath.Ball_Clock.Q[5] ));
 sg13g2_o21ai_1 _4490_ (.B1(_1933_),
    .Y(_1633_),
    .A1(_0114_),
    .A2(_1930_));
 sg13g2_nand3_1 _4491_ (.B(\Pong.datapath.Ball_Clock.Q[15] ),
    .C(_1633_),
    .A(\Pong.datapath.Ball_Clock.Q[16] ),
    .Y(_1634_));
 sg13g2_and2_2 _4492_ (.A(_1632_),
    .B(_1634_),
    .X(_1635_));
 sg13g2_nor2_2 _4493_ (.A(net653),
    .B(_1635_),
    .Y(_1636_));
 sg13g2_or2_1 _4494_ (.X(_1637_),
    .B(_1635_),
    .A(net653));
 sg13g2_o21ai_1 _4495_ (.B1(net744),
    .Y(_1638_),
    .A1(net351),
    .A2(_1635_));
 sg13g2_a21oi_1 _4496_ (.A1(net351),
    .A2(_1637_),
    .Y(_0259_),
    .B1(_1638_));
 sg13g2_a21oi_1 _4497_ (.A1(\Pong.datapath.Ball_Clock.Q[0] ),
    .A2(_1637_),
    .Y(_1639_),
    .B1(net334));
 sg13g2_and3_1 _4498_ (.X(_1640_),
    .A(net334),
    .B(net351),
    .C(_1635_));
 sg13g2_nor3_1 _4499_ (.A(net737),
    .B(net335),
    .C(_1640_),
    .Y(_0260_));
 sg13g2_nand2_1 _4500_ (.Y(_1641_),
    .A(\Pong.datapath.Ball_Clock.Q[2] ),
    .B(\Pong.datapath.Ball_Clock.Q[1] ));
 sg13g2_and2_1 _4501_ (.A(net465),
    .B(_1640_),
    .X(_1642_));
 sg13g2_o21ai_1 _4502_ (.B1(net744),
    .Y(_1643_),
    .A1(net465),
    .A2(_1640_));
 sg13g2_nor2_1 _4503_ (.A(_1642_),
    .B(_1643_),
    .Y(_0261_));
 sg13g2_xnor2_1 _4504_ (.Y(_1644_),
    .A(net442),
    .B(_1642_));
 sg13g2_nor2_1 _4505_ (.A(net737),
    .B(net443),
    .Y(_0262_));
 sg13g2_a21oi_1 _4506_ (.A1(\Pong.datapath.Ball_Clock.Q[3] ),
    .A2(_1642_),
    .Y(_1645_),
    .B1(net330));
 sg13g2_and3_1 _4507_ (.X(_1646_),
    .A(net330),
    .B(net442),
    .C(_1642_));
 sg13g2_nor3_1 _4508_ (.A(net737),
    .B(net331),
    .C(_1646_),
    .Y(_0263_));
 sg13g2_nand2b_2 _4509_ (.Y(_1647_),
    .B(net744),
    .A_N(net653));
 sg13g2_xnor2_1 _4510_ (.Y(_1648_),
    .A(net454),
    .B(_1646_));
 sg13g2_nor2_1 _4511_ (.A(_1647_),
    .B(_1648_),
    .Y(_0264_));
 sg13g2_a21oi_1 _4512_ (.A1(\Pong.datapath.Ball_Clock.Q[5] ),
    .A2(_1646_),
    .Y(_1649_),
    .B1(net315));
 sg13g2_nand4_1 _4513_ (.B(\Pong.datapath.Ball_Clock.Q[5] ),
    .C(\Pong.datapath.Ball_Clock.Q[4] ),
    .A(\Pong.datapath.Ball_Clock.Q[6] ),
    .Y(_1650_),
    .D(\Pong.datapath.Ball_Clock.Q[3] ));
 sg13g2_nor3_2 _4514_ (.A(_1779_),
    .B(_1641_),
    .C(_1650_),
    .Y(_1651_));
 sg13g2_a21oi_1 _4515_ (.A1(_1637_),
    .A2(_1651_),
    .Y(_1652_),
    .B1(net737));
 sg13g2_nor2b_1 _4516_ (.A(net316),
    .B_N(_1652_),
    .Y(_0265_));
 sg13g2_and2_1 _4517_ (.A(\Pong.datapath.Ball_Clock.Q[7] ),
    .B(_1651_),
    .X(_1653_));
 sg13g2_xor2_1 _4518_ (.B(_1651_),
    .A(net401),
    .X(_1654_));
 sg13g2_a22oi_1 _4519_ (.Y(_1655_),
    .B1(_1654_),
    .B2(_1635_),
    .A2(_1636_),
    .A1(net401));
 sg13g2_nor2_1 _4520_ (.A(net737),
    .B(_1655_),
    .Y(_0266_));
 sg13g2_xnor2_1 _4521_ (.Y(_1656_),
    .A(_0114_),
    .B(_1653_));
 sg13g2_a22oi_1 _4522_ (.Y(_1657_),
    .B1(_1656_),
    .B2(_1635_),
    .A2(_1636_),
    .A1(net431));
 sg13g2_nor2_1 _4523_ (.A(net737),
    .B(net432),
    .Y(_0267_));
 sg13g2_nand3_1 _4524_ (.B(\Pong.datapath.Ball_Clock.Q[8] ),
    .C(_1653_),
    .A(net354),
    .Y(_1658_));
 sg13g2_a21oi_1 _4525_ (.A1(\Pong.datapath.Ball_Clock.Q[8] ),
    .A2(_1653_),
    .Y(_1659_),
    .B1(net354));
 sg13g2_a22oi_1 _4526_ (.Y(_1660_),
    .B1(_1658_),
    .B2(_1635_),
    .A2(_1636_),
    .A1(net354));
 sg13g2_nor3_1 _4527_ (.A(net737),
    .B(net355),
    .C(_1660_),
    .Y(_0268_));
 sg13g2_nor2_1 _4528_ (.A(_1636_),
    .B(_1658_),
    .Y(_1661_));
 sg13g2_nor2_1 _4529_ (.A(net371),
    .B(_1661_),
    .Y(_1662_));
 sg13g2_and2_1 _4530_ (.A(net371),
    .B(_1661_),
    .X(_1663_));
 sg13g2_nor3_1 _4531_ (.A(_1647_),
    .B(net372),
    .C(_1663_),
    .Y(_0269_));
 sg13g2_and2_1 _4532_ (.A(net458),
    .B(_1663_),
    .X(_1664_));
 sg13g2_o21ai_1 _4533_ (.B1(net744),
    .Y(_1665_),
    .A1(net458),
    .A2(_1663_));
 sg13g2_nor2_1 _4534_ (.A(_1664_),
    .B(_1665_),
    .Y(_0270_));
 sg13g2_nor2_1 _4535_ (.A(net416),
    .B(_1664_),
    .Y(_1666_));
 sg13g2_and2_1 _4536_ (.A(net416),
    .B(_1664_),
    .X(_1667_));
 sg13g2_nor3_1 _4537_ (.A(net737),
    .B(net417),
    .C(_1667_),
    .Y(_0271_));
 sg13g2_o21ai_1 _4538_ (.B1(net744),
    .Y(_1668_),
    .A1(net390),
    .A2(_1667_));
 sg13g2_a21oi_1 _4539_ (.A1(net390),
    .A2(_1667_),
    .Y(_0272_),
    .B1(_1668_));
 sg13g2_a21oi_1 _4540_ (.A1(\Pong.datapath.Ball_Clock.Q[13] ),
    .A2(_1667_),
    .Y(_1669_),
    .B1(net343));
 sg13g2_nand4_1 _4541_ (.B(\Pong.datapath.Ball_Clock.Q[13] ),
    .C(\Pong.datapath.Ball_Clock.Q[12] ),
    .A(\Pong.datapath.Ball_Clock.Q[14] ),
    .Y(_1670_),
    .D(\Pong.datapath.Ball_Clock.Q[11] ));
 sg13g2_nor2_1 _4542_ (.A(_1930_),
    .B(_1670_),
    .Y(_1671_));
 sg13g2_nand3_1 _4543_ (.B(_1653_),
    .C(_1671_),
    .A(\Pong.datapath.Ball_Clock.Q[8] ),
    .Y(_1672_));
 sg13g2_inv_1 _4544_ (.Y(_1673_),
    .A(_1672_));
 sg13g2_o21ai_1 _4545_ (.B1(net744),
    .Y(_1674_),
    .A1(_1636_),
    .A2(_1672_));
 sg13g2_nor2_1 _4546_ (.A(net344),
    .B(_1674_),
    .Y(_0273_));
 sg13g2_xor2_1 _4547_ (.B(_1672_),
    .A(net490),
    .X(_1675_));
 sg13g2_a21oi_1 _4548_ (.A1(_1637_),
    .A2(_1675_),
    .Y(_0274_),
    .B1(_1647_));
 sg13g2_a21oi_1 _4549_ (.A1(\Pong.datapath.Ball_Clock.Q[15] ),
    .A2(_1673_),
    .Y(_1676_),
    .B1(net274));
 sg13g2_nor2_1 _4550_ (.A(_1647_),
    .B(net275),
    .Y(_0275_));
 sg13g2_nand2_1 _4551_ (.Y(_1677_),
    .A(\Pong.control_unit.state_ballMovement[2] ),
    .B(_0110_));
 sg13g2_nand2_1 _4552_ (.Y(_1678_),
    .A(_1800_),
    .B(\Pong.control_unit.state_ballMovement[1] ));
 sg13g2_o21ai_1 _4553_ (.B1(_0110_),
    .Y(_1679_),
    .A1(\Pong.control_unit.state_ballMovement[2] ),
    .A2(_1678_));
 sg13g2_inv_1 _4554_ (.Y(_1680_),
    .A(_1679_));
 sg13g2_nor2_2 _4555_ (.A(\Pong.control_unit.state_ballMovement[3] ),
    .B(\Pong.control_unit.state_ballMovement[0] ),
    .Y(_1681_));
 sg13g2_nand2_2 _4556_ (.Y(_1682_),
    .A(_1799_),
    .B(_1800_));
 sg13g2_nor2_2 _4557_ (.A(_1679_),
    .B(_1682_),
    .Y(_1683_));
 sg13g2_nand2_1 _4558_ (.Y(_1684_),
    .A(_1677_),
    .B(_1681_));
 sg13g2_nand2_1 _4559_ (.Y(_1685_),
    .A(_1677_),
    .B(net638));
 sg13g2_or2_1 _4560_ (.X(_1686_),
    .B(_1685_),
    .A(net631));
 sg13g2_nor2_1 _4561_ (.A(_1799_),
    .B(_1679_),
    .Y(_1687_));
 sg13g2_nand2_1 _4562_ (.Y(_1688_),
    .A(\Pong.control_unit.state_ballMovement[3] ),
    .B(_1680_));
 sg13g2_o21ai_1 _4563_ (.B1(_1684_),
    .Y(_1689_),
    .A1(_0108_),
    .A2(net635));
 sg13g2_o21ai_1 _4564_ (.B1(net733),
    .Y(_1690_),
    .A1(net631),
    .A2(net578));
 sg13g2_a21oi_1 _4565_ (.A1(_1686_),
    .A2(_1689_),
    .Y(_0276_),
    .B1(_1690_));
 sg13g2_o21ai_1 _4566_ (.B1(net578),
    .Y(_1691_),
    .A1(_0632_),
    .A2(_1681_));
 sg13g2_a21oi_1 _4567_ (.A1(_0632_),
    .A2(net638),
    .Y(_1692_),
    .B1(_1691_));
 sg13g2_o21ai_1 _4568_ (.B1(net734),
    .Y(_1693_),
    .A1(net628),
    .A2(net578));
 sg13g2_nor2_1 _4569_ (.A(_1692_),
    .B(_1693_),
    .Y(_0277_));
 sg13g2_xnor2_1 _4570_ (.Y(_1694_),
    .A(_0067_),
    .B(_1950_));
 sg13g2_nor3_1 _4571_ (.A(_1681_),
    .B(net636),
    .C(_1694_),
    .Y(_1695_));
 sg13g2_nand2_1 _4572_ (.Y(_1696_),
    .A(_0670_),
    .B(net638));
 sg13g2_o21ai_1 _4573_ (.B1(_1696_),
    .Y(_1697_),
    .A1(net625),
    .A2(net578));
 sg13g2_o21ai_1 _4574_ (.B1(net733),
    .Y(_0278_),
    .A1(_1695_),
    .A2(_1697_));
 sg13g2_xnor2_1 _4575_ (.Y(_1698_),
    .A(_0068_),
    .B(_0664_));
 sg13g2_xor2_1 _4576_ (.B(_1955_),
    .A(_0068_),
    .X(_1699_));
 sg13g2_a221oi_1 _4577_ (.B2(_1682_),
    .C1(net636),
    .B1(_1699_),
    .A1(net638),
    .Y(_1700_),
    .A2(_1698_));
 sg13g2_a21oi_1 _4578_ (.A1(net624),
    .A2(net636),
    .Y(_1701_),
    .B1(_1700_));
 sg13g2_nand2_1 _4579_ (.Y(_0279_),
    .A(net734),
    .B(_1701_));
 sg13g2_xnor2_1 _4580_ (.Y(_1702_),
    .A(net621),
    .B(_0665_));
 sg13g2_a21oi_1 _4581_ (.A1(net621),
    .A2(_1956_),
    .Y(_1703_),
    .B1(_1681_));
 sg13g2_o21ai_1 _4582_ (.B1(_1703_),
    .Y(_1704_),
    .A1(net621),
    .A2(_1956_));
 sg13g2_a21oi_1 _4583_ (.A1(net638),
    .A2(_1702_),
    .Y(_1705_),
    .B1(net634));
 sg13g2_a22oi_1 _4584_ (.Y(_1706_),
    .B1(_1704_),
    .B2(_1705_),
    .A2(net636),
    .A1(net623));
 sg13g2_nand2_1 _4585_ (.Y(_0280_),
    .A(net733),
    .B(_1706_));
 sg13g2_xnor2_1 _4586_ (.Y(_1707_),
    .A(net619),
    .B(_1958_));
 sg13g2_nor3_1 _4587_ (.A(_1681_),
    .B(net634),
    .C(_1707_),
    .Y(_1708_));
 sg13g2_a221oi_1 _4588_ (.B2(net620),
    .C1(_1708_),
    .B1(net634),
    .A1(_0667_),
    .Y(_1709_),
    .A2(net638));
 sg13g2_nor2b_1 _4589_ (.A(_1709_),
    .B_N(net733),
    .Y(_0281_));
 sg13g2_o21ai_1 _4590_ (.B1(_1682_),
    .Y(_1710_),
    .A1(net616),
    .A2(_0614_));
 sg13g2_a21o_1 _4591_ (.A2(_0614_),
    .A1(net616),
    .B1(_1710_),
    .X(_1711_));
 sg13g2_xor2_1 _4592_ (.B(_0675_),
    .A(net616),
    .X(_1712_));
 sg13g2_a21oi_1 _4593_ (.A1(_1683_),
    .A2(_1712_),
    .Y(_1713_),
    .B1(net635));
 sg13g2_a22oi_1 _4594_ (.Y(_1714_),
    .B1(_1711_),
    .B2(_1713_),
    .A2(net634),
    .A1(net618));
 sg13g2_nand2_1 _4595_ (.Y(_0282_),
    .A(net733),
    .B(_1714_));
 sg13g2_xnor2_1 _4596_ (.Y(_1715_),
    .A(_1833_),
    .B(_0684_));
 sg13g2_o21ai_1 _4597_ (.B1(_1682_),
    .Y(_1716_),
    .A1(_0097_),
    .A2(_0615_));
 sg13g2_a21o_1 _4598_ (.A2(_0615_),
    .A1(_0097_),
    .B1(_1716_),
    .X(_1717_));
 sg13g2_a21oi_1 _4599_ (.A1(net638),
    .A2(_1715_),
    .Y(_1718_),
    .B1(net634));
 sg13g2_a22oi_1 _4600_ (.Y(_1719_),
    .B1(_1717_),
    .B2(_1718_),
    .A2(net634),
    .A1(net615));
 sg13g2_nand2_1 _4601_ (.Y(_0283_),
    .A(net734),
    .B(_1719_));
 sg13g2_a21oi_1 _4602_ (.A1(net610),
    .A2(_0620_),
    .Y(_1720_),
    .B1(_1681_));
 sg13g2_o21ai_1 _4603_ (.B1(_1720_),
    .Y(_1721_),
    .A1(net610),
    .A2(_0620_));
 sg13g2_xnor2_1 _4604_ (.Y(_1722_),
    .A(net610),
    .B(_0677_));
 sg13g2_a21oi_1 _4605_ (.A1(net638),
    .A2(_1722_),
    .Y(_1723_),
    .B1(net634));
 sg13g2_o21ai_1 _4606_ (.B1(net734),
    .Y(_1724_),
    .A1(net612),
    .A2(net578));
 sg13g2_a21oi_1 _4607_ (.A1(_1721_),
    .A2(_1723_),
    .Y(_0284_),
    .B1(_1724_));
 sg13g2_a21oi_1 _4608_ (.A1(_0113_),
    .A2(_0646_),
    .Y(_1725_),
    .B1(_1681_));
 sg13g2_o21ai_1 _4609_ (.B1(_1725_),
    .Y(_1726_),
    .A1(_0113_),
    .A2(_0646_));
 sg13g2_xnor2_1 _4610_ (.Y(_1727_),
    .A(_0113_),
    .B(_0679_));
 sg13g2_a21oi_1 _4611_ (.A1(_1683_),
    .A2(_1727_),
    .Y(_1728_),
    .B1(net634));
 sg13g2_o21ai_1 _4612_ (.B1(net734),
    .Y(_1729_),
    .A1(net608),
    .A2(net578));
 sg13g2_a21oi_1 _4613_ (.A1(_1726_),
    .A2(_1728_),
    .Y(_0285_),
    .B1(_1729_));
 sg13g2_or2_1 _4614_ (.X(_1730_),
    .B(_1685_),
    .A(\Pong.datapath.ballFunction.ball_center_x[0] ));
 sg13g2_o21ai_1 _4615_ (.B1(_1684_),
    .Y(_1731_),
    .A1(_0107_),
    .A2(net635));
 sg13g2_o21ai_1 _4616_ (.B1(net733),
    .Y(_1732_),
    .A1(\Pong.datapath.ballFunction.ball_center_x[0] ),
    .A2(net577));
 sg13g2_a21oi_1 _4617_ (.A1(_1730_),
    .A2(_1731_),
    .Y(_0286_),
    .B1(_1732_));
 sg13g2_a21oi_2 _4618_ (.B1(\Pong.control_unit.state_ballMovement[3] ),
    .Y(_1733_),
    .A2(_1677_),
    .A1(_1800_));
 sg13g2_nor2_1 _4619_ (.A(_1680_),
    .B(_1682_),
    .Y(_1734_));
 sg13g2_nor3_1 _4620_ (.A(net633),
    .B(net654),
    .C(_1734_),
    .Y(_1735_));
 sg13g2_nand2_1 _4621_ (.Y(_1736_),
    .A(_0872_),
    .B(net574));
 sg13g2_nor2b_1 _4622_ (.A(_0872_),
    .B_N(net654),
    .Y(_1737_));
 sg13g2_nor2_1 _4623_ (.A(net633),
    .B(_1737_),
    .Y(_1738_));
 sg13g2_o21ai_1 _4624_ (.B1(net732),
    .Y(_1739_),
    .A1(net606),
    .A2(net577));
 sg13g2_a21oi_1 _4625_ (.A1(_1736_),
    .A2(_1738_),
    .Y(_0287_),
    .B1(_1739_));
 sg13g2_a221oi_1 _4626_ (.B2(_0898_),
    .C1(net633),
    .B1(net574),
    .A1(_0876_),
    .Y(_1740_),
    .A2(net654));
 sg13g2_o21ai_1 _4627_ (.B1(net732),
    .Y(_1741_),
    .A1(net604),
    .A2(net577));
 sg13g2_nor2_1 _4628_ (.A(_1740_),
    .B(_1741_),
    .Y(_0288_));
 sg13g2_xnor2_1 _4629_ (.Y(_1742_),
    .A(_0100_),
    .B(_2163_));
 sg13g2_xnor2_1 _4630_ (.Y(_1743_),
    .A(_0100_),
    .B(_0896_));
 sg13g2_a221oi_1 _4631_ (.B2(_1735_),
    .C1(net633),
    .B1(_1743_),
    .A1(_1733_),
    .Y(_1744_),
    .A2(_1742_));
 sg13g2_o21ai_1 _4632_ (.B1(net733),
    .Y(_1745_),
    .A1(net601),
    .A2(net578));
 sg13g2_nor2_1 _4633_ (.A(_1744_),
    .B(_1745_),
    .Y(_0289_));
 sg13g2_nand2b_1 _4634_ (.Y(_1746_),
    .B(net574),
    .A_N(_0916_));
 sg13g2_a21oi_1 _4635_ (.A1(net599),
    .A2(_2152_),
    .Y(_1747_),
    .B1(_1746_));
 sg13g2_o21ai_1 _4636_ (.B1(net654),
    .Y(_1748_),
    .A1(net599),
    .A2(_0864_));
 sg13g2_a21oi_1 _4637_ (.A1(net599),
    .A2(_0864_),
    .Y(_1749_),
    .B1(_1748_));
 sg13g2_nor3_1 _4638_ (.A(net637),
    .B(_1747_),
    .C(_1749_),
    .Y(_1750_));
 sg13g2_o21ai_1 _4639_ (.B1(net732),
    .Y(_1751_),
    .A1(net600),
    .A2(net577));
 sg13g2_nor2_1 _4640_ (.A(_1750_),
    .B(_1751_),
    .Y(_0290_));
 sg13g2_a22oi_1 _4641_ (.Y(_1752_),
    .B1(net574),
    .B2(_0916_),
    .A2(_1733_),
    .A1(_0865_));
 sg13g2_inv_1 _4642_ (.Y(_1753_),
    .A(_1752_));
 sg13g2_o21ai_1 _4643_ (.B1(net654),
    .Y(_1754_),
    .A1(_2162_),
    .A2(_0708_));
 sg13g2_a21oi_1 _4644_ (.A1(_1746_),
    .A2(_1754_),
    .Y(_1755_),
    .B1(_0102_));
 sg13g2_a221oi_1 _4645_ (.B2(_0102_),
    .C1(_1755_),
    .B1(_1753_),
    .A1(net598),
    .Y(_1756_),
    .A2(net637));
 sg13g2_nor2b_1 _4646_ (.A(_1756_),
    .B_N(net732),
    .Y(_0291_));
 sg13g2_xnor2_1 _4647_ (.Y(_1757_),
    .A(_0103_),
    .B(_0866_));
 sg13g2_xnor2_1 _4648_ (.Y(_1758_),
    .A(_0103_),
    .B(_0891_));
 sg13g2_a221oi_1 _4649_ (.B2(net574),
    .C1(net633),
    .B1(_1758_),
    .A1(net654),
    .Y(_1759_),
    .A2(_1757_));
 sg13g2_a21oi_1 _4650_ (.A1(net596),
    .A2(net633),
    .Y(_1760_),
    .B1(_1759_));
 sg13g2_nand2_1 _4651_ (.Y(_0292_),
    .A(net732),
    .B(_1760_));
 sg13g2_xor2_1 _4652_ (.B(_0868_),
    .A(_0104_),
    .X(_1761_));
 sg13g2_xnor2_1 _4653_ (.Y(_1762_),
    .A(_0104_),
    .B(_0892_));
 sg13g2_a22oi_1 _4654_ (.Y(_1763_),
    .B1(_1762_),
    .B2(net574),
    .A2(_1761_),
    .A1(net654));
 sg13g2_o21ai_1 _4655_ (.B1(net732),
    .Y(_1764_),
    .A1(net595),
    .A2(net577));
 sg13g2_a21oi_1 _4656_ (.A1(net577),
    .A2(_1763_),
    .Y(_0293_),
    .B1(_1764_));
 sg13g2_xor2_1 _4657_ (.B(_0867_),
    .A(_0105_),
    .X(_1765_));
 sg13g2_o21ai_1 _4658_ (.B1(_0105_),
    .Y(_1766_),
    .A1(net591),
    .A2(_0748_));
 sg13g2_nand2b_1 _4659_ (.Y(_1767_),
    .B(_1766_),
    .A_N(_0899_));
 sg13g2_a221oi_1 _4660_ (.B2(net574),
    .C1(net633),
    .B1(_1767_),
    .A1(net654),
    .Y(_1768_),
    .A2(_1765_));
 sg13g2_a21oi_1 _4661_ (.A1(net594),
    .A2(net633),
    .Y(_1769_),
    .B1(_1768_));
 sg13g2_nand2_1 _4662_ (.Y(_0294_),
    .A(net732),
    .B(_1769_));
 sg13g2_xnor2_1 _4663_ (.Y(_1770_),
    .A(_0106_),
    .B(_0869_));
 sg13g2_xnor2_1 _4664_ (.Y(_1771_),
    .A(_0106_),
    .B(_0899_));
 sg13g2_a22oi_1 _4665_ (.Y(_1772_),
    .B1(_1771_),
    .B2(net574),
    .A2(_1770_),
    .A1(_1733_));
 sg13g2_o21ai_1 _4666_ (.B1(net732),
    .Y(_1773_),
    .A1(\Pong.datapath.ballFunction.ball_center_x[9] ),
    .A2(net577));
 sg13g2_a21oi_1 _4667_ (.A1(net577),
    .A2(_1772_),
    .Y(_0295_),
    .B1(_1773_));
 sg13g2_dfrbp_1 _4668_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net14),
    .D(_0131_),
    .Q_N(_2301_),
    .Q(\Pong.datapath.score_flag ));
 sg13g2_dfrbp_1 _4669_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net15),
    .D(_0000_),
    .Q_N(_0115_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[0] ));
 sg13g2_dfrbp_1 _4670_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net16),
    .D(_0010_),
    .Q_N(_2302_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[1] ));
 sg13g2_dfrbp_1 _4671_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net17),
    .D(_0011_),
    .Q_N(_0118_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[2] ));
 sg13g2_dfrbp_1 _4672_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net18),
    .D(_0012_),
    .Q_N(_2303_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ));
 sg13g2_dfrbp_1 _4673_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net19),
    .D(_0013_),
    .Q_N(_0120_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ));
 sg13g2_dfrbp_1 _4674_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net20),
    .D(_0014_),
    .Q_N(_2304_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[5] ));
 sg13g2_dfrbp_1 _4675_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net21),
    .D(_0015_),
    .Q_N(_2305_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[6] ));
 sg13g2_dfrbp_1 _4676_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net22),
    .D(_0016_),
    .Q_N(_0123_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ));
 sg13g2_dfrbp_1 _4677_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net23),
    .D(_0017_),
    .Q_N(_2306_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[8] ));
 sg13g2_dfrbp_1 _4678_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net24),
    .D(_0018_),
    .Q_N(_2307_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ));
 sg13g2_dfrbp_1 _4679_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net25),
    .D(_0001_),
    .Q_N(_2308_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[10] ));
 sg13g2_dfrbp_1 _4680_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net26),
    .D(_0002_),
    .Q_N(_2309_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[11] ));
 sg13g2_dfrbp_1 _4681_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net27),
    .D(_0003_),
    .Q_N(_0122_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ));
 sg13g2_dfrbp_1 _4682_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net28),
    .D(_0004_),
    .Q_N(_2310_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[13] ));
 sg13g2_dfrbp_1 _4683_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net29),
    .D(_0005_),
    .Q_N(_0121_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[14] ));
 sg13g2_dfrbp_1 _4684_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net30),
    .D(_0006_),
    .Q_N(_2311_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ));
 sg13g2_dfrbp_1 _4685_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net31),
    .D(_0007_),
    .Q_N(_0119_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ));
 sg13g2_dfrbp_1 _4686_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net36),
    .D(_0008_),
    .Q_N(_0117_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[17] ));
 sg13g2_dfrbp_1 _4687_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net13),
    .D(_0009_),
    .Q_N(_2300_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[18] ));
 sg13g2_dfrbp_1 _4688_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net177),
    .D(_0132_),
    .Q_N(_0052_),
    .Q(\Pong.datapath.NES_wire_Right[2] ));
 sg13g2_dfrbp_1 _4689_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net175),
    .D(_0133_),
    .Q_N(_0051_),
    .Q(\Pong.datapath.NES_wire_Left[5] ));
 sg13g2_dfrbp_1 _4690_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net173),
    .D(_0134_),
    .Q_N(_0050_),
    .Q(\Pong.datapath.NES_wire_Left[4] ));
 sg13g2_dfrbp_1 _4691_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net37),
    .D(_0135_),
    .Q_N(_0049_),
    .Q(\Pong.datapath.NES_wire_Left[3] ));
 sg13g2_dfrbp_1 _4692_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net38),
    .D(_0043_),
    .Q_N(_2312_),
    .Q(\Pong.datapath.sw_ballMovement_reg[0] ));
 sg13g2_dfrbp_1 _4693_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net39),
    .D(_0044_),
    .Q_N(_2313_),
    .Q(\Pong.datapath.sw_ballMovement_reg[2] ));
 sg13g2_dfrbp_1 _4694_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net40),
    .D(_0045_),
    .Q_N(_2314_),
    .Q(\Pong.datapath.sw_ballMovement_reg[3] ));
 sg13g2_dfrbp_1 _4695_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net41),
    .D(_0046_),
    .Q_N(_2315_),
    .Q(\Pong.datapath.sw_ballMovement_reg[4] ));
 sg13g2_dfrbp_1 _4696_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net42),
    .D(_0047_),
    .Q_N(_2316_),
    .Q(\Pong.datapath.sw_ballMovement_reg[5] ));
 sg13g2_dfrbp_1 _4697_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net43),
    .D(net404),
    .Q_N(_2317_),
    .Q(\Pong.control_unit.state_ballMovement[0] ));
 sg13g2_dfrbp_1 _4698_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net44),
    .D(net258),
    .Q_N(_2318_),
    .Q(\Pong.control_unit.state_ballMovement[1] ));
 sg13g2_dfrbp_1 _4699_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net45),
    .D(net441),
    .Q_N(_2319_),
    .Q(\Pong.control_unit.state_ballMovement[2] ));
 sg13g2_dfrbp_1 _4700_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net50),
    .D(net448),
    .Q_N(_0110_),
    .Q(\Pong.control_unit.state_ballMovement[3] ));
 sg13g2_dfrbp_1 _4701_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net171),
    .D(net420),
    .Q_N(_2299_),
    .Q(\Pong.control_unit.state_ballMovement[4] ));
 sg13g2_dfrbp_1 _4702_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net169),
    .D(_0136_),
    .Q_N(_0048_),
    .Q(\Pong.datapath.NES_wire_Left[2] ));
 sg13g2_dfrbp_1 _4703_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net167),
    .D(_0137_),
    .Q_N(_0053_),
    .Q(\Pong.datapath.NES_wire_Right[3] ));
 sg13g2_dfrbp_1 _4704_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net165),
    .D(_0138_),
    .Q_N(_0054_),
    .Q(\Pong.datapath.NES_wire_Right[4] ));
 sg13g2_dfrbp_1 _4705_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net51),
    .D(_0139_),
    .Q_N(_0055_),
    .Q(\Pong.datapath.NES_wire_Right[5] ));
 sg13g2_dfrbp_1 _4706_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net52),
    .D(net434),
    .Q_N(_0116_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[0] ));
 sg13g2_dfrbp_1 _4707_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net53),
    .D(_0029_),
    .Q_N(_2320_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ));
 sg13g2_dfrbp_1 _4708_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net54),
    .D(_0030_),
    .Q_N(_0125_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[2] ));
 sg13g2_dfrbp_1 _4709_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net55),
    .D(_0031_),
    .Q_N(_2321_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ));
 sg13g2_dfrbp_1 _4710_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net56),
    .D(_0032_),
    .Q_N(_0127_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[4] ));
 sg13g2_dfrbp_1 _4711_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net57),
    .D(_0033_),
    .Q_N(_2322_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[5] ));
 sg13g2_dfrbp_1 _4712_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net58),
    .D(_0034_),
    .Q_N(_2323_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[6] ));
 sg13g2_dfrbp_1 _4713_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net59),
    .D(_0035_),
    .Q_N(_0130_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[7] ));
 sg13g2_dfrbp_1 _4714_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net60),
    .D(_0036_),
    .Q_N(_2324_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[8] ));
 sg13g2_dfrbp_1 _4715_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net61),
    .D(_0037_),
    .Q_N(_2325_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[9] ));
 sg13g2_dfrbp_1 _4716_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net62),
    .D(net290),
    .Q_N(_2326_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[10] ));
 sg13g2_dfrbp_1 _4717_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net63),
    .D(_0021_),
    .Q_N(_2327_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[11] ));
 sg13g2_dfrbp_1 _4718_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net64),
    .D(_0022_),
    .Q_N(_0129_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[12] ));
 sg13g2_dfrbp_1 _4719_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net65),
    .D(_0023_),
    .Q_N(_2328_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[13] ));
 sg13g2_dfrbp_1 _4720_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net66),
    .D(_0024_),
    .Q_N(_0128_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[14] ));
 sg13g2_dfrbp_1 _4721_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net67),
    .D(_0025_),
    .Q_N(_2329_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ));
 sg13g2_dfrbp_1 _4722_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net68),
    .D(_0026_),
    .Q_N(_0126_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[16] ));
 sg13g2_dfrbp_1 _4723_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net186),
    .D(_0027_),
    .Q_N(_0124_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ));
 sg13g2_dfrbp_1 _4724_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net163),
    .D(_0028_),
    .Q_N(_2298_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ));
 sg13g2_dfrbp_1 _4725_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net161),
    .D(net488),
    .Q_N(_2297_),
    .Q(\Pong.datapath.scoreRight[0] ));
 sg13g2_dfrbp_1 _4726_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net160),
    .D(_0141_),
    .Q_N(_2296_),
    .Q(\Pong.datapath.scoreRight[1] ));
 sg13g2_dfrbp_1 _4727_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net159),
    .D(_0142_),
    .Q_N(_2295_),
    .Q(\Pong.datapath.scoreRight[2] ));
 sg13g2_dfrbp_1 _4728_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net158),
    .D(net427),
    .Q_N(_2294_),
    .Q(\Pong.datapath.scoreRight[3] ));
 sg13g2_dfrbp_1 _4729_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net157),
    .D(_0144_),
    .Q_N(_2293_),
    .Q(\Pong.datapath.scoreLeft[0] ));
 sg13g2_dfrbp_1 _4730_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net156),
    .D(_0145_),
    .Q_N(_2292_),
    .Q(\Pong.datapath.scoreLeft[1] ));
 sg13g2_dfrbp_1 _4731_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net155),
    .D(net423),
    .Q_N(_2291_),
    .Q(\Pong.datapath.scoreLeft[2] ));
 sg13g2_dfrbp_1 _4732_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net154),
    .D(net374),
    .Q_N(_2290_),
    .Q(\Pong.datapath.scoreLeft[3] ));
 sg13g2_dfrbp_1 _4733_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net153),
    .D(_0148_),
    .Q_N(_2289_),
    .Q(\Pong.datapath.ballFunction.reset_n ));
 sg13g2_dfrbp_1 _4734_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net152),
    .D(_0149_),
    .Q_N(_2288_),
    .Q(\Pong.datapath.rightPaddle[0] ));
 sg13g2_dfrbp_1 _4735_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net151),
    .D(_0150_),
    .Q_N(_2287_),
    .Q(\Pong.datapath.rightPaddle[1] ));
 sg13g2_dfrbp_1 _4736_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net150),
    .D(_0151_),
    .Q_N(_0077_),
    .Q(\Pong.datapath.rightPaddle[2] ));
 sg13g2_dfrbp_1 _4737_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net149),
    .D(_0152_),
    .Q_N(_0066_),
    .Q(\Pong.datapath.rightPaddle[3] ));
 sg13g2_dfrbp_1 _4738_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net148),
    .D(_0153_),
    .Q_N(_0065_),
    .Q(\Pong.datapath.rightPaddle[4] ));
 sg13g2_dfrbp_1 _4739_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net147),
    .D(_0154_),
    .Q_N(_0061_),
    .Q(\Pong.datapath.rightPaddle[5] ));
 sg13g2_dfrbp_1 _4740_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net146),
    .D(_0155_),
    .Q_N(_0060_),
    .Q(\Pong.datapath.rightPaddle[6] ));
 sg13g2_dfrbp_1 _4741_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net145),
    .D(net464),
    .Q_N(_0059_),
    .Q(\Pong.datapath.rightPaddle[7] ));
 sg13g2_dfrbp_1 _4742_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net144),
    .D(_0157_),
    .Q_N(_0058_),
    .Q(\Pong.datapath.rightPaddle[8] ));
 sg13g2_dfrbp_1 _4743_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net143),
    .D(net456),
    .Q_N(_0056_),
    .Q(\Pong.datapath.rightPaddle[9] ));
 sg13g2_dfrbp_1 _4744_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net142),
    .D(_0159_),
    .Q_N(_2286_),
    .Q(\Pong.datapath.old_NES_Right[2] ));
 sg13g2_dfrbp_1 _4745_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net141),
    .D(_0160_),
    .Q_N(_2285_),
    .Q(\Pong.datapath.old_NES_Right[3] ));
 sg13g2_dfrbp_1 _4746_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net140),
    .D(_0161_),
    .Q_N(_2284_),
    .Q(\Pong.datapath.old_NES_Right[4] ));
 sg13g2_dfrbp_1 _4747_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net139),
    .D(_0162_),
    .Q_N(_2283_),
    .Q(\Pong.datapath.old_NES_Right[5] ));
 sg13g2_dfrbp_1 _4748_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net138),
    .D(net241),
    .Q_N(_2282_),
    .Q(\Pong.datapath.NES_activity_Right[2] ));
 sg13g2_dfrbp_1 _4749_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net137),
    .D(net250),
    .Q_N(_2281_),
    .Q(\Pong.datapath.NES_activity_Right[3] ));
 sg13g2_dfrbp_1 _4750_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net136),
    .D(net237),
    .Q_N(_2280_),
    .Q(\Pong.datapath.NES_activity_Right[4] ));
 sg13g2_dfrbp_1 _4751_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net135),
    .D(net243),
    .Q_N(_0076_),
    .Q(\Pong.datapath.NES_activity_Right[5] ));
 sg13g2_dfrbp_1 _4752_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net134),
    .D(net353),
    .Q_N(_0078_),
    .Q(\Pong.datapath.leftPaddle[0] ));
 sg13g2_dfrbp_1 _4753_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net133),
    .D(net254),
    .Q_N(_0080_),
    .Q(\Pong.datapath.leftPaddle[1] ));
 sg13g2_dfrbp_1 _4754_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net132),
    .D(net511),
    .Q_N(_0079_),
    .Q(\Pong.datapath.leftPaddle[2] ));
 sg13g2_dfrbp_1 _4755_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net131),
    .D(_0170_),
    .Q_N(_0075_),
    .Q(\Pong.datapath.leftPaddle[3] ));
 sg13g2_dfrbp_1 _4756_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net130),
    .D(_0171_),
    .Q_N(_0074_),
    .Q(\Pong.datapath.leftPaddle[4] ));
 sg13g2_dfrbp_1 _4757_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net129),
    .D(net520),
    .Q_N(_0073_),
    .Q(\Pong.datapath.leftPaddle[5] ));
 sg13g2_dfrbp_1 _4758_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net128),
    .D(_0173_),
    .Q_N(_0072_),
    .Q(\Pong.datapath.leftPaddle[6] ));
 sg13g2_dfrbp_1 _4759_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net127),
    .D(net513),
    .Q_N(_0071_),
    .Q(\Pong.datapath.leftPaddle[7] ));
 sg13g2_dfrbp_1 _4760_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net126),
    .D(net532),
    .Q_N(_0070_),
    .Q(\Pong.datapath.leftPaddle[8] ));
 sg13g2_dfrbp_1 _4761_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net125),
    .D(_0176_),
    .Q_N(_0069_),
    .Q(\Pong.datapath.leftPaddle[9] ));
 sg13g2_dfrbp_1 _4762_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net124),
    .D(net248),
    .Q_N(_2279_),
    .Q(\Pong.datapath.NES_activity_Left[2] ));
 sg13g2_dfrbp_1 _4763_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net123),
    .D(net252),
    .Q_N(_2278_),
    .Q(\Pong.datapath.NES_activity_Left[3] ));
 sg13g2_dfrbp_1 _4764_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net122),
    .D(net239),
    .Q_N(_2277_),
    .Q(\Pong.datapath.NES_activity_Left[4] ));
 sg13g2_dfrbp_1 _4765_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net121),
    .D(net246),
    .Q_N(_2276_),
    .Q(\Pong.datapath.NES_activity_Left[5] ));
 sg13g2_dfrbp_1 _4766_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net120),
    .D(_0181_),
    .Q_N(_2275_),
    .Q(\Pong.datapath.old_NES_Left[2] ));
 sg13g2_dfrbp_1 _4767_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net119),
    .D(_0182_),
    .Q_N(_2274_),
    .Q(\Pong.datapath.old_NES_Left[3] ));
 sg13g2_dfrbp_1 _4768_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net118),
    .D(_0183_),
    .Q_N(_2273_),
    .Q(\Pong.datapath.old_NES_Left[4] ));
 sg13g2_dfrbp_1 _4769_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net117),
    .D(_0184_),
    .Q_N(_2272_),
    .Q(\Pong.datapath.old_NES_Left[5] ));
 sg13g2_dfrbp_1 _4770_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net116),
    .D(_0185_),
    .Q_N(_2271_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[0] ));
 sg13g2_dfrbp_1 _4771_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net114),
    .D(_0186_),
    .Q_N(_0096_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[1] ));
 sg13g2_dfrbp_1 _4772_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net112),
    .D(_0187_),
    .Q_N(_0081_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[2] ));
 sg13g2_dfrbp_1 _4773_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net110),
    .D(_0188_),
    .Q_N(_0082_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[3] ));
 sg13g2_dfrbp_1 _4774_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net108),
    .D(_0189_),
    .Q_N(_0083_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[4] ));
 sg13g2_dfrbp_1 _4775_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net106),
    .D(_0190_),
    .Q_N(_0084_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[5] ));
 sg13g2_dfrbp_1 _4776_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net104),
    .D(_0191_),
    .Q_N(_0085_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[6] ));
 sg13g2_dfrbp_1 _4777_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net102),
    .D(_0192_),
    .Q_N(_0086_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[7] ));
 sg13g2_dfrbp_1 _4778_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net100),
    .D(_0193_),
    .Q_N(_0087_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[8] ));
 sg13g2_dfrbp_1 _4779_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net98),
    .D(_0194_),
    .Q_N(_0088_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[9] ));
 sg13g2_dfrbp_1 _4780_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net96),
    .D(_0195_),
    .Q_N(_2270_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[0] ));
 sg13g2_dfrbp_1 _4781_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net94),
    .D(_0196_),
    .Q_N(_0098_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[1] ));
 sg13g2_dfrbp_1 _4782_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net92),
    .D(_0197_),
    .Q_N(_0089_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[2] ));
 sg13g2_dfrbp_1 _4783_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net90),
    .D(_0198_),
    .Q_N(_0090_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[3] ));
 sg13g2_dfrbp_1 _4784_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net88),
    .D(_0199_),
    .Q_N(_0091_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[4] ));
 sg13g2_dfrbp_1 _4785_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net86),
    .D(_0200_),
    .Q_N(_0092_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[5] ));
 sg13g2_dfrbp_1 _4786_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net84),
    .D(_0201_),
    .Q_N(_0093_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[6] ));
 sg13g2_dfrbp_1 _4787_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net82),
    .D(_0202_),
    .Q_N(_0094_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[7] ));
 sg13g2_dfrbp_1 _4788_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net80),
    .D(_0203_),
    .Q_N(_0109_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[8] ));
 sg13g2_dfrbp_1 _4789_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net78),
    .D(_0204_),
    .Q_N(_0095_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[9] ));
 sg13g2_dfrbp_1 _4790_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net76),
    .D(net474),
    .Q_N(_2269_),
    .Q(\Pong.datapath.NES_counter_left.Q[0] ));
 sg13g2_dfrbp_1 _4791_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net74),
    .D(_0206_),
    .Q_N(_2268_),
    .Q(\Pong.datapath.NES_counter_left.Q[1] ));
 sg13g2_dfrbp_1 _4792_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net72),
    .D(net319),
    .Q_N(_2267_),
    .Q(\Pong.datapath.NES_counter_left.Q[2] ));
 sg13g2_dfrbp_1 _4793_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net70),
    .D(_0208_),
    .Q_N(_2266_),
    .Q(\Pong.datapath.NES_counter_left.Q[3] ));
 sg13g2_dfrbp_1 _4794_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net49),
    .D(_0209_),
    .Q_N(_2265_),
    .Q(\Pong.datapath.NES_counter_left.Q[4] ));
 sg13g2_dfrbp_1 _4795_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net47),
    .D(_0210_),
    .Q_N(_2264_),
    .Q(\Pong.datapath.NES_counter_left.Q[5] ));
 sg13g2_dfrbp_1 _4796_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net35),
    .D(_0211_),
    .Q_N(_2263_),
    .Q(\Pong.datapath.NES_counter_left.Q[6] ));
 sg13g2_dfrbp_1 _4797_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net33),
    .D(_0212_),
    .Q_N(_2262_),
    .Q(\Pong.datapath.NES_counter_left.Q[7] ));
 sg13g2_dfrbp_1 _4798_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net12),
    .D(net484),
    .Q_N(_2261_),
    .Q(\Pong.datapath.NES_counter_right.Q[0] ));
 sg13g2_dfrbp_1 _4799_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net223),
    .D(_0214_),
    .Q_N(_2260_),
    .Q(\Pong.datapath.NES_counter_right.Q[1] ));
 sg13g2_dfrbp_1 _4800_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net221),
    .D(net359),
    .Q_N(_2259_),
    .Q(\Pong.datapath.NES_counter_right.Q[2] ));
 sg13g2_dfrbp_1 _4801_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net219),
    .D(net406),
    .Q_N(_2258_),
    .Q(\Pong.datapath.NES_counter_right.Q[3] ));
 sg13g2_dfrbp_1 _4802_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net217),
    .D(net379),
    .Q_N(_2257_),
    .Q(\Pong.datapath.NES_counter_right.Q[4] ));
 sg13g2_dfrbp_1 _4803_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net215),
    .D(_0218_),
    .Q_N(_2256_),
    .Q(\Pong.datapath.NES_counter_right.Q[5] ));
 sg13g2_dfrbp_1 _4804_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net213),
    .D(net376),
    .Q_N(_2255_),
    .Q(\Pong.datapath.NES_counter_right.Q[6] ));
 sg13g2_dfrbp_1 _4805_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net211),
    .D(net367),
    .Q_N(_2254_),
    .Q(\Pong.datapath.NES_counter_right.Q[7] ));
 sg13g2_dfrbp_1 _4806_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net209),
    .D(_0221_),
    .Q_N(_2253_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[0] ));
 sg13g2_dfrbp_1 _4807_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net207),
    .D(net288),
    .Q_N(_2252_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[1] ));
 sg13g2_dfrbp_1 _4808_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net205),
    .D(_0223_),
    .Q_N(_2251_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[2] ));
 sg13g2_dfrbp_1 _4809_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net203),
    .D(_0224_),
    .Q_N(_2250_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[3] ));
 sg13g2_dfrbp_1 _4810_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net201),
    .D(_0225_),
    .Q_N(_2249_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[4] ));
 sg13g2_dfrbp_1 _4811_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net199),
    .D(net308),
    .Q_N(_2248_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[5] ));
 sg13g2_dfrbp_1 _4812_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net197),
    .D(net327),
    .Q_N(_2247_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[6] ));
 sg13g2_dfrbp_1 _4813_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net195),
    .D(_0228_),
    .Q_N(_2246_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[7] ));
 sg13g2_dfrbp_1 _4814_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net193),
    .D(_0229_),
    .Q_N(_2245_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[8] ));
 sg13g2_dfrbp_1 _4815_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net191),
    .D(_0230_),
    .Q_N(_2244_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[9] ));
 sg13g2_dfrbp_1 _4816_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net189),
    .D(net300),
    .Q_N(_2243_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[10] ));
 sg13g2_dfrbp_1 _4817_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net187),
    .D(_0232_),
    .Q_N(_0112_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[11] ));
 sg13g2_dfrbp_1 _4818_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net185),
    .D(_0233_),
    .Q_N(_2242_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[12] ));
 sg13g2_dfrbp_1 _4819_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net183),
    .D(_0234_),
    .Q_N(_2241_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[13] ));
 sg13g2_dfrbp_1 _4820_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net181),
    .D(net461),
    .Q_N(_2240_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[14] ));
 sg13g2_dfrbp_1 _4821_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net179),
    .D(_0236_),
    .Q_N(_2239_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[15] ));
 sg13g2_dfrbp_1 _4822_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net176),
    .D(net515),
    .Q_N(_2238_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[16] ));
 sg13g2_dfrbp_1 _4823_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net172),
    .D(net350),
    .Q_N(_2237_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[17] ));
 sg13g2_dfrbp_1 _4824_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net168),
    .D(_0239_),
    .Q_N(_2236_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[18] ));
 sg13g2_dfrbp_1 _4825_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net164),
    .D(_0240_),
    .Q_N(_2235_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[0] ));
 sg13g2_dfrbp_1 _4826_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net115),
    .D(_0241_),
    .Q_N(_2234_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[1] ));
 sg13g2_dfrbp_1 _4827_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net111),
    .D(_0242_),
    .Q_N(_2233_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[2] ));
 sg13g2_dfrbp_1 _4828_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net107),
    .D(net269),
    .Q_N(_2232_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[3] ));
 sg13g2_dfrbp_1 _4829_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net103),
    .D(_0244_),
    .Q_N(_2231_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[4] ));
 sg13g2_dfrbp_1 _4830_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net99),
    .D(_0245_),
    .Q_N(_2230_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[5] ));
 sg13g2_dfrbp_1 _4831_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net95),
    .D(_0246_),
    .Q_N(_2229_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[6] ));
 sg13g2_dfrbp_1 _4832_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net91),
    .D(_0247_),
    .Q_N(_2228_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[7] ));
 sg13g2_dfrbp_1 _4833_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net87),
    .D(_0248_),
    .Q_N(_2227_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[8] ));
 sg13g2_dfrbp_1 _4834_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net83),
    .D(net364),
    .Q_N(_2226_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[9] ));
 sg13g2_dfrbp_1 _4835_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net79),
    .D(_0250_),
    .Q_N(_2225_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[10] ));
 sg13g2_dfrbp_1 _4836_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net75),
    .D(_0251_),
    .Q_N(_0111_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[11] ));
 sg13g2_dfrbp_1 _4837_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net71),
    .D(_0252_),
    .Q_N(_2224_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[12] ));
 sg13g2_dfrbp_1 _4838_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net48),
    .D(_0253_),
    .Q_N(_2223_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[13] ));
 sg13g2_dfrbp_1 _4839_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net34),
    .D(net285),
    .Q_N(_2222_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[14] ));
 sg13g2_dfrbp_1 _4840_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net224),
    .D(_0255_),
    .Q_N(_2221_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[15] ));
 sg13g2_dfrbp_1 _4841_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net220),
    .D(_0256_),
    .Q_N(_2220_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[16] ));
 sg13g2_dfrbp_1 _4842_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net216),
    .D(net329),
    .Q_N(_2219_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[17] ));
 sg13g2_dfrbp_1 _4843_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net212),
    .D(_0258_),
    .Q_N(_2218_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[18] ));
 sg13g2_dfrbp_1 _4844_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net208),
    .D(_0259_),
    .Q_N(_2217_),
    .Q(\Pong.datapath.Ball_Clock.Q[0] ));
 sg13g2_dfrbp_1 _4845_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net204),
    .D(net336),
    .Q_N(_2216_),
    .Q(\Pong.datapath.Ball_Clock.Q[1] ));
 sg13g2_dfrbp_1 _4846_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net200),
    .D(_0261_),
    .Q_N(_2215_),
    .Q(\Pong.datapath.Ball_Clock.Q[2] ));
 sg13g2_dfrbp_1 _4847_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net196),
    .D(_0262_),
    .Q_N(_2214_),
    .Q(\Pong.datapath.Ball_Clock.Q[3] ));
 sg13g2_dfrbp_1 _4848_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net192),
    .D(net332),
    .Q_N(_2213_),
    .Q(\Pong.datapath.Ball_Clock.Q[4] ));
 sg13g2_dfrbp_1 _4849_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net188),
    .D(_0264_),
    .Q_N(_2212_),
    .Q(\Pong.datapath.Ball_Clock.Q[5] ));
 sg13g2_dfrbp_1 _4850_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net184),
    .D(_0265_),
    .Q_N(_2211_),
    .Q(\Pong.datapath.Ball_Clock.Q[6] ));
 sg13g2_dfrbp_1 _4851_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net180),
    .D(_0266_),
    .Q_N(_2210_),
    .Q(\Pong.datapath.Ball_Clock.Q[7] ));
 sg13g2_dfrbp_1 _4852_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net174),
    .D(_0267_),
    .Q_N(_0114_),
    .Q(\Pong.datapath.Ball_Clock.Q[8] ));
 sg13g2_dfrbp_1 _4853_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net166),
    .D(net356),
    .Q_N(_2209_),
    .Q(\Pong.datapath.Ball_Clock.Q[9] ));
 sg13g2_dfrbp_1 _4854_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net113),
    .D(_0269_),
    .Q_N(_2208_),
    .Q(\Pong.datapath.Ball_Clock.Q[10] ));
 sg13g2_dfrbp_1 _4855_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net105),
    .D(_0270_),
    .Q_N(_2207_),
    .Q(\Pong.datapath.Ball_Clock.Q[11] ));
 sg13g2_dfrbp_1 _4856_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net97),
    .D(_0271_),
    .Q_N(_2206_),
    .Q(\Pong.datapath.Ball_Clock.Q[12] ));
 sg13g2_dfrbp_1 _4857_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net89),
    .D(net391),
    .Q_N(_2205_),
    .Q(\Pong.datapath.Ball_Clock.Q[13] ));
 sg13g2_dfrbp_1 _4858_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net81),
    .D(_0273_),
    .Q_N(_2204_),
    .Q(\Pong.datapath.Ball_Clock.Q[14] ));
 sg13g2_dfrbp_1 _4859_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net73),
    .D(_0274_),
    .Q_N(_2203_),
    .Q(\Pong.datapath.Ball_Clock.Q[15] ));
 sg13g2_dfrbp_1 _4860_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net46),
    .D(_0275_),
    .Q_N(_2202_),
    .Q(\Pong.datapath.Ball_Clock.Q[16] ));
 sg13g2_dfrbp_1 _4861_ (.CLK(net651),
    .RESET_B(net222),
    .D(_0276_),
    .Q_N(_0108_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[0] ));
 sg13g2_dfrbp_1 _4862_ (.CLK(net652),
    .RESET_B(net214),
    .D(_0277_),
    .Q_N(_2201_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[1] ));
 sg13g2_dfrbp_1 _4863_ (.CLK(net652),
    .RESET_B(net206),
    .D(_0278_),
    .Q_N(_0067_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[2] ));
 sg13g2_dfrbp_1 _4864_ (.CLK(net652),
    .RESET_B(net198),
    .D(_0279_),
    .Q_N(_0068_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[3] ));
 sg13g2_dfrbp_1 _4865_ (.CLK(net652),
    .RESET_B(net190),
    .D(_0280_),
    .Q_N(_0064_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[4] ));
 sg13g2_dfrbp_1 _4866_ (.CLK(net652),
    .RESET_B(net182),
    .D(_0281_),
    .Q_N(_0063_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[5] ));
 sg13g2_dfrbp_1 _4867_ (.CLK(net652),
    .RESET_B(net170),
    .D(_0282_),
    .Q_N(_0062_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[6] ));
 sg13g2_dfrbp_1 _4868_ (.CLK(net651),
    .RESET_B(net109),
    .D(_0283_),
    .Q_N(_0097_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[7] ));
 sg13g2_dfrbp_1 _4869_ (.CLK(net651),
    .RESET_B(net93),
    .D(_0284_),
    .Q_N(_0057_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[8] ));
 sg13g2_dfrbp_1 _4870_ (.CLK(net651),
    .RESET_B(net77),
    .D(_0285_),
    .Q_N(_0113_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[9] ));
 sg13g2_dfrbp_1 _4871_ (.CLK(net651),
    .RESET_B(net32),
    .D(_0286_),
    .Q_N(_0107_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[0] ));
 sg13g2_dfrbp_1 _4872_ (.CLK(net652),
    .RESET_B(net210),
    .D(_0287_),
    .Q_N(_2200_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[1] ));
 sg13g2_dfrbp_1 _4873_ (.CLK(net653),
    .RESET_B(net194),
    .D(_0288_),
    .Q_N(_0099_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[2] ));
 sg13g2_dfrbp_1 _4874_ (.CLK(net651),
    .RESET_B(net178),
    .D(_0289_),
    .Q_N(_0100_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[3] ));
 sg13g2_dfrbp_1 _4875_ (.CLK(net651),
    .RESET_B(net101),
    .D(_0290_),
    .Q_N(_0101_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[4] ));
 sg13g2_dfrbp_1 _4876_ (.CLK(net651),
    .RESET_B(net69),
    .D(_0291_),
    .Q_N(_0102_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[5] ));
 sg13g2_dfrbp_1 _4877_ (.CLK(net653),
    .RESET_B(net202),
    .D(_0292_),
    .Q_N(_0103_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[6] ));
 sg13g2_dfrbp_1 _4878_ (.CLK(net653),
    .RESET_B(net162),
    .D(_0293_),
    .Q_N(_0104_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[7] ));
 sg13g2_dfrbp_1 _4879_ (.CLK(net653),
    .RESET_B(net218),
    .D(_0294_),
    .Q_N(_0105_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[8] ));
 sg13g2_dfrbp_1 _4880_ (.CLK(net653),
    .RESET_B(net85),
    .D(_0295_),
    .Q_N(_0106_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[9] ));
 sg13g2_tiehi _4687__13 (.L_HI(net13));
 sg13g2_tiehi _4668__14 (.L_HI(net14));
 sg13g2_tiehi _4669__15 (.L_HI(net15));
 sg13g2_tiehi _4670__16 (.L_HI(net16));
 sg13g2_tiehi _4671__17 (.L_HI(net17));
 sg13g2_tiehi _4672__18 (.L_HI(net18));
 sg13g2_tiehi _4673__19 (.L_HI(net19));
 sg13g2_tiehi _4674__20 (.L_HI(net20));
 sg13g2_tiehi _4675__21 (.L_HI(net21));
 sg13g2_tiehi _4676__22 (.L_HI(net22));
 sg13g2_tiehi _4677__23 (.L_HI(net23));
 sg13g2_tiehi _4678__24 (.L_HI(net24));
 sg13g2_tiehi _4679__25 (.L_HI(net25));
 sg13g2_tiehi _4680__26 (.L_HI(net26));
 sg13g2_tiehi _4681__27 (.L_HI(net27));
 sg13g2_tiehi _4682__28 (.L_HI(net28));
 sg13g2_tiehi _4683__29 (.L_HI(net29));
 sg13g2_tiehi _4684__30 (.L_HI(net30));
 sg13g2_tiehi _4685__31 (.L_HI(net31));
 sg13g2_tiehi _4871__32 (.L_HI(net32));
 sg13g2_tiehi _4797__33 (.L_HI(net33));
 sg13g2_tiehi _4839__34 (.L_HI(net34));
 sg13g2_tiehi _4796__35 (.L_HI(net35));
 sg13g2_tiehi _4686__36 (.L_HI(net36));
 sg13g2_tiehi _4691__37 (.L_HI(net37));
 sg13g2_tiehi _4692__38 (.L_HI(net38));
 sg13g2_tiehi _4693__39 (.L_HI(net39));
 sg13g2_tiehi _4694__40 (.L_HI(net40));
 sg13g2_tiehi _4695__41 (.L_HI(net41));
 sg13g2_tiehi _4696__42 (.L_HI(net42));
 sg13g2_tiehi _4697__43 (.L_HI(net43));
 sg13g2_tiehi _4698__44 (.L_HI(net44));
 sg13g2_tiehi _4699__45 (.L_HI(net45));
 sg13g2_tiehi _4860__46 (.L_HI(net46));
 sg13g2_tiehi _4795__47 (.L_HI(net47));
 sg13g2_tiehi _4838__48 (.L_HI(net48));
 sg13g2_tiehi _4794__49 (.L_HI(net49));
 sg13g2_tiehi _4700__50 (.L_HI(net50));
 sg13g2_tiehi _4705__51 (.L_HI(net51));
 sg13g2_tiehi _4706__52 (.L_HI(net52));
 sg13g2_tiehi _4707__53 (.L_HI(net53));
 sg13g2_tiehi _4708__54 (.L_HI(net54));
 sg13g2_tiehi _4709__55 (.L_HI(net55));
 sg13g2_tiehi _4710__56 (.L_HI(net56));
 sg13g2_tiehi _4711__57 (.L_HI(net57));
 sg13g2_tiehi _4712__58 (.L_HI(net58));
 sg13g2_tiehi _4713__59 (.L_HI(net59));
 sg13g2_tiehi _4714__60 (.L_HI(net60));
 sg13g2_tiehi _4715__61 (.L_HI(net61));
 sg13g2_tiehi _4716__62 (.L_HI(net62));
 sg13g2_tiehi _4717__63 (.L_HI(net63));
 sg13g2_tiehi _4718__64 (.L_HI(net64));
 sg13g2_tiehi _4719__65 (.L_HI(net65));
 sg13g2_tiehi _4720__66 (.L_HI(net66));
 sg13g2_tiehi _4721__67 (.L_HI(net67));
 sg13g2_tiehi _4722__68 (.L_HI(net68));
 sg13g2_tiehi _4876__69 (.L_HI(net69));
 sg13g2_tiehi _4793__70 (.L_HI(net70));
 sg13g2_tiehi _4837__71 (.L_HI(net71));
 sg13g2_tiehi _4792__72 (.L_HI(net72));
 sg13g2_tiehi _4859__73 (.L_HI(net73));
 sg13g2_tiehi _4791__74 (.L_HI(net74));
 sg13g2_tiehi _4836__75 (.L_HI(net75));
 sg13g2_tiehi _4790__76 (.L_HI(net76));
 sg13g2_tiehi _4870__77 (.L_HI(net77));
 sg13g2_tiehi _4789__78 (.L_HI(net78));
 sg13g2_tiehi _4835__79 (.L_HI(net79));
 sg13g2_tiehi _4788__80 (.L_HI(net80));
 sg13g2_tiehi _4858__81 (.L_HI(net81));
 sg13g2_tiehi _4787__82 (.L_HI(net82));
 sg13g2_tiehi _4834__83 (.L_HI(net83));
 sg13g2_tiehi _4786__84 (.L_HI(net84));
 sg13g2_tiehi _4880__85 (.L_HI(net85));
 sg13g2_tiehi _4785__86 (.L_HI(net86));
 sg13g2_tiehi _4833__87 (.L_HI(net87));
 sg13g2_tiehi _4784__88 (.L_HI(net88));
 sg13g2_tiehi _4857__89 (.L_HI(net89));
 sg13g2_tiehi _4783__90 (.L_HI(net90));
 sg13g2_tiehi _4832__91 (.L_HI(net91));
 sg13g2_tiehi _4782__92 (.L_HI(net92));
 sg13g2_tiehi _4869__93 (.L_HI(net93));
 sg13g2_tiehi _4781__94 (.L_HI(net94));
 sg13g2_tiehi _4831__95 (.L_HI(net95));
 sg13g2_tiehi _4780__96 (.L_HI(net96));
 sg13g2_tiehi _4856__97 (.L_HI(net97));
 sg13g2_tiehi _4779__98 (.L_HI(net98));
 sg13g2_tiehi _4830__99 (.L_HI(net99));
 sg13g2_tiehi _4778__100 (.L_HI(net100));
 sg13g2_tiehi _4875__101 (.L_HI(net101));
 sg13g2_tiehi _4777__102 (.L_HI(net102));
 sg13g2_tiehi _4829__103 (.L_HI(net103));
 sg13g2_tiehi _4776__104 (.L_HI(net104));
 sg13g2_tiehi _4855__105 (.L_HI(net105));
 sg13g2_tiehi _4775__106 (.L_HI(net106));
 sg13g2_tiehi _4828__107 (.L_HI(net107));
 sg13g2_tiehi _4774__108 (.L_HI(net108));
 sg13g2_tiehi _4868__109 (.L_HI(net109));
 sg13g2_tiehi _4773__110 (.L_HI(net110));
 sg13g2_tiehi _4827__111 (.L_HI(net111));
 sg13g2_tiehi _4772__112 (.L_HI(net112));
 sg13g2_tiehi _4854__113 (.L_HI(net113));
 sg13g2_tiehi _4771__114 (.L_HI(net114));
 sg13g2_tiehi _4826__115 (.L_HI(net115));
 sg13g2_tiehi _4770__116 (.L_HI(net116));
 sg13g2_tiehi _4769__117 (.L_HI(net117));
 sg13g2_tiehi _4768__118 (.L_HI(net118));
 sg13g2_tiehi _4767__119 (.L_HI(net119));
 sg13g2_tiehi _4766__120 (.L_HI(net120));
 sg13g2_tiehi _4765__121 (.L_HI(net121));
 sg13g2_tiehi _4764__122 (.L_HI(net122));
 sg13g2_tiehi _4763__123 (.L_HI(net123));
 sg13g2_tiehi _4762__124 (.L_HI(net124));
 sg13g2_tiehi _4761__125 (.L_HI(net125));
 sg13g2_tiehi _4760__126 (.L_HI(net126));
 sg13g2_tiehi _4759__127 (.L_HI(net127));
 sg13g2_tiehi _4758__128 (.L_HI(net128));
 sg13g2_tiehi _4757__129 (.L_HI(net129));
 sg13g2_tiehi _4756__130 (.L_HI(net130));
 sg13g2_tiehi _4755__131 (.L_HI(net131));
 sg13g2_tiehi _4754__132 (.L_HI(net132));
 sg13g2_tiehi _4753__133 (.L_HI(net133));
 sg13g2_tiehi _4752__134 (.L_HI(net134));
 sg13g2_tiehi _4751__135 (.L_HI(net135));
 sg13g2_tiehi _4750__136 (.L_HI(net136));
 sg13g2_tiehi _4749__137 (.L_HI(net137));
 sg13g2_tiehi _4748__138 (.L_HI(net138));
 sg13g2_tiehi _4747__139 (.L_HI(net139));
 sg13g2_tiehi _4746__140 (.L_HI(net140));
 sg13g2_tiehi _4745__141 (.L_HI(net141));
 sg13g2_tiehi _4744__142 (.L_HI(net142));
 sg13g2_tiehi _4743__143 (.L_HI(net143));
 sg13g2_tiehi _4742__144 (.L_HI(net144));
 sg13g2_tiehi _4741__145 (.L_HI(net145));
 sg13g2_tiehi _4740__146 (.L_HI(net146));
 sg13g2_tiehi _4739__147 (.L_HI(net147));
 sg13g2_tiehi _4738__148 (.L_HI(net148));
 sg13g2_tiehi _4737__149 (.L_HI(net149));
 sg13g2_tiehi _4736__150 (.L_HI(net150));
 sg13g2_tiehi _4735__151 (.L_HI(net151));
 sg13g2_tiehi _4734__152 (.L_HI(net152));
 sg13g2_tiehi _4733__153 (.L_HI(net153));
 sg13g2_tiehi _4732__154 (.L_HI(net154));
 sg13g2_tiehi _4731__155 (.L_HI(net155));
 sg13g2_tiehi _4730__156 (.L_HI(net156));
 sg13g2_tiehi _4729__157 (.L_HI(net157));
 sg13g2_tiehi _4728__158 (.L_HI(net158));
 sg13g2_tiehi _4727__159 (.L_HI(net159));
 sg13g2_tiehi _4726__160 (.L_HI(net160));
 sg13g2_tiehi _4725__161 (.L_HI(net161));
 sg13g2_tiehi _4878__162 (.L_HI(net162));
 sg13g2_tiehi _4724__163 (.L_HI(net163));
 sg13g2_tiehi _4825__164 (.L_HI(net164));
 sg13g2_tiehi _4704__165 (.L_HI(net165));
 sg13g2_tiehi _4853__166 (.L_HI(net166));
 sg13g2_tiehi _4703__167 (.L_HI(net167));
 sg13g2_tiehi _4824__168 (.L_HI(net168));
 sg13g2_tiehi _4702__169 (.L_HI(net169));
 sg13g2_tiehi _4867__170 (.L_HI(net170));
 sg13g2_tiehi _4701__171 (.L_HI(net171));
 sg13g2_tiehi _4823__172 (.L_HI(net172));
 sg13g2_tiehi _4690__173 (.L_HI(net173));
 sg13g2_tiehi _4852__174 (.L_HI(net174));
 sg13g2_tiehi _4689__175 (.L_HI(net175));
 sg13g2_tiehi _4822__176 (.L_HI(net176));
 sg13g2_tiehi _4688__177 (.L_HI(net177));
 sg13g2_tiehi _4874__178 (.L_HI(net178));
 sg13g2_tiehi _4821__179 (.L_HI(net179));
 sg13g2_tiehi _4851__180 (.L_HI(net180));
 sg13g2_tiehi _4820__181 (.L_HI(net181));
 sg13g2_tiehi _4866__182 (.L_HI(net182));
 sg13g2_tiehi _4819__183 (.L_HI(net183));
 sg13g2_tiehi _4850__184 (.L_HI(net184));
 sg13g2_tiehi _4818__185 (.L_HI(net185));
 sg13g2_tiehi _4723__186 (.L_HI(net186));
 sg13g2_tiehi _4817__187 (.L_HI(net187));
 sg13g2_tiehi _4849__188 (.L_HI(net188));
 sg13g2_tiehi _4816__189 (.L_HI(net189));
 sg13g2_tiehi _4865__190 (.L_HI(net190));
 sg13g2_tiehi _4815__191 (.L_HI(net191));
 sg13g2_tiehi _4848__192 (.L_HI(net192));
 sg13g2_tiehi _4814__193 (.L_HI(net193));
 sg13g2_tiehi _4873__194 (.L_HI(net194));
 sg13g2_tiehi _4813__195 (.L_HI(net195));
 sg13g2_tiehi _4847__196 (.L_HI(net196));
 sg13g2_tiehi _4812__197 (.L_HI(net197));
 sg13g2_tiehi _4864__198 (.L_HI(net198));
 sg13g2_tiehi _4811__199 (.L_HI(net199));
 sg13g2_tiehi _4846__200 (.L_HI(net200));
 sg13g2_tiehi _4810__201 (.L_HI(net201));
 sg13g2_tiehi _4877__202 (.L_HI(net202));
 sg13g2_tiehi _4809__203 (.L_HI(net203));
 sg13g2_tiehi _4845__204 (.L_HI(net204));
 sg13g2_tiehi _4808__205 (.L_HI(net205));
 sg13g2_tiehi _4863__206 (.L_HI(net206));
 sg13g2_tiehi _4807__207 (.L_HI(net207));
 sg13g2_tiehi _4844__208 (.L_HI(net208));
 sg13g2_tiehi _4806__209 (.L_HI(net209));
 sg13g2_tiehi _4872__210 (.L_HI(net210));
 sg13g2_tiehi _4805__211 (.L_HI(net211));
 sg13g2_tiehi _4843__212 (.L_HI(net212));
 sg13g2_tiehi _4804__213 (.L_HI(net213));
 sg13g2_tiehi _4862__214 (.L_HI(net214));
 sg13g2_tiehi _4803__215 (.L_HI(net215));
 sg13g2_tiehi _4842__216 (.L_HI(net216));
 sg13g2_tiehi _4802__217 (.L_HI(net217));
 sg13g2_tiehi _4879__218 (.L_HI(net218));
 sg13g2_tiehi _4801__219 (.L_HI(net219));
 sg13g2_tiehi _4841__220 (.L_HI(net220));
 sg13g2_tiehi _4800__221 (.L_HI(net221));
 sg13g2_tiehi _4861__222 (.L_HI(net222));
 sg13g2_tiehi _4799__223 (.L_HI(net223));
 sg13g2_tiehi _4840__224 (.L_HI(net224));
 sg13g2_tiehi tt_um_brandonramos_VGA_Pong_with_NES_Controllers_225 (.L_HI(net225));
 sg13g2_tiehi tt_um_brandonramos_VGA_Pong_with_NES_Controllers_226 (.L_HI(net226));
 sg13g2_tiehi tt_um_brandonramos_VGA_Pong_with_NES_Controllers_227 (.L_HI(net227));
 sg13g2_tiehi tt_um_brandonramos_VGA_Pong_with_NES_Controllers_228 (.L_HI(net228));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_brandonramos_VGA_Pong_with_NES_Controllers_5 (.L_LO(net5));
 sg13g2_tielo tt_um_brandonramos_VGA_Pong_with_NES_Controllers_6 (.L_LO(net6));
 sg13g2_tielo tt_um_brandonramos_VGA_Pong_with_NES_Controllers_7 (.L_LO(net7));
 sg13g2_tielo tt_um_brandonramos_VGA_Pong_with_NES_Controllers_8 (.L_LO(net8));
 sg13g2_tielo tt_um_brandonramos_VGA_Pong_with_NES_Controllers_9 (.L_LO(net9));
 sg13g2_tielo tt_um_brandonramos_VGA_Pong_with_NES_Controllers_10 (.L_LO(net10));
 sg13g2_tielo tt_um_brandonramos_VGA_Pong_with_NES_Controllers_11 (.L_LO(net11));
 sg13g2_tiehi _4798__12 (.L_HI(net12));
 sg13g2_buf_4 _5106_ (.X(uo_out[0]),
    .A(\Pong.datapath.h_sync ));
 sg13g2_buf_4 _5107_ (.X(uo_out[1]),
    .A(\Pong.b ));
 sg13g2_buf_4 _5108_ (.X(uo_out[2]),
    .A(\Pong.b ));
 sg13g2_buf_4 _5109_ (.X(uo_out[3]),
    .A(\Pong.b ));
 sg13g2_buf_4 _5110_ (.X(uo_out[4]),
    .A(\Pong.datapath.v_sync ));
 sg13g2_buf_4 _5111_ (.X(uo_out[5]),
    .A(\Pong.b ));
 sg13g2_buf_4 _5112_ (.X(uo_out[6]),
    .A(\Pong.b ));
 sg13g2_buf_4 _5113_ (.X(uo_out[7]),
    .A(\Pong.b ));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(_1372_));
 sg13g2_buf_2 fanout572 (.A(_1250_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_1250_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_1735_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_1366_),
    .X(net575));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(_0747_));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(_1688_));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(_0725_));
 sg13g2_buf_2 fanout580 (.A(_0722_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_0719_),
    .X(net581));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(_0643_));
 sg13g2_buf_1 fanout583 (.A(_0643_),
    .X(net583));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(_0635_));
 sg13g2_buf_4 fanout585 (.X(net585),
    .A(_0630_));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(_0627_));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(_0611_));
 sg13g2_buf_2 fanout588 (.A(_0611_),
    .X(net588));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(_0609_));
 sg13g2_buf_2 fanout590 (.A(_2162_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_2150_),
    .X(net591));
 sg13g2_buf_1 fanout592 (.A(_2150_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_1951_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(\Pong.datapath.ballFunction.ball_center_x[8] ),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(\Pong.datapath.ballFunction.ball_center_x[7] ));
 sg13g2_buf_2 fanout596 (.A(\Pong.datapath.ballFunction.ball_center_x[6] ),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(\Pong.datapath.ballFunction.ball_center_x[6] ),
    .X(net597));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(\Pong.datapath.ballFunction.ball_center_x[5] ));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(_0101_));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(\Pong.datapath.ballFunction.ball_center_x[4] ));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(\Pong.datapath.ballFunction.ball_center_x[3] ));
 sg13g2_buf_1 fanout602 (.A(\Pong.datapath.ballFunction.ball_center_x[3] ),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(\Pong.datapath.ballFunction.ball_center_x[2] ));
 sg13g2_buf_2 fanout605 (.A(net607),
    .X(net605));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(\Pong.datapath.ballFunction.ball_center_x[1] ));
 sg13g2_buf_2 fanout607 (.A(\Pong.datapath.ballFunction.ball_center_x[1] ),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(\Pong.datapath.ballFunction.ball_center_y[9] ));
 sg13g2_buf_2 fanout609 (.A(\Pong.datapath.ballFunction.ball_center_y[9] ),
    .X(net609));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(net611));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(_0057_));
 sg13g2_buf_2 fanout612 (.A(net613),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(\Pong.datapath.ballFunction.ball_center_y[8] ),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(\Pong.datapath.ballFunction.ball_center_y[7] ),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_4 fanout617 (.X(net617),
    .A(_0062_));
 sg13g2_buf_4 fanout618 (.X(net618),
    .A(\Pong.datapath.ballFunction.ball_center_y[6] ));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(_0063_));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(\Pong.datapath.ballFunction.ball_center_y[5] ));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(_0064_));
 sg13g2_buf_2 fanout622 (.A(_0064_),
    .X(net622));
 sg13g2_buf_4 fanout623 (.X(net623),
    .A(\Pong.datapath.ballFunction.ball_center_y[4] ));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(\Pong.datapath.ballFunction.ball_center_y[3] ));
 sg13g2_buf_2 fanout625 (.A(net626),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(\Pong.datapath.ballFunction.ball_center_y[2] ));
 sg13g2_buf_4 fanout628 (.X(net628),
    .A(net630));
 sg13g2_buf_1 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(\Pong.datapath.ballFunction.ball_center_y[1] ));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(net632));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(\Pong.datapath.ballFunction.ball_center_y[0] ));
 sg13g2_buf_2 fanout633 (.A(net637),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_1 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_1 fanout637 (.A(_1687_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_1683_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_1435_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_1434_),
    .X(net640));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(net642));
 sg13g2_buf_2 fanout642 (.A(_1872_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_1871_),
    .X(net644));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(net647));
 sg13g2_buf_2 fanout646 (.A(net647),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_1840_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(net650),
    .X(net648));
 sg13g2_buf_1 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_1839_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_4 fanout652 (.X(net652),
    .A(\Pong.datapath.Ball_Clock.roll ));
 sg13g2_buf_2 fanout653 (.A(\Pong.datapath.Ball_Clock.roll ),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_1733_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_1826_),
    .X(net655));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(_1808_));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(_0095_));
 sg13g2_buf_2 fanout658 (.A(net659),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(\Pong.datapath.vga.Column_Counter.Q[9] ),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(net494),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(net498),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net479),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(net534),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(net503),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(net492),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net495),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(\Pong.datapath.vga.Column_Counter.Q[1] ),
    .X(net673));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net388));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_0088_));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(net525));
 sg13g2_buf_2 fanout677 (.A(\Pong.datapath.vga.Row_Counter.Q[9] ),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(_0087_));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(net524));
 sg13g2_buf_2 fanout680 (.A(\Pong.datapath.vga.Row_Counter.Q[7] ),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(\Pong.datapath.vga.Row_Counter.Q[7] ),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(_0085_));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(net505));
 sg13g2_buf_2 fanout684 (.A(\Pong.datapath.vga.Row_Counter.Q[6] ),
    .X(net684));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(_0084_));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_1 fanout687 (.A(net530),
    .X(net687));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(_0083_));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(net521),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(\Pong.datapath.vga.Row_Counter.Q[3] ));
 sg13g2_buf_8 fanout694 (.A(_0081_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(\Pong.datapath.vga.Row_Counter.Q[2] ));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(\Pong.datapath.vga.Row_Counter.Q[1] ));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(net491));
 sg13g2_buf_2 fanout699 (.A(\Pong.datapath.vga.Row_Counter.Q[0] ),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(net702),
    .X(net700));
 sg13g2_buf_1 fanout701 (.A(net702),
    .X(net701));
 sg13g2_buf_1 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net471),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(\Pong.datapath.NES_activity_Left[3] ));
 sg13g2_buf_2 fanout705 (.A(net531),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(net536));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(net509));
 sg13g2_buf_2 fanout708 (.A(net709),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(\Pong.datapath.leftPaddle[5] ),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(\Pong.datapath.leftPaddle[4] ),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(net522),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(\Pong.datapath.leftPaddle[3] ),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(\Pong.datapath.leftPaddle[2] ),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(net510),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(\Pong.datapath.leftPaddle[1] ));
 sg13g2_buf_2 fanout717 (.A(\Pong.datapath.leftPaddle[0] ),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(\Pong.datapath.leftPaddle[0] ),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net721),
    .X(net720));
 sg13g2_buf_1 fanout721 (.A(\Pong.datapath.NES_activity_Right[4] ),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net478),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net478),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(\Pong.datapath.rightPaddle[7] ),
    .X(net724));
 sg13g2_buf_1 fanout725 (.A(\Pong.datapath.rightPaddle[7] ),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(\Pong.datapath.rightPaddle[6] ));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(\Pong.datapath.rightPaddle[2] ));
 sg13g2_buf_2 fanout728 (.A(net729),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net489),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(\Pong.datapath.rightPaddle[0] ),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(\Pong.datapath.rightPaddle[0] ),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(net734),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(\Pong.datapath.ballFunction.reset_n ),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(net739),
    .X(net736));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net739));
 sg13g2_buf_4 fanout738 (.X(net738),
    .A(net739));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(_1796_));
 sg13g2_buf_2 fanout740 (.A(net741),
    .X(net740));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net742));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(_1796_));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(net744));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(net745));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(net1));
 sg13g2_buf_2 fanout746 (.A(net748),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net750),
    .X(net748));
 sg13g2_buf_4 fanout749 (.X(net749),
    .A(net750));
 sg13g2_buf_2 fanout750 (.A(net1),
    .X(net750));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_2 input2 (.A(uio_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(uio_in[3]),
    .X(net3));
 sg13g2_tielo tt_um_brandonramos_VGA_Pong_with_NES_Controllers_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0052_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0054_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0051_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0053_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0048_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0049_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0050_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold8 (.A(\Pong.datapath.old_NES_Right[4] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0165_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold10 (.A(\Pong.datapath.old_NES_Left[4] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0179_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold12 (.A(\Pong.datapath.old_NES_Right[2] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0163_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold14 (.A(\Pong.datapath.old_NES_Right[5] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0166_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0055_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold17 (.A(\Pong.datapath.old_NES_Left[5] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0180_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold19 (.A(\Pong.datapath.old_NES_Left[2] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0177_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold21 (.A(\Pong.datapath.old_NES_Right[3] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0164_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold23 (.A(\Pong.datapath.old_NES_Left[3] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0178_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0080_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0168_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold27 (.A(\Pong.datapath.NES_delay_counter_right.Q[18] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold28 (.A(_1631_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold29 (.A(\Pong.datapath.sw_ballMovement_reg[5] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0039_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold31 (.A(\Pong.datapath.NES_delay_counter_left.Q[18] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold32 (.A(_1581_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold33 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[10] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold34 (.A(_1843_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold35 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[7] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold36 (.A(_1875_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold37 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[11] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold38 (.A(_1896_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold39 (.A(\Pong.datapath.NES_delay_counter_right.Q[3] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold40 (.A(_1597_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0243_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold42 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[1] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold43 (.A(_1841_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold44 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[14] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold45 (.A(_1899_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold46 (.A(\Pong.datapath.Ball_Clock.Q[16] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold47 (.A(_1676_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold48 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[12] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold49 (.A(_1897_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold50 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[9] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold51 (.A(\Pong.datapath.NES_delay_counter_left.Q[7] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold52 (.A(_1553_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold53 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[5] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold54 (.A(_1946_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold55 (.A(\Pong.datapath.NES_delay_counter_right.Q[14] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold56 (.A(_1621_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0254_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold58 (.A(\Pong.datapath.NES_delay_counter_left.Q[1] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold59 (.A(_1543_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0222_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold61 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[10] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0020_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold63 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold64 (.A(_1941_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold65 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[11] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold66 (.A(_1847_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold67 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[14] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold68 (.A(_1864_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold69 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[5] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold70 (.A(\Pong.datapath.NES_delay_counter_left.Q[10] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold71 (.A(_1560_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0231_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold73 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold74 (.A(_1943_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold75 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold76 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[2] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1940_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold78 (.A(\Pong.datapath.NES_delay_counter_left.Q[5] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold79 (.A(_1550_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0226_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold81 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold82 (.A(_1945_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold83 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold84 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold85 (.A(_1938_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold86 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[18] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold87 (.A(\Pong.datapath.Ball_Clock.Q[6] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold88 (.A(_1649_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold89 (.A(\Pong.datapath.NES_counter_left.Q[2] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold90 (.A(_1500_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0207_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold92 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold93 (.A(_1937_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold94 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[2] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold95 (.A(_1949_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold96 (.A(\Pong.datapath.NES_delay_counter_right.Q[7] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold97 (.A(_1605_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold98 (.A(\Pong.datapath.NES_delay_counter_left.Q[6] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0227_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold100 (.A(\Pong.datapath.NES_delay_counter_right.Q[17] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0257_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold102 (.A(\Pong.datapath.Ball_Clock.Q[4] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold103 (.A(_1645_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0263_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold105 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold106 (.A(\Pong.datapath.Ball_Clock.Q[1] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold107 (.A(_1639_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0260_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold109 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[0] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold110 (.A(_1859_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold111 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[17] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold112 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[16] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold113 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[6] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold114 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold115 (.A(\Pong.datapath.Ball_Clock.Q[14] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold116 (.A(_1669_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold117 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold118 (.A(_1846_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold119 (.A(\Pong.datapath.NES_delay_counter_right.Q[12] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold120 (.A(_1618_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold121 (.A(\Pong.datapath.NES_delay_counter_left.Q[17] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0238_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold123 (.A(\Pong.datapath.Ball_Clock.Q[0] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0078_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0167_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold126 (.A(\Pong.datapath.Ball_Clock.Q[9] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold127 (.A(_1659_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0268_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold129 (.A(\Pong.datapath.NES_counter_right.Q[2] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold130 (.A(_1521_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0215_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold132 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[13] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold133 (.A(_1898_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold134 (.A(\Pong.datapath.NES_delay_counter_right.Q[9] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold135 (.A(_1610_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0249_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold137 (.A(\Pong.datapath.NES_counter_right.Q[7] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold138 (.A(_1531_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0220_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold140 (.A(\Pong.datapath.NES_delay_counter_right.Q[4] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold141 (.A(_1599_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold142 (.A(\Pong.datapath.NES_delay_counter_right.Q[0] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold143 (.A(\Pong.datapath.Ball_Clock.Q[10] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold144 (.A(_1662_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold145 (.A(\Pong.datapath.scoreLeft[3] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0147_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold147 (.A(\Pong.datapath.NES_counter_right.Q[6] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0219_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold149 (.A(\Pong.datapath.NES_counter_right.Q[4] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold150 (.A(_1526_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0217_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold152 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold153 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[8] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold154 (.A(\Pong.datapath.NES_counter_left.Q[6] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold155 (.A(_1510_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold156 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[13] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold157 (.A(\Pong.datapath.NES_delay_counter_right.Q[10] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold158 (.A(_1611_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold159 (.A(\Pong.datapath.NES_wire_Right[2] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold160 (.A(\Pong.datapath.vga.Column_Counter.Q[0] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold161 (.A(\Pong.datapath.NES_wire_Right[4] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold162 (.A(\Pong.datapath.Ball_Clock.Q[13] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0272_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold164 (.A(\Pong.datapath.NES_counter_left.Q[5] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold165 (.A(_1507_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold166 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[8] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold167 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold168 (.A(\Pong.datapath.NES_delay_counter_left.Q[11] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold169 (.A(_1567_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold170 (.A(\Pong.datapath.NES_wire_Left[5] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold171 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold172 (.A(\Pong.datapath.NES_wire_Right[3] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold173 (.A(\Pong.datapath.Ball_Clock.Q[7] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold174 (.A(\Pong.control_unit.state_ballMovement[1] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold175 (.A(_1917_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0038_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold177 (.A(\Pong.datapath.NES_counter_right.Q[3] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0216_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold179 (.A(\Pong.datapath.NES_delay_counter_right.Q[5] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold180 (.A(\Pong.datapath.NES_delay_counter_right.Q[1] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold181 (.A(\Pong.datapath.NES_delay_counter_left.Q[8] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold182 (.A(\Pong.datapath.NES_counter_left.Q[4] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold183 (.A(_1505_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0111_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold185 (.A(_1615_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0112_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold187 (.A(\Pong.datapath.NES_wire_Right[5] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold188 (.A(\Pong.datapath.Ball_Clock.Q[12] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1666_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold190 (.A(\Pong.control_unit.state_ballMovement[4] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold191 (.A(_1927_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0042_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold193 (.A(\Pong.datapath.scoreLeft[2] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold194 (.A(_1204_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0146_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold196 (.A(\Pong.datapath.NES_counter_left.Q[1] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold197 (.A(_1499_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold198 (.A(\Pong.datapath.scoreRight[3] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0143_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold200 (.A(\Pong.datapath.NES_delay_counter_left.Q[2] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold201 (.A(_1546_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold202 (.A(\Pong.datapath.NES_counter_left.Q[3] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold203 (.A(\Pong.datapath.Ball_Clock.Q[8] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold204 (.A(_1657_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold205 (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[0] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0019_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold207 (.A(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold208 (.A(_1549_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold209 (.A(\Pong.datapath.NES_delay_counter_right.Q[13] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold210 (.A(_1619_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold211 (.A(\Pong.datapath.sw_ballMovement_reg[0] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold212 (.A(_1913_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0040_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold214 (.A(\Pong.datapath.Ball_Clock.Q[3] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold215 (.A(_1644_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold216 (.A(\Pong.datapath.NES_delay_counter_left.Q[0] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold217 (.A(\Pong.datapath.NES_delay_counter_left.Q[3] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold218 (.A(\Pong.datapath.NES_counter_right.Q[5] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold219 (.A(\Pong.datapath.sw_ballMovement_reg[2] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0041_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold221 (.A(\Pong.datapath.NES_counter_right.Q[1] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold222 (.A(_1520_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold223 (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[6] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold224 (.A(_1863_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold225 (.A(\Pong.datapath.NES_delay_counter_left.Q[9] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold226 (.A(\Pong.datapath.Ball_Clock.Q[5] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0076_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0158_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold229 (.A(\Pong.datapath.NES_delay_counter_right.Q[2] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold230 (.A(\Pong.datapath.Ball_Clock.Q[11] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold231 (.A(\Pong.datapath.NES_delay_counter_left.Q[14] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold232 (.A(_1572_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0235_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold234 (.A(\Pong.datapath.NES_delay_counter_right.Q[6] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold235 (.A(\Pong.datapath.NES_activity_Right[5] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0156_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold237 (.A(\Pong.datapath.Ball_Clock.Q[2] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold238 (.A(\Pong.datapath.NES_delay_counter_right.Q[8] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold239 (.A(\Pong.datapath.NES_delay_counter_left.Q[15] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold240 (.A(_1575_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold241 (.A(\Pong.datapath.scoreRight[2] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold242 (.A(_1195_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold243 (.A(\Pong.datapath.NES_activity_Left[4] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold244 (.A(_1210_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold245 (.A(\Pong.datapath.NES_counter_left.Q[0] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0205_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0086_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold248 (.A(_1456_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold249 (.A(\Pong.datapath.NES_activity_Left[5] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold250 (.A(\Pong.datapath.NES_activity_Right[3] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold251 (.A(\Pong.datapath.vga.Column_Counter.Q[6] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold252 (.A(_1483_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold253 (.A(\Pong.datapath.scoreRight[1] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold254 (.A(\Pong.datapath.NES_counter_right.Q[0] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold255 (.A(_1518_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0213_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold257 (.A(\Pong.datapath.scoreLeft[1] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold258 (.A(_1203_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold259 (.A(\Pong.datapath.scoreRight[0] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0140_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold261 (.A(\Pong.datapath.rightPaddle[1] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold262 (.A(\Pong.datapath.Ball_Clock.Q[15] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold263 (.A(\Pong.datapath.vga.Row_Counter.Q[0] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold264 (.A(\Pong.datapath.vga.Column_Counter.Q[3] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold265 (.A(_1474_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold266 (.A(\Pong.datapath.vga.Column_Counter.Q[8] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold267 (.A(\Pong.datapath.vga.Column_Counter.Q[2] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold268 (.A(_1472_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold269 (.A(\Pong.datapath.NES_wire_Left[4] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold270 (.A(\Pong.datapath.vga.Column_Counter.Q[7] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold271 (.A(_1485_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold272 (.A(\Pong.datapath.NES_wire_Left[2] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold273 (.A(\Pong.datapath.NES_wire_Left[3] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold274 (.A(\Pong.datapath.NES_activity_Left[5] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold275 (.A(\Pong.datapath.vga.Column_Counter.Q[4] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold276 (.A(_1477_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold277 (.A(\Pong.datapath.vga.Row_Counter.Q[6] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold278 (.A(\Pong.datapath.NES_delay_counter_left.Q[13] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold279 (.A(_1571_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold280 (.A(\Pong.datapath.NES_activity_Right[2] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold281 (.A(\Pong.datapath.leftPaddle[6] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold282 (.A(\Pong.datapath.leftPaddle[2] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0169_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold284 (.A(\Pong.datapath.leftPaddle[7] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0174_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold286 (.A(\Pong.datapath.NES_delay_counter_left.Q[16] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0237_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0082_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold289 (.A(\Pong.datapath.NES_delay_counter_right.Q[16] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold290 (.A(_1625_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0073_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0172_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold293 (.A(\Pong.datapath.vga.Row_Counter.Q[4] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold294 (.A(\Pong.datapath.leftPaddle[3] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold295 (.A(\Pong.datapath.scoreLeft[0] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold296 (.A(\Pong.datapath.vga.Row_Counter.Q[8] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold297 (.A(\Pong.datapath.vga.Row_Counter.Q[9] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold298 (.A(\Pong.datapath.NES_activity_Right[5] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold299 (.A(_1078_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold300 (.A(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold301 (.A(\Pong.datapath.leftPaddle[9] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold302 (.A(\Pong.datapath.vga.Row_Counter.Q[5] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold303 (.A(\Pong.datapath.NES_activity_Left[3] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0175_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0095_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold306 (.A(\Pong.datapath.vga.Column_Counter.Q[5] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold307 (.A(_1479_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0069_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold309 (.A(\Pong.datapath.NES_delay_counter_left.Q[16] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold310 (.A(_1862_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold311 (.A(\Pong.datapath.NES_delay_counter_left.Q[3] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold312 (.A(_1853_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold313 (.A(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .X(net541));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_4 FILLER_0_196 ();
 sg13g2_fill_2 FILLER_0_204 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_fill_2 FILLER_1_126 ();
 sg13g2_fill_1 FILLER_1_128 ();
 sg13g2_decap_8 FILLER_1_134 ();
 sg13g2_decap_8 FILLER_1_141 ();
 sg13g2_decap_8 FILLER_1_148 ();
 sg13g2_decap_8 FILLER_1_155 ();
 sg13g2_decap_8 FILLER_1_162 ();
 sg13g2_decap_8 FILLER_1_169 ();
 sg13g2_decap_8 FILLER_1_176 ();
 sg13g2_decap_8 FILLER_1_183 ();
 sg13g2_decap_4 FILLER_1_190 ();
 sg13g2_fill_1 FILLER_1_194 ();
 sg13g2_fill_2 FILLER_1_221 ();
 sg13g2_fill_2 FILLER_1_228 ();
 sg13g2_decap_8 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_267 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_decap_8 FILLER_1_288 ();
 sg13g2_decap_8 FILLER_1_295 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_4 FILLER_2_112 ();
 sg13g2_fill_2 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_4 FILLER_2_172 ();
 sg13g2_fill_1 FILLER_2_176 ();
 sg13g2_fill_1 FILLER_2_203 ();
 sg13g2_fill_2 FILLER_2_209 ();
 sg13g2_fill_1 FILLER_2_211 ();
 sg13g2_decap_8 FILLER_2_253 ();
 sg13g2_decap_8 FILLER_2_260 ();
 sg13g2_decap_8 FILLER_2_267 ();
 sg13g2_decap_8 FILLER_2_274 ();
 sg13g2_decap_8 FILLER_2_281 ();
 sg13g2_decap_8 FILLER_2_288 ();
 sg13g2_decap_8 FILLER_2_295 ();
 sg13g2_decap_8 FILLER_2_302 ();
 sg13g2_decap_8 FILLER_2_309 ();
 sg13g2_decap_8 FILLER_2_316 ();
 sg13g2_decap_8 FILLER_2_323 ();
 sg13g2_decap_8 FILLER_2_330 ();
 sg13g2_decap_8 FILLER_2_337 ();
 sg13g2_decap_8 FILLER_2_344 ();
 sg13g2_decap_8 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_4 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_95 ();
 sg13g2_fill_2 FILLER_3_122 ();
 sg13g2_decap_8 FILLER_3_155 ();
 sg13g2_decap_8 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_169 ();
 sg13g2_decap_4 FILLER_3_176 ();
 sg13g2_fill_2 FILLER_3_180 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_4 FILLER_4_91 ();
 sg13g2_fill_1 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_fill_2 FILLER_4_179 ();
 sg13g2_fill_1 FILLER_4_181 ();
 sg13g2_fill_2 FILLER_4_196 ();
 sg13g2_fill_1 FILLER_4_198 ();
 sg13g2_fill_2 FILLER_4_207 ();
 sg13g2_fill_1 FILLER_4_217 ();
 sg13g2_fill_2 FILLER_4_223 ();
 sg13g2_fill_1 FILLER_4_231 ();
 sg13g2_fill_2 FILLER_4_254 ();
 sg13g2_fill_1 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_262 ();
 sg13g2_decap_8 FILLER_4_269 ();
 sg13g2_decap_8 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_fill_2 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_fill_2 FILLER_5_91 ();
 sg13g2_fill_2 FILLER_5_129 ();
 sg13g2_fill_2 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_173 ();
 sg13g2_fill_2 FILLER_5_180 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_189 ();
 sg13g2_fill_1 FILLER_5_198 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_8 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_fill_2 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_fill_1 FILLER_5_298 ();
 sg13g2_fill_1 FILLER_5_313 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_98 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_2 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_fill_1 FILLER_6_207 ();
 sg13g2_fill_2 FILLER_6_212 ();
 sg13g2_decap_8 FILLER_6_219 ();
 sg13g2_decap_4 FILLER_6_226 ();
 sg13g2_fill_2 FILLER_6_236 ();
 sg13g2_fill_2 FILLER_6_243 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_fill_2 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_159 ();
 sg13g2_fill_1 FILLER_7_186 ();
 sg13g2_fill_2 FILLER_7_207 ();
 sg13g2_fill_1 FILLER_7_209 ();
 sg13g2_fill_2 FILLER_7_215 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_fill_2 FILLER_7_235 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_fill_2 FILLER_7_280 ();
 sg13g2_fill_1 FILLER_7_310 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_369 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_98 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_fill_1 FILLER_8_162 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_fill_1 FILLER_8_218 ();
 sg13g2_fill_1 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_252 ();
 sg13g2_decap_4 FILLER_8_266 ();
 sg13g2_fill_1 FILLER_8_270 ();
 sg13g2_fill_1 FILLER_8_297 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_fill_2 FILLER_9_124 ();
 sg13g2_fill_1 FILLER_9_126 ();
 sg13g2_fill_2 FILLER_9_136 ();
 sg13g2_fill_1 FILLER_9_138 ();
 sg13g2_fill_2 FILLER_9_164 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_175 ();
 sg13g2_fill_1 FILLER_9_177 ();
 sg13g2_fill_2 FILLER_9_191 ();
 sg13g2_fill_1 FILLER_9_193 ();
 sg13g2_fill_2 FILLER_9_200 ();
 sg13g2_fill_1 FILLER_9_202 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_224 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_fill_2 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_235 ();
 sg13g2_fill_2 FILLER_9_252 ();
 sg13g2_decap_4 FILLER_9_275 ();
 sg13g2_fill_2 FILLER_9_279 ();
 sg13g2_fill_2 FILLER_9_293 ();
 sg13g2_fill_1 FILLER_9_295 ();
 sg13g2_fill_2 FILLER_9_306 ();
 sg13g2_fill_1 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_fill_2 FILLER_10_98 ();
 sg13g2_fill_1 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_118 ();
 sg13g2_fill_2 FILLER_10_129 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_fill_1 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_213 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_fill_1 FILLER_10_221 ();
 sg13g2_fill_2 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_250 ();
 sg13g2_fill_1 FILLER_10_256 ();
 sg13g2_fill_2 FILLER_10_272 ();
 sg13g2_fill_1 FILLER_10_304 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_fill_1 FILLER_10_312 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_fill_2 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_180 ();
 sg13g2_fill_2 FILLER_11_187 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_decap_4 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_fill_2 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_239 ();
 sg13g2_decap_4 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_265 ();
 sg13g2_decap_8 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_279 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_fill_1 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_fill_2 FILLER_12_105 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_fill_2 FILLER_12_206 ();
 sg13g2_fill_2 FILLER_12_251 ();
 sg13g2_decap_4 FILLER_12_275 ();
 sg13g2_fill_1 FILLER_12_279 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_fill_1 FILLER_12_332 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_fill_2 FILLER_13_187 ();
 sg13g2_fill_1 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_fill_2 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_227 ();
 sg13g2_fill_2 FILLER_13_243 ();
 sg13g2_fill_1 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_278 ();
 sg13g2_decap_4 FILLER_13_285 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_4 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_209 ();
 sg13g2_fill_2 FILLER_14_215 ();
 sg13g2_decap_4 FILLER_14_222 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_fill_2 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_288 ();
 sg13g2_decap_8 FILLER_14_295 ();
 sg13g2_fill_2 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_4 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_129 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_171 ();
 sg13g2_fill_1 FILLER_15_173 ();
 sg13g2_decap_8 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_228 ();
 sg13g2_fill_2 FILLER_15_235 ();
 sg13g2_fill_2 FILLER_15_247 ();
 sg13g2_decap_4 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_257 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_fill_2 FILLER_15_270 ();
 sg13g2_fill_1 FILLER_15_272 ();
 sg13g2_decap_4 FILLER_15_299 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_decap_4 FILLER_15_320 ();
 sg13g2_decap_4 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_fill_1 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_decap_4 FILLER_16_142 ();
 sg13g2_fill_1 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_213 ();
 sg13g2_fill_1 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_fill_2 FILLER_16_265 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_325 ();
 sg13g2_fill_2 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_fill_2 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_114 ();
 sg13g2_decap_4 FILLER_17_157 ();
 sg13g2_decap_4 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_174 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_fill_2 FILLER_17_205 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_fill_2 FILLER_17_318 ();
 sg13g2_fill_1 FILLER_17_320 ();
 sg13g2_fill_2 FILLER_17_326 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_fill_2 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_decap_4 FILLER_18_326 ();
 sg13g2_fill_2 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_fill_2 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_170 ();
 sg13g2_decap_8 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_decap_4 FILLER_19_206 ();
 sg13g2_fill_2 FILLER_19_262 ();
 sg13g2_fill_1 FILLER_19_264 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_decap_4 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_341 ();
 sg13g2_decap_4 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_119 ();
 sg13g2_fill_2 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_174 ();
 sg13g2_decap_4 FILLER_20_181 ();
 sg13g2_fill_2 FILLER_20_185 ();
 sg13g2_decap_8 FILLER_20_195 ();
 sg13g2_fill_2 FILLER_20_202 ();
 sg13g2_fill_1 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_fill_2 FILLER_20_242 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_275 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_4 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_decap_4 FILLER_21_211 ();
 sg13g2_decap_4 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_4 FILLER_21_249 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_273 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_fill_2 FILLER_21_363 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_4 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_decap_4 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_decap_4 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_decap_4 FILLER_22_310 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_324 ();
 sg13g2_decap_4 FILLER_22_334 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_fill_2 FILLER_22_354 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_4 FILLER_23_126 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_4 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_302 ();
 sg13g2_decap_4 FILLER_23_330 ();
 sg13g2_decap_4 FILLER_23_352 ();
 sg13g2_fill_2 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_128 ();
 sg13g2_fill_2 FILLER_24_146 ();
 sg13g2_fill_2 FILLER_24_156 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_decap_4 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_251 ();
 sg13g2_fill_2 FILLER_24_284 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_decap_4 FILLER_24_310 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_357 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_126 ();
 sg13g2_fill_1 FILLER_25_128 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_192 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_decap_4 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_336 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_fill_2 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_fill_2 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_4 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_241 ();
 sg13g2_decap_8 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_fill_1 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_decap_4 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_fill_2 FILLER_26_298 ();
 sg13g2_fill_1 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_fill_2 FILLER_26_344 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_fill_2 FILLER_26_352 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_220 ();
 sg13g2_decap_8 FILLER_27_227 ();
 sg13g2_decap_4 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_decap_8 FILLER_27_271 ();
 sg13g2_decap_8 FILLER_27_278 ();
 sg13g2_decap_8 FILLER_27_285 ();
 sg13g2_decap_8 FILLER_27_292 ();
 sg13g2_decap_4 FILLER_27_299 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_decap_4 FILLER_27_327 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_decap_4 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_decap_4 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_fill_2 FILLER_27_374 ();
 sg13g2_fill_1 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_decap_4 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_fill_1 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_357 ();
 sg13g2_fill_2 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_4 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_166 ();
 sg13g2_fill_1 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_decap_4 FILLER_29_265 ();
 sg13g2_fill_2 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_decap_4 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_370 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_decap_4 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_290 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_fill_2 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_4 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_341 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_fill_2 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_4 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_251 ();
 sg13g2_decap_4 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_278 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_decap_4 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_32_323 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_196 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_decap_4 FILLER_33_300 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_decap_4 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_fill_2 FILLER_34_143 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_decap_4 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_309 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_357 ();
 sg13g2_decap_4 FILLER_34_365 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_4 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_decap_4 FILLER_35_347 ();
 sg13g2_decap_8 FILLER_35_356 ();
 sg13g2_decap_8 FILLER_35_363 ();
 sg13g2_decap_4 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_74 ();
 sg13g2_decap_8 FILLER_36_81 ();
 sg13g2_decap_8 FILLER_36_88 ();
 sg13g2_decap_4 FILLER_36_95 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_2 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_fill_2 FILLER_36_211 ();
 sg13g2_fill_1 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_decap_4 FILLER_36_362 ();
 sg13g2_fill_2 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_85 ();
 sg13g2_decap_8 FILLER_37_92 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_fill_2 FILLER_37_106 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_fill_1 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_fill_2 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_4 FILLER_37_298 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_decap_4 FILLER_37_318 ();
 sg13g2_fill_2 FILLER_37_322 ();
 sg13g2_decap_4 FILLER_37_328 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_71 ();
 sg13g2_decap_8 FILLER_38_94 ();
 sg13g2_decap_4 FILLER_38_101 ();
 sg13g2_decap_4 FILLER_38_109 ();
 sg13g2_fill_2 FILLER_38_113 ();
 sg13g2_fill_2 FILLER_38_154 ();
 sg13g2_fill_2 FILLER_38_191 ();
 sg13g2_fill_2 FILLER_38_203 ();
 sg13g2_fill_1 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_decap_4 FILLER_38_238 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_253 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_305 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_362 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_55 ();
 sg13g2_decap_4 FILLER_39_88 ();
 sg13g2_fill_1 FILLER_39_92 ();
 sg13g2_fill_2 FILLER_39_201 ();
 sg13g2_fill_1 FILLER_39_203 ();
 sg13g2_fill_2 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_270 ();
 sg13g2_fill_1 FILLER_39_272 ();
 sg13g2_fill_2 FILLER_39_353 ();
 sg13g2_fill_2 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_4 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_194 ();
 sg13g2_fill_2 FILLER_40_211 ();
 sg13g2_fill_1 FILLER_40_228 ();
 sg13g2_fill_1 FILLER_40_235 ();
 sg13g2_fill_2 FILLER_40_323 ();
 sg13g2_fill_2 FILLER_40_333 ();
 sg13g2_fill_1 FILLER_40_340 ();
 sg13g2_fill_2 FILLER_40_366 ();
 sg13g2_fill_2 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_374 ();
 sg13g2_decap_8 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_398 ();
 sg13g2_decap_4 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_47 ();
 sg13g2_fill_1 FILLER_41_57 ();
 sg13g2_decap_8 FILLER_41_76 ();
 sg13g2_decap_4 FILLER_41_83 ();
 sg13g2_fill_2 FILLER_41_87 ();
 sg13g2_fill_1 FILLER_41_135 ();
 sg13g2_fill_2 FILLER_41_154 ();
 sg13g2_fill_2 FILLER_41_206 ();
 sg13g2_decap_8 FILLER_41_229 ();
 sg13g2_fill_2 FILLER_41_236 ();
 sg13g2_fill_1 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_256 ();
 sg13g2_decap_8 FILLER_41_271 ();
 sg13g2_fill_2 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_285 ();
 sg13g2_fill_2 FILLER_41_336 ();
 sg13g2_fill_2 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_345 ();
 sg13g2_fill_2 FILLER_41_368 ();
 sg13g2_fill_1 FILLER_41_370 ();
 sg13g2_decap_8 FILLER_41_387 ();
 sg13g2_decap_8 FILLER_41_394 ();
 sg13g2_decap_8 FILLER_41_401 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_21 ();
 sg13g2_fill_1 FILLER_42_23 ();
 sg13g2_fill_1 FILLER_42_55 ();
 sg13g2_fill_2 FILLER_42_65 ();
 sg13g2_fill_1 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_72 ();
 sg13g2_fill_2 FILLER_42_79 ();
 sg13g2_fill_2 FILLER_42_111 ();
 sg13g2_fill_2 FILLER_42_150 ();
 sg13g2_decap_8 FILLER_42_172 ();
 sg13g2_decap_8 FILLER_42_179 ();
 sg13g2_decap_4 FILLER_42_186 ();
 sg13g2_decap_8 FILLER_42_195 ();
 sg13g2_decap_8 FILLER_42_202 ();
 sg13g2_decap_4 FILLER_42_209 ();
 sg13g2_decap_8 FILLER_42_222 ();
 sg13g2_decap_8 FILLER_42_229 ();
 sg13g2_decap_4 FILLER_42_236 ();
 sg13g2_fill_2 FILLER_42_240 ();
 sg13g2_fill_2 FILLER_42_246 ();
 sg13g2_decap_4 FILLER_42_253 ();
 sg13g2_decap_8 FILLER_42_263 ();
 sg13g2_decap_8 FILLER_42_270 ();
 sg13g2_fill_2 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_fill_2 FILLER_42_301 ();
 sg13g2_fill_1 FILLER_42_303 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_fill_1 FILLER_42_327 ();
 sg13g2_fill_2 FILLER_42_337 ();
 sg13g2_fill_1 FILLER_42_351 ();
 sg13g2_fill_1 FILLER_42_365 ();
 sg13g2_decap_8 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_4 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_4 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_84 ();
 sg13g2_fill_1 FILLER_43_127 ();
 sg13g2_fill_2 FILLER_43_133 ();
 sg13g2_fill_1 FILLER_43_140 ();
 sg13g2_fill_2 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_165 ();
 sg13g2_decap_4 FILLER_43_174 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_4 FILLER_43_189 ();
 sg13g2_fill_2 FILLER_43_193 ();
 sg13g2_decap_4 FILLER_43_199 ();
 sg13g2_fill_2 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_fill_2 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_fill_2 FILLER_43_238 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_fill_1 FILLER_43_274 ();
 sg13g2_decap_8 FILLER_43_291 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_decap_8 FILLER_43_305 ();
 sg13g2_fill_2 FILLER_43_312 ();
 sg13g2_fill_1 FILLER_43_314 ();
 sg13g2_decap_8 FILLER_43_323 ();
 sg13g2_decap_8 FILLER_43_330 ();
 sg13g2_decap_8 FILLER_43_337 ();
 sg13g2_fill_1 FILLER_43_344 ();
 sg13g2_fill_1 FILLER_43_349 ();
 sg13g2_fill_2 FILLER_43_354 ();
 sg13g2_decap_8 FILLER_43_361 ();
 sg13g2_fill_1 FILLER_43_368 ();
 sg13g2_decap_8 FILLER_43_373 ();
 sg13g2_decap_8 FILLER_43_380 ();
 sg13g2_decap_8 FILLER_43_387 ();
 sg13g2_decap_8 FILLER_43_394 ();
 sg13g2_decap_8 FILLER_43_401 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_9 ();
 sg13g2_fill_2 FILLER_44_36 ();
 sg13g2_fill_2 FILLER_44_115 ();
 sg13g2_fill_1 FILLER_44_117 ();
 sg13g2_fill_1 FILLER_44_151 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_fill_2 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_257 ();
 sg13g2_fill_2 FILLER_44_265 ();
 sg13g2_fill_1 FILLER_44_267 ();
 sg13g2_fill_2 FILLER_44_276 ();
 sg13g2_decap_4 FILLER_44_298 ();
 sg13g2_fill_2 FILLER_44_302 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_decap_4 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_342 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_355 ();
 sg13g2_decap_8 FILLER_44_362 ();
 sg13g2_fill_2 FILLER_44_369 ();
 sg13g2_fill_1 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_381 ();
 sg13g2_decap_8 FILLER_44_388 ();
 sg13g2_decap_8 FILLER_44_395 ();
 sg13g2_decap_8 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_11 ();
 sg13g2_fill_2 FILLER_45_50 ();
 sg13g2_fill_1 FILLER_45_90 ();
 sg13g2_fill_1 FILLER_45_193 ();
 sg13g2_fill_2 FILLER_45_209 ();
 sg13g2_fill_2 FILLER_45_222 ();
 sg13g2_fill_2 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_261 ();
 sg13g2_fill_1 FILLER_45_263 ();
 sg13g2_fill_2 FILLER_45_271 ();
 sg13g2_fill_1 FILLER_45_273 ();
 sg13g2_fill_1 FILLER_45_292 ();
 sg13g2_fill_2 FILLER_45_348 ();
 sg13g2_fill_1 FILLER_45_350 ();
 sg13g2_fill_2 FILLER_45_377 ();
 sg13g2_fill_1 FILLER_45_379 ();
 sg13g2_decap_8 FILLER_45_384 ();
 sg13g2_decap_8 FILLER_45_391 ();
 sg13g2_decap_8 FILLER_45_398 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_9 ();
 sg13g2_fill_2 FILLER_46_51 ();
 sg13g2_fill_2 FILLER_46_96 ();
 sg13g2_fill_2 FILLER_46_169 ();
 sg13g2_fill_2 FILLER_46_180 ();
 sg13g2_fill_2 FILLER_46_229 ();
 sg13g2_fill_1 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_332 ();
 sg13g2_fill_2 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_391 ();
 sg13g2_decap_8 FILLER_46_398 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_60 ();
 sg13g2_fill_1 FILLER_47_130 ();
 sg13g2_fill_2 FILLER_47_174 ();
 sg13g2_fill_1 FILLER_47_199 ();
 sg13g2_fill_1 FILLER_47_208 ();
 sg13g2_fill_2 FILLER_47_214 ();
 sg13g2_fill_1 FILLER_47_216 ();
 sg13g2_fill_2 FILLER_47_242 ();
 sg13g2_decap_8 FILLER_47_263 ();
 sg13g2_decap_8 FILLER_47_270 ();
 sg13g2_decap_8 FILLER_47_277 ();
 sg13g2_decap_8 FILLER_47_284 ();
 sg13g2_decap_4 FILLER_47_291 ();
 sg13g2_decap_8 FILLER_47_299 ();
 sg13g2_fill_1 FILLER_47_306 ();
 sg13g2_fill_2 FILLER_47_327 ();
 sg13g2_fill_1 FILLER_47_329 ();
 sg13g2_fill_2 FILLER_47_377 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_fill_2 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_1 FILLER_48_29 ();
 sg13g2_fill_1 FILLER_48_51 ();
 sg13g2_fill_2 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_228 ();
 sg13g2_decap_4 FILLER_48_235 ();
 sg13g2_fill_2 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_258 ();
 sg13g2_decap_8 FILLER_48_267 ();
 sg13g2_decap_4 FILLER_48_286 ();
 sg13g2_fill_1 FILLER_48_290 ();
 sg13g2_fill_2 FILLER_48_317 ();
 sg13g2_decap_8 FILLER_48_333 ();
 sg13g2_decap_8 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_347 ();
 sg13g2_decap_8 FILLER_48_352 ();
 sg13g2_fill_1 FILLER_48_359 ();
 sg13g2_fill_2 FILLER_48_370 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_28 ();
 sg13g2_fill_1 FILLER_49_70 ();
 sg13g2_fill_1 FILLER_49_85 ();
 sg13g2_fill_2 FILLER_49_141 ();
 sg13g2_fill_1 FILLER_49_143 ();
 sg13g2_fill_2 FILLER_49_165 ();
 sg13g2_fill_1 FILLER_49_167 ();
 sg13g2_fill_2 FILLER_49_178 ();
 sg13g2_fill_2 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_218 ();
 sg13g2_decap_8 FILLER_49_225 ();
 sg13g2_decap_8 FILLER_49_232 ();
 sg13g2_decap_8 FILLER_49_239 ();
 sg13g2_decap_8 FILLER_49_246 ();
 sg13g2_fill_1 FILLER_49_253 ();
 sg13g2_fill_2 FILLER_49_272 ();
 sg13g2_decap_4 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_338 ();
 sg13g2_fill_2 FILLER_49_362 ();
 sg13g2_fill_1 FILLER_49_364 ();
 sg13g2_fill_1 FILLER_49_369 ();
 sg13g2_decap_8 FILLER_49_388 ();
 sg13g2_decap_8 FILLER_49_395 ();
 sg13g2_decap_8 FILLER_49_402 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_4 ();
 sg13g2_fill_2 FILLER_50_50 ();
 sg13g2_fill_1 FILLER_50_71 ();
 sg13g2_fill_2 FILLER_50_89 ();
 sg13g2_fill_1 FILLER_50_91 ();
 sg13g2_fill_1 FILLER_50_118 ();
 sg13g2_fill_1 FILLER_50_150 ();
 sg13g2_fill_2 FILLER_50_159 ();
 sg13g2_fill_1 FILLER_50_196 ();
 sg13g2_fill_1 FILLER_50_204 ();
 sg13g2_decap_4 FILLER_50_214 ();
 sg13g2_decap_8 FILLER_50_222 ();
 sg13g2_decap_8 FILLER_50_229 ();
 sg13g2_decap_8 FILLER_50_236 ();
 sg13g2_fill_1 FILLER_50_270 ();
 sg13g2_fill_1 FILLER_50_301 ();
 sg13g2_fill_2 FILLER_50_306 ();
 sg13g2_decap_8 FILLER_50_312 ();
 sg13g2_fill_1 FILLER_50_341 ();
 sg13g2_decap_8 FILLER_50_368 ();
 sg13g2_decap_8 FILLER_50_387 ();
 sg13g2_decap_8 FILLER_50_394 ();
 sg13g2_decap_8 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_27 ();
 sg13g2_fill_1 FILLER_51_59 ();
 sg13g2_fill_2 FILLER_51_86 ();
 sg13g2_fill_1 FILLER_51_88 ();
 sg13g2_decap_4 FILLER_51_158 ();
 sg13g2_fill_2 FILLER_51_162 ();
 sg13g2_fill_1 FILLER_51_181 ();
 sg13g2_decap_4 FILLER_51_232 ();
 sg13g2_fill_2 FILLER_51_236 ();
 sg13g2_fill_1 FILLER_51_266 ();
 sg13g2_fill_1 FILLER_51_287 ();
 sg13g2_fill_2 FILLER_51_292 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_388 ();
 sg13g2_decap_8 FILLER_51_395 ();
 sg13g2_decap_8 FILLER_51_402 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_27 ();
 sg13g2_fill_1 FILLER_52_44 ();
 sg13g2_fill_2 FILLER_52_80 ();
 sg13g2_fill_1 FILLER_52_117 ();
 sg13g2_fill_1 FILLER_52_137 ();
 sg13g2_decap_8 FILLER_52_164 ();
 sg13g2_fill_2 FILLER_52_195 ();
 sg13g2_fill_2 FILLER_52_205 ();
 sg13g2_decap_4 FILLER_52_239 ();
 sg13g2_fill_2 FILLER_52_243 ();
 sg13g2_decap_4 FILLER_52_260 ();
 sg13g2_fill_2 FILLER_52_272 ();
 sg13g2_fill_1 FILLER_52_274 ();
 sg13g2_fill_2 FILLER_52_280 ();
 sg13g2_fill_1 FILLER_52_282 ();
 sg13g2_decap_8 FILLER_52_292 ();
 sg13g2_decap_8 FILLER_52_299 ();
 sg13g2_decap_8 FILLER_52_310 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_fill_1 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_fill_1 FILLER_52_350 ();
 sg13g2_decap_4 FILLER_52_369 ();
 sg13g2_fill_1 FILLER_52_373 ();
 sg13g2_fill_1 FILLER_52_379 ();
 sg13g2_decap_8 FILLER_52_384 ();
 sg13g2_decap_8 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_398 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_fill_2 FILLER_53_47 ();
 sg13g2_fill_1 FILLER_53_49 ();
 sg13g2_fill_1 FILLER_53_55 ();
 sg13g2_fill_2 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_126 ();
 sg13g2_fill_1 FILLER_53_141 ();
 sg13g2_fill_1 FILLER_53_200 ();
 sg13g2_fill_2 FILLER_53_206 ();
 sg13g2_decap_4 FILLER_53_238 ();
 sg13g2_decap_8 FILLER_53_258 ();
 sg13g2_decap_4 FILLER_53_265 ();
 sg13g2_fill_1 FILLER_53_277 ();
 sg13g2_decap_8 FILLER_53_303 ();
 sg13g2_fill_1 FILLER_53_310 ();
 sg13g2_decap_8 FILLER_53_342 ();
 sg13g2_decap_8 FILLER_53_349 ();
 sg13g2_fill_2 FILLER_53_356 ();
 sg13g2_decap_8 FILLER_53_362 ();
 sg13g2_fill_1 FILLER_53_369 ();
 sg13g2_decap_8 FILLER_53_390 ();
 sg13g2_decap_8 FILLER_53_397 ();
 sg13g2_decap_4 FILLER_53_404 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_fill_1 FILLER_54_103 ();
 sg13g2_fill_1 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_187 ();
 sg13g2_fill_2 FILLER_54_230 ();
 sg13g2_decap_8 FILLER_54_270 ();
 sg13g2_fill_1 FILLER_54_277 ();
 sg13g2_fill_1 FILLER_54_297 ();
 sg13g2_fill_2 FILLER_54_313 ();
 sg13g2_fill_1 FILLER_54_315 ();
 sg13g2_fill_1 FILLER_54_327 ();
 sg13g2_fill_1 FILLER_54_336 ();
 sg13g2_decap_4 FILLER_54_358 ();
 sg13g2_fill_1 FILLER_54_362 ();
 sg13g2_decap_8 FILLER_54_402 ();
 sg13g2_fill_2 FILLER_55_42 ();
 sg13g2_fill_1 FILLER_55_58 ();
 sg13g2_fill_1 FILLER_55_74 ();
 sg13g2_fill_2 FILLER_55_189 ();
 sg13g2_fill_1 FILLER_55_191 ();
 sg13g2_fill_2 FILLER_55_224 ();
 sg13g2_fill_1 FILLER_55_226 ();
 sg13g2_decap_4 FILLER_55_321 ();
 sg13g2_fill_1 FILLER_55_325 ();
 sg13g2_decap_4 FILLER_55_362 ();
 sg13g2_fill_1 FILLER_55_366 ();
 sg13g2_fill_1 FILLER_55_372 ();
 sg13g2_decap_8 FILLER_55_390 ();
 sg13g2_decap_8 FILLER_55_397 ();
 sg13g2_decap_4 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_15 ();
 sg13g2_fill_1 FILLER_56_17 ();
 sg13g2_fill_1 FILLER_56_65 ();
 sg13g2_fill_2 FILLER_56_78 ();
 sg13g2_fill_1 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_119 ();
 sg13g2_fill_1 FILLER_56_121 ();
 sg13g2_fill_2 FILLER_56_137 ();
 sg13g2_fill_1 FILLER_56_191 ();
 sg13g2_decap_8 FILLER_56_227 ();
 sg13g2_fill_2 FILLER_56_234 ();
 sg13g2_fill_2 FILLER_56_245 ();
 sg13g2_fill_1 FILLER_56_260 ();
 sg13g2_decap_4 FILLER_56_283 ();
 sg13g2_fill_2 FILLER_56_287 ();
 sg13g2_fill_2 FILLER_56_312 ();
 sg13g2_fill_2 FILLER_56_322 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_decap_8 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_decap_8 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_1 FILLER_57_38 ();
 sg13g2_fill_1 FILLER_57_113 ();
 sg13g2_fill_2 FILLER_57_147 ();
 sg13g2_fill_2 FILLER_57_165 ();
 sg13g2_fill_2 FILLER_57_184 ();
 sg13g2_fill_1 FILLER_57_186 ();
 sg13g2_fill_1 FILLER_57_205 ();
 sg13g2_decap_8 FILLER_57_237 ();
 sg13g2_fill_2 FILLER_57_248 ();
 sg13g2_fill_1 FILLER_57_250 ();
 sg13g2_decap_4 FILLER_57_289 ();
 sg13g2_fill_2 FILLER_57_293 ();
 sg13g2_decap_8 FILLER_57_299 ();
 sg13g2_decap_8 FILLER_57_306 ();
 sg13g2_fill_2 FILLER_57_313 ();
 sg13g2_decap_8 FILLER_57_318 ();
 sg13g2_decap_4 FILLER_57_325 ();
 sg13g2_fill_2 FILLER_57_329 ();
 sg13g2_decap_4 FILLER_57_345 ();
 sg13g2_fill_2 FILLER_57_349 ();
 sg13g2_decap_4 FILLER_57_355 ();
 sg13g2_fill_2 FILLER_57_359 ();
 sg13g2_decap_8 FILLER_57_379 ();
 sg13g2_decap_8 FILLER_57_386 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_51 ();
 sg13g2_fill_1 FILLER_58_79 ();
 sg13g2_fill_2 FILLER_58_85 ();
 sg13g2_fill_2 FILLER_58_125 ();
 sg13g2_decap_4 FILLER_58_166 ();
 sg13g2_fill_1 FILLER_58_170 ();
 sg13g2_decap_4 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_179 ();
 sg13g2_fill_2 FILLER_58_206 ();
 sg13g2_fill_1 FILLER_58_208 ();
 sg13g2_decap_4 FILLER_58_235 ();
 sg13g2_fill_2 FILLER_58_239 ();
 sg13g2_fill_2 FILLER_58_252 ();
 sg13g2_fill_1 FILLER_58_254 ();
 sg13g2_fill_2 FILLER_58_266 ();
 sg13g2_fill_2 FILLER_58_272 ();
 sg13g2_fill_1 FILLER_58_274 ();
 sg13g2_decap_8 FILLER_58_279 ();
 sg13g2_decap_4 FILLER_58_286 ();
 sg13g2_fill_2 FILLER_58_290 ();
 sg13g2_decap_4 FILLER_58_305 ();
 sg13g2_fill_2 FILLER_58_309 ();
 sg13g2_fill_1 FILLER_58_346 ();
 sg13g2_fill_1 FILLER_58_351 ();
 sg13g2_decap_4 FILLER_58_359 ();
 sg13g2_fill_1 FILLER_58_363 ();
 sg13g2_fill_2 FILLER_58_369 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_1 FILLER_59_26 ();
 sg13g2_fill_2 FILLER_59_31 ();
 sg13g2_fill_1 FILLER_59_39 ();
 sg13g2_fill_1 FILLER_59_66 ();
 sg13g2_fill_2 FILLER_59_85 ();
 sg13g2_fill_2 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_133 ();
 sg13g2_fill_2 FILLER_59_186 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_decap_8 FILLER_59_233 ();
 sg13g2_decap_8 FILLER_59_276 ();
 sg13g2_fill_2 FILLER_59_283 ();
 sg13g2_fill_1 FILLER_59_303 ();
 sg13g2_fill_2 FILLER_59_333 ();
 sg13g2_fill_1 FILLER_59_335 ();
 sg13g2_fill_1 FILLER_59_353 ();
 sg13g2_fill_2 FILLER_59_370 ();
 sg13g2_fill_1 FILLER_59_372 ();
 sg13g2_decap_8 FILLER_59_397 ();
 sg13g2_decap_4 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_29 ();
 sg13g2_fill_1 FILLER_60_31 ();
 sg13g2_fill_2 FILLER_60_217 ();
 sg13g2_fill_2 FILLER_60_224 ();
 sg13g2_fill_1 FILLER_60_226 ();
 sg13g2_fill_1 FILLER_60_240 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_fill_1 FILLER_60_287 ();
 sg13g2_decap_4 FILLER_60_307 ();
 sg13g2_fill_1 FILLER_60_316 ();
 sg13g2_fill_1 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_328 ();
 sg13g2_fill_1 FILLER_60_339 ();
 sg13g2_fill_2 FILLER_60_368 ();
 sg13g2_fill_1 FILLER_60_370 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_decap_8 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_63 ();
 sg13g2_fill_2 FILLER_61_89 ();
 sg13g2_fill_1 FILLER_61_106 ();
 sg13g2_fill_1 FILLER_61_205 ();
 sg13g2_decap_4 FILLER_61_243 ();
 sg13g2_fill_2 FILLER_61_247 ();
 sg13g2_fill_1 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_291 ();
 sg13g2_decap_8 FILLER_61_298 ();
 sg13g2_decap_8 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_312 ();
 sg13g2_decap_8 FILLER_61_328 ();
 sg13g2_fill_2 FILLER_61_344 ();
 sg13g2_fill_1 FILLER_61_346 ();
 sg13g2_decap_4 FILLER_61_355 ();
 sg13g2_fill_1 FILLER_61_359 ();
 sg13g2_decap_4 FILLER_61_365 ();
 sg13g2_fill_1 FILLER_61_369 ();
 sg13g2_decap_8 FILLER_61_376 ();
 sg13g2_decap_8 FILLER_61_383 ();
 sg13g2_decap_8 FILLER_61_390 ();
 sg13g2_decap_8 FILLER_61_397 ();
 sg13g2_decap_4 FILLER_61_404 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_2 FILLER_62_22 ();
 sg13g2_fill_1 FILLER_62_24 ();
 sg13g2_fill_2 FILLER_62_67 ();
 sg13g2_fill_1 FILLER_62_94 ();
 sg13g2_fill_1 FILLER_62_100 ();
 sg13g2_fill_1 FILLER_62_128 ();
 sg13g2_fill_2 FILLER_62_211 ();
 sg13g2_decap_8 FILLER_62_241 ();
 sg13g2_decap_8 FILLER_62_248 ();
 sg13g2_fill_2 FILLER_62_265 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_decap_8 FILLER_62_299 ();
 sg13g2_fill_2 FILLER_62_306 ();
 sg13g2_fill_2 FILLER_62_335 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_decap_8 FILLER_62_342 ();
 sg13g2_decap_4 FILLER_62_349 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_decap_8 FILLER_62_402 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_30 ();
 sg13g2_fill_1 FILLER_63_46 ();
 sg13g2_fill_2 FILLER_63_77 ();
 sg13g2_fill_2 FILLER_63_117 ();
 sg13g2_fill_1 FILLER_63_119 ();
 sg13g2_decap_4 FILLER_63_255 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_fill_2 FILLER_63_273 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_fill_2 FILLER_63_284 ();
 sg13g2_fill_2 FILLER_63_299 ();
 sg13g2_decap_8 FILLER_63_348 ();
 sg13g2_fill_2 FILLER_63_355 ();
 sg13g2_fill_1 FILLER_63_357 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_fill_1 FILLER_63_368 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_fill_1 FILLER_64_66 ();
 sg13g2_fill_1 FILLER_64_159 ();
 sg13g2_fill_1 FILLER_64_169 ();
 sg13g2_fill_2 FILLER_64_237 ();
 sg13g2_fill_1 FILLER_64_263 ();
 sg13g2_fill_2 FILLER_64_276 ();
 sg13g2_fill_1 FILLER_64_278 ();
 sg13g2_fill_2 FILLER_64_291 ();
 sg13g2_fill_1 FILLER_64_302 ();
 sg13g2_decap_4 FILLER_64_329 ();
 sg13g2_fill_2 FILLER_64_333 ();
 sg13g2_fill_2 FILLER_64_357 ();
 sg13g2_fill_1 FILLER_64_359 ();
 sg13g2_fill_2 FILLER_64_378 ();
 sg13g2_fill_1 FILLER_64_380 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_1 FILLER_65_25 ();
 sg13g2_fill_2 FILLER_65_94 ();
 sg13g2_fill_1 FILLER_65_104 ();
 sg13g2_fill_2 FILLER_65_254 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_decap_4 FILLER_65_261 ();
 sg13g2_decap_4 FILLER_65_269 ();
 sg13g2_fill_2 FILLER_65_282 ();
 sg13g2_fill_1 FILLER_65_284 ();
 sg13g2_fill_1 FILLER_65_292 ();
 sg13g2_decap_4 FILLER_65_321 ();
 sg13g2_fill_1 FILLER_65_330 ();
 sg13g2_decap_4 FILLER_65_341 ();
 sg13g2_fill_2 FILLER_65_345 ();
 sg13g2_fill_2 FILLER_65_352 ();
 sg13g2_fill_1 FILLER_65_366 ();
 sg13g2_decap_8 FILLER_65_374 ();
 sg13g2_decap_8 FILLER_65_381 ();
 sg13g2_decap_8 FILLER_65_388 ();
 sg13g2_decap_8 FILLER_65_395 ();
 sg13g2_decap_8 FILLER_65_402 ();
 sg13g2_fill_2 FILLER_66_155 ();
 sg13g2_decap_4 FILLER_66_170 ();
 sg13g2_fill_2 FILLER_66_178 ();
 sg13g2_fill_2 FILLER_66_184 ();
 sg13g2_fill_2 FILLER_66_225 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_decap_8 FILLER_66_271 ();
 sg13g2_fill_2 FILLER_66_278 ();
 sg13g2_fill_1 FILLER_66_280 ();
 sg13g2_fill_2 FILLER_66_289 ();
 sg13g2_fill_1 FILLER_66_291 ();
 sg13g2_decap_8 FILLER_66_314 ();
 sg13g2_fill_1 FILLER_66_356 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_decap_8 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_393 ();
 sg13g2_decap_8 FILLER_66_400 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_176 ();
 sg13g2_decap_8 FILLER_67_183 ();
 sg13g2_decap_8 FILLER_67_190 ();
 sg13g2_fill_2 FILLER_67_197 ();
 sg13g2_decap_4 FILLER_67_204 ();
 sg13g2_fill_1 FILLER_67_217 ();
 sg13g2_fill_2 FILLER_67_228 ();
 sg13g2_fill_1 FILLER_67_230 ();
 sg13g2_fill_2 FILLER_67_236 ();
 sg13g2_fill_1 FILLER_67_242 ();
 sg13g2_decap_8 FILLER_67_257 ();
 sg13g2_decap_8 FILLER_67_264 ();
 sg13g2_fill_2 FILLER_67_271 ();
 sg13g2_decap_8 FILLER_67_306 ();
 sg13g2_decap_8 FILLER_67_313 ();
 sg13g2_decap_4 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_346 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_61 ();
 sg13g2_fill_2 FILLER_68_107 ();
 sg13g2_decap_8 FILLER_68_178 ();
 sg13g2_decap_8 FILLER_68_185 ();
 sg13g2_decap_8 FILLER_68_192 ();
 sg13g2_decap_4 FILLER_68_199 ();
 sg13g2_fill_2 FILLER_68_203 ();
 sg13g2_fill_2 FILLER_68_210 ();
 sg13g2_fill_1 FILLER_68_212 ();
 sg13g2_fill_2 FILLER_68_226 ();
 sg13g2_fill_2 FILLER_68_243 ();
 sg13g2_decap_4 FILLER_68_257 ();
 sg13g2_fill_2 FILLER_68_261 ();
 sg13g2_fill_2 FILLER_68_268 ();
 sg13g2_decap_8 FILLER_68_303 ();
 sg13g2_decap_4 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_2 FILLER_68_334 ();
 sg13g2_decap_8 FILLER_68_361 ();
 sg13g2_fill_1 FILLER_68_368 ();
 sg13g2_decap_8 FILLER_68_373 ();
 sg13g2_fill_2 FILLER_68_380 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_decap_8 FILLER_68_393 ();
 sg13g2_decap_8 FILLER_68_400 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_fill_1 FILLER_69_26 ();
 sg13g2_fill_1 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_146 ();
 sg13g2_fill_1 FILLER_69_222 ();
 sg13g2_fill_2 FILLER_69_237 ();
 sg13g2_decap_4 FILLER_69_246 ();
 sg13g2_fill_2 FILLER_69_267 ();
 sg13g2_fill_2 FILLER_69_295 ();
 sg13g2_decap_8 FILLER_69_389 ();
 sg13g2_decap_8 FILLER_69_396 ();
 sg13g2_decap_4 FILLER_69_403 ();
 sg13g2_fill_2 FILLER_69_407 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_20 ();
 sg13g2_fill_1 FILLER_70_49 ();
 sg13g2_fill_1 FILLER_70_74 ();
 sg13g2_fill_1 FILLER_70_146 ();
 sg13g2_fill_1 FILLER_70_168 ();
 sg13g2_fill_2 FILLER_70_199 ();
 sg13g2_fill_1 FILLER_70_258 ();
 sg13g2_fill_2 FILLER_70_273 ();
 sg13g2_decap_4 FILLER_70_289 ();
 sg13g2_decap_8 FILLER_70_313 ();
 sg13g2_decap_4 FILLER_70_324 ();
 sg13g2_fill_1 FILLER_70_328 ();
 sg13g2_fill_1 FILLER_70_333 ();
 sg13g2_decap_4 FILLER_70_343 ();
 sg13g2_fill_1 FILLER_70_365 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_fill_2 FILLER_70_406 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_42 ();
 sg13g2_fill_2 FILLER_71_63 ();
 sg13g2_fill_1 FILLER_71_104 ();
 sg13g2_fill_1 FILLER_71_122 ();
 sg13g2_fill_2 FILLER_71_139 ();
 sg13g2_fill_2 FILLER_71_211 ();
 sg13g2_fill_1 FILLER_71_213 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_fill_1 FILLER_71_271 ();
 sg13g2_fill_2 FILLER_71_293 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_2 FILLER_71_320 ();
 sg13g2_decap_4 FILLER_71_333 ();
 sg13g2_fill_2 FILLER_71_350 ();
 sg13g2_fill_1 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_394 ();
 sg13g2_decap_8 FILLER_71_401 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_fill_1 FILLER_72_89 ();
 sg13g2_fill_2 FILLER_72_113 ();
 sg13g2_fill_2 FILLER_72_152 ();
 sg13g2_fill_1 FILLER_72_174 ();
 sg13g2_fill_2 FILLER_72_184 ();
 sg13g2_fill_2 FILLER_72_205 ();
 sg13g2_fill_1 FILLER_72_220 ();
 sg13g2_fill_1 FILLER_72_226 ();
 sg13g2_fill_2 FILLER_72_255 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_fill_2 FILLER_72_270 ();
 sg13g2_fill_1 FILLER_72_272 ();
 sg13g2_fill_2 FILLER_72_285 ();
 sg13g2_decap_8 FILLER_72_292 ();
 sg13g2_decap_4 FILLER_72_299 ();
 sg13g2_fill_1 FILLER_72_303 ();
 sg13g2_fill_1 FILLER_72_338 ();
 sg13g2_fill_1 FILLER_72_363 ();
 sg13g2_fill_2 FILLER_72_374 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_fill_2 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_fill_2 FILLER_73_13 ();
 sg13g2_fill_2 FILLER_73_28 ();
 sg13g2_fill_2 FILLER_73_110 ();
 sg13g2_fill_1 FILLER_73_147 ();
 sg13g2_fill_2 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_171 ();
 sg13g2_fill_2 FILLER_73_198 ();
 sg13g2_fill_1 FILLER_73_200 ();
 sg13g2_decap_4 FILLER_73_218 ();
 sg13g2_decap_4 FILLER_73_227 ();
 sg13g2_fill_1 FILLER_73_274 ();
 sg13g2_decap_4 FILLER_73_308 ();
 sg13g2_fill_2 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_318 ();
 sg13g2_fill_2 FILLER_73_329 ();
 sg13g2_fill_2 FILLER_73_363 ();
 sg13g2_fill_1 FILLER_73_365 ();
 sg13g2_decap_8 FILLER_73_390 ();
 sg13g2_decap_8 FILLER_73_397 ();
 sg13g2_decap_4 FILLER_73_404 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_fill_1 FILLER_74_85 ();
 sg13g2_fill_1 FILLER_74_148 ();
 sg13g2_fill_2 FILLER_74_164 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_fill_1 FILLER_74_182 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_1 FILLER_74_262 ();
 sg13g2_fill_2 FILLER_74_269 ();
 sg13g2_fill_1 FILLER_74_271 ();
 sg13g2_fill_2 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_287 ();
 sg13g2_fill_2 FILLER_74_304 ();
 sg13g2_fill_1 FILLER_74_306 ();
 sg13g2_fill_2 FILLER_74_320 ();
 sg13g2_fill_1 FILLER_74_322 ();
 sg13g2_fill_1 FILLER_74_328 ();
 sg13g2_fill_2 FILLER_74_342 ();
 sg13g2_fill_1 FILLER_74_344 ();
 sg13g2_fill_1 FILLER_74_373 ();
 sg13g2_decap_8 FILLER_74_387 ();
 sg13g2_decap_8 FILLER_74_394 ();
 sg13g2_decap_8 FILLER_74_401 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_8 ();
 sg13g2_fill_1 FILLER_75_57 ();
 sg13g2_fill_1 FILLER_75_81 ();
 sg13g2_fill_2 FILLER_75_120 ();
 sg13g2_decap_4 FILLER_75_204 ();
 sg13g2_fill_1 FILLER_75_208 ();
 sg13g2_fill_2 FILLER_75_235 ();
 sg13g2_fill_1 FILLER_75_237 ();
 sg13g2_fill_2 FILLER_75_242 ();
 sg13g2_fill_2 FILLER_75_268 ();
 sg13g2_decap_4 FILLER_75_298 ();
 sg13g2_fill_1 FILLER_75_302 ();
 sg13g2_fill_2 FILLER_75_329 ();
 sg13g2_fill_2 FILLER_75_340 ();
 sg13g2_fill_2 FILLER_75_356 ();
 sg13g2_fill_1 FILLER_75_358 ();
 sg13g2_fill_2 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_388 ();
 sg13g2_decap_8 FILLER_75_395 ();
 sg13g2_decap_8 FILLER_75_402 ();
 sg13g2_decap_4 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_4 ();
 sg13g2_fill_1 FILLER_76_16 ();
 sg13g2_fill_2 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_167 ();
 sg13g2_decap_4 FILLER_76_200 ();
 sg13g2_decap_4 FILLER_76_208 ();
 sg13g2_fill_1 FILLER_76_212 ();
 sg13g2_fill_2 FILLER_76_227 ();
 sg13g2_fill_1 FILLER_76_229 ();
 sg13g2_decap_8 FILLER_76_293 ();
 sg13g2_decap_8 FILLER_76_300 ();
 sg13g2_decap_8 FILLER_76_307 ();
 sg13g2_decap_4 FILLER_76_314 ();
 sg13g2_fill_2 FILLER_76_318 ();
 sg13g2_fill_2 FILLER_76_348 ();
 sg13g2_fill_1 FILLER_76_350 ();
 sg13g2_fill_1 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_386 ();
 sg13g2_decap_8 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_77 ();
 sg13g2_fill_1 FILLER_77_144 ();
 sg13g2_fill_2 FILLER_77_175 ();
 sg13g2_fill_1 FILLER_77_186 ();
 sg13g2_fill_2 FILLER_77_283 ();
 sg13g2_fill_1 FILLER_77_311 ();
 sg13g2_fill_1 FILLER_77_324 ();
 sg13g2_fill_2 FILLER_77_343 ();
 sg13g2_fill_1 FILLER_77_345 ();
 sg13g2_decap_4 FILLER_77_358 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_275 ();
 sg13g2_fill_1 FILLER_78_316 ();
 sg13g2_fill_2 FILLER_78_334 ();
 sg13g2_fill_1 FILLER_78_336 ();
 sg13g2_fill_1 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_14 ();
 sg13g2_fill_2 FILLER_79_53 ();
 sg13g2_fill_2 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_155 ();
 sg13g2_decap_4 FILLER_79_240 ();
 sg13g2_decap_4 FILLER_79_258 ();
 sg13g2_fill_1 FILLER_79_262 ();
 sg13g2_fill_2 FILLER_79_289 ();
 sg13g2_fill_1 FILLER_79_291 ();
 sg13g2_fill_2 FILLER_79_300 ();
 sg13g2_fill_2 FILLER_79_328 ();
 sg13g2_fill_1 FILLER_79_330 ();
 sg13g2_fill_1 FILLER_79_357 ();
 sg13g2_fill_1 FILLER_79_363 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_4 FILLER_80_7 ();
 sg13g2_fill_2 FILLER_80_11 ();
 sg13g2_fill_2 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_96 ();
 sg13g2_fill_1 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_132 ();
 sg13g2_fill_2 FILLER_80_137 ();
 sg13g2_fill_2 FILLER_80_150 ();
 sg13g2_fill_2 FILLER_80_173 ();
 sg13g2_fill_1 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_fill_2 FILLER_80_208 ();
 sg13g2_fill_1 FILLER_80_210 ();
 sg13g2_fill_1 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_fill_2 FILLER_80_227 ();
 sg13g2_fill_1 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_233 ();
 sg13g2_decap_8 FILLER_80_240 ();
 sg13g2_decap_8 FILLER_80_247 ();
 sg13g2_decap_8 FILLER_80_254 ();
 sg13g2_decap_8 FILLER_80_261 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_fill_1 FILLER_80_299 ();
 sg13g2_fill_2 FILLER_80_309 ();
 sg13g2_fill_1 FILLER_80_311 ();
 sg13g2_fill_2 FILLER_80_321 ();
 sg13g2_fill_1 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_346 ();
 sg13g2_decap_8 FILLER_80_353 ();
 sg13g2_decap_8 FILLER_80_360 ();
 sg13g2_decap_8 FILLER_80_367 ();
 sg13g2_fill_2 FILLER_80_374 ();
 sg13g2_decap_8 FILLER_80_384 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_4 FILLER_80_405 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net225;
 assign uio_oe[2] = net226;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net227;
 assign uio_oe[5] = net228;
 assign uio_oe[6] = net6;
 assign uio_oe[7] = net7;
 assign uio_out[0] = net8;
 assign uio_out[3] = net9;
 assign uio_out[6] = net10;
 assign uio_out[7] = net11;
endmodule

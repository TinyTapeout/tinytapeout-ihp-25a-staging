module tt_um_silice (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire \main._w_demo_audio1 ;
 wire \main._w_demo_video_hs ;
 wire \main._w_demo_video_vs ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[0] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[10] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[5] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[8] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[9] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[5] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[5] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[0] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[1] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[2] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[3] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[4] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[5] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[0] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[1] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[2] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_l[0] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_l[1] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[9] ;
 wire \main.demo._d_prev_b[0] ;
 wire \main.demo._d_prev_b[1] ;
 wire \main.demo._d_prev_b[2] ;
 wire \main.demo._d_prev_b[3] ;
 wire \main.demo._d_prev_b[4] ;
 wire \main.demo._d_prev_b[5] ;
 wire \main.demo._d_prev_b[6] ;
 wire \main.demo._d_prev_b[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[0] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[10] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[1] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[2] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[3] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[4] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[5] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[6] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[8] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[9] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[0] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[10] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[1] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[2] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[3] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[4] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[5] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[6] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[8] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[9] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[0] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[10] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[5] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[8] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[9] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[0] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[10] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[5] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[8] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[9] ;
 wire \main.demo._q_effect[0] ;
 wire \main.demo._q_effect[1] ;
 wire \main.demo._q_frame[0] ;
 wire \main.demo._q_frame[10] ;
 wire \main.demo._q_frame[11] ;
 wire \main.demo._q_frame[12] ;
 wire \main.demo._q_frame[13] ;
 wire \main.demo._q_frame[14] ;
 wire \main.demo._q_frame[1] ;
 wire \main.demo._q_frame[2] ;
 wire \main.demo._q_frame[3] ;
 wire \main.demo._q_frame[4] ;
 wire \main.demo._q_frame[5] ;
 wire \main.demo._q_frame[6] ;
 wire \main.demo._q_frame[7] ;
 wire \main.demo._q_frame[8] ;
 wire \main.demo._q_frame[9] ;
 wire \main.demo._q_go ;
 wire \main.demo._q_prev_b[6] ;
 wire \main.demo._q_prev_b[7] ;
 wire \main.demo._q_prev_vs ;
 wire \main.demo._q_rot_en ;
 wire \main.demo._q_speed[0] ;
 wire \main.demo._q_speed[10] ;
 wire \main.demo._q_speed[11] ;
 wire \main.demo._q_speed[12] ;
 wire \main.demo._q_speed[13] ;
 wire \main.demo._q_speed[14] ;
 wire \main.demo._q_speed[15] ;
 wire \main.demo._q_speed[1] ;
 wire \main.demo._q_speed[2] ;
 wire \main.demo._q_speed[3] ;
 wire \main.demo._q_speed[4] ;
 wire \main.demo._q_speed[5] ;
 wire \main.demo._q_speed[6] ;
 wire \main.demo._q_speed[7] ;
 wire \main.demo._q_speed[8] ;
 wire \main.demo._q_speed[9] ;
 wire \main.demo._q_th[0] ;
 wire \main.demo._q_th[1] ;
 wire \main.demo._q_th[2] ;
 wire \main.demo._q_th[3] ;
 wire \main.demo._q_th[4] ;
 wire \main.demo._q_th[5] ;
 wire \main.demo._q_th[6] ;
 wire \main.demo._q_th[7] ;
 wire \main.demo._q_th[8] ;
 wire \main.demo._t___block_68_frag[0] ;
 wire \main.demo._t___block_68_frag[1] ;
 wire \main.demo._t___block_68_frag[2] ;
 wire \main.demo._t___block_68_frag[3] ;
 wire \main.demo._t___block_68_frag[4] ;
 wire \main.demo._t___block_68_frag[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_a[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_a[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[0] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[10] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[1] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[2] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[3] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[4] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[8] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[9] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[0] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[10] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[1] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[2] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[3] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[4] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[8] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[9] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[0] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[1] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[2] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_l[0] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_l[1] ;
 wire \main.demo._t___stage___block_3_x[0] ;
 wire \main.demo._t___stage___block_3_x[1] ;
 wire \main.demo._t___stage___block_3_x[2] ;
 wire \main.demo._t___stage___block_3_y[0] ;
 wire \main.demo._t___stage___block_3_y[1] ;
 wire \main.demo._t___stage___block_3_y[2] ;
 wire \main.demo._w_vga_active ;
 wire \main.demo._w_vga_vga_x[10] ;
 wire \main.demo._w_vga_vga_x[3] ;
 wire \main.demo._w_vga_vga_x[4] ;
 wire \main.demo._w_vga_vga_x[5] ;
 wire \main.demo._w_vga_vga_x[6] ;
 wire \main.demo._w_vga_vga_x[7] ;
 wire \main.demo._w_vga_vga_x[8] ;
 wire \main.demo._w_vga_vga_x[9] ;
 wire \main.demo._w_vga_vga_y[10] ;
 wire \main.demo._w_vga_vga_y[3] ;
 wire \main.demo._w_vga_vga_y[4] ;
 wire \main.demo._w_vga_vga_y[5] ;
 wire \main.demo._w_vga_vga_y[6] ;
 wire \main.demo._w_vga_vga_y[7] ;
 wire \main.demo._w_vga_vga_y[8] ;
 wire \main.demo.vga._d_active ;
 wire \main.demo.vga._d_vblank ;
 wire \main.demo.vga._q_active_h ;
 wire \main.demo.vga._q_active_v ;
 wire \main.demo.vga._q_xcount[0] ;
 wire \main.demo.vga._q_xcount[10] ;
 wire \main.demo.vga._q_xcount[1] ;
 wire \main.demo.vga._q_xcount[2] ;
 wire \main.demo.vga._q_xcount[3] ;
 wire \main.demo.vga._q_xcount[4] ;
 wire \main.demo.vga._q_xcount[5] ;
 wire \main.demo.vga._q_xcount[6] ;
 wire \main.demo.vga._q_xcount[7] ;
 wire \main.demo.vga._q_xcount[8] ;
 wire \main.demo.vga._q_xcount[9] ;
 wire \main.demo.vga._q_ycount[0] ;
 wire \main.demo.vga._q_ycount[1] ;
 wire \main.demo.vga._q_ycount[2] ;
 wire \main.demo.vga._q_ycount[3] ;
 wire \main.demo.vga._q_ycount[4] ;
 wire \main.demo.vga._q_ycount[5] ;
 wire \main.demo.vga._q_ycount[6] ;
 wire \main.demo.vga._q_ycount[7] ;
 wire \main.demo.vga._q_ycount[8] ;
 wire \main.demo.zic._q_clock_count[0] ;
 wire \main.demo.zic._q_clock_count[1] ;
 wire \main.demo.zic._q_clock_count[2] ;
 wire \main.demo.zic._q_clock_count[3] ;
 wire \main.demo.zic._q_clock_count[4] ;
 wire \main.demo.zic._q_clock_count[5] ;
 wire \main.demo.zic._q_clock_count[6] ;
 wire \main.demo.zic._q_clock_count[7] ;
 wire \main.demo.zic._q_clock_count[8] ;
 wire \main.demo.zic._q_drum_inc[0] ;
 wire \main.demo.zic._q_drum_inc[1] ;
 wire \main.demo.zic._q_drum_inc[2] ;
 wire \main.demo.zic._q_drum_inc[3] ;
 wire \main.demo.zic._q_idx[0] ;
 wire \main.demo.zic._q_idx[1] ;
 wire \main.demo.zic._q_idx[2] ;
 wire \main.demo.zic._q_idx[3] ;
 wire \main.demo.zic._q_idx[4] ;
 wire \main.demo.zic._q_idx[5] ;
 wire \main.demo.zic._q_idx[6] ;
 wire \main.demo.zic._q_qpos[0] ;
 wire \main.demo.zic._q_qpos[10] ;
 wire \main.demo.zic._q_qpos[11] ;
 wire \main.demo.zic._q_qpos[12] ;
 wire \main.demo.zic._q_qpos[1] ;
 wire \main.demo.zic._q_qpos[2] ;
 wire \main.demo.zic._q_qpos[3] ;
 wire \main.demo.zic._q_qpos[4] ;
 wire \main.demo.zic._q_qpos[5] ;
 wire \main.demo.zic._q_qpos[6] ;
 wire \main.demo.zic._q_qpos[7] ;
 wire \main.demo.zic._q_qpos[8] ;
 wire \main.demo.zic._q_qpos[9] ;
 wire \main.demo.zic._q_rythm_count[0] ;
 wire \main.demo.zic._q_rythm_count[10] ;
 wire \main.demo.zic._q_rythm_count[11] ;
 wire \main.demo.zic._q_rythm_count[12] ;
 wire \main.demo.zic._q_rythm_count[1] ;
 wire \main.demo.zic._q_rythm_count[2] ;
 wire \main.demo.zic._q_rythm_count[3] ;
 wire \main.demo.zic._q_rythm_count[4] ;
 wire \main.demo.zic._q_rythm_count[5] ;
 wire \main.demo.zic._q_rythm_count[6] ;
 wire \main.demo.zic._q_rythm_count[7] ;
 wire \main.demo.zic._q_rythm_count[8] ;
 wire \main.demo.zic._q_rythm_count[9] ;
 wire \main.demo.zic._q_squ_env[0] ;
 wire \main.demo.zic._q_squ_env[1] ;
 wire \main.demo.zic._q_squ_env[2] ;
 wire \main.demo.zic._q_squ_env[3] ;
 wire \main.demo.zic._q_squ_env[4] ;
 wire \main.demo.zic._q_squ_env[5] ;
 wire \main.demo.zic._q_tpos[0] ;
 wire \main.demo.zic._q_tpos[10] ;
 wire \main.demo.zic._q_tpos[11] ;
 wire \main.demo.zic._q_tpos[1] ;
 wire \main.demo.zic._q_tpos[2] ;
 wire \main.demo.zic._q_tpos[3] ;
 wire \main.demo.zic._q_tpos[4] ;
 wire \main.demo.zic._q_tpos[5] ;
 wire \main.demo.zic._q_tpos[6] ;
 wire \main.demo.zic._q_tpos[7] ;
 wire \main.demo.zic._q_tpos[8] ;
 wire \main.demo.zic._q_tpos[9] ;
 wire rst_n_q;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_leaf_0_clk;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;

 sg13g2_inv_1 _3783_ (.Y(_2902_),
    .A(net564));
 sg13g2_inv_1 _3784_ (.Y(_2903_),
    .A(net535));
 sg13g2_inv_1 _3785_ (.Y(_2904_),
    .A(net522));
 sg13g2_inv_1 _3786_ (.Y(_2905_),
    .A(net534));
 sg13g2_inv_1 _3787_ (.Y(_2906_),
    .A(\main.demo.zic._q_rythm_count[10] ));
 sg13g2_inv_1 _3788_ (.Y(_2907_),
    .A(net334));
 sg13g2_inv_1 _3789_ (.Y(_2908_),
    .A(net524));
 sg13g2_inv_2 _3790_ (.Y(_2909_),
    .A(\main.demo._q_th[6] ));
 sg13g2_inv_2 _3791_ (.Y(_2910_),
    .A(\main.demo._q_th[3] ));
 sg13g2_inv_1 _3792_ (.Y(_2911_),
    .A(\main.demo._q_th[2] ));
 sg13g2_inv_1 _3793_ (.Y(_2912_),
    .A(net474));
 sg13g2_inv_2 _3794_ (.Y(_2913_),
    .A(net478));
 sg13g2_inv_1 _3795_ (.Y(_2914_),
    .A(net463));
 sg13g2_inv_1 _3796_ (.Y(_2915_),
    .A(net483));
 sg13g2_inv_1 _3797_ (.Y(_2916_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_inv_4 _3798_ (.A(net499),
    .Y(_2917_));
 sg13g2_inv_1 _3799_ (.Y(_2918_),
    .A(_0040_));
 sg13g2_inv_1 _3800_ (.Y(_2919_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ));
 sg13g2_inv_1 _3801_ (.Y(_2920_),
    .A(_0046_));
 sg13g2_inv_1 _3802_ (.Y(_2921_),
    .A(_0047_));
 sg13g2_inv_1 _3803_ (.Y(_2922_),
    .A(_0048_));
 sg13g2_inv_1 _3804_ (.Y(_2923_),
    .A(_0049_));
 sg13g2_inv_1 _3805_ (.Y(_2924_),
    .A(_0050_));
 sg13g2_inv_2 _3806_ (.Y(_2925_),
    .A(net491));
 sg13g2_inv_1 _3807_ (.Y(_2926_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ));
 sg13g2_inv_1 _3808_ (.Y(_2927_),
    .A(\main.demo._w_vga_vga_x[8] ));
 sg13g2_inv_1 _3809_ (.Y(_2928_),
    .A(net467));
 sg13g2_inv_1 _3810_ (.Y(_2929_),
    .A(net653));
 sg13g2_inv_1 _3811_ (.Y(_2930_),
    .A(\main.demo._q_frame[4] ));
 sg13g2_inv_1 _3812_ (.Y(_2931_),
    .A(net471));
 sg13g2_inv_1 _3813_ (.Y(_2932_),
    .A(\main.demo._q_frame[3] ));
 sg13g2_inv_1 _3814_ (.Y(_2933_),
    .A(\main.demo._w_vga_vga_x[3] ));
 sg13g2_inv_1 _3815_ (.Y(_2934_),
    .A(_0061_));
 sg13g2_inv_1 _3816_ (.Y(_2935_),
    .A(\main.demo._w_vga_vga_y[5] ));
 sg13g2_inv_1 _3817_ (.Y(_2936_),
    .A(net506));
 sg13g2_inv_1 _3818_ (.Y(_2937_),
    .A(\main.demo.vga._q_active_h ));
 sg13g2_inv_2 _3819_ (.Y(_2938_),
    .A(\main.demo._t___stage___block_3_y[0] ));
 sg13g2_inv_1 _3820_ (.Y(_2939_),
    .A(\main.demo._t___stage___block_3_x[0] ));
 sg13g2_inv_1 _3821_ (.Y(_2940_),
    .A(\main.demo._t___stage___block_3_y[1] ));
 sg13g2_inv_1 _3822_ (.Y(_2941_),
    .A(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_inv_1 _3823_ (.Y(_2942_),
    .A(\main.demo._t___stage___block_3_y[2] ));
 sg13g2_inv_2 _3824_ (.Y(_2943_),
    .A(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_inv_1 _3825_ (.Y(_2944_),
    .A(\main.demo._q_frame[13] ));
 sg13g2_inv_2 _3826_ (.Y(_2945_),
    .A(net654));
 sg13g2_inv_1 _3827_ (.Y(_2946_),
    .A(net634));
 sg13g2_inv_2 _3828_ (.Y(_2947_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ));
 sg13g2_inv_1 _3829_ (.Y(_2948_),
    .A(net488));
 sg13g2_inv_2 _3830_ (.Y(_2949_),
    .A(_0008_));
 sg13g2_inv_2 _3831_ (.Y(_2950_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ));
 sg13g2_inv_1 _3832_ (.Y(_2951_),
    .A(_0014_));
 sg13g2_inv_1 _3833_ (.Y(_2952_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ));
 sg13g2_inv_1 _3834_ (.Y(_2953_),
    .A(_0017_));
 sg13g2_inv_1 _3835_ (.Y(_2954_),
    .A(_0019_));
 sg13g2_inv_1 _3836_ (.Y(_2955_),
    .A(_0020_));
 sg13g2_inv_1 _3837_ (.Y(_2956_),
    .A(_0021_));
 sg13g2_inv_1 _3838_ (.Y(_2957_),
    .A(_0024_));
 sg13g2_inv_1 _3839_ (.Y(_2958_),
    .A(net635));
 sg13g2_inv_1 _3840_ (.Y(_2959_),
    .A(net614));
 sg13g2_inv_1 _3841_ (.Y(_2960_),
    .A(net577));
 sg13g2_inv_1 _3842_ (.Y(_2961_),
    .A(net558));
 sg13g2_inv_1 _3843_ (.Y(_2962_),
    .A(_0030_));
 sg13g2_inv_1 _3844_ (.Y(_2963_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_inv_1 _3845_ (.Y(_2964_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[3] ));
 sg13g2_inv_1 _3846_ (.Y(_2965_),
    .A(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ));
 sg13g2_inv_1 _3847_ (.Y(_2966_),
    .A(\main.demo._d___pip_58_1_4___stage___block_3_cx[3] ));
 sg13g2_inv_1 _3848_ (.Y(_2967_),
    .A(net285));
 sg13g2_nor2_1 _3849_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .Y(_2968_));
 sg13g2_or2_1 _3850_ (.X(_2969_),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ));
 sg13g2_nand2_2 _3851_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ),
    .A(net297),
    .B(net453));
 sg13g2_inv_1 _3852_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .A(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ));
 sg13g2_nor2b_1 _3853_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ),
    .B_N(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .Y(_2970_));
 sg13g2_xor2_1 _3854_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ),
    .X(_2971_));
 sg13g2_nor3_1 _3855_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ),
    .Y(_2972_));
 sg13g2_nand2b_1 _3856_ (.Y(_2973_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ),
    .A_N(_2972_));
 sg13g2_nand2b_1 _3857_ (.Y(_2974_),
    .B(_2972_),
    .A_N(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_nand3_1 _3858_ (.B(_2973_),
    .C(_2974_),
    .A(_2917_),
    .Y(_2975_));
 sg13g2_o21ai_1 _3859_ (.B1(_2975_),
    .Y(_2976_),
    .A1(_2917_),
    .A2(_0039_));
 sg13g2_nand2b_1 _3860_ (.Y(_2977_),
    .B(_2976_),
    .A_N(_0038_));
 sg13g2_o21ai_1 _3861_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ),
    .Y(_2978_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_nor2_1 _3862_ (.A(net497),
    .B(_2972_),
    .Y(_2979_));
 sg13g2_a22oi_1 _3863_ (.Y(_2980_),
    .B1(_2978_),
    .B2(_2979_),
    .A2(_2918_),
    .A1(net497));
 sg13g2_nor2b_1 _3864_ (.A(_2980_),
    .B_N(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ),
    .Y(_2981_));
 sg13g2_xnor2_1 _3865_ (.Y(_2982_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_mux2_1 _3866_ (.A0(_0041_),
    .A1(_2982_),
    .S(_2917_),
    .X(_2983_));
 sg13g2_nand2_1 _3867_ (.Y(_2984_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ));
 sg13g2_xnor2_1 _3868_ (.Y(_2985_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ),
    .B(_2983_));
 sg13g2_nand2b_1 _3869_ (.Y(_2986_),
    .B(_2985_),
    .A_N(_2984_));
 sg13g2_o21ai_1 _3870_ (.B1(_2986_),
    .Y(_2987_),
    .A1(_2919_),
    .A2(_2983_));
 sg13g2_xnor2_1 _3871_ (.Y(_2988_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ),
    .B(_2980_));
 sg13g2_a21oi_1 _3872_ (.A1(_2987_),
    .A2(_2988_),
    .Y(_2989_),
    .B1(_2981_));
 sg13g2_xor2_1 _3873_ (.B(_2976_),
    .A(_0038_),
    .X(_2990_));
 sg13g2_o21ai_1 _3874_ (.B1(_2977_),
    .Y(_2991_),
    .A1(_2989_),
    .A2(_2990_));
 sg13g2_nand2_1 _3875_ (.Y(_2992_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ),
    .B(_2974_));
 sg13g2_or2_2 _3876_ (.X(_2993_),
    .B(_2974_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ));
 sg13g2_a21oi_1 _3877_ (.A1(_2992_),
    .A2(_2993_),
    .Y(_2994_),
    .B1(net495));
 sg13g2_a21oi_1 _3878_ (.A1(_0037_),
    .A2(net495),
    .Y(_2995_),
    .B1(_2994_));
 sg13g2_xor2_1 _3879_ (.B(_2995_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ),
    .X(_2996_));
 sg13g2_xnor2_1 _3880_ (.Y(_2997_),
    .A(_2991_),
    .B(_2996_));
 sg13g2_nor2_1 _3881_ (.A(_2971_),
    .B(_2997_),
    .Y(_2998_));
 sg13g2_inv_1 _3882_ (.Y(_2999_),
    .A(_2998_));
 sg13g2_xnor2_1 _3883_ (.Y(_3000_),
    .A(_2971_),
    .B(_2997_));
 sg13g2_a22oi_1 _3884_ (.Y(_3001_),
    .B1(_2996_),
    .B2(_2991_),
    .A2(_2995_),
    .A1(_2924_));
 sg13g2_inv_1 _3885_ (.Y(_3002_),
    .A(_3001_));
 sg13g2_a21oi_1 _3886_ (.A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .A2(_2993_),
    .Y(_3003_),
    .B1(net496));
 sg13g2_o21ai_1 _3887_ (.B1(_3003_),
    .Y(_3004_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .A2(_2993_));
 sg13g2_o21ai_1 _3888_ (.B1(_3004_),
    .Y(_3005_),
    .A1(_2917_),
    .A2(_0044_));
 sg13g2_xor2_1 _3889_ (.B(_3005_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ),
    .X(_3006_));
 sg13g2_xor2_1 _3890_ (.B(_3006_),
    .A(_3001_),
    .X(_3007_));
 sg13g2_nor2_1 _3891_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ),
    .Y(_3008_));
 sg13g2_nor3_1 _3892_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ),
    .Y(_3009_));
 sg13g2_nor2b_1 _3893_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ),
    .B_N(_3009_),
    .Y(_3010_));
 sg13g2_nand2b_2 _3894_ (.Y(_3011_),
    .B(_3010_),
    .A_N(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ));
 sg13g2_nand2_1 _3895_ (.Y(_3012_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ),
    .B(_3011_));
 sg13g2_nor2_2 _3896_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ),
    .B(_3011_),
    .Y(_3013_));
 sg13g2_nor2_1 _3897_ (.A(net495),
    .B(_3013_),
    .Y(_3014_));
 sg13g2_a22oi_1 _3898_ (.Y(_3015_),
    .B1(_3012_),
    .B2(_3014_),
    .A2(_2920_),
    .A1(net495));
 sg13g2_nand2b_1 _3899_ (.Y(_3016_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ),
    .A_N(_3010_));
 sg13g2_a21oi_1 _3900_ (.A1(_3011_),
    .A2(_3016_),
    .Y(_3017_),
    .B1(net495));
 sg13g2_a21oi_2 _3901_ (.B1(_3017_),
    .Y(_3018_),
    .A2(_0047_),
    .A1(net495));
 sg13g2_nand2b_1 _3902_ (.Y(_3019_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ),
    .A_N(_3009_));
 sg13g2_nor2_1 _3903_ (.A(net496),
    .B(_3010_),
    .Y(_3020_));
 sg13g2_a22oi_1 _3904_ (.Y(_3021_),
    .B1(_3019_),
    .B2(_3020_),
    .A2(_2922_),
    .A1(net496));
 sg13g2_o21ai_1 _3905_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ),
    .Y(_3022_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ));
 sg13g2_nor2_1 _3906_ (.A(net497),
    .B(_3009_),
    .Y(_3023_));
 sg13g2_a22oi_1 _3907_ (.Y(_3024_),
    .B1(_3022_),
    .B2(_3023_),
    .A2(_2923_),
    .A1(net497));
 sg13g2_nand2_1 _3908_ (.Y(_3025_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ));
 sg13g2_nor2_1 _3909_ (.A(net497),
    .B(_3008_),
    .Y(_3026_));
 sg13g2_a22oi_1 _3910_ (.Y(_3027_),
    .B1(_3025_),
    .B2(_3026_),
    .A2(_2924_),
    .A1(net497));
 sg13g2_nand2_1 _3911_ (.Y(_3028_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[1] ),
    .B(_3027_));
 sg13g2_xnor2_1 _3912_ (.Y(_3029_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[1] ),
    .B(_3027_));
 sg13g2_o21ai_1 _3913_ (.B1(_3028_),
    .Y(_3030_),
    .A1(_2970_),
    .A2(_3029_));
 sg13g2_xnor2_1 _3914_ (.Y(_3031_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ),
    .B(_3024_));
 sg13g2_nor2b_1 _3915_ (.A(_3031_),
    .B_N(_3030_),
    .Y(_3032_));
 sg13g2_a21o_1 _3916_ (.A2(_3024_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ),
    .B1(_3032_),
    .X(_3033_));
 sg13g2_xnor2_1 _3917_ (.Y(_3034_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B(_3021_));
 sg13g2_nor2b_1 _3918_ (.A(_3034_),
    .B_N(_3033_),
    .Y(_3035_));
 sg13g2_a21o_1 _3919_ (.A2(_3021_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B1(_3035_),
    .X(_3036_));
 sg13g2_xor2_1 _3920_ (.B(_3018_),
    .A(_0041_),
    .X(_3037_));
 sg13g2_nand2_1 _3921_ (.Y(_3038_),
    .A(_3036_),
    .B(_3037_));
 sg13g2_o21ai_1 _3922_ (.B1(_3038_),
    .Y(_3039_),
    .A1(_2916_),
    .A2(_3018_));
 sg13g2_xnor2_1 _3923_ (.Y(_3040_),
    .A(_0040_),
    .B(_3015_));
 sg13g2_a22oi_1 _3924_ (.Y(_3041_),
    .B1(_3039_),
    .B2(_3040_),
    .A2(_3015_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ));
 sg13g2_xnor2_1 _3925_ (.Y(_3042_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .B(_3013_));
 sg13g2_nand2_1 _3926_ (.Y(_3043_),
    .A(net495),
    .B(_0045_));
 sg13g2_o21ai_1 _3927_ (.B1(_3043_),
    .Y(_3044_),
    .A1(net495),
    .A2(_3042_));
 sg13g2_xnor2_1 _3928_ (.Y(_3045_),
    .A(_0039_),
    .B(_3044_));
 sg13g2_nor2b_1 _3929_ (.A(_3041_),
    .B_N(_3045_),
    .Y(_3046_));
 sg13g2_a21o_1 _3930_ (.A2(_3044_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ),
    .B1(_3046_),
    .X(_3047_));
 sg13g2_nand3_1 _3931_ (.B(_0045_),
    .C(_3013_),
    .A(_0043_),
    .Y(_3048_));
 sg13g2_xor2_1 _3932_ (.B(_3048_),
    .A(_0037_),
    .X(_3049_));
 sg13g2_nand2_1 _3933_ (.Y(_3050_),
    .A(_3047_),
    .B(_3049_));
 sg13g2_nand4_1 _3934_ (.B(_0043_),
    .C(_0045_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ),
    .Y(_3051_),
    .D(_3013_));
 sg13g2_nor4_2 _3935_ (.A(net496),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ),
    .Y(_3052_),
    .D(_3011_));
 sg13g2_nand2_2 _3936_ (.Y(_3053_),
    .A(_0043_),
    .B(_3052_));
 sg13g2_xnor2_1 _3937_ (.Y(_3054_),
    .A(_0044_),
    .B(_3053_));
 sg13g2_a21o_1 _3938_ (.A2(_3051_),
    .A1(_3050_),
    .B1(_3054_),
    .X(_3055_));
 sg13g2_nand3_1 _3939_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .C(_3052_),
    .A(_0043_),
    .Y(_3056_));
 sg13g2_xnor2_1 _3940_ (.Y(_3057_),
    .A(_0042_),
    .B(_3053_));
 sg13g2_a21oi_2 _3941_ (.B1(_3057_),
    .Y(_3058_),
    .A2(_3056_),
    .A1(_3055_));
 sg13g2_nand3_1 _3942_ (.B(_3056_),
    .C(_3057_),
    .A(_3055_),
    .Y(_3059_));
 sg13g2_nor2b_2 _3943_ (.A(_3058_),
    .B_N(_3059_),
    .Y(_3060_));
 sg13g2_inv_1 _3944_ (.Y(_3061_),
    .A(_3060_));
 sg13g2_nand3_1 _3945_ (.B(_3051_),
    .C(_3054_),
    .A(_3050_),
    .Y(_3062_));
 sg13g2_nand2_2 _3946_ (.Y(_3063_),
    .A(_3055_),
    .B(_3062_));
 sg13g2_xnor2_1 _3947_ (.Y(_3064_),
    .A(_3041_),
    .B(_3045_));
 sg13g2_xor2_1 _3948_ (.B(_3040_),
    .A(_3039_),
    .X(_3065_));
 sg13g2_xnor2_1 _3949_ (.Y(_3066_),
    .A(_3036_),
    .B(_3037_));
 sg13g2_nor2b_1 _3950_ (.A(_3065_),
    .B_N(_3066_),
    .Y(_3067_));
 sg13g2_nand2b_1 _3951_ (.Y(_3068_),
    .B(_3067_),
    .A_N(_3064_));
 sg13g2_xor2_1 _3952_ (.B(_3049_),
    .A(_3047_),
    .X(_3069_));
 sg13g2_nor2_1 _3953_ (.A(_3068_),
    .B(_3069_),
    .Y(_3070_));
 sg13g2_nand2_1 _3954_ (.Y(_3071_),
    .A(_3063_),
    .B(_3070_));
 sg13g2_or3_1 _3955_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .C(_2993_),
    .X(_3072_));
 sg13g2_nor2_1 _3956_ (.A(net499),
    .B(_3072_),
    .Y(_3073_));
 sg13g2_nor2_1 _3957_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ),
    .B(_3073_),
    .Y(_3074_));
 sg13g2_nand2_1 _3958_ (.Y(_3075_),
    .A(_2917_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ));
 sg13g2_a21oi_1 _3959_ (.A1(net499),
    .A2(_0051_),
    .Y(_3076_),
    .B1(_3073_));
 sg13g2_nand2_2 _3960_ (.Y(_3077_),
    .A(_3075_),
    .B(_3076_));
 sg13g2_o21ai_1 _3961_ (.B1(_3077_),
    .Y(_3078_),
    .A1(_3072_),
    .A2(_3075_));
 sg13g2_o21ai_1 _3962_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .Y(_3079_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .A2(_2993_));
 sg13g2_a21oi_1 _3963_ (.A1(_3072_),
    .A2(_3079_),
    .Y(_3080_),
    .B1(net496));
 sg13g2_a21oi_1 _3964_ (.A1(net496),
    .A2(_0042_),
    .Y(_3081_),
    .B1(_3080_));
 sg13g2_a22oi_1 _3965_ (.Y(_3082_),
    .B1(_3006_),
    .B2(_3002_),
    .A2(_3005_),
    .A1(_2923_));
 sg13g2_inv_1 _3966_ (.Y(_3083_),
    .A(_3082_));
 sg13g2_xor2_1 _3967_ (.B(_3081_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ),
    .X(_3084_));
 sg13g2_a22oi_1 _3968_ (.Y(_3085_),
    .B1(_3083_),
    .B2(_3084_),
    .A2(_3081_),
    .A1(_2922_));
 sg13g2_inv_1 _3969_ (.Y(_3086_),
    .A(_3085_));
 sg13g2_xor2_1 _3970_ (.B(_3078_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ),
    .X(_3087_));
 sg13g2_a22oi_1 _3971_ (.Y(_3088_),
    .B1(_3086_),
    .B2(_3087_),
    .A2(_3078_),
    .A1(_2921_));
 sg13g2_xor2_1 _3972_ (.B(_3077_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ),
    .X(_3089_));
 sg13g2_or2_1 _3973_ (.X(_3090_),
    .B(_3089_),
    .A(_3088_));
 sg13g2_xor2_1 _3974_ (.B(_3077_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .X(_3091_));
 sg13g2_o21ai_1 _3975_ (.B1(_0045_),
    .Y(_3092_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .A2(_0046_));
 sg13g2_nand3_1 _3976_ (.B(_3076_),
    .C(_3092_),
    .A(_3075_),
    .Y(_3093_));
 sg13g2_o21ai_1 _3977_ (.B1(_3093_),
    .Y(_3094_),
    .A1(_3090_),
    .A2(_3091_));
 sg13g2_xor2_1 _3978_ (.B(_3094_),
    .A(_3074_),
    .X(_3095_));
 sg13g2_inv_2 _3979_ (.Y(_3096_),
    .A(net406));
 sg13g2_a21oi_1 _3980_ (.A1(_3063_),
    .A2(_3070_),
    .Y(_3097_),
    .B1(net404));
 sg13g2_xnor2_1 _3981_ (.Y(_3098_),
    .A(_3060_),
    .B(_3097_));
 sg13g2_nor2_1 _3982_ (.A(_3007_),
    .B(_3098_),
    .Y(_3099_));
 sg13g2_xor2_1 _3983_ (.B(_3098_),
    .A(_3007_),
    .X(_3100_));
 sg13g2_nor2_1 _3984_ (.A(_3070_),
    .B(net404),
    .Y(_3101_));
 sg13g2_xor2_1 _3985_ (.B(_3101_),
    .A(_3063_),
    .X(_3102_));
 sg13g2_nor2_1 _3986_ (.A(_3066_),
    .B(net404),
    .Y(_3103_));
 sg13g2_nor2_1 _3987_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ),
    .Y(_3104_));
 sg13g2_nor2_1 _3988_ (.A(_3066_),
    .B(_3104_),
    .Y(_3105_));
 sg13g2_a21o_1 _3989_ (.A2(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B1(_2985_),
    .X(_3106_));
 sg13g2_o21ai_1 _3990_ (.B1(_2986_),
    .Y(_3107_),
    .A1(_3105_),
    .A2(_3106_));
 sg13g2_a21oi_1 _3991_ (.A1(_3065_),
    .A2(_3103_),
    .Y(_3108_),
    .B1(_3107_));
 sg13g2_o21ai_1 _3992_ (.B1(_3108_),
    .Y(_3109_),
    .A1(_3065_),
    .A2(_3103_));
 sg13g2_nand3_1 _3993_ (.B(_2985_),
    .C(_3105_),
    .A(_2984_),
    .Y(_3110_));
 sg13g2_xnor2_1 _3994_ (.Y(_3111_),
    .A(_2987_),
    .B(_2988_));
 sg13g2_nor2_1 _3995_ (.A(_3067_),
    .B(net404),
    .Y(_3112_));
 sg13g2_xnor2_1 _3996_ (.Y(_3113_),
    .A(_3064_),
    .B(_3112_));
 sg13g2_a22oi_1 _3997_ (.Y(_3114_),
    .B1(_3111_),
    .B2(_3113_),
    .A2(_3110_),
    .A1(_3109_));
 sg13g2_xnor2_1 _3998_ (.Y(_3115_),
    .A(_2989_),
    .B(_2990_));
 sg13g2_nor2b_1 _3999_ (.A(net404),
    .B_N(_3068_),
    .Y(_3116_));
 sg13g2_xnor2_1 _4000_ (.Y(_3117_),
    .A(_3069_),
    .B(_3116_));
 sg13g2_or2_1 _4001_ (.X(_3118_),
    .B(_3117_),
    .A(_3115_));
 sg13g2_o21ai_1 _4002_ (.B1(_3118_),
    .Y(_3119_),
    .A1(_3111_),
    .A2(_3113_));
 sg13g2_a22oi_1 _4003_ (.Y(_3120_),
    .B1(_3115_),
    .B2(_3117_),
    .A2(_3102_),
    .A1(_2997_));
 sg13g2_o21ai_1 _4004_ (.B1(_3120_),
    .Y(_3121_),
    .A1(_3114_),
    .A2(_3119_));
 sg13g2_o21ai_1 _4005_ (.B1(_3121_),
    .Y(_3122_),
    .A1(_2997_),
    .A2(_3102_));
 sg13g2_xnor2_1 _4006_ (.Y(_3123_),
    .A(_3100_),
    .B(_3122_));
 sg13g2_inv_1 _4007_ (.Y(_3124_),
    .A(_3123_));
 sg13g2_nor2_1 _4008_ (.A(_3000_),
    .B(_3123_),
    .Y(_3125_));
 sg13g2_xnor2_1 _4009_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[0] ),
    .A(_3000_),
    .B(_3123_));
 sg13g2_nand2b_1 _4010_ (.Y(_3126_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ));
 sg13g2_nor2b_1 _4011_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ),
    .Y(_3127_));
 sg13g2_nand2b_1 _4012_ (.Y(_3128_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ));
 sg13g2_nand2b_1 _4013_ (.Y(_3129_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ));
 sg13g2_nand2_2 _4014_ (.Y(_3130_),
    .A(_3128_),
    .B(_3129_));
 sg13g2_nor2b_1 _4015_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ),
    .Y(_3131_));
 sg13g2_nand2b_1 _4016_ (.Y(_3132_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ));
 sg13g2_nand2b_1 _4017_ (.Y(_3133_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ));
 sg13g2_xor2_1 _4018_ (.B(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ),
    .X(_3134_));
 sg13g2_nor2b_1 _4019_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ),
    .Y(_3135_));
 sg13g2_nand2b_1 _4020_ (.Y(_3136_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ));
 sg13g2_nand2b_1 _4021_ (.Y(_3137_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ));
 sg13g2_nand2b_1 _4022_ (.Y(_3138_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ));
 sg13g2_nand2_2 _4023_ (.Y(_3139_),
    .A(_3137_),
    .B(_3138_));
 sg13g2_nor2b_1 _4024_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ),
    .Y(_3140_));
 sg13g2_nor2b_1 _4025_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ),
    .Y(_3141_));
 sg13g2_nand2b_1 _4026_ (.Y(_3142_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ));
 sg13g2_xnor2_1 _4027_ (.Y(_3143_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ));
 sg13g2_nand2b_1 _4028_ (.Y(_3144_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ));
 sg13g2_nand2b_1 _4029_ (.Y(_3145_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ));
 sg13g2_nand3b_1 _4030_ (.B(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ),
    .C(_3145_),
    .Y(_3146_),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ));
 sg13g2_and2_1 _4031_ (.A(_3144_),
    .B(_3146_),
    .X(_3147_));
 sg13g2_nand2_1 _4032_ (.Y(_3148_),
    .A(_3143_),
    .B(_3147_));
 sg13g2_a21oi_1 _4033_ (.A1(_3142_),
    .A2(_3148_),
    .Y(_3149_),
    .B1(_3140_));
 sg13g2_nor2_1 _4034_ (.A(_3141_),
    .B(_3149_),
    .Y(_3150_));
 sg13g2_o21ai_1 _4035_ (.B1(_3137_),
    .Y(_3151_),
    .A1(_3139_),
    .A2(_3150_));
 sg13g2_o21ai_1 _4036_ (.B1(_3136_),
    .Y(_3152_),
    .A1(_3135_),
    .A2(_3151_));
 sg13g2_nor2_1 _4037_ (.A(_3134_),
    .B(_3152_),
    .Y(_3153_));
 sg13g2_a21oi_1 _4038_ (.A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ),
    .A2(_2926_),
    .Y(_3154_),
    .B1(_3153_));
 sg13g2_o21ai_1 _4039_ (.B1(_3132_),
    .Y(_3155_),
    .A1(_3131_),
    .A2(_3154_));
 sg13g2_inv_1 _4040_ (.Y(_3156_),
    .A(_3155_));
 sg13g2_o21ai_1 _4041_ (.B1(_3128_),
    .Y(_3157_),
    .A1(_3130_),
    .A2(_3156_));
 sg13g2_a21oi_1 _4042_ (.A1(_3126_),
    .A2(_3157_),
    .Y(_3158_),
    .B1(_3127_));
 sg13g2_xnor2_1 _4043_ (.Y(_3159_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ));
 sg13g2_nor2b_1 _4044_ (.A(_3135_),
    .B_N(_3136_),
    .Y(_3160_));
 sg13g2_inv_1 _4045_ (.Y(_3161_),
    .A(_3160_));
 sg13g2_nand3b_1 _4046_ (.B(_3144_),
    .C(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .Y(_3162_),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_and2_1 _4047_ (.A(_3145_),
    .B(_3162_),
    .X(_3163_));
 sg13g2_nand2_1 _4048_ (.Y(_3164_),
    .A(_3143_),
    .B(_3163_));
 sg13g2_a21o_1 _4049_ (.A2(_3164_),
    .A1(_3149_),
    .B1(_3141_),
    .X(_3165_));
 sg13g2_nor2_1 _4050_ (.A(_3139_),
    .B(_3165_),
    .Y(_3166_));
 sg13g2_nor3_1 _4051_ (.A(_3139_),
    .B(_3161_),
    .C(_3165_),
    .Y(_3167_));
 sg13g2_nand2b_2 _4052_ (.Y(_3168_),
    .B(_3132_),
    .A_N(_3131_));
 sg13g2_nor2_1 _4053_ (.A(_3134_),
    .B(_3168_),
    .Y(_3169_));
 sg13g2_a21oi_1 _4054_ (.A1(_3167_),
    .A2(_3169_),
    .Y(_3170_),
    .B1(_3156_));
 sg13g2_nor2_1 _4055_ (.A(_3130_),
    .B(_3170_),
    .Y(_3171_));
 sg13g2_a21oi_1 _4056_ (.A1(_3159_),
    .A2(_3171_),
    .Y(_3172_),
    .B1(_3158_));
 sg13g2_nor2_1 _4057_ (.A(net490),
    .B(_3172_),
    .Y(_3173_));
 sg13g2_and2_1 _4058_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ),
    .X(_3174_));
 sg13g2_and2_1 _4059_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ),
    .X(_3175_));
 sg13g2_and2_1 _4060_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ),
    .X(_3176_));
 sg13g2_and2_1 _4061_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ),
    .X(_3177_));
 sg13g2_and2_1 _4062_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ),
    .X(_3178_));
 sg13g2_and2_1 _4063_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ),
    .X(_3179_));
 sg13g2_nor2_1 _4064_ (.A(_3140_),
    .B(_3141_),
    .Y(_3180_));
 sg13g2_inv_1 _4065_ (.Y(_3181_),
    .A(_3180_));
 sg13g2_nand2_1 _4066_ (.Y(_3182_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_a21oi_1 _4067_ (.A1(_3144_),
    .A2(_3145_),
    .Y(_3183_),
    .B1(_3182_));
 sg13g2_a21o_1 _4068_ (.A2(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ),
    .A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ),
    .B1(_3183_),
    .X(_3184_));
 sg13g2_nor2b_1 _4069_ (.A(_3143_),
    .B_N(_3184_),
    .Y(_3185_));
 sg13g2_a21o_1 _4070_ (.A2(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ),
    .A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ),
    .B1(_3185_),
    .X(_3186_));
 sg13g2_a21o_1 _4071_ (.A2(_3186_),
    .A1(_3181_),
    .B1(_3179_),
    .X(_3187_));
 sg13g2_a21o_1 _4072_ (.A2(_3187_),
    .A1(_3139_),
    .B1(_3178_),
    .X(_3188_));
 sg13g2_a21o_1 _4073_ (.A2(_3188_),
    .A1(_3161_),
    .B1(_3177_),
    .X(_3189_));
 sg13g2_a21o_1 _4074_ (.A2(_3189_),
    .A1(_3134_),
    .B1(_3176_),
    .X(_3190_));
 sg13g2_a21o_1 _4075_ (.A2(_3190_),
    .A1(_3168_),
    .B1(_3175_),
    .X(_3191_));
 sg13g2_a21o_1 _4076_ (.A2(_3191_),
    .A1(_3130_),
    .B1(_3174_),
    .X(_3192_));
 sg13g2_nor2b_1 _4077_ (.A(_3159_),
    .B_N(_3192_),
    .Y(_3193_));
 sg13g2_a21o_1 _4078_ (.A2(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ),
    .A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ),
    .B1(_3193_),
    .X(_3194_));
 sg13g2_a21oi_1 _4079_ (.A1(net490),
    .A2(_3194_),
    .Y(_3195_),
    .B1(_3173_));
 sg13g2_xor2_1 _4080_ (.B(_3195_),
    .A(net628),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ));
 sg13g2_inv_2 _4081_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .A(net402));
 sg13g2_xnor2_1 _4082_ (.Y(_3196_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_nand3_1 _4083_ (.B(_3145_),
    .C(_3182_),
    .A(_3144_),
    .Y(_3197_));
 sg13g2_nand2b_1 _4084_ (.Y(_3198_),
    .B(_3197_),
    .A_N(_3183_));
 sg13g2_nor2b_1 _4085_ (.A(net494),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .Y(_3199_));
 sg13g2_xnor2_1 _4086_ (.Y(_3200_),
    .A(_3198_),
    .B(_3199_));
 sg13g2_inv_1 _4087_ (.Y(_3201_),
    .A(_3200_));
 sg13g2_nand2_1 _4088_ (.Y(_3202_),
    .A(_3196_),
    .B(_3200_));
 sg13g2_xor2_1 _4089_ (.B(_3200_),
    .A(_3196_),
    .X(_3203_));
 sg13g2_nand2_1 _4090_ (.Y(_3204_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ),
    .B(net494));
 sg13g2_xor2_1 _4091_ (.B(_3204_),
    .A(_3198_),
    .X(_3205_));
 sg13g2_inv_1 _4092_ (.Y(_3206_),
    .A(_3205_));
 sg13g2_nand2_1 _4093_ (.Y(_3207_),
    .A(net396),
    .B(_3205_));
 sg13g2_xor2_1 _4094_ (.B(_3184_),
    .A(_3143_),
    .X(_3208_));
 sg13g2_inv_1 _4095_ (.Y(_3209_),
    .A(_3208_));
 sg13g2_xnor2_1 _4096_ (.Y(_3210_),
    .A(_3143_),
    .B(_3147_));
 sg13g2_nor2_1 _4097_ (.A(_2925_),
    .B(_3210_),
    .Y(_3211_));
 sg13g2_a21oi_2 _4098_ (.B1(_3211_),
    .Y(_3212_),
    .A2(_3209_),
    .A1(_2925_));
 sg13g2_xnor2_1 _4099_ (.Y(_3213_),
    .A(_3207_),
    .B(_3212_));
 sg13g2_nor2_1 _4100_ (.A(_3201_),
    .B(_3213_),
    .Y(_3214_));
 sg13g2_nand2b_1 _4101_ (.Y(_3215_),
    .B(_3205_),
    .A_N(_3196_));
 sg13g2_inv_1 _4102_ (.Y(_3216_),
    .A(_3215_));
 sg13g2_xnor2_1 _4103_ (.Y(_3217_),
    .A(_3200_),
    .B(_3213_));
 sg13g2_a21oi_1 _4104_ (.A1(_3216_),
    .A2(_3217_),
    .Y(_3218_),
    .B1(_3214_));
 sg13g2_inv_1 _4105_ (.Y(_3219_),
    .A(_3218_));
 sg13g2_or2_1 _4106_ (.X(_3220_),
    .B(_3163_),
    .A(_3143_));
 sg13g2_a21oi_1 _4107_ (.A1(_3143_),
    .A2(_3163_),
    .Y(_3221_),
    .B1(net493));
 sg13g2_a22oi_1 _4108_ (.Y(_3222_),
    .B1(_3220_),
    .B2(_3221_),
    .A2(_3209_),
    .A1(net493));
 sg13g2_nand2_1 _4109_ (.Y(_3223_),
    .A(_3206_),
    .B(_3212_));
 sg13g2_nand2_1 _4110_ (.Y(_3224_),
    .A(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .B(_3223_));
 sg13g2_nor2_1 _4111_ (.A(net493),
    .B(_3186_),
    .Y(_3225_));
 sg13g2_a21oi_1 _4112_ (.A1(_3142_),
    .A2(_3148_),
    .Y(_3226_),
    .B1(_2925_));
 sg13g2_nor2_1 _4113_ (.A(_3225_),
    .B(_3226_),
    .Y(_3227_));
 sg13g2_xnor2_1 _4114_ (.Y(_3228_),
    .A(_3180_),
    .B(_3227_));
 sg13g2_inv_1 _4115_ (.Y(_3229_),
    .A(_3228_));
 sg13g2_xnor2_1 _4116_ (.Y(_3230_),
    .A(_3224_),
    .B(_3229_));
 sg13g2_nor2_1 _4117_ (.A(_3222_),
    .B(_3230_),
    .Y(_3231_));
 sg13g2_xor2_1 _4118_ (.B(_3230_),
    .A(_3222_),
    .X(_3232_));
 sg13g2_xnor2_1 _4119_ (.Y(_3233_),
    .A(_3218_),
    .B(_3232_));
 sg13g2_nand2_1 _4120_ (.Y(_3234_),
    .A(_3203_),
    .B(_3233_));
 sg13g2_xnor2_1 _4121_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[0] ),
    .A(_3203_),
    .B(_3233_));
 sg13g2_nand2_2 _4122_ (.Y(_3235_),
    .A(net478),
    .B(\main.demo._q_frame[6] ));
 sg13g2_nor2_1 _4123_ (.A(_0059_),
    .B(_3235_),
    .Y(_3236_));
 sg13g2_and2_1 _4124_ (.A(\main.demo._q_frame[6] ),
    .B(\main.demo._q_frame[5] ),
    .X(_3237_));
 sg13g2_xor2_1 _4125_ (.B(\main.demo._q_frame[5] ),
    .A(\main.demo._q_frame[6] ),
    .X(_3238_));
 sg13g2_a21oi_1 _4126_ (.A1(\main.demo._q_frame[4] ),
    .A2(net447),
    .Y(_3239_),
    .B1(_2913_));
 sg13g2_o21ai_1 _4127_ (.B1(_3239_),
    .Y(_3240_),
    .A1(\main.demo._q_frame[4] ),
    .A2(net447));
 sg13g2_nor2_1 _4128_ (.A(_0060_),
    .B(_3240_),
    .Y(_3241_));
 sg13g2_xor2_1 _4129_ (.B(_3235_),
    .A(\main.demo._w_vga_vga_y[8] ),
    .X(_3242_));
 sg13g2_nand2_1 _4130_ (.Y(_3243_),
    .A(_3241_),
    .B(_3242_));
 sg13g2_xnor2_1 _4131_ (.Y(_3244_),
    .A(_3241_),
    .B(_3242_));
 sg13g2_a21oi_1 _4132_ (.A1(net501),
    .A2(net447),
    .Y(_3245_),
    .B1(_2913_));
 sg13g2_o21ai_1 _4133_ (.B1(_3245_),
    .Y(_3246_),
    .A1(net501),
    .A2(net447));
 sg13g2_nand2b_1 _4134_ (.Y(_3247_),
    .B(_2934_),
    .A_N(_3246_));
 sg13g2_xnor2_1 _4135_ (.Y(_3248_),
    .A(_2934_),
    .B(_3246_));
 sg13g2_a21oi_1 _4136_ (.A1(net502),
    .A2(net447),
    .Y(_3249_),
    .B1(_2913_));
 sg13g2_o21ai_1 _4137_ (.B1(_3249_),
    .Y(_3250_),
    .A1(net502),
    .A2(net447));
 sg13g2_nor2_1 _4138_ (.A(_0062_),
    .B(_3250_),
    .Y(_3251_));
 sg13g2_xnor2_1 _4139_ (.Y(_3252_),
    .A(_3248_),
    .B(_3251_));
 sg13g2_xor2_1 _4140_ (.B(net447),
    .A(\main.demo._q_frame[1] ),
    .X(_3253_));
 sg13g2_a21oi_2 _4141_ (.B1(\main.demo._w_vga_vga_y[4] ),
    .Y(_3254_),
    .A2(_3253_),
    .A1(net478));
 sg13g2_xor2_1 _4142_ (.B(_3250_),
    .A(_0062_),
    .X(_3255_));
 sg13g2_inv_1 _4143_ (.Y(_3256_),
    .A(_3255_));
 sg13g2_a21oi_1 _4144_ (.A1(\main.demo._q_frame[0] ),
    .A2(net448),
    .Y(_3257_),
    .B1(_2913_));
 sg13g2_o21ai_1 _4145_ (.B1(_3257_),
    .Y(_3258_),
    .A1(\main.demo._q_frame[0] ),
    .A2(net448));
 sg13g2_nor2_1 _4146_ (.A(net638),
    .B(_3258_),
    .Y(_3259_));
 sg13g2_nand3_1 _4147_ (.B(\main.demo._w_vga_vga_y[4] ),
    .C(_3253_),
    .A(\main.demo._q_rot_en ),
    .Y(_3260_));
 sg13g2_nand2b_1 _4148_ (.Y(_3261_),
    .B(_3260_),
    .A_N(_3254_));
 sg13g2_nand2_1 _4149_ (.Y(_3262_),
    .A(_3259_),
    .B(_3261_));
 sg13g2_xor2_1 _4150_ (.B(_3261_),
    .A(_3259_),
    .X(_3263_));
 sg13g2_xnor2_1 _4151_ (.Y(_3264_),
    .A(_3254_),
    .B(_3255_));
 sg13g2_xnor2_1 _4152_ (.Y(_3265_),
    .A(_3262_),
    .B(_3264_));
 sg13g2_or2_1 _4153_ (.X(_3266_),
    .B(_3265_),
    .A(_3263_));
 sg13g2_o21ai_1 _4154_ (.B1(_3266_),
    .Y(_3267_),
    .A1(_3254_),
    .A2(_3256_));
 sg13g2_nor2b_1 _4155_ (.A(_3252_),
    .B_N(_3267_),
    .Y(_3268_));
 sg13g2_xor2_1 _4156_ (.B(_3240_),
    .A(_0060_),
    .X(_3269_));
 sg13g2_a21o_1 _4157_ (.A2(_3251_),
    .A1(_3248_),
    .B1(_3268_),
    .X(_3270_));
 sg13g2_nand2_1 _4158_ (.Y(_3271_),
    .A(_3269_),
    .B(_3270_));
 sg13g2_nand2_1 _4159_ (.Y(_3272_),
    .A(_3247_),
    .B(_3271_));
 sg13g2_o21ai_1 _4160_ (.B1(_3272_),
    .Y(_3273_),
    .A1(_3268_),
    .A2(_3269_));
 sg13g2_xor2_1 _4161_ (.B(_3273_),
    .A(_3244_),
    .X(_3274_));
 sg13g2_o21ai_1 _4162_ (.B1(_3243_),
    .Y(_3275_),
    .A1(_3244_),
    .A2(_3273_));
 sg13g2_a21oi_1 _4163_ (.A1(\main.demo._w_vga_vga_y[8] ),
    .A2(_3235_),
    .Y(_3276_),
    .B1(\main.demo._w_vga_vga_y[10] ));
 sg13g2_nand3_1 _4164_ (.B(\main.demo._w_vga_vga_y[8] ),
    .C(_3235_),
    .A(\main.demo._w_vga_vga_y[10] ),
    .Y(_3277_));
 sg13g2_nand2b_1 _4165_ (.Y(_3278_),
    .B(_3277_),
    .A_N(_3276_));
 sg13g2_xor2_1 _4166_ (.B(_3278_),
    .A(_3275_),
    .X(_3279_));
 sg13g2_nor2_1 _4167_ (.A(_3274_),
    .B(_3279_),
    .Y(_3280_));
 sg13g2_a22oi_1 _4168_ (.Y(_3281_),
    .B1(_3243_),
    .B2(_3276_),
    .A2(_3235_),
    .A1(\main.demo._w_vga_vga_y[10] ));
 sg13g2_nor2_1 _4169_ (.A(_3280_),
    .B(_3281_),
    .Y(_3282_));
 sg13g2_xnor2_1 _4170_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ),
    .A(_3236_),
    .B(_3282_));
 sg13g2_nand2_1 _4171_ (.Y(_3283_),
    .A(net478),
    .B(net500));
 sg13g2_nor2_1 _4172_ (.A(_0053_),
    .B(_3283_),
    .Y(_3284_));
 sg13g2_xor2_1 _4173_ (.B(_3283_),
    .A(_0053_),
    .X(_3285_));
 sg13g2_a21oi_1 _4174_ (.A1(net500),
    .A2(net447),
    .Y(_3286_),
    .B1(_2913_));
 sg13g2_o21ai_1 _4175_ (.B1(_3286_),
    .Y(_3287_),
    .A1(net500),
    .A2(net448));
 sg13g2_nand2_1 _4176_ (.Y(_3288_),
    .A(_0054_),
    .B(_3287_));
 sg13g2_and2_1 _4177_ (.A(_3285_),
    .B(_3288_),
    .X(_3289_));
 sg13g2_xor2_1 _4178_ (.B(\main.demo._q_frame[6] ),
    .A(net500),
    .X(_3290_));
 sg13g2_a21oi_1 _4179_ (.A1(\main.demo._q_frame[4] ),
    .A2(_3290_),
    .Y(_3291_),
    .B1(_2913_));
 sg13g2_o21ai_1 _4180_ (.B1(_3291_),
    .Y(_3292_),
    .A1(\main.demo._q_frame[4] ),
    .A2(_3290_));
 sg13g2_nand2_1 _4181_ (.Y(_3293_),
    .A(_0055_),
    .B(_3292_));
 sg13g2_xnor2_1 _4182_ (.Y(_3294_),
    .A(_2928_),
    .B(_3287_));
 sg13g2_nand2_1 _4183_ (.Y(_3295_),
    .A(_3293_),
    .B(_3294_));
 sg13g2_xor2_1 _4184_ (.B(_3294_),
    .A(_3293_),
    .X(_3296_));
 sg13g2_inv_1 _4185_ (.Y(_3297_),
    .A(_3296_));
 sg13g2_a21oi_1 _4186_ (.A1(net501),
    .A2(_3290_),
    .Y(_3298_),
    .B1(_2913_));
 sg13g2_o21ai_1 _4187_ (.B1(_3298_),
    .Y(_3299_),
    .A1(net501),
    .A2(_3290_));
 sg13g2_o21ai_1 _4188_ (.B1(net478),
    .Y(_3300_),
    .A1(net502),
    .A2(_3290_));
 sg13g2_a21oi_1 _4189_ (.A1(net502),
    .A2(_3290_),
    .Y(_3301_),
    .B1(_3300_));
 sg13g2_nand2b_1 _4190_ (.Y(_3302_),
    .B(_3301_),
    .A_N(_0057_));
 sg13g2_o21ai_1 _4191_ (.B1(net478),
    .Y(_3303_),
    .A1(\main.demo._q_frame[1] ),
    .A2(_3290_));
 sg13g2_a21oi_1 _4192_ (.A1(\main.demo._q_frame[1] ),
    .A2(_3290_),
    .Y(_3304_),
    .B1(_3303_));
 sg13g2_nor2b_1 _4193_ (.A(_0058_),
    .B_N(_3304_),
    .Y(_3305_));
 sg13g2_xnor2_1 _4194_ (.Y(_3306_),
    .A(_0057_),
    .B(_3301_));
 sg13g2_nand2_1 _4195_ (.Y(_3307_),
    .A(_3305_),
    .B(_3306_));
 sg13g2_xnor2_1 _4196_ (.Y(_3308_),
    .A(_0056_),
    .B(_3299_));
 sg13g2_a21o_1 _4197_ (.A2(_3307_),
    .A1(_3302_),
    .B1(_3308_),
    .X(_3309_));
 sg13g2_o21ai_1 _4198_ (.B1(_3309_),
    .Y(_3310_),
    .A1(_0056_),
    .A2(_3299_));
 sg13g2_xor2_1 _4199_ (.B(_3292_),
    .A(\main.demo._w_vga_vga_x[6] ),
    .X(_3311_));
 sg13g2_nand2_1 _4200_ (.Y(_3312_),
    .A(_3310_),
    .B(_3311_));
 sg13g2_o21ai_1 _4201_ (.B1(_3295_),
    .Y(_3313_),
    .A1(_3297_),
    .A2(_3312_));
 sg13g2_xor2_1 _4202_ (.B(_3288_),
    .A(_3285_),
    .X(_3314_));
 sg13g2_a21o_1 _4203_ (.A2(_3314_),
    .A1(_3313_),
    .B1(_3289_),
    .X(_3315_));
 sg13g2_nand3_1 _4204_ (.B(net500),
    .C(_0053_),
    .A(net478),
    .Y(_3316_));
 sg13g2_xor2_1 _4205_ (.B(_3316_),
    .A(\main.demo._w_vga_vga_x[9] ),
    .X(_3317_));
 sg13g2_a22oi_1 _4206_ (.Y(_3318_),
    .B1(_3315_),
    .B2(_3317_),
    .A2(_3284_),
    .A1(\main.demo._w_vga_vga_x[9] ));
 sg13g2_a21oi_1 _4207_ (.A1(net478),
    .A2(net500),
    .Y(_3319_),
    .B1(_0052_));
 sg13g2_xor2_1 _4208_ (.B(_3319_),
    .A(\main.demo._w_vga_vga_x[10] ),
    .X(_3320_));
 sg13g2_xnor2_1 _4209_ (.Y(_3321_),
    .A(_3318_),
    .B(_3320_));
 sg13g2_nor2b_2 _4210_ (.A(net397),
    .B_N(_3321_),
    .Y(_3322_));
 sg13g2_inv_2 _4211_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .A(net395));
 sg13g2_nor2_1 _4212_ (.A(\main.demo.vga._q_xcount[5] ),
    .B(\main.demo.vga._q_xcount[4] ),
    .Y(_3323_));
 sg13g2_and2_1 _4213_ (.A(\main.demo.vga._q_xcount[7] ),
    .B(_3323_),
    .X(_3324_));
 sg13g2_nor2_1 _4214_ (.A(net319),
    .B(net317),
    .Y(_3325_));
 sg13g2_nor4_2 _4215_ (.A(\main.demo.vga._q_xcount[1] ),
    .B(\main.demo.vga._q_xcount[0] ),
    .C(\main.demo.vga._q_xcount[3] ),
    .Y(_3326_),
    .D(\main.demo.vga._q_xcount[2] ));
 sg13g2_inv_1 _4216_ (.Y(_3327_),
    .A(_3326_));
 sg13g2_nor2_1 _4217_ (.A(\main.demo.vga._q_xcount[6] ),
    .B(\main.demo.vga._q_xcount[10] ),
    .Y(_0229_));
 sg13g2_nor2b_1 _4218_ (.A(\main.demo.vga._q_xcount[8] ),
    .B_N(\main.demo.vga._q_xcount[9] ),
    .Y(_0230_));
 sg13g2_and4_1 _4219_ (.A(_3324_),
    .B(_3326_),
    .C(_0229_),
    .D(_0230_),
    .X(_0231_));
 sg13g2_nor3_1 _4220_ (.A(\main.demo.vga._q_xcount[7] ),
    .B(\main.demo.vga._q_xcount[9] ),
    .C(\main.demo.vga._q_xcount[8] ),
    .Y(_0232_));
 sg13g2_nand4_1 _4221_ (.B(_3326_),
    .C(_0229_),
    .A(_3323_),
    .Y(_0233_),
    .D(_0232_));
 sg13g2_o21ai_1 _4222_ (.B1(_0233_),
    .Y(_0234_),
    .A1(_2937_),
    .A2(_0231_));
 sg13g2_inv_1 _4223_ (.Y(_0235_),
    .A(net422));
 sg13g2_and3_1 _4224_ (.X(_0236_),
    .A(net320),
    .B(\main.demo.vga._q_ycount[7] ),
    .C(net593));
 sg13g2_nor4_2 _4225_ (.A(net364),
    .B(\main.demo.vga._q_ycount[2] ),
    .C(net514),
    .Y(_0237_),
    .D(net527));
 sg13g2_nor2_1 _4226_ (.A(\main.demo.vga._q_ycount[4] ),
    .B(\main.demo.vga._d_vblank ),
    .Y(_0238_));
 sg13g2_and2_1 _4227_ (.A(net334),
    .B(_0238_),
    .X(_0239_));
 sg13g2_nand3_1 _4228_ (.B(_0237_),
    .C(_0239_),
    .A(_0236_),
    .Y(_0240_));
 sg13g2_nor4_1 _4229_ (.A(\main.demo.vga._q_ycount[8] ),
    .B(\main.demo.vga._q_ycount[7] ),
    .C(\main.demo.vga._q_ycount[6] ),
    .D(\main.demo.vga._q_ycount[5] ),
    .Y(_0241_));
 sg13g2_and2_1 _4230_ (.A(_0238_),
    .B(_0241_),
    .X(_0242_));
 sg13g2_a22oi_1 _4231_ (.Y(_0243_),
    .B1(_0242_),
    .B2(_0237_),
    .A2(_0240_),
    .A1(net314));
 sg13g2_nor2_1 _4232_ (.A(_0235_),
    .B(net421),
    .Y(\main.demo.vga._d_active ));
 sg13g2_nor2_1 _4233_ (.A(net644),
    .B(net401),
    .Y(_0244_));
 sg13g2_a21oi_1 _4234_ (.A1(_2939_),
    .A2(net401),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[0] ),
    .B1(_0244_));
 sg13g2_xor2_1 _4235_ (.B(\main.demo._t___stage___block_3_x[1] ),
    .A(\main.demo._t___stage___block_3_x[0] ),
    .X(_0245_));
 sg13g2_nand2_1 _4236_ (.Y(_0246_),
    .A(net401),
    .B(_0245_));
 sg13g2_nor2_1 _4237_ (.A(_2938_),
    .B(_3321_),
    .Y(_0247_));
 sg13g2_xnor2_1 _4238_ (.Y(_0248_),
    .A(net643),
    .B(_0247_));
 sg13g2_o21ai_1 _4239_ (.B1(_0246_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[1] ),
    .A1(net401),
    .A2(_0248_));
 sg13g2_nor3_2 _4240_ (.A(\main.demo._t___stage___block_3_x[0] ),
    .B(\main.demo._t___stage___block_3_x[1] ),
    .C(\main.demo._t___stage___block_3_x[2] ),
    .Y(_0249_));
 sg13g2_o21ai_1 _4241_ (.B1(\main.demo._t___stage___block_3_x[2] ),
    .Y(_0250_),
    .A1(\main.demo._t___stage___block_3_x[0] ),
    .A2(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_nor2b_1 _4242_ (.A(_0249_),
    .B_N(_0250_),
    .Y(_0251_));
 sg13g2_nand2_1 _4243_ (.Y(_0252_),
    .A(net400),
    .B(_0251_));
 sg13g2_nor2_1 _4244_ (.A(\main.demo._t___stage___block_3_y[0] ),
    .B(\main.demo._t___stage___block_3_y[1] ),
    .Y(_0253_));
 sg13g2_nor2_1 _4245_ (.A(_3321_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_xor2_1 _4246_ (.B(_0254_),
    .A(net588),
    .X(_0255_));
 sg13g2_o21ai_1 _4247_ (.B1(_0252_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[2] ),
    .A1(net400),
    .A2(_0255_));
 sg13g2_xnor2_1 _4248_ (.Y(_0256_),
    .A(_0058_),
    .B(_3304_));
 sg13g2_nor2b_1 _4249_ (.A(_0256_),
    .B_N(_0249_),
    .Y(_0257_));
 sg13g2_xnor2_1 _4250_ (.Y(_0258_),
    .A(_0249_),
    .B(_0256_));
 sg13g2_xor2_1 _4251_ (.B(_3258_),
    .A(net626),
    .X(_0259_));
 sg13g2_a21oi_1 _4252_ (.A1(_2942_),
    .A2(_0253_),
    .Y(_0260_),
    .B1(_3321_));
 sg13g2_xor2_1 _4253_ (.B(_0260_),
    .A(_0259_),
    .X(_0261_));
 sg13g2_mux2_1 _4254_ (.A0(_0261_),
    .A1(_0258_),
    .S(net400),
    .X(\main.demo._t___pip_58_1_0___stage___block_3_cy[3] ));
 sg13g2_xor2_1 _4255_ (.B(_3306_),
    .A(_3305_),
    .X(_0262_));
 sg13g2_nand2b_1 _4256_ (.Y(_0263_),
    .B(_0257_),
    .A_N(_0262_));
 sg13g2_xnor2_1 _4257_ (.Y(_0264_),
    .A(_0257_),
    .B(_0262_));
 sg13g2_nand2_1 _4258_ (.Y(_0265_),
    .A(net398),
    .B(_0264_));
 sg13g2_nand3b_1 _4259_ (.B(_0253_),
    .C(net588),
    .Y(_0266_),
    .A_N(_0259_));
 sg13g2_nor2b_1 _4260_ (.A(_3321_),
    .B_N(_0266_),
    .Y(_0267_));
 sg13g2_xnor2_1 _4261_ (.Y(_0268_),
    .A(_3263_),
    .B(_0267_));
 sg13g2_o21ai_1 _4262_ (.B1(_0265_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[4] ),
    .A1(net399),
    .A2(_0268_));
 sg13g2_o21ai_1 _4263_ (.B1(_3265_),
    .Y(_0269_),
    .A1(_3263_),
    .A2(_0266_));
 sg13g2_nor2_1 _4264_ (.A(_3266_),
    .B(_0266_),
    .Y(_0270_));
 sg13g2_nor2_1 _4265_ (.A(_3321_),
    .B(_0270_),
    .Y(_0271_));
 sg13g2_nand2_1 _4266_ (.Y(_0272_),
    .A(_0269_),
    .B(_0271_));
 sg13g2_nand3_1 _4267_ (.B(_3307_),
    .C(_3308_),
    .A(_3302_),
    .Y(_0273_));
 sg13g2_and2_1 _4268_ (.A(_3309_),
    .B(_0273_),
    .X(_0274_));
 sg13g2_nor2_1 _4269_ (.A(_0263_),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_xor2_1 _4270_ (.B(_0274_),
    .A(_0263_),
    .X(_0276_));
 sg13g2_nor2_1 _4271_ (.A(net397),
    .B(_3321_),
    .Y(_0277_));
 sg13g2_inv_1 _4272_ (.Y(_0278_),
    .A(net393));
 sg13g2_a22oi_1 _4273_ (.Y(_0279_),
    .B1(_0276_),
    .B2(net398),
    .A2(_3322_),
    .A1(_3265_));
 sg13g2_o21ai_1 _4274_ (.B1(_0279_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[5] ),
    .A1(net398),
    .A2(_0272_));
 sg13g2_xnor2_1 _4275_ (.Y(_0280_),
    .A(_3310_),
    .B(_3311_));
 sg13g2_nand2_1 _4276_ (.Y(_0281_),
    .A(_0275_),
    .B(_0280_));
 sg13g2_xor2_1 _4277_ (.B(_0280_),
    .A(_0275_),
    .X(_0282_));
 sg13g2_xor2_1 _4278_ (.B(_3267_),
    .A(_3252_),
    .X(_0283_));
 sg13g2_inv_1 _4279_ (.Y(_0284_),
    .A(_0283_));
 sg13g2_xnor2_1 _4280_ (.Y(_0285_),
    .A(_0271_),
    .B(_0284_));
 sg13g2_nand2_1 _4281_ (.Y(_0286_),
    .A(net398),
    .B(_0282_));
 sg13g2_o21ai_1 _4282_ (.B1(_0286_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[6] ),
    .A1(net398),
    .A2(_0285_));
 sg13g2_xnor2_1 _4283_ (.Y(_0287_),
    .A(_3247_),
    .B(_3269_));
 sg13g2_xnor2_1 _4284_ (.Y(_0288_),
    .A(_3270_),
    .B(_0287_));
 sg13g2_inv_1 _4285_ (.Y(_0289_),
    .A(_0288_));
 sg13g2_nand3_1 _4286_ (.B(_0283_),
    .C(_0288_),
    .A(_0270_),
    .Y(_0290_));
 sg13g2_inv_1 _4287_ (.Y(_0291_),
    .A(_0290_));
 sg13g2_a21oi_1 _4288_ (.A1(_0270_),
    .A2(_0283_),
    .Y(_0292_),
    .B1(_0288_));
 sg13g2_nand2b_1 _4289_ (.Y(_0293_),
    .B(net393),
    .A_N(_0292_));
 sg13g2_xnor2_1 _4290_ (.Y(_0294_),
    .A(_3297_),
    .B(_3312_));
 sg13g2_nor2b_1 _4291_ (.A(_0281_),
    .B_N(_0294_),
    .Y(_0295_));
 sg13g2_xnor2_1 _4292_ (.Y(_0296_),
    .A(_0281_),
    .B(_0294_));
 sg13g2_a22oi_1 _4293_ (.Y(_0297_),
    .B1(_0296_),
    .B2(net399),
    .A2(_0289_),
    .A1(net395));
 sg13g2_o21ai_1 _4294_ (.B1(_0297_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[7] ),
    .A1(_0291_),
    .A2(_0293_));
 sg13g2_xnor2_1 _4295_ (.Y(_0298_),
    .A(_3274_),
    .B(_0290_));
 sg13g2_xor2_1 _4296_ (.B(_3314_),
    .A(_3313_),
    .X(_0299_));
 sg13g2_nor2b_1 _4297_ (.A(_0299_),
    .B_N(_0295_),
    .Y(_0300_));
 sg13g2_xnor2_1 _4298_ (.Y(_0301_),
    .A(_0295_),
    .B(_0299_));
 sg13g2_a22oi_1 _4299_ (.Y(_0302_),
    .B1(_0301_),
    .B2(net397),
    .A2(net395),
    .A1(_3274_));
 sg13g2_o21ai_1 _4300_ (.B1(_0302_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[8] ),
    .A1(_0278_),
    .A2(_0298_));
 sg13g2_o21ai_1 _4301_ (.B1(_3279_),
    .Y(_0303_),
    .A1(_3274_),
    .A2(_0290_));
 sg13g2_a21oi_1 _4302_ (.A1(_3280_),
    .A2(_0291_),
    .Y(_0304_),
    .B1(_0278_));
 sg13g2_xor2_1 _4303_ (.B(_3317_),
    .A(_3315_),
    .X(_0305_));
 sg13g2_nand2b_1 _4304_ (.Y(_0306_),
    .B(_0300_),
    .A_N(_0305_));
 sg13g2_xnor2_1 _4305_ (.Y(_0307_),
    .A(_0300_),
    .B(_0305_));
 sg13g2_nand2_1 _4306_ (.Y(_0308_),
    .A(net397),
    .B(_0307_));
 sg13g2_a22oi_1 _4307_ (.Y(_0309_),
    .B1(_0303_),
    .B2(_0304_),
    .A2(net395),
    .A1(_3279_));
 sg13g2_nand2_1 _4308_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[9] ),
    .A(_0308_),
    .B(_0309_));
 sg13g2_xor2_1 _4309_ (.B(_0306_),
    .A(_3321_),
    .X(_0310_));
 sg13g2_a21oi_1 _4310_ (.A1(net397),
    .A2(_0310_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[10] ),
    .B1(_0304_));
 sg13g2_nor2_1 _4311_ (.A(net648),
    .B(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .Y(_0311_));
 sg13g2_a221oi_1 _4312_ (.B2(\main.demo._t___stage___block_3_x[0] ),
    .C1(_0311_),
    .B1(net394),
    .A1(\main.demo._t___stage___block_3_y[0] ),
    .Y(_0312_),
    .A2(net400));
 sg13g2_inv_1 _4313_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[0] ),
    .A(_0312_));
 sg13g2_a22oi_1 _4314_ (.Y(_0313_),
    .B1(_0245_),
    .B2(net394),
    .A2(net400),
    .A1(\main.demo._t___stage___block_3_y[1] ));
 sg13g2_o21ai_1 _4315_ (.B1(_0313_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[1] ),
    .A1(net323),
    .A2(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ));
 sg13g2_nand2_1 _4316_ (.Y(_0314_),
    .A(net567),
    .B(net400));
 sg13g2_a22oi_1 _4317_ (.Y(_0315_),
    .B1(_0251_),
    .B2(net394),
    .A2(net395),
    .A1(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_nand2_1 _4318_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[2] ),
    .A(_0314_),
    .B(_0315_));
 sg13g2_nand2_1 _4319_ (.Y(_0316_),
    .A(net400),
    .B(_0259_));
 sg13g2_a22oi_1 _4320_ (.Y(_0317_),
    .B1(_0258_),
    .B2(net393),
    .A2(_0256_),
    .A1(_3322_));
 sg13g2_nand2_1 _4321_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[3] ),
    .A(_0316_),
    .B(_0317_));
 sg13g2_nand2_1 _4322_ (.Y(_0318_),
    .A(_3263_),
    .B(net398));
 sg13g2_a22oi_1 _4323_ (.Y(_0319_),
    .B1(_0264_),
    .B2(net394),
    .A2(_0262_),
    .A1(net395));
 sg13g2_nand2_1 _4324_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[4] ),
    .A(_0318_),
    .B(_0319_));
 sg13g2_nand2_1 _4325_ (.Y(_0320_),
    .A(_3265_),
    .B(net398));
 sg13g2_a22oi_1 _4326_ (.Y(_0321_),
    .B1(_0276_),
    .B2(net393),
    .A2(_0274_),
    .A1(_3322_));
 sg13g2_nand2_1 _4327_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[5] ),
    .A(_0320_),
    .B(_0321_));
 sg13g2_a22oi_1 _4328_ (.Y(_0322_),
    .B1(_0284_),
    .B2(net398),
    .A2(_0282_),
    .A1(net393));
 sg13g2_o21ai_1 _4329_ (.B1(_0322_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[6] ),
    .A1(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .A2(_0280_));
 sg13g2_a22oi_1 _4330_ (.Y(_0323_),
    .B1(_0296_),
    .B2(net393),
    .A2(_0289_),
    .A1(net397));
 sg13g2_o21ai_1 _4331_ (.B1(_0323_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[7] ),
    .A1(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .A2(_0294_));
 sg13g2_nand2_1 _4332_ (.Y(_0324_),
    .A(_3274_),
    .B(net397));
 sg13g2_a22oi_1 _4333_ (.Y(_0325_),
    .B1(_0301_),
    .B2(net393),
    .A2(_0299_),
    .A1(net395));
 sg13g2_nand2_1 _4334_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[8] ),
    .A(_0324_),
    .B(_0325_));
 sg13g2_nand2_1 _4335_ (.Y(_0326_),
    .A(_3279_),
    .B(net397));
 sg13g2_a22oi_1 _4336_ (.Y(_0327_),
    .B1(_0307_),
    .B2(net393),
    .A2(_0305_),
    .A1(net395));
 sg13g2_nand2_1 _4337_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[9] ),
    .A(_0326_),
    .B(_0327_));
 sg13g2_nor2_1 _4338_ (.A(_0278_),
    .B(_0306_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[10] ));
 sg13g2_nor2_1 _4339_ (.A(_3223_),
    .B(_3228_),
    .Y(_0328_));
 sg13g2_xnor2_1 _4340_ (.Y(_0329_),
    .A(_3139_),
    .B(_3187_));
 sg13g2_inv_1 _4341_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_nor2_1 _4342_ (.A(net493),
    .B(_0329_),
    .Y(_0331_));
 sg13g2_xor2_1 _4343_ (.B(_3150_),
    .A(_3139_),
    .X(_0332_));
 sg13g2_a21oi_2 _4344_ (.B1(_0331_),
    .Y(_0333_),
    .A2(_0332_),
    .A1(net493));
 sg13g2_nand2_1 _4345_ (.Y(_0334_),
    .A(_0328_),
    .B(_0333_));
 sg13g2_nor2_1 _4346_ (.A(net492),
    .B(_3188_),
    .Y(_0335_));
 sg13g2_a21oi_1 _4347_ (.A1(net492),
    .A2(_3151_),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_xnor2_1 _4348_ (.Y(_0337_),
    .A(_3160_),
    .B(_0336_));
 sg13g2_inv_1 _4349_ (.Y(_0338_),
    .A(_0337_));
 sg13g2_nor2_1 _4350_ (.A(_0334_),
    .B(_0337_),
    .Y(_0339_));
 sg13g2_xnor2_1 _4351_ (.Y(_0340_),
    .A(_3134_),
    .B(_3189_));
 sg13g2_inv_1 _4352_ (.Y(_0341_),
    .A(_0340_));
 sg13g2_nand2_1 _4353_ (.Y(_0342_),
    .A(_3134_),
    .B(_3152_));
 sg13g2_nor2_1 _4354_ (.A(_2925_),
    .B(_3153_),
    .Y(_0343_));
 sg13g2_a22oi_1 _4355_ (.Y(_0344_),
    .B1(_0342_),
    .B2(_0343_),
    .A2(_0341_),
    .A1(_2925_));
 sg13g2_nand2_1 _4356_ (.Y(_0345_),
    .A(_0339_),
    .B(_0344_));
 sg13g2_mux2_1 _4357_ (.A0(_3154_),
    .A1(_3190_),
    .S(_2925_),
    .X(_0346_));
 sg13g2_xor2_1 _4358_ (.B(_0346_),
    .A(_3168_),
    .X(_0347_));
 sg13g2_inv_1 _4359_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_nor2_1 _4360_ (.A(_0345_),
    .B(_0347_),
    .Y(_0349_));
 sg13g2_xor2_1 _4361_ (.B(_3191_),
    .A(_3130_),
    .X(_0350_));
 sg13g2_and2_1 _4362_ (.A(_2925_),
    .B(_0350_),
    .X(_0351_));
 sg13g2_xnor2_1 _4363_ (.Y(_0352_),
    .A(_3130_),
    .B(_3155_));
 sg13g2_a21oi_2 _4364_ (.B1(_0351_),
    .Y(_0353_),
    .A2(_0352_),
    .A1(net491));
 sg13g2_nand2_1 _4365_ (.Y(_0354_),
    .A(_0349_),
    .B(_0353_));
 sg13g2_nor2_1 _4366_ (.A(net490),
    .B(_3192_),
    .Y(_0355_));
 sg13g2_a21oi_1 _4367_ (.A1(net490),
    .A2(_3157_),
    .Y(_0356_),
    .B1(_0355_));
 sg13g2_xnor2_1 _4368_ (.Y(_0357_),
    .A(_3159_),
    .B(_0356_));
 sg13g2_nor2_1 _4369_ (.A(_0354_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_nor2_1 _4370_ (.A(net490),
    .B(_3194_),
    .Y(_0359_));
 sg13g2_a21oi_1 _4371_ (.A1(net490),
    .A2(_3158_),
    .Y(_0360_),
    .B1(_0359_));
 sg13g2_xor2_1 _4372_ (.B(_0360_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ),
    .X(_0361_));
 sg13g2_a21oi_2 _4373_ (.B1(_0361_),
    .Y(_0362_),
    .A2(_0358_),
    .A1(net396));
 sg13g2_nor2_1 _4374_ (.A(net490),
    .B(_3171_),
    .Y(_0363_));
 sg13g2_a22oi_1 _4375_ (.Y(_0364_),
    .B1(_0363_),
    .B2(_3129_),
    .A2(_3192_),
    .A1(net490));
 sg13g2_xnor2_1 _4376_ (.Y(_0365_),
    .A(_3159_),
    .B(_0364_));
 sg13g2_nor2_1 _4377_ (.A(net402),
    .B(_0358_),
    .Y(_0366_));
 sg13g2_xnor2_1 _4378_ (.Y(_0367_),
    .A(_0361_),
    .B(_0366_));
 sg13g2_xor2_1 _4379_ (.B(_0367_),
    .A(_0365_),
    .X(_0368_));
 sg13g2_nand2_1 _4380_ (.Y(_0369_),
    .A(_3130_),
    .B(_3170_));
 sg13g2_a22oi_1 _4381_ (.Y(_0370_),
    .B1(_0363_),
    .B2(_0369_),
    .A2(_0350_),
    .A1(net491));
 sg13g2_nand2_1 _4382_ (.Y(_0371_),
    .A(net396),
    .B(_0354_));
 sg13g2_xor2_1 _4383_ (.B(_0371_),
    .A(_0357_),
    .X(_0372_));
 sg13g2_nor2_1 _4384_ (.A(_0370_),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_nor2_1 _4385_ (.A(_3152_),
    .B(_3167_),
    .Y(_0374_));
 sg13g2_nor2_1 _4386_ (.A(_3134_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_nor2_1 _4387_ (.A(net492),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_a22oi_1 _4388_ (.Y(_0377_),
    .B1(_0376_),
    .B2(_3133_),
    .A2(_3190_),
    .A1(net491));
 sg13g2_xnor2_1 _4389_ (.Y(_0378_),
    .A(_3168_),
    .B(_0377_));
 sg13g2_nor2_1 _4390_ (.A(net402),
    .B(_0349_),
    .Y(_0379_));
 sg13g2_xnor2_1 _4391_ (.Y(_0380_),
    .A(_0353_),
    .B(_0379_));
 sg13g2_nand2_1 _4392_ (.Y(_0381_),
    .A(_3134_),
    .B(_0374_));
 sg13g2_a22oi_1 _4393_ (.Y(_0382_),
    .B1(_0376_),
    .B2(_0381_),
    .A2(_0341_),
    .A1(net492));
 sg13g2_nand2_1 _4394_ (.Y(_0383_),
    .A(net396),
    .B(_0345_));
 sg13g2_xnor2_1 _4395_ (.Y(_0384_),
    .A(_0348_),
    .B(_0383_));
 sg13g2_nor2_1 _4396_ (.A(_0382_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_xnor2_1 _4397_ (.Y(_0386_),
    .A(_0382_),
    .B(_0384_));
 sg13g2_inv_1 _4398_ (.Y(_0387_),
    .A(_0386_));
 sg13g2_nor2_1 _4399_ (.A(net492),
    .B(_3166_),
    .Y(_0388_));
 sg13g2_a22oi_1 _4400_ (.Y(_0389_),
    .B1(_0388_),
    .B2(_3138_),
    .A2(_3188_),
    .A1(net492));
 sg13g2_xnor2_1 _4401_ (.Y(_0390_),
    .A(_3161_),
    .B(_0389_));
 sg13g2_nor2_1 _4402_ (.A(net403),
    .B(_0339_),
    .Y(_0391_));
 sg13g2_xnor2_1 _4403_ (.Y(_0392_),
    .A(_0344_),
    .B(_0391_));
 sg13g2_nand2_1 _4404_ (.Y(_0393_),
    .A(_3139_),
    .B(_3165_));
 sg13g2_a22oi_1 _4405_ (.Y(_0394_),
    .B1(_0388_),
    .B2(_0393_),
    .A2(_0330_),
    .A1(net492));
 sg13g2_nand2_1 _4406_ (.Y(_0395_),
    .A(net396),
    .B(_0334_));
 sg13g2_xnor2_1 _4407_ (.Y(_0396_),
    .A(_0338_),
    .B(_0395_));
 sg13g2_nor2_1 _4408_ (.A(_0394_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_nand2b_1 _4409_ (.Y(_0398_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ));
 sg13g2_a22oi_1 _4410_ (.Y(_0399_),
    .B1(_3221_),
    .B2(_0398_),
    .A2(_3186_),
    .A1(net493));
 sg13g2_xnor2_1 _4411_ (.Y(_0400_),
    .A(_3181_),
    .B(_0399_));
 sg13g2_nor2_1 _4412_ (.A(net402),
    .B(_0328_),
    .Y(_0401_));
 sg13g2_xnor2_1 _4413_ (.Y(_0402_),
    .A(_0333_),
    .B(_0401_));
 sg13g2_a21oi_1 _4414_ (.A1(_3219_),
    .A2(_3232_),
    .Y(_0403_),
    .B1(_3231_));
 sg13g2_xor2_1 _4415_ (.B(_0402_),
    .A(_0400_),
    .X(_0404_));
 sg13g2_nor2b_1 _4416_ (.A(_0403_),
    .B_N(_0404_),
    .Y(_0405_));
 sg13g2_a21o_1 _4417_ (.A2(_0402_),
    .A1(_0400_),
    .B1(_0405_),
    .X(_0406_));
 sg13g2_xor2_1 _4418_ (.B(_0396_),
    .A(_0394_),
    .X(_0407_));
 sg13g2_a21oi_1 _4419_ (.A1(_0406_),
    .A2(_0407_),
    .Y(_0408_),
    .B1(_0397_));
 sg13g2_xor2_1 _4420_ (.B(_0392_),
    .A(_0390_),
    .X(_0409_));
 sg13g2_nor2b_1 _4421_ (.A(_0408_),
    .B_N(_0409_),
    .Y(_0410_));
 sg13g2_a21o_1 _4422_ (.A2(_0392_),
    .A1(_0390_),
    .B1(_0410_),
    .X(_0411_));
 sg13g2_a21oi_1 _4423_ (.A1(_0387_),
    .A2(_0411_),
    .Y(_0412_),
    .B1(_0385_));
 sg13g2_xor2_1 _4424_ (.B(_0380_),
    .A(_0378_),
    .X(_0413_));
 sg13g2_nor2b_1 _4425_ (.A(_0412_),
    .B_N(_0413_),
    .Y(_0414_));
 sg13g2_a21o_1 _4426_ (.A2(_0380_),
    .A1(_0378_),
    .B1(_0414_),
    .X(_0415_));
 sg13g2_xor2_1 _4427_ (.B(_0372_),
    .A(_0370_),
    .X(_0416_));
 sg13g2_and2_1 _4428_ (.A(_0415_),
    .B(_0416_),
    .X(_0417_));
 sg13g2_o21ai_1 _4429_ (.B1(_0368_),
    .Y(_0418_),
    .A1(_0373_),
    .A2(_0417_));
 sg13g2_o21ai_1 _4430_ (.B1(_0418_),
    .Y(_0419_),
    .A1(_0365_),
    .A2(_0367_));
 sg13g2_xor2_1 _4431_ (.B(_0419_),
    .A(_0362_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ));
 sg13g2_inv_1 _4432_ (.Y(_0420_),
    .A(net388));
 sg13g2_nand2_2 _4433_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .A(net482),
    .B(net453));
 sg13g2_and2_1 _4434_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .X(_0421_));
 sg13g2_nand2_2 _4435_ (.Y(_0422_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ));
 sg13g2_or2_1 _4436_ (.X(_0423_),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .A(net483));
 sg13g2_a21oi_1 _4437_ (.A1(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .A2(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ),
    .Y(_0424_),
    .B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ));
 sg13g2_a21o_2 _4438_ (.A2(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ),
    .A1(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .X(_0425_));
 sg13g2_o21ai_1 _4439_ (.B1(_0425_),
    .Y(_0426_),
    .A1(_0421_),
    .A2(_0423_));
 sg13g2_and2_1 _4440_ (.A(net481),
    .B(_0426_),
    .X(_0427_));
 sg13g2_nand2_2 _4441_ (.Y(_0428_),
    .A(net481),
    .B(_0426_));
 sg13g2_nor2_2 _4442_ (.A(_0422_),
    .B(_0425_),
    .Y(_0429_));
 sg13g2_nand3_1 _4443_ (.B(_0421_),
    .C(_0424_),
    .A(net483),
    .Y(_0430_));
 sg13g2_a21o_2 _4444_ (.A2(_0426_),
    .A1(net481),
    .B1(_0430_),
    .X(_0431_));
 sg13g2_nand3_1 _4445_ (.B(_0426_),
    .C(_0430_),
    .A(net481),
    .Y(_0432_));
 sg13g2_and2_1 _4446_ (.A(_0431_),
    .B(_0432_),
    .X(_0433_));
 sg13g2_a21oi_2 _4447_ (.B1(_0425_),
    .Y(_0434_),
    .A2(_0422_),
    .A1(_2915_));
 sg13g2_and2_2 _4448_ (.A(_0430_),
    .B(_0434_),
    .X(_0435_));
 sg13g2_nand2_1 _4449_ (.Y(_0436_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .B(_2947_));
 sg13g2_nand2_1 _4450_ (.Y(_0437_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .B(_0426_));
 sg13g2_a21oi_2 _4451_ (.B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .Y(_0438_),
    .A2(_0425_),
    .A1(_0423_));
 sg13g2_nand2_2 _4452_ (.Y(_0439_),
    .A(_0426_),
    .B(_0436_));
 sg13g2_a221oi_1 _4453_ (.B2(_0426_),
    .C1(_0435_),
    .B1(_0436_),
    .A1(_0431_),
    .Y(_0440_),
    .A2(_0432_));
 sg13g2_nand2_1 _4454_ (.Y(_0441_),
    .A(net449),
    .B(_0440_));
 sg13g2_o21ai_1 _4455_ (.B1(_0426_),
    .Y(_0442_),
    .A1(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ),
    .A2(net482));
 sg13g2_nor4_2 _4456_ (.A(net483),
    .B(net481),
    .C(_0422_),
    .Y(_0443_),
    .D(_0425_));
 sg13g2_o21ai_1 _4457_ (.B1(net449),
    .Y(_0444_),
    .A1(_0440_),
    .A2(_0443_));
 sg13g2_and2_1 _4458_ (.A(_2947_),
    .B(_0438_),
    .X(_0445_));
 sg13g2_nand2_1 _4459_ (.Y(_0446_),
    .A(_2947_),
    .B(_0438_));
 sg13g2_a221oi_1 _4460_ (.B2(_0430_),
    .C1(_0446_),
    .B1(_0434_),
    .A1(_0431_),
    .Y(_0447_),
    .A2(_0432_));
 sg13g2_nand2_1 _4461_ (.Y(_0448_),
    .A(net449),
    .B(_0447_));
 sg13g2_nand2_1 _4462_ (.Y(_0449_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .B(_0438_));
 sg13g2_a221oi_1 _4463_ (.B2(_0430_),
    .C1(_0449_),
    .B1(_0434_),
    .A1(_0431_),
    .Y(_0450_),
    .A2(_0432_));
 sg13g2_nor2_1 _4464_ (.A(net450),
    .B(_0431_),
    .Y(_0451_));
 sg13g2_or2_1 _4465_ (.X(_0452_),
    .B(_0431_),
    .A(net449));
 sg13g2_xnor2_1 _4466_ (.Y(_0453_),
    .A(net450),
    .B(_0431_));
 sg13g2_nand2_1 _4467_ (.Y(_0454_),
    .A(_0450_),
    .B(_0453_));
 sg13g2_a22oi_1 _4468_ (.Y(_0455_),
    .B1(_0450_),
    .B2(_0453_),
    .A2(_0447_),
    .A1(net449));
 sg13g2_and2_1 _4469_ (.A(_0442_),
    .B(_0445_),
    .X(_0456_));
 sg13g2_nand2_1 _4470_ (.Y(_0457_),
    .A(net449),
    .B(_0456_));
 sg13g2_nor4_2 _4471_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .B(_0427_),
    .C(_0435_),
    .Y(_0458_),
    .D(_0437_));
 sg13g2_or4_1 _4472_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .B(_0427_),
    .C(_0435_),
    .D(_0437_),
    .X(_0459_));
 sg13g2_o21ai_1 _4473_ (.B1(_2969_),
    .Y(_0460_),
    .A1(_0456_),
    .A2(_0458_));
 sg13g2_and3_1 _4474_ (.X(_0461_),
    .A(net450),
    .B(_0439_),
    .C(_0442_));
 sg13g2_nand3_1 _4475_ (.B(_0439_),
    .C(_0442_),
    .A(net450),
    .Y(_0462_));
 sg13g2_nand3_1 _4476_ (.B(net482),
    .C(_0424_),
    .A(net483),
    .Y(_0463_));
 sg13g2_nor2_2 _4477_ (.A(net451),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_nand2b_1 _4478_ (.Y(_0465_),
    .B(net450),
    .A_N(_0463_));
 sg13g2_nor4_2 _4479_ (.A(net483),
    .B(net451),
    .C(_0422_),
    .Y(_0466_),
    .D(_0428_));
 sg13g2_nor3_1 _4480_ (.A(_0461_),
    .B(_0464_),
    .C(_0466_),
    .Y(_0467_));
 sg13g2_and2_1 _4481_ (.A(_0460_),
    .B(_0467_),
    .X(_0468_));
 sg13g2_nand4_1 _4482_ (.B(_0455_),
    .C(_0460_),
    .A(_0444_),
    .Y(_0469_),
    .D(_0467_));
 sg13g2_and2_1 _4483_ (.A(net452),
    .B(_0450_),
    .X(_0470_));
 sg13g2_nand2_2 _4484_ (.Y(_0471_),
    .A(net452),
    .B(_0450_));
 sg13g2_nand2_2 _4485_ (.Y(_0472_),
    .A(net452),
    .B(_0440_));
 sg13g2_o21ai_1 _4486_ (.B1(net452),
    .Y(_0473_),
    .A1(_0440_),
    .A2(_0450_));
 sg13g2_nand4_1 _4487_ (.B(net481),
    .C(net453),
    .A(_2915_),
    .Y(_0474_),
    .D(_0421_));
 sg13g2_nand4_1 _4488_ (.B(net481),
    .C(net451),
    .A(net483),
    .Y(_0475_),
    .D(_0439_));
 sg13g2_nor2_1 _4489_ (.A(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .B(_0430_),
    .Y(_0476_));
 sg13g2_or2_2 _4490_ (.X(_0477_),
    .B(_0430_),
    .A(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ));
 sg13g2_nand4_1 _4491_ (.B(_0474_),
    .C(_0475_),
    .A(_0473_),
    .Y(_0478_),
    .D(_0477_));
 sg13g2_and2_1 _4492_ (.A(net452),
    .B(_0456_),
    .X(_0479_));
 sg13g2_nand3_1 _4493_ (.B(_0442_),
    .C(_0445_),
    .A(net451),
    .Y(_0480_));
 sg13g2_nand2_2 _4494_ (.Y(_0481_),
    .A(net451),
    .B(_0443_));
 sg13g2_nand2_1 _4495_ (.Y(_0482_),
    .A(net452),
    .B(_0458_));
 sg13g2_nand3_1 _4496_ (.B(_0439_),
    .C(_0442_),
    .A(net451),
    .Y(_0483_));
 sg13g2_nand2_1 _4497_ (.Y(_0484_),
    .A(_0482_),
    .B(_0483_));
 sg13g2_o21ai_1 _4498_ (.B1(_0480_),
    .Y(_0485_),
    .A1(net450),
    .A2(_0459_));
 sg13g2_nand2_1 _4499_ (.Y(_0486_),
    .A(_0481_),
    .B(_0483_));
 sg13g2_nand4_1 _4500_ (.B(_0428_),
    .C(_0435_),
    .A(net451),
    .Y(_0487_),
    .D(_0439_));
 sg13g2_nand2_1 _4501_ (.Y(_0488_),
    .A(_0452_),
    .B(_0487_));
 sg13g2_nand4_1 _4502_ (.B(_0428_),
    .C(_0435_),
    .A(net451),
    .Y(_0489_),
    .D(_0438_));
 sg13g2_nand2_1 _4503_ (.Y(_0490_),
    .A(_0463_),
    .B(_0489_));
 sg13g2_or4_1 _4504_ (.A(_0485_),
    .B(_0486_),
    .C(_0488_),
    .D(_0490_),
    .X(_0491_));
 sg13g2_nor3_2 _4505_ (.A(_0469_),
    .B(_0478_),
    .C(_0491_),
    .Y(_0492_));
 sg13g2_or3_2 _4506_ (.A(_0469_),
    .B(_0478_),
    .C(_0491_),
    .X(_0493_));
 sg13g2_or2_1 _4507_ (.X(_0494_),
    .B(_0489_),
    .A(_2947_));
 sg13g2_nand2_2 _4508_ (.Y(_0495_),
    .A(_0487_),
    .B(_0494_));
 sg13g2_nand4_1 _4509_ (.B(net481),
    .C(net453),
    .A(net483),
    .Y(_0496_),
    .D(_0438_));
 sg13g2_nand2b_2 _4510_ (.Y(_0497_),
    .B(_2947_),
    .A_N(_0496_));
 sg13g2_or2_1 _4511_ (.X(_0498_),
    .B(_0466_),
    .A(_0451_));
 sg13g2_nand2_1 _4512_ (.Y(_0499_),
    .A(_0429_),
    .B(_0464_));
 sg13g2_nand2_1 _4513_ (.Y(_0500_),
    .A(_0462_),
    .B(_0497_));
 sg13g2_nor2_1 _4514_ (.A(_0466_),
    .B(_0488_),
    .Y(_0501_));
 sg13g2_o21ai_1 _4515_ (.B1(_0481_),
    .Y(_0502_),
    .A1(_0449_),
    .A2(_0465_));
 sg13g2_nor2_1 _4516_ (.A(_0500_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_nand4_1 _4517_ (.B(_0474_),
    .C(_0499_),
    .A(_0448_),
    .Y(_0504_),
    .D(_0503_));
 sg13g2_nor4_1 _4518_ (.A(_0492_),
    .B(_0495_),
    .C(_0498_),
    .D(_0504_),
    .Y(_0505_));
 sg13g2_nand2_1 _4519_ (.Y(_0506_),
    .A(_0472_),
    .B(_0474_));
 sg13g2_nand2b_1 _4520_ (.Y(_0507_),
    .B(_0464_),
    .A_N(_0429_));
 sg13g2_nand3_1 _4521_ (.B(_0435_),
    .C(_0445_),
    .A(_0428_),
    .Y(_0508_));
 sg13g2_nor2_1 _4522_ (.A(net449),
    .B(_0508_),
    .Y(_0509_));
 sg13g2_nand3_1 _4523_ (.B(_0496_),
    .C(_0507_),
    .A(_0481_),
    .Y(_0510_));
 sg13g2_nor4_1 _4524_ (.A(_0485_),
    .B(_0506_),
    .C(_0509_),
    .D(_0510_),
    .Y(_0511_));
 sg13g2_nand3_1 _4525_ (.B(_0501_),
    .C(_0511_),
    .A(_0493_),
    .Y(_0512_));
 sg13g2_and2_1 _4526_ (.A(_0452_),
    .B(_0455_),
    .X(_0513_));
 sg13g2_and3_1 _4527_ (.X(_0514_),
    .A(_0441_),
    .B(_0452_),
    .C(_0455_));
 sg13g2_nand2_1 _4528_ (.Y(_0515_),
    .A(_0468_),
    .B(_0514_));
 sg13g2_and3_2 _4529_ (.X(_0516_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .B(_0468_),
    .C(_0514_));
 sg13g2_nand3_1 _4530_ (.B(_0468_),
    .C(_0514_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .Y(_0517_));
 sg13g2_nor2_1 _4531_ (.A(_0440_),
    .B(_0470_),
    .Y(_0518_));
 sg13g2_a21oi_1 _4532_ (.A1(_0445_),
    .A2(_0464_),
    .Y(_0519_),
    .B1(_0466_));
 sg13g2_a21oi_1 _4533_ (.A1(_0438_),
    .A2(_0464_),
    .Y(_0520_),
    .B1(_0466_));
 sg13g2_and4_1 _4534_ (.A(_0474_),
    .B(_0481_),
    .C(_0483_),
    .D(_0520_),
    .X(_0521_));
 sg13g2_nand3_1 _4535_ (.B(_0518_),
    .C(_0521_),
    .A(_0497_),
    .Y(_0522_));
 sg13g2_nand3_1 _4536_ (.B(_0480_),
    .C(_0497_),
    .A(_0477_),
    .Y(_0523_));
 sg13g2_nor4_2 _4537_ (.A(_0495_),
    .B(_0516_),
    .C(_0522_),
    .Y(_0524_),
    .D(_0523_));
 sg13g2_nor2_1 _4538_ (.A(_0512_),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_xnor2_1 _4539_ (.Y(_0526_),
    .A(_0512_),
    .B(_0524_));
 sg13g2_and2_1 _4540_ (.A(_0475_),
    .B(_0477_),
    .X(_0527_));
 sg13g2_nand4_1 _4541_ (.B(_0487_),
    .C(_0519_),
    .A(_0471_),
    .Y(_0528_),
    .D(_0527_));
 sg13g2_nor2_1 _4542_ (.A(_2947_),
    .B(_0496_),
    .Y(_0529_));
 sg13g2_a21oi_2 _4543_ (.B1(_0529_),
    .Y(_0530_),
    .A2(_0464_),
    .A1(_0429_));
 sg13g2_nand2_1 _4544_ (.Y(_0531_),
    .A(_0460_),
    .B(_0530_));
 sg13g2_nand4_1 _4545_ (.B(_0481_),
    .C(_0482_),
    .A(_0455_),
    .Y(_0532_),
    .D(_0483_));
 sg13g2_or4_2 _4546_ (.A(_0492_),
    .B(_0528_),
    .C(_0531_),
    .D(_0532_),
    .X(_0533_));
 sg13g2_nand2_1 _4547_ (.Y(_0534_),
    .A(_0475_),
    .B(_0496_));
 sg13g2_and4_1 _4548_ (.A(net450),
    .B(_0427_),
    .C(_0435_),
    .D(_0439_),
    .X(_0535_));
 sg13g2_nor4_1 _4549_ (.A(_0479_),
    .B(_0498_),
    .C(_0534_),
    .D(_0535_),
    .Y(_0536_));
 sg13g2_nor4_2 _4550_ (.A(_0433_),
    .B(_0435_),
    .C(_0446_),
    .Y(_0537_),
    .D(_0453_));
 sg13g2_inv_1 _4551_ (.Y(_0538_),
    .A(_0537_));
 sg13g2_nand4_1 _4552_ (.B(_0494_),
    .C(_0536_),
    .A(_0441_),
    .Y(_0539_),
    .D(_0538_));
 sg13g2_nand3_1 _4553_ (.B(_0457_),
    .C(_0499_),
    .A(_0448_),
    .Y(_0540_));
 sg13g2_or2_1 _4554_ (.X(_0541_),
    .B(_0540_),
    .A(_0484_));
 sg13g2_nor3_1 _4555_ (.A(_0516_),
    .B(_0539_),
    .C(_0541_),
    .Y(_0542_));
 sg13g2_and2_1 _4556_ (.A(_0533_),
    .B(_0542_),
    .X(_0543_));
 sg13g2_nand4_1 _4557_ (.B(_0475_),
    .C(_0477_),
    .A(_0444_),
    .Y(_0544_),
    .D(_0497_));
 sg13g2_nor3_2 _4558_ (.A(_0492_),
    .B(_0541_),
    .C(_0544_),
    .Y(_0545_));
 sg13g2_nand3_1 _4559_ (.B(_0462_),
    .C(_0475_),
    .A(_0454_),
    .Y(_0546_));
 sg13g2_nor4_1 _4560_ (.A(_0451_),
    .B(_0485_),
    .C(_0535_),
    .D(_0546_),
    .Y(_0547_));
 sg13g2_and4_1 _4561_ (.A(_0474_),
    .B(_0517_),
    .C(_0530_),
    .D(_0547_),
    .X(_0548_));
 sg13g2_nand2b_1 _4562_ (.Y(_0549_),
    .B(_0545_),
    .A_N(_0548_));
 sg13g2_and2_1 _4563_ (.A(_0473_),
    .B(_0493_),
    .X(_0550_));
 sg13g2_nand4_1 _4564_ (.B(_0475_),
    .C(_0482_),
    .A(_0457_),
    .Y(_0551_),
    .D(_0507_));
 sg13g2_nor4_1 _4565_ (.A(_0495_),
    .B(_0498_),
    .C(_0500_),
    .D(_0551_),
    .Y(_0552_));
 sg13g2_and3_2 _4566_ (.X(_0553_),
    .A(_0473_),
    .B(_0493_),
    .C(_0552_));
 sg13g2_nor2_1 _4567_ (.A(_0470_),
    .B(_0537_),
    .Y(_0554_));
 sg13g2_a21oi_1 _4568_ (.A1(net449),
    .A2(_0458_),
    .Y(_0555_),
    .B1(_0509_));
 sg13g2_and4_1 _4569_ (.A(_0441_),
    .B(_0487_),
    .C(_0494_),
    .D(_0555_),
    .X(_0556_));
 sg13g2_and4_1 _4570_ (.A(_0474_),
    .B(_0480_),
    .C(_0520_),
    .D(_0530_),
    .X(_0557_));
 sg13g2_nand4_1 _4571_ (.B(_0554_),
    .C(_0556_),
    .A(_0517_),
    .Y(_0558_),
    .D(_0557_));
 sg13g2_nor2_1 _4572_ (.A(_0553_),
    .B(_0558_),
    .Y(_0559_));
 sg13g2_nor2b_1 _4573_ (.A(_0545_),
    .B_N(_0548_),
    .Y(_0560_));
 sg13g2_xnor2_1 _4574_ (.Y(_0561_),
    .A(_0545_),
    .B(_0548_));
 sg13g2_o21ai_1 _4575_ (.B1(_0549_),
    .Y(_0562_),
    .A1(_0559_),
    .A2(_0560_));
 sg13g2_o21ai_1 _4576_ (.B1(_0483_),
    .Y(_0563_),
    .A1(_0446_),
    .A2(_0465_));
 sg13g2_nor4_1 _4577_ (.A(_0451_),
    .B(_0506_),
    .C(_0535_),
    .D(_0563_),
    .Y(_0564_));
 sg13g2_nand3_1 _4578_ (.B(_0556_),
    .C(_0564_),
    .A(_0517_),
    .Y(_0565_));
 sg13g2_nand2_1 _4579_ (.Y(_0566_),
    .A(net413),
    .B(_0565_));
 sg13g2_inv_1 _4580_ (.Y(_0567_),
    .A(_0566_));
 sg13g2_xor2_1 _4581_ (.B(_0565_),
    .A(net413),
    .X(_0568_));
 sg13g2_or2_1 _4582_ (.X(_0569_),
    .B(_0542_),
    .A(_0533_));
 sg13g2_nand2_1 _4583_ (.Y(_0570_),
    .A(_0566_),
    .B(_0569_));
 sg13g2_a21oi_1 _4584_ (.A1(_0562_),
    .A2(_0568_),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_nor3_1 _4585_ (.A(_0526_),
    .B(_0543_),
    .C(_0571_),
    .Y(_0572_));
 sg13g2_or3_1 _4586_ (.A(_0526_),
    .B(_0543_),
    .C(_0571_),
    .X(_0573_));
 sg13g2_o21ai_1 _4587_ (.B1(_0526_),
    .Y(_0574_),
    .A1(_0543_),
    .A2(_0571_));
 sg13g2_and2_2 _4588_ (.A(_0573_),
    .B(_0574_),
    .X(_0575_));
 sg13g2_nor2b_1 _4589_ (.A(_0543_),
    .B_N(_0569_),
    .Y(_0576_));
 sg13g2_a21oi_1 _4590_ (.A1(_0562_),
    .A2(_0568_),
    .Y(_0577_),
    .B1(_0567_));
 sg13g2_xnor2_1 _4591_ (.Y(_0578_),
    .A(_0576_),
    .B(_0577_));
 sg13g2_nand2_2 _4592_ (.Y(_0579_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .B(_0578_));
 sg13g2_xor2_1 _4593_ (.B(_0568_),
    .A(_0562_),
    .X(_0580_));
 sg13g2_nand2_2 _4594_ (.Y(_0581_),
    .A(net489),
    .B(_0580_));
 sg13g2_nand2_2 _4595_ (.Y(_0582_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .B(_0580_));
 sg13g2_nand2_2 _4596_ (.Y(_0583_),
    .A(net489),
    .B(_0578_));
 sg13g2_or2_1 _4597_ (.X(_0584_),
    .B(_0583_),
    .A(_0582_));
 sg13g2_nor2_1 _4598_ (.A(_0575_),
    .B(_0584_),
    .Y(_0585_));
 sg13g2_nand3_1 _4599_ (.B(_0573_),
    .C(_0574_),
    .A(net489),
    .Y(_0586_));
 sg13g2_nor2_2 _4600_ (.A(_0579_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_xor2_1 _4601_ (.B(_0586_),
    .A(_0579_),
    .X(_0588_));
 sg13g2_mux2_1 _4602_ (.A0(_0575_),
    .A1(_0588_),
    .S(_0584_),
    .X(_0589_));
 sg13g2_nand2_2 _4603_ (.Y(_0590_),
    .A(net488),
    .B(_0580_));
 sg13g2_xnor2_1 _4604_ (.Y(_0591_),
    .A(_0559_),
    .B(_0561_));
 sg13g2_nor2b_1 _4605_ (.A(_0010_),
    .B_N(_0591_),
    .Y(_0592_));
 sg13g2_xor2_1 _4606_ (.B(_0558_),
    .A(_0553_),
    .X(_0593_));
 sg13g2_nor2_1 _4607_ (.A(_0009_),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_nand2_1 _4608_ (.Y(_0595_),
    .A(_0592_),
    .B(_0594_));
 sg13g2_xnor2_1 _4609_ (.Y(_0596_),
    .A(_0592_),
    .B(_0594_));
 sg13g2_xor2_1 _4610_ (.B(_0596_),
    .A(_0590_),
    .X(_0597_));
 sg13g2_a21oi_2 _4611_ (.B1(_0585_),
    .Y(_0598_),
    .A2(_0597_),
    .A1(_0589_));
 sg13g2_nand2_2 _4612_ (.Y(_0599_),
    .A(net487),
    .B(_0578_));
 sg13g2_nand2_1 _4613_ (.Y(_0600_),
    .A(net484),
    .B(_0580_));
 sg13g2_nand2_1 _4614_ (.Y(_0601_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .B(_0591_));
 sg13g2_nor2_1 _4615_ (.A(_0600_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_xor2_1 _4616_ (.B(_0601_),
    .A(_0600_),
    .X(_0603_));
 sg13g2_nand2b_1 _4617_ (.Y(_0604_),
    .B(_0603_),
    .A_N(_0599_));
 sg13g2_xnor2_1 _4618_ (.Y(_0605_),
    .A(_0599_),
    .B(_0603_));
 sg13g2_nor3_1 _4619_ (.A(_0476_),
    .B(_0484_),
    .C(_0488_),
    .Y(_0606_));
 sg13g2_and4_1 _4620_ (.A(_0496_),
    .B(_0514_),
    .C(_0550_),
    .D(_0606_),
    .X(_0607_));
 sg13g2_nand3_1 _4621_ (.B(_0475_),
    .C(_0497_),
    .A(_0474_),
    .Y(_0608_));
 sg13g2_nor3_1 _4622_ (.A(_0485_),
    .B(_0495_),
    .C(_0608_),
    .Y(_0609_));
 sg13g2_nand4_1 _4623_ (.B(_0517_),
    .C(_0554_),
    .A(_0513_),
    .Y(_0610_),
    .D(_0609_));
 sg13g2_nand2_1 _4624_ (.Y(_0611_),
    .A(net412),
    .B(_0610_));
 sg13g2_xor2_1 _4625_ (.B(_0610_),
    .A(net412),
    .X(_0612_));
 sg13g2_o21ai_1 _4626_ (.B1(_0612_),
    .Y(_0613_),
    .A1(_0525_),
    .A2(_0572_));
 sg13g2_or3_1 _4627_ (.A(_0525_),
    .B(_0572_),
    .C(_0612_),
    .X(_0614_));
 sg13g2_and2_2 _4628_ (.A(_0613_),
    .B(_0614_),
    .X(_0615_));
 sg13g2_nand3_1 _4629_ (.B(_0613_),
    .C(_0614_),
    .A(net489),
    .Y(_0616_));
 sg13g2_nand3_1 _4630_ (.B(_0573_),
    .C(_0574_),
    .A(_2949_),
    .Y(_0617_));
 sg13g2_xor2_1 _4631_ (.B(_0617_),
    .A(_0616_),
    .X(_0618_));
 sg13g2_xnor2_1 _4632_ (.Y(_0619_),
    .A(_0587_),
    .B(_0618_));
 sg13g2_nor2b_1 _4633_ (.A(_0619_),
    .B_N(_0605_),
    .Y(_0620_));
 sg13g2_xnor2_1 _4634_ (.Y(_0621_),
    .A(_0605_),
    .B(_0619_));
 sg13g2_nor2b_1 _4635_ (.A(_0598_),
    .B_N(_0621_),
    .Y(_0622_));
 sg13g2_o21ai_1 _4636_ (.B1(_0595_),
    .Y(_0623_),
    .A1(_0590_),
    .A2(_0596_));
 sg13g2_xnor2_1 _4637_ (.Y(_0624_),
    .A(_0598_),
    .B(_0621_));
 sg13g2_a21oi_2 _4638_ (.B1(_0622_),
    .Y(_0625_),
    .A2(_0624_),
    .A1(_0623_));
 sg13g2_nand2b_2 _4639_ (.Y(_0626_),
    .B(_0604_),
    .A_N(_0602_));
 sg13g2_nand2b_2 _4640_ (.Y(_0627_),
    .B(_0615_),
    .A_N(_0011_));
 sg13g2_nor2_2 _4641_ (.A(_0617_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_xor2_1 _4642_ (.B(_0627_),
    .A(_0617_),
    .X(_0629_));
 sg13g2_a21o_1 _4643_ (.A2(_0629_),
    .A1(_0587_),
    .B1(_0620_),
    .X(_0630_));
 sg13g2_nand2_1 _4644_ (.Y(_0631_),
    .A(net484),
    .B(_0578_));
 sg13g2_nand2_1 _4645_ (.Y(_0632_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .B(_0580_));
 sg13g2_or2_1 _4646_ (.X(_0633_),
    .B(_0632_),
    .A(_0631_));
 sg13g2_xor2_1 _4647_ (.B(_0632_),
    .A(_0631_),
    .X(_0634_));
 sg13g2_nand2_1 _4648_ (.Y(_0635_),
    .A(net487),
    .B(_0575_));
 sg13g2_nand3_1 _4649_ (.B(_0575_),
    .C(_0634_),
    .A(net487),
    .Y(_0636_));
 sg13g2_xor2_1 _4650_ (.B(_0635_),
    .A(_0634_),
    .X(_0637_));
 sg13g2_nor4_1 _4651_ (.A(_0469_),
    .B(_0488_),
    .C(_0506_),
    .D(_0523_),
    .Y(_0638_));
 sg13g2_nand2_2 _4652_ (.Y(_0639_),
    .A(_0493_),
    .B(_0638_));
 sg13g2_nor4_2 _4653_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .B(_0478_),
    .C(_0495_),
    .Y(_0640_),
    .D(_0515_));
 sg13g2_nor2_1 _4654_ (.A(_0639_),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_xnor2_1 _4655_ (.Y(_0642_),
    .A(_0639_),
    .B(_0640_));
 sg13g2_a21oi_2 _4656_ (.B1(_0642_),
    .Y(_0643_),
    .A2(_0613_),
    .A1(_0611_));
 sg13g2_nor2_1 _4657_ (.A(_0537_),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_or3_2 _4658_ (.A(_0008_),
    .B(_0537_),
    .C(_0643_),
    .X(_0645_));
 sg13g2_nor3_2 _4659_ (.A(_2950_),
    .B(_0537_),
    .C(_0643_),
    .Y(_0646_));
 sg13g2_and2_1 _4660_ (.A(_2949_),
    .B(_0615_),
    .X(_0647_));
 sg13g2_nor2_2 _4661_ (.A(_0616_),
    .B(_0645_),
    .Y(_0648_));
 sg13g2_xnor2_1 _4662_ (.Y(_0649_),
    .A(_0646_),
    .B(_0647_));
 sg13g2_or3_1 _4663_ (.A(_0617_),
    .B(_0627_),
    .C(_0649_),
    .X(_0650_));
 sg13g2_xor2_1 _4664_ (.B(_0649_),
    .A(_0628_),
    .X(_0651_));
 sg13g2_xor2_1 _4665_ (.B(_0651_),
    .A(_0637_),
    .X(_0652_));
 sg13g2_xnor2_1 _4666_ (.Y(_0653_),
    .A(_0630_),
    .B(_0652_));
 sg13g2_nor2b_1 _4667_ (.A(_0653_),
    .B_N(_0626_),
    .Y(_0654_));
 sg13g2_xor2_1 _4668_ (.B(_0653_),
    .A(_0626_),
    .X(_0655_));
 sg13g2_or2_1 _4669_ (.X(_0656_),
    .B(_0655_),
    .A(_0625_));
 sg13g2_and2_1 _4670_ (.A(_0625_),
    .B(_0655_),
    .X(_0657_));
 sg13g2_xor2_1 _4671_ (.B(_0655_),
    .A(_0625_),
    .X(_0658_));
 sg13g2_xnor2_1 _4672_ (.Y(_0659_),
    .A(_0623_),
    .B(_0624_));
 sg13g2_xor2_1 _4673_ (.B(_0583_),
    .A(_0582_),
    .X(_0660_));
 sg13g2_nand2_2 _4674_ (.Y(_0661_),
    .A(_2949_),
    .B(_0591_));
 sg13g2_nor2_2 _4675_ (.A(_0581_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_and2_1 _4676_ (.A(_0660_),
    .B(_0662_),
    .X(_0663_));
 sg13g2_nand2b_2 _4677_ (.Y(_0664_),
    .B(net486),
    .A_N(_0593_));
 sg13g2_inv_1 _4678_ (.Y(_0665_),
    .A(_0664_));
 sg13g2_nand2_2 _4679_ (.Y(_0666_),
    .A(net488),
    .B(_0591_));
 sg13g2_nor2_2 _4680_ (.A(_0664_),
    .B(_0666_),
    .Y(_0667_));
 sg13g2_xnor2_1 _4681_ (.Y(_0668_),
    .A(_0665_),
    .B(_0666_));
 sg13g2_xor2_1 _4682_ (.B(_0662_),
    .A(_0660_),
    .X(_0669_));
 sg13g2_a21o_1 _4683_ (.A2(_0669_),
    .A1(_0668_),
    .B1(_0663_),
    .X(_0670_));
 sg13g2_xnor2_1 _4684_ (.Y(_0671_),
    .A(_0589_),
    .B(_0597_));
 sg13g2_nor2b_1 _4685_ (.A(_0671_),
    .B_N(_0670_),
    .Y(_0672_));
 sg13g2_xnor2_1 _4686_ (.Y(_0673_),
    .A(_0670_),
    .B(_0671_));
 sg13g2_and2_1 _4687_ (.A(_0667_),
    .B(_0673_),
    .X(_0674_));
 sg13g2_or2_1 _4688_ (.X(_0675_),
    .B(_0661_),
    .A(_0011_));
 sg13g2_nor3_1 _4689_ (.A(_2948_),
    .B(_0593_),
    .C(_0675_),
    .Y(_0676_));
 sg13g2_inv_1 _4690_ (.Y(_0677_),
    .A(_0676_));
 sg13g2_a21oi_1 _4691_ (.A1(_2948_),
    .A2(_0675_),
    .Y(_0678_),
    .B1(_0593_));
 sg13g2_xor2_1 _4692_ (.B(_0661_),
    .A(_0581_),
    .X(_0679_));
 sg13g2_a21o_1 _4693_ (.A2(_0679_),
    .A1(_0678_),
    .B1(_0676_),
    .X(_0680_));
 sg13g2_xnor2_1 _4694_ (.Y(_0681_),
    .A(_0668_),
    .B(_0669_));
 sg13g2_o21ai_1 _4695_ (.B1(_0680_),
    .Y(_0682_),
    .A1(_0667_),
    .A2(_0673_));
 sg13g2_nor3_1 _4696_ (.A(_0674_),
    .B(_0681_),
    .C(_0682_),
    .Y(_0683_));
 sg13g2_or3_1 _4697_ (.A(_0672_),
    .B(_0674_),
    .C(_0683_),
    .X(_0684_));
 sg13g2_nand2b_1 _4698_ (.Y(_0685_),
    .B(_0684_),
    .A_N(_0659_));
 sg13g2_o21ai_1 _4699_ (.B1(_0656_),
    .Y(_0686_),
    .A1(_0657_),
    .A2(_0685_));
 sg13g2_a21oi_2 _4700_ (.B1(_0654_),
    .Y(_0687_),
    .A2(_0652_),
    .A1(_0630_));
 sg13g2_nand2_2 _4701_ (.Y(_0688_),
    .A(_0633_),
    .B(_0636_));
 sg13g2_o21ai_1 _4702_ (.B1(_0650_),
    .Y(_0689_),
    .A1(_0637_),
    .A2(_0651_));
 sg13g2_nand2_2 _4703_ (.Y(_0690_),
    .A(net487),
    .B(_0615_));
 sg13g2_nand2_1 _4704_ (.Y(_0691_),
    .A(net484),
    .B(_0575_));
 sg13g2_nor2b_1 _4705_ (.A(_0009_),
    .B_N(_0578_),
    .Y(_0692_));
 sg13g2_nand3_1 _4706_ (.B(_0575_),
    .C(_0692_),
    .A(net484),
    .Y(_0693_));
 sg13g2_xnor2_1 _4707_ (.Y(_0694_),
    .A(_0691_),
    .B(_0692_));
 sg13g2_nand2b_1 _4708_ (.Y(_0695_),
    .B(_0694_),
    .A_N(_0690_));
 sg13g2_xnor2_1 _4709_ (.Y(_0696_),
    .A(_0690_),
    .B(_0694_));
 sg13g2_inv_1 _4710_ (.Y(_0697_),
    .A(_0696_));
 sg13g2_nor3_1 _4711_ (.A(_0476_),
    .B(_0485_),
    .C(_0486_),
    .Y(_0698_));
 sg13g2_nand4_1 _4712_ (.B(_0475_),
    .C(_0508_),
    .A(_0472_),
    .Y(_0699_),
    .D(_0698_));
 sg13g2_nor3_1 _4713_ (.A(_0516_),
    .B(_0537_),
    .C(_0699_),
    .Y(_0700_));
 sg13g2_and3_1 _4714_ (.X(_0701_),
    .A(_0471_),
    .B(_0474_),
    .C(_0493_));
 sg13g2_nand3_1 _4715_ (.B(_0698_),
    .C(_0701_),
    .A(_0489_),
    .Y(_0702_));
 sg13g2_xor2_1 _4716_ (.B(_0702_),
    .A(_0700_),
    .X(_0703_));
 sg13g2_o21ai_1 _4717_ (.B1(_0703_),
    .Y(_0704_),
    .A1(_0641_),
    .A2(_0643_));
 sg13g2_and2_2 _4718_ (.A(_0472_),
    .B(net408),
    .X(_0705_));
 sg13g2_inv_1 _4719_ (.Y(_0706_),
    .A(_0705_));
 sg13g2_nand2_1 _4720_ (.Y(_0707_),
    .A(_0648_),
    .B(_0706_));
 sg13g2_nand2_1 _4721_ (.Y(_0708_),
    .A(net489),
    .B(_0704_));
 sg13g2_inv_1 _4722_ (.Y(_0709_),
    .A(_0708_));
 sg13g2_nand3_1 _4723_ (.B(_0472_),
    .C(net408),
    .A(net489),
    .Y(_0710_));
 sg13g2_or2_2 _4724_ (.X(_0711_),
    .B(_0710_),
    .A(_0645_));
 sg13g2_xnor2_1 _4725_ (.Y(_0712_),
    .A(_0645_),
    .B(_0710_));
 sg13g2_mux2_1 _4726_ (.A0(_0712_),
    .A1(_0706_),
    .S(_0648_),
    .X(_0713_));
 sg13g2_xnor2_1 _4727_ (.Y(_0714_),
    .A(_0697_),
    .B(_0713_));
 sg13g2_nand2b_1 _4728_ (.Y(_0715_),
    .B(_0689_),
    .A_N(_0714_));
 sg13g2_xor2_1 _4729_ (.B(_0714_),
    .A(_0689_),
    .X(_0716_));
 sg13g2_nand2b_1 _4730_ (.Y(_0717_),
    .B(_0688_),
    .A_N(_0716_));
 sg13g2_xor2_1 _4731_ (.B(_0716_),
    .A(_0688_),
    .X(_0718_));
 sg13g2_nor2_1 _4732_ (.A(_0687_),
    .B(_0718_),
    .Y(_0719_));
 sg13g2_xor2_1 _4733_ (.B(_0718_),
    .A(_0687_),
    .X(_0720_));
 sg13g2_xor2_1 _4734_ (.B(_0720_),
    .A(_0686_),
    .X(_0721_));
 sg13g2_nand2b_1 _4735_ (.Y(_0722_),
    .B(_0721_),
    .A_N(_0505_));
 sg13g2_nor2b_1 _4736_ (.A(_0721_),
    .B_N(net413),
    .Y(_0723_));
 sg13g2_xnor2_1 _4737_ (.Y(_0724_),
    .A(net413),
    .B(_0721_));
 sg13g2_nand2_1 _4738_ (.Y(_0725_),
    .A(_0597_),
    .B(_0667_));
 sg13g2_xor2_1 _4739_ (.B(_0667_),
    .A(_0597_),
    .X(_0726_));
 sg13g2_nand2_1 _4740_ (.Y(_0727_),
    .A(_0588_),
    .B(_0726_));
 sg13g2_nand2_1 _4741_ (.Y(_0728_),
    .A(_0725_),
    .B(_0727_));
 sg13g2_or2_1 _4742_ (.X(_0729_),
    .B(_0623_),
    .A(_0605_));
 sg13g2_and2_1 _4743_ (.A(_0605_),
    .B(_0623_),
    .X(_0730_));
 sg13g2_xor2_1 _4744_ (.B(_0623_),
    .A(_0605_),
    .X(_0731_));
 sg13g2_xnor2_1 _4745_ (.Y(_0732_),
    .A(_0618_),
    .B(_0731_));
 sg13g2_a21oi_1 _4746_ (.A1(_0725_),
    .A2(_0727_),
    .Y(_0733_),
    .B1(_0732_));
 sg13g2_xor2_1 _4747_ (.B(_0732_),
    .A(_0728_),
    .X(_0734_));
 sg13g2_inv_1 _4748_ (.Y(_0735_),
    .A(_0734_));
 sg13g2_xor2_1 _4749_ (.B(_0734_),
    .A(_0587_),
    .X(_0736_));
 sg13g2_nand2_1 _4750_ (.Y(_0737_),
    .A(_0660_),
    .B(_0668_));
 sg13g2_xnor2_1 _4751_ (.Y(_0738_),
    .A(_0588_),
    .B(_0726_));
 sg13g2_nor2_1 _4752_ (.A(_0737_),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_xnor2_1 _4753_ (.Y(_0740_),
    .A(_0737_),
    .B(_0738_));
 sg13g2_or2_1 _4754_ (.X(_0741_),
    .B(_0740_),
    .A(_0584_));
 sg13g2_nor2b_1 _4755_ (.A(_0739_),
    .B_N(_0741_),
    .Y(_0742_));
 sg13g2_or2_1 _4756_ (.X(_0743_),
    .B(_0742_),
    .A(_0736_));
 sg13g2_xnor2_1 _4757_ (.Y(_0744_),
    .A(_0736_),
    .B(_0742_));
 sg13g2_nand2_1 _4758_ (.Y(_0745_),
    .A(_0584_),
    .B(_0740_));
 sg13g2_xor2_1 _4759_ (.B(_0666_),
    .A(_0582_),
    .X(_0746_));
 sg13g2_nand2b_1 _4760_ (.Y(_0747_),
    .B(_0746_),
    .A_N(_0583_));
 sg13g2_xnor2_1 _4761_ (.Y(_0748_),
    .A(_0583_),
    .B(_0746_));
 sg13g2_xnor2_1 _4762_ (.Y(_0749_),
    .A(_0664_),
    .B(_0748_));
 sg13g2_o21ai_1 _4763_ (.B1(_0749_),
    .Y(_0750_),
    .A1(_0662_),
    .A2(_0680_));
 sg13g2_o21ai_1 _4764_ (.B1(_0750_),
    .Y(_0751_),
    .A1(_0581_),
    .A2(_0677_));
 sg13g2_nand3_1 _4765_ (.B(_0745_),
    .C(_0751_),
    .A(_0741_),
    .Y(_0752_));
 sg13g2_xnor2_1 _4766_ (.Y(_0753_),
    .A(_0744_),
    .B(_0752_));
 sg13g2_nor2_1 _4767_ (.A(_0553_),
    .B(_0753_),
    .Y(_0754_));
 sg13g2_or2_2 _4768_ (.X(_0755_),
    .B(_0753_),
    .A(_0553_));
 sg13g2_nand2_1 _4769_ (.Y(_0756_),
    .A(_0545_),
    .B(_0755_));
 sg13g2_nor2_1 _4770_ (.A(_0545_),
    .B(_0755_),
    .Y(_0757_));
 sg13g2_xnor2_1 _4771_ (.Y(_0758_),
    .A(_0658_),
    .B(_0685_));
 sg13g2_a21oi_1 _4772_ (.A1(_0756_),
    .A2(_0758_),
    .Y(_0759_),
    .B1(_0757_));
 sg13g2_o21ai_1 _4773_ (.B1(_0722_),
    .Y(_0760_),
    .A1(_0723_),
    .A2(_0759_));
 sg13g2_a21oi_1 _4774_ (.A1(_0686_),
    .A2(_0720_),
    .Y(_0761_),
    .B1(_0719_));
 sg13g2_nand2_1 _4775_ (.Y(_0762_),
    .A(_0715_),
    .B(_0717_));
 sg13g2_and2_2 _4776_ (.A(_0693_),
    .B(_0695_),
    .X(_0763_));
 sg13g2_o21ai_1 _4777_ (.B1(_0707_),
    .Y(_0764_),
    .A1(_0697_),
    .A2(_0713_));
 sg13g2_nand2_2 _4778_ (.Y(_0765_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .B(_0615_));
 sg13g2_nand2_1 _4779_ (.Y(_0766_),
    .A(net484),
    .B(_0615_));
 sg13g2_nand2_1 _4780_ (.Y(_0767_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .B(_0575_));
 sg13g2_nor2_2 _4781_ (.A(_0691_),
    .B(_0765_),
    .Y(_0768_));
 sg13g2_xor2_1 _4782_ (.B(_0767_),
    .A(_0766_),
    .X(_0769_));
 sg13g2_nor3_2 _4783_ (.A(_2948_),
    .B(_0537_),
    .C(_0643_),
    .Y(_0770_));
 sg13g2_xnor2_1 _4784_ (.Y(_0771_),
    .A(_0769_),
    .B(_0770_));
 sg13g2_and2_2 _4785_ (.A(_0471_),
    .B(net408),
    .X(_0772_));
 sg13g2_nand2_2 _4786_ (.Y(_0773_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .B(_0772_));
 sg13g2_nand2_2 _4787_ (.Y(_0774_),
    .A(net489),
    .B(_0772_));
 sg13g2_nand3_1 _4788_ (.B(_0472_),
    .C(net408),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .Y(_0775_));
 sg13g2_nor2_1 _4789_ (.A(_0710_),
    .B(_0773_),
    .Y(_0776_));
 sg13g2_xor2_1 _4790_ (.B(_0775_),
    .A(_0774_),
    .X(_0777_));
 sg13g2_nor2b_1 _4791_ (.A(_0711_),
    .B_N(_0777_),
    .Y(_0778_));
 sg13g2_xnor2_1 _4792_ (.Y(_0779_),
    .A(_0711_),
    .B(_0777_));
 sg13g2_nor2b_1 _4793_ (.A(_0771_),
    .B_N(_0779_),
    .Y(_0780_));
 sg13g2_xnor2_1 _4794_ (.Y(_0781_),
    .A(_0771_),
    .B(_0779_));
 sg13g2_nand2_1 _4795_ (.Y(_0782_),
    .A(_0764_),
    .B(_0781_));
 sg13g2_xnor2_1 _4796_ (.Y(_0783_),
    .A(_0764_),
    .B(_0781_));
 sg13g2_xor2_1 _4797_ (.B(_0783_),
    .A(_0763_),
    .X(_0784_));
 sg13g2_nand2_1 _4798_ (.Y(_0785_),
    .A(_0762_),
    .B(_0784_));
 sg13g2_xnor2_1 _4799_ (.Y(_0786_),
    .A(_0762_),
    .B(_0784_));
 sg13g2_xor2_1 _4800_ (.B(_0786_),
    .A(_0761_),
    .X(_0787_));
 sg13g2_and2_1 _4801_ (.A(_0533_),
    .B(_0787_),
    .X(_0788_));
 sg13g2_xor2_1 _4802_ (.B(_0787_),
    .A(_0533_),
    .X(_0789_));
 sg13g2_xnor2_1 _4803_ (.Y(_0790_),
    .A(_0760_),
    .B(_0789_));
 sg13g2_nor2_1 _4804_ (.A(_0015_),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_xnor2_1 _4805_ (.Y(_0792_),
    .A(_0724_),
    .B(_0759_));
 sg13g2_and2_1 _4806_ (.A(\main.demo._q_speed[0] ),
    .B(_0792_),
    .X(_0793_));
 sg13g2_xor2_1 _4807_ (.B(_0790_),
    .A(_0015_),
    .X(_0794_));
 sg13g2_a21o_1 _4808_ (.A2(_0794_),
    .A1(_0793_),
    .B1(_0791_),
    .X(_0795_));
 sg13g2_a21oi_1 _4809_ (.A1(_0760_),
    .A2(_0789_),
    .Y(_0796_),
    .B1(_0788_));
 sg13g2_o21ai_1 _4810_ (.B1(_0785_),
    .Y(_0797_),
    .A1(_0761_),
    .A2(_0786_));
 sg13g2_o21ai_1 _4811_ (.B1(_0782_),
    .Y(_0798_),
    .A1(_0763_),
    .A2(_0783_));
 sg13g2_a21oi_2 _4812_ (.B1(_0768_),
    .Y(_0799_),
    .A2(_0770_),
    .A1(_0769_));
 sg13g2_and2_1 _4813_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .B(_0644_),
    .X(_0800_));
 sg13g2_nand2_1 _4814_ (.Y(_0801_),
    .A(net485),
    .B(_0644_));
 sg13g2_nor2_1 _4815_ (.A(_0765_),
    .B(_0801_),
    .Y(_0802_));
 sg13g2_inv_1 _4816_ (.Y(_0803_),
    .A(_0802_));
 sg13g2_xor2_1 _4817_ (.B(_0801_),
    .A(_0765_),
    .X(_0804_));
 sg13g2_nand2_1 _4818_ (.Y(_0805_),
    .A(net488),
    .B(net408));
 sg13g2_inv_1 _4819_ (.Y(_0806_),
    .A(_0805_));
 sg13g2_nand2_1 _4820_ (.Y(_0807_),
    .A(net487),
    .B(_0705_));
 sg13g2_nand3_1 _4821_ (.B(_0705_),
    .C(_0804_),
    .A(net487),
    .Y(_0808_));
 sg13g2_xor2_1 _4822_ (.B(_0807_),
    .A(_0804_),
    .X(_0809_));
 sg13g2_nand3_1 _4823_ (.B(net489),
    .C(_0772_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .Y(_0810_));
 sg13g2_inv_1 _4824_ (.Y(_0811_),
    .A(_0810_));
 sg13g2_xnor2_1 _4825_ (.Y(_0812_),
    .A(_0709_),
    .B(_0773_));
 sg13g2_nor2_1 _4826_ (.A(_0776_),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_or2_1 _4827_ (.X(_0814_),
    .B(_0813_),
    .A(_0809_));
 sg13g2_xnor2_1 _4828_ (.Y(_0815_),
    .A(_0809_),
    .B(_0813_));
 sg13g2_nor2_1 _4829_ (.A(_0778_),
    .B(_0780_),
    .Y(_0816_));
 sg13g2_nor2_1 _4830_ (.A(_0815_),
    .B(_0816_),
    .Y(_0817_));
 sg13g2_xnor2_1 _4831_ (.Y(_0818_),
    .A(_0815_),
    .B(_0816_));
 sg13g2_nor2_1 _4832_ (.A(_0799_),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_xor2_1 _4833_ (.B(_0818_),
    .A(_0799_),
    .X(_0820_));
 sg13g2_and2_1 _4834_ (.A(_0798_),
    .B(_0820_),
    .X(_0821_));
 sg13g2_or2_1 _4835_ (.X(_0822_),
    .B(_0820_),
    .A(_0798_));
 sg13g2_xnor2_1 _4836_ (.Y(_0823_),
    .A(_0798_),
    .B(_0820_));
 sg13g2_xnor2_1 _4837_ (.Y(_0824_),
    .A(_0797_),
    .B(_0823_));
 sg13g2_nand2_1 _4838_ (.Y(_0825_),
    .A(_0512_),
    .B(_0824_));
 sg13g2_xnor2_1 _4839_ (.Y(_0826_),
    .A(_0512_),
    .B(_0824_));
 sg13g2_xnor2_1 _4840_ (.Y(_0827_),
    .A(_0796_),
    .B(_0826_));
 sg13g2_xnor2_1 _4841_ (.Y(_0828_),
    .A(\main.demo._q_speed[2] ),
    .B(_0827_));
 sg13g2_xor2_1 _4842_ (.B(_0828_),
    .A(_0795_),
    .X(_0829_));
 sg13g2_inv_1 _4843_ (.Y(_0830_),
    .A(_0829_));
 sg13g2_a21oi_1 _4844_ (.A1(_0797_),
    .A2(_0822_),
    .Y(_0831_),
    .B1(_0821_));
 sg13g2_nor2_1 _4845_ (.A(_0817_),
    .B(_0819_),
    .Y(_0832_));
 sg13g2_nand2_2 _4846_ (.Y(_0833_),
    .A(_0803_),
    .B(_0808_));
 sg13g2_nand2_2 _4847_ (.Y(_0834_),
    .A(net487),
    .B(_0772_));
 sg13g2_nand2_1 _4848_ (.Y(_0835_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .B(_0705_));
 sg13g2_nand3_1 _4849_ (.B(_0705_),
    .C(_0800_),
    .A(net485),
    .Y(_0836_));
 sg13g2_a21o_1 _4850_ (.A2(_0705_),
    .A1(net485),
    .B1(_0800_),
    .X(_0837_));
 sg13g2_nand2_2 _4851_ (.Y(_0838_),
    .A(_0836_),
    .B(_0837_));
 sg13g2_xor2_1 _4852_ (.B(_0838_),
    .A(_0834_),
    .X(_0839_));
 sg13g2_nor2_2 _4853_ (.A(_2950_),
    .B(_0516_),
    .Y(_0840_));
 sg13g2_nor2_2 _4854_ (.A(_0008_),
    .B(_0516_),
    .Y(_0841_));
 sg13g2_nor3_2 _4855_ (.A(_0008_),
    .B(_2950_),
    .C(_0516_),
    .Y(_0842_));
 sg13g2_inv_1 _4856_ (.Y(_0843_),
    .A(_0842_));
 sg13g2_and2_1 _4857_ (.A(_2949_),
    .B(net408),
    .X(_0844_));
 sg13g2_o21ai_1 _4858_ (.B1(_0843_),
    .Y(_0845_),
    .A1(_0840_),
    .A2(_0844_));
 sg13g2_nor2_1 _4859_ (.A(_0810_),
    .B(_0845_),
    .Y(_0846_));
 sg13g2_xor2_1 _4860_ (.B(_0845_),
    .A(_0810_),
    .X(_0847_));
 sg13g2_and2_1 _4861_ (.A(_0839_),
    .B(_0847_),
    .X(_0848_));
 sg13g2_xnor2_1 _4862_ (.Y(_0849_),
    .A(_0839_),
    .B(_0847_));
 sg13g2_nor2_1 _4863_ (.A(_0814_),
    .B(_0849_),
    .Y(_0850_));
 sg13g2_xor2_1 _4864_ (.B(_0849_),
    .A(_0814_),
    .X(_0851_));
 sg13g2_xnor2_1 _4865_ (.Y(_0852_),
    .A(_0833_),
    .B(_0851_));
 sg13g2_or2_1 _4866_ (.X(_0853_),
    .B(_0852_),
    .A(_0832_));
 sg13g2_xnor2_1 _4867_ (.Y(_0854_),
    .A(_0832_),
    .B(_0852_));
 sg13g2_xnor2_1 _4868_ (.Y(_0855_),
    .A(_0831_),
    .B(_0854_));
 sg13g2_nor2_1 _4869_ (.A(_0607_),
    .B(_0855_),
    .Y(_0856_));
 sg13g2_o21ai_1 _4870_ (.B1(_0825_),
    .Y(_0857_),
    .A1(_0796_),
    .A2(_0826_));
 sg13g2_xor2_1 _4871_ (.B(_0855_),
    .A(net412),
    .X(_0858_));
 sg13g2_a21oi_1 _4872_ (.A1(_0857_),
    .A2(_0858_),
    .Y(_0859_),
    .B1(_0856_));
 sg13g2_o21ai_1 _4873_ (.B1(_0853_),
    .Y(_0860_),
    .A1(_0831_),
    .A2(_0854_));
 sg13g2_a21oi_1 _4874_ (.A1(_0833_),
    .A2(_0851_),
    .Y(_0861_),
    .B1(_0850_));
 sg13g2_o21ai_1 _4875_ (.B1(_0836_),
    .Y(_0862_),
    .A1(_0834_),
    .A2(_0838_));
 sg13g2_nor2_2 _4876_ (.A(_0840_),
    .B(_0841_),
    .Y(_0863_));
 sg13g2_nand2_1 _4877_ (.Y(_0864_),
    .A(net484),
    .B(_0772_));
 sg13g2_nor2_2 _4878_ (.A(_0835_),
    .B(_0864_),
    .Y(_0865_));
 sg13g2_xor2_1 _4879_ (.B(_0864_),
    .A(_0835_),
    .X(_0866_));
 sg13g2_xnor2_1 _4880_ (.Y(_0867_),
    .A(_0805_),
    .B(_0866_));
 sg13g2_xnor2_1 _4881_ (.Y(_0868_),
    .A(_0863_),
    .B(_0867_));
 sg13g2_o21ai_1 _4882_ (.B1(_0868_),
    .Y(_0869_),
    .A1(_0846_),
    .A2(_0848_));
 sg13g2_inv_1 _4883_ (.Y(_0870_),
    .A(_0869_));
 sg13g2_nor3_1 _4884_ (.A(_0846_),
    .B(_0848_),
    .C(_0868_),
    .Y(_0871_));
 sg13g2_nor2_1 _4885_ (.A(_0870_),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_xnor2_1 _4886_ (.Y(_0873_),
    .A(_0862_),
    .B(_0872_));
 sg13g2_nor2_1 _4887_ (.A(_0861_),
    .B(_0873_),
    .Y(_0874_));
 sg13g2_xor2_1 _4888_ (.B(_0873_),
    .A(_0861_),
    .X(_0875_));
 sg13g2_xor2_1 _4889_ (.B(_0875_),
    .A(_0860_),
    .X(_0876_));
 sg13g2_nand2_1 _4890_ (.Y(_0877_),
    .A(_0639_),
    .B(_0876_));
 sg13g2_xnor2_1 _4891_ (.Y(_0878_),
    .A(_0639_),
    .B(_0876_));
 sg13g2_xnor2_1 _4892_ (.Y(_0879_),
    .A(_0859_),
    .B(_0878_));
 sg13g2_nor2_1 _4893_ (.A(_0012_),
    .B(_0879_),
    .Y(_0880_));
 sg13g2_xnor2_1 _4894_ (.Y(_0881_),
    .A(_0857_),
    .B(_0858_));
 sg13g2_or2_1 _4895_ (.X(_0882_),
    .B(_0881_),
    .A(_0013_));
 sg13g2_nor2_1 _4896_ (.A(_0014_),
    .B(_0827_),
    .Y(_0883_));
 sg13g2_a21oi_1 _4897_ (.A1(_0795_),
    .A2(_0828_),
    .Y(_0884_),
    .B1(_0883_));
 sg13g2_xnor2_1 _4898_ (.Y(_0885_),
    .A(_0013_),
    .B(_0881_));
 sg13g2_o21ai_1 _4899_ (.B1(_0882_),
    .Y(_0886_),
    .A1(_0884_),
    .A2(_0885_));
 sg13g2_xor2_1 _4900_ (.B(_0879_),
    .A(_0012_),
    .X(_0887_));
 sg13g2_a21oi_1 _4901_ (.A1(_0886_),
    .A2(_0887_),
    .Y(_0888_),
    .B1(_0880_));
 sg13g2_o21ai_1 _4902_ (.B1(_0877_),
    .Y(_0889_),
    .A1(_0859_),
    .A2(_0878_));
 sg13g2_a21oi_1 _4903_ (.A1(_0860_),
    .A2(_0875_),
    .Y(_0890_),
    .B1(_0874_));
 sg13g2_a21oi_1 _4904_ (.A1(_0862_),
    .A2(_0872_),
    .Y(_0891_),
    .B1(_0870_));
 sg13g2_inv_1 _4905_ (.Y(_0892_),
    .A(_0891_));
 sg13g2_a21oi_2 _4906_ (.B1(_0865_),
    .Y(_0893_),
    .A2(_0866_),
    .A1(_0806_));
 sg13g2_nand2_2 _4907_ (.Y(_0894_),
    .A(net487),
    .B(_0517_));
 sg13g2_inv_1 _4908_ (.Y(_0895_),
    .A(_0894_));
 sg13g2_nor2b_1 _4909_ (.A(_0009_),
    .B_N(net408),
    .Y(_0896_));
 sg13g2_nor2b_1 _4910_ (.A(_0009_),
    .B_N(_0772_),
    .Y(_0897_));
 sg13g2_nand2b_1 _4911_ (.Y(_0898_),
    .B(net408),
    .A_N(_0010_));
 sg13g2_nor2b_2 _4912_ (.A(_0010_),
    .B_N(_0897_),
    .Y(_0899_));
 sg13g2_xnor2_1 _4913_ (.Y(_0900_),
    .A(_0897_),
    .B(_0898_));
 sg13g2_xnor2_1 _4914_ (.Y(_0901_),
    .A(_0895_),
    .B(_0900_));
 sg13g2_nor2_1 _4915_ (.A(_0863_),
    .B(_0867_),
    .Y(_0902_));
 sg13g2_nor2b_1 _4916_ (.A(_0863_),
    .B_N(_0901_),
    .Y(_0903_));
 sg13g2_xor2_1 _4917_ (.B(_0902_),
    .A(_0901_),
    .X(_0904_));
 sg13g2_nor2_1 _4918_ (.A(_0893_),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_xor2_1 _4919_ (.B(_0904_),
    .A(_0893_),
    .X(_0906_));
 sg13g2_xnor2_1 _4920_ (.Y(_0907_),
    .A(_0891_),
    .B(_0906_));
 sg13g2_nor2b_1 _4921_ (.A(_0890_),
    .B_N(_0907_),
    .Y(_0908_));
 sg13g2_xnor2_1 _4922_ (.Y(_0909_),
    .A(_0890_),
    .B(_0907_));
 sg13g2_xnor2_1 _4923_ (.Y(_0910_),
    .A(_0702_),
    .B(_0909_));
 sg13g2_nor2b_1 _4924_ (.A(_0910_),
    .B_N(_0889_),
    .Y(_0911_));
 sg13g2_xor2_1 _4925_ (.B(_0910_),
    .A(_0889_),
    .X(_0912_));
 sg13g2_nor2_1 _4926_ (.A(_0007_),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_xor2_1 _4927_ (.B(_0912_),
    .A(_0007_),
    .X(_0914_));
 sg13g2_nor2b_1 _4928_ (.A(_0888_),
    .B_N(_0914_),
    .Y(_0915_));
 sg13g2_xnor2_1 _4929_ (.Y(_0916_),
    .A(_0888_),
    .B(_0914_));
 sg13g2_inv_1 _4930_ (.Y(_0917_),
    .A(_0916_));
 sg13g2_nor2_1 _4931_ (.A(net472),
    .B(net476),
    .Y(_0918_));
 sg13g2_or2_1 _4932_ (.X(_0919_),
    .B(net476),
    .A(net472));
 sg13g2_nor2_2 _4933_ (.A(_2945_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_nand2_2 _4934_ (.Y(_0921_),
    .A(\main.demo._q_speed[1] ),
    .B(net445));
 sg13g2_o21ai_1 _4935_ (.B1(net445),
    .Y(_0922_),
    .A1(\main.demo._q_speed[1] ),
    .A2(\main.demo._q_speed[2] ));
 sg13g2_nand2b_1 _4936_ (.Y(_0923_),
    .B(_0921_),
    .A_N(_0920_));
 sg13g2_a21oi_1 _4937_ (.A1(\main.demo._q_speed[1] ),
    .A2(_0920_),
    .Y(_0924_),
    .B1(_0922_));
 sg13g2_mux2_1 _4938_ (.A0(_0920_),
    .A1(_0924_),
    .S(_0916_),
    .X(_0925_));
 sg13g2_nand2_1 _4939_ (.Y(_0926_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ),
    .B(_0925_));
 sg13g2_xnor2_1 _4940_ (.Y(_0927_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ),
    .B(_0925_));
 sg13g2_inv_1 _4941_ (.Y(_0928_),
    .A(_0927_));
 sg13g2_o21ai_1 _4942_ (.B1(_0926_),
    .Y(_0929_),
    .A1(_0921_),
    .A2(_0927_));
 sg13g2_nand2_1 _4943_ (.Y(_0930_),
    .A(\main.demo._q_speed[3] ),
    .B(net445));
 sg13g2_nand2_1 _4944_ (.Y(_0931_),
    .A(_0916_),
    .B(_0923_));
 sg13g2_xor2_1 _4945_ (.B(_0931_),
    .A(_0930_),
    .X(_0932_));
 sg13g2_xor2_1 _4946_ (.B(_0932_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ),
    .X(_0933_));
 sg13g2_xor2_1 _4947_ (.B(_0933_),
    .A(_0929_),
    .X(_0934_));
 sg13g2_and2_2 _4948_ (.A(net472),
    .B(net476),
    .X(_0935_));
 sg13g2_nand2_2 _4949_ (.Y(_0936_),
    .A(net475),
    .B(net477));
 sg13g2_o21ai_1 _4950_ (.B1(net477),
    .Y(_0937_),
    .A1(net475),
    .A2(_0934_));
 sg13g2_nor2_1 _4951_ (.A(_0830_),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_nor2_1 _4952_ (.A(_0927_),
    .B(_0936_),
    .Y(_0939_));
 sg13g2_nor2b_1 _4953_ (.A(net472),
    .B_N(net476),
    .Y(_0940_));
 sg13g2_nand2_2 _4954_ (.Y(_0941_),
    .A(net460),
    .B(net477));
 sg13g2_nor2b_1 _4955_ (.A(_0018_),
    .B_N(_0932_),
    .Y(_0942_));
 sg13g2_a21o_1 _4956_ (.A2(_0933_),
    .A1(_0929_),
    .B1(_0942_),
    .X(_0943_));
 sg13g2_nand2_2 _4957_ (.Y(_0944_),
    .A(\main.demo._q_speed[4] ),
    .B(net444));
 sg13g2_o21ai_1 _4958_ (.B1(net444),
    .Y(_0945_),
    .A1(\main.demo._q_speed[2] ),
    .A2(\main.demo._q_speed[3] ));
 sg13g2_nand2_1 _4959_ (.Y(_0946_),
    .A(_0921_),
    .B(_0945_));
 sg13g2_nand2_1 _4960_ (.Y(_0947_),
    .A(_0916_),
    .B(_0946_));
 sg13g2_xnor2_1 _4961_ (.Y(_0948_),
    .A(_0944_),
    .B(_0947_));
 sg13g2_nor2_1 _4962_ (.A(_0017_),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_nand2_1 _4963_ (.Y(_0950_),
    .A(_0017_),
    .B(_0948_));
 sg13g2_nand2b_1 _4964_ (.Y(_0951_),
    .B(_0950_),
    .A_N(_0949_));
 sg13g2_xnor2_1 _4965_ (.Y(_0952_),
    .A(_0943_),
    .B(_0951_));
 sg13g2_nand2_1 _4966_ (.Y(_0953_),
    .A(net441),
    .B(_0952_));
 sg13g2_xnor2_1 _4967_ (.Y(_0954_),
    .A(_0884_),
    .B(_0885_));
 sg13g2_inv_1 _4968_ (.Y(_0955_),
    .A(_0954_));
 sg13g2_xnor2_1 _4969_ (.Y(_0956_),
    .A(_0953_),
    .B(_0955_));
 sg13g2_nand4_1 _4970_ (.B(net476),
    .C(_0928_),
    .A(net472),
    .Y(_0957_),
    .D(_0955_));
 sg13g2_xnor2_1 _4971_ (.Y(_0958_),
    .A(_0939_),
    .B(_0956_));
 sg13g2_or3_1 _4972_ (.A(_0830_),
    .B(_0937_),
    .C(_0958_),
    .X(_0959_));
 sg13g2_nor2_2 _4973_ (.A(net459),
    .B(net476),
    .Y(_0960_));
 sg13g2_nand2b_2 _4974_ (.Y(_0961_),
    .B(net472),
    .A_N(net476));
 sg13g2_o21ai_1 _4975_ (.B1(_0957_),
    .Y(_0962_),
    .A1(_0953_),
    .A2(_0954_));
 sg13g2_inv_1 _4976_ (.Y(_0963_),
    .A(_0962_));
 sg13g2_a21oi_1 _4977_ (.A1(_0943_),
    .A2(_0950_),
    .Y(_0964_),
    .B1(_0949_));
 sg13g2_nand2_2 _4978_ (.Y(_0965_),
    .A(\main.demo._q_speed[5] ),
    .B(net444));
 sg13g2_nand2_1 _4979_ (.Y(_0966_),
    .A(_0944_),
    .B(_0945_));
 sg13g2_nand3_1 _4980_ (.B(_0944_),
    .C(_0945_),
    .A(_0922_),
    .Y(_0967_));
 sg13g2_nand2_1 _4981_ (.Y(_0968_),
    .A(_0916_),
    .B(_0967_));
 sg13g2_xor2_1 _4982_ (.B(_0968_),
    .A(_0965_),
    .X(_0969_));
 sg13g2_nand2b_1 _4983_ (.Y(_0970_),
    .B(_0969_),
    .A_N(_0016_));
 sg13g2_xnor2_1 _4984_ (.Y(_0971_),
    .A(_0016_),
    .B(_0969_));
 sg13g2_inv_1 _4985_ (.Y(_0972_),
    .A(_0971_));
 sg13g2_xnor2_1 _4986_ (.Y(_0973_),
    .A(_0964_),
    .B(_0971_));
 sg13g2_xor2_1 _4987_ (.B(_0887_),
    .A(_0886_),
    .X(_0974_));
 sg13g2_nand3_1 _4988_ (.B(_0973_),
    .C(_0974_),
    .A(net441),
    .Y(_0975_));
 sg13g2_a21o_1 _4989_ (.A2(_0973_),
    .A1(net441),
    .B1(_0974_),
    .X(_0976_));
 sg13g2_nand4_1 _4990_ (.B(net477),
    .C(_0934_),
    .A(net472),
    .Y(_0977_),
    .D(_0974_));
 sg13g2_inv_1 _4991_ (.Y(_0978_),
    .A(_0977_));
 sg13g2_a22oi_1 _4992_ (.Y(_0979_),
    .B1(_0975_),
    .B2(_0976_),
    .A2(_0935_),
    .A1(_0934_));
 sg13g2_nor3_1 _4993_ (.A(_0963_),
    .B(_0978_),
    .C(_0979_),
    .Y(_0980_));
 sg13g2_or3_1 _4994_ (.A(_0963_),
    .B(_0978_),
    .C(_0979_),
    .X(_0981_));
 sg13g2_o21ai_1 _4995_ (.B1(_0963_),
    .Y(_0982_),
    .A1(_0978_),
    .A2(_0979_));
 sg13g2_and3_1 _4996_ (.X(_0983_),
    .A(_0960_),
    .B(_0981_),
    .C(_0982_));
 sg13g2_a21oi_1 _4997_ (.A1(_0981_),
    .A2(_0982_),
    .Y(_0984_),
    .B1(_0960_));
 sg13g2_nor3_1 _4998_ (.A(_0959_),
    .B(_0983_),
    .C(_0984_),
    .Y(_0985_));
 sg13g2_xnor2_1 _4999_ (.Y(_0986_),
    .A(_0830_),
    .B(_0937_));
 sg13g2_nor2_2 _5000_ (.A(_0927_),
    .B(_0941_),
    .Y(_0987_));
 sg13g2_xor2_1 _5001_ (.B(_0794_),
    .A(_0793_),
    .X(_0988_));
 sg13g2_nand2_1 _5002_ (.Y(_0989_),
    .A(_0987_),
    .B(_0988_));
 sg13g2_nor2_1 _5003_ (.A(_0986_),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_nor2b_1 _5004_ (.A(_0958_),
    .B_N(_0990_),
    .Y(_0991_));
 sg13g2_xnor2_1 _5005_ (.Y(_0992_),
    .A(_0987_),
    .B(_0988_));
 sg13g2_o21ai_1 _5006_ (.B1(net442),
    .Y(_0993_),
    .A1(\main.demo._q_speed[0] ),
    .A2(_0792_));
 sg13g2_nor2_2 _5007_ (.A(_0793_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_nor2b_1 _5008_ (.A(_0992_),
    .B_N(_0994_),
    .Y(_0995_));
 sg13g2_nor2b_1 _5009_ (.A(_0986_),
    .B_N(_0995_),
    .Y(_0996_));
 sg13g2_nor2_1 _5010_ (.A(_0938_),
    .B(_0990_),
    .Y(_0997_));
 sg13g2_xor2_1 _5011_ (.B(_0997_),
    .A(_0958_),
    .X(_0998_));
 sg13g2_a21o_1 _5012_ (.A2(_0998_),
    .A1(_0996_),
    .B1(_0991_),
    .X(_0999_));
 sg13g2_o21ai_1 _5013_ (.B1(_0959_),
    .Y(_1000_),
    .A1(_0983_),
    .A2(_0984_));
 sg13g2_nor2b_1 _5014_ (.A(_0985_),
    .B_N(_1000_),
    .Y(_1001_));
 sg13g2_a21oi_1 _5015_ (.A1(_0999_),
    .A2(_1000_),
    .Y(_1002_),
    .B1(_0985_));
 sg13g2_or2_1 _5016_ (.X(_1003_),
    .B(_0983_),
    .A(_0980_));
 sg13g2_nor2_2 _5017_ (.A(_0927_),
    .B(_0961_),
    .Y(_1004_));
 sg13g2_nand2_1 _5018_ (.Y(_1005_),
    .A(_0928_),
    .B(_0960_));
 sg13g2_nand2_1 _5019_ (.Y(_1006_),
    .A(_0975_),
    .B(_0977_));
 sg13g2_nand2_1 _5020_ (.Y(_1007_),
    .A(_0935_),
    .B(_0952_));
 sg13g2_o21ai_1 _5021_ (.B1(_0970_),
    .Y(_1008_),
    .A1(_0964_),
    .A2(_0972_));
 sg13g2_nand2_2 _5022_ (.Y(_1009_),
    .A(\main.demo._q_speed[6] ),
    .B(net444));
 sg13g2_nand3_1 _5023_ (.B(_0945_),
    .C(_0965_),
    .A(_0944_),
    .Y(_1010_));
 sg13g2_o21ai_1 _5024_ (.B1(_0916_),
    .Y(_1011_),
    .A1(_0923_),
    .A2(_1010_));
 sg13g2_xor2_1 _5025_ (.B(_1011_),
    .A(_1009_),
    .X(_1012_));
 sg13g2_xor2_1 _5026_ (.B(_1012_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[5] ),
    .X(_1013_));
 sg13g2_xor2_1 _5027_ (.B(_1013_),
    .A(_1008_),
    .X(_1014_));
 sg13g2_xnor2_1 _5028_ (.Y(_1015_),
    .A(_1008_),
    .B(_1013_));
 sg13g2_nand2_1 _5029_ (.Y(_1016_),
    .A(net442),
    .B(_1014_));
 sg13g2_nor3_1 _5030_ (.A(_0917_),
    .B(_0941_),
    .C(_1015_),
    .Y(_1017_));
 sg13g2_a21oi_1 _5031_ (.A1(net441),
    .A2(_1014_),
    .Y(_1018_),
    .B1(_0916_));
 sg13g2_nand4_1 _5032_ (.B(net477),
    .C(_0916_),
    .A(net472),
    .Y(_1019_),
    .D(_0952_));
 sg13g2_o21ai_1 _5033_ (.B1(_1007_),
    .Y(_1020_),
    .A1(_1017_),
    .A2(_1018_));
 sg13g2_nand3_1 _5034_ (.B(_1019_),
    .C(_1020_),
    .A(_1006_),
    .Y(_1021_));
 sg13g2_a21o_1 _5035_ (.A2(_1020_),
    .A1(_1019_),
    .B1(_1006_),
    .X(_1022_));
 sg13g2_nand3_1 _5036_ (.B(_1021_),
    .C(_1022_),
    .A(_1004_),
    .Y(_1023_));
 sg13g2_a21o_1 _5037_ (.A2(_1022_),
    .A1(_1021_),
    .B1(_1004_),
    .X(_1024_));
 sg13g2_and3_1 _5038_ (.X(_1025_),
    .A(_1003_),
    .B(_1023_),
    .C(_1024_));
 sg13g2_nand3_1 _5039_ (.B(_1023_),
    .C(_1024_),
    .A(_1003_),
    .Y(_1026_));
 sg13g2_a21oi_1 _5040_ (.A1(_1023_),
    .A2(_1024_),
    .Y(_1027_),
    .B1(_1003_));
 sg13g2_nor3_1 _5041_ (.A(_1002_),
    .B(_1025_),
    .C(_1027_),
    .Y(_1028_));
 sg13g2_o21ai_1 _5042_ (.B1(_1002_),
    .Y(_1029_),
    .A1(_1025_),
    .A2(_1027_));
 sg13g2_nor2b_1 _5043_ (.A(_1028_),
    .B_N(_1029_),
    .Y(_1030_));
 sg13g2_nor2_1 _5044_ (.A(net443),
    .B(_1015_),
    .Y(_1031_));
 sg13g2_xnor2_1 _5045_ (.Y(_1032_),
    .A(_1030_),
    .B(_1031_));
 sg13g2_nor2_1 _5046_ (.A(_0582_),
    .B(_0599_),
    .Y(_1033_));
 sg13g2_xor2_1 _5047_ (.B(_0590_),
    .A(_0579_),
    .X(_1034_));
 sg13g2_nor2b_1 _5048_ (.A(_0586_),
    .B_N(_1034_),
    .Y(_1035_));
 sg13g2_nor2_1 _5049_ (.A(_1033_),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_xnor2_1 _5050_ (.Y(_1037_),
    .A(_0586_),
    .B(_1034_));
 sg13g2_nand2b_1 _5051_ (.Y(_1038_),
    .B(_1037_),
    .A_N(_0596_));
 sg13g2_nor2b_1 _5052_ (.A(_0595_),
    .B_N(_0603_),
    .Y(_1039_));
 sg13g2_xnor2_1 _5053_ (.Y(_1040_),
    .A(_0595_),
    .B(_0603_));
 sg13g2_xor2_1 _5054_ (.B(_0617_),
    .A(_0599_),
    .X(_1041_));
 sg13g2_xnor2_1 _5055_ (.Y(_1042_),
    .A(_0616_),
    .B(_1041_));
 sg13g2_xor2_1 _5056_ (.B(_1042_),
    .A(_1040_),
    .X(_1043_));
 sg13g2_nand2b_1 _5057_ (.Y(_1044_),
    .B(_1043_),
    .A_N(_1038_));
 sg13g2_xor2_1 _5058_ (.B(_1043_),
    .A(_1038_),
    .X(_1045_));
 sg13g2_xor2_1 _5059_ (.B(_1037_),
    .A(_0596_),
    .X(_1046_));
 sg13g2_o21ai_1 _5060_ (.B1(_0747_),
    .Y(_1047_),
    .A1(_0582_),
    .A2(_0666_));
 sg13g2_nand3_1 _5061_ (.B(_0748_),
    .C(_1047_),
    .A(_0665_),
    .Y(_1048_));
 sg13g2_a21oi_1 _5062_ (.A1(_0665_),
    .A2(_0748_),
    .Y(_1049_),
    .B1(_1047_));
 sg13g2_a21oi_1 _5063_ (.A1(_1046_),
    .A2(_1048_),
    .Y(_1050_),
    .B1(_1049_));
 sg13g2_o21ai_1 _5064_ (.B1(_1050_),
    .Y(_1051_),
    .A1(_1036_),
    .A2(_1045_));
 sg13g2_a21o_1 _5065_ (.A2(_1045_),
    .A1(_1036_),
    .B1(_1051_),
    .X(_1052_));
 sg13g2_o21ai_1 _5066_ (.B1(_1052_),
    .Y(_1053_),
    .A1(_0744_),
    .A2(_0752_));
 sg13g2_o21ai_1 _5067_ (.B1(_1044_),
    .Y(_1054_),
    .A1(_1036_),
    .A2(_1045_));
 sg13g2_a21oi_1 _5068_ (.A1(_1040_),
    .A2(_1042_),
    .Y(_1055_),
    .B1(_1039_));
 sg13g2_nand2_1 _5069_ (.Y(_1056_),
    .A(_0602_),
    .B(_0634_));
 sg13g2_xnor2_1 _5070_ (.Y(_1057_),
    .A(_0602_),
    .B(_0634_));
 sg13g2_nand3_1 _5071_ (.B(_0613_),
    .C(_0614_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .Y(_1058_));
 sg13g2_xor2_1 _5072_ (.B(_1058_),
    .A(_0635_),
    .X(_1059_));
 sg13g2_nand2_1 _5073_ (.Y(_1060_),
    .A(_0646_),
    .B(_1059_));
 sg13g2_xnor2_1 _5074_ (.Y(_1061_),
    .A(_0646_),
    .B(_1059_));
 sg13g2_xor2_1 _5075_ (.B(_1061_),
    .A(_1057_),
    .X(_1062_));
 sg13g2_nand2b_1 _5076_ (.Y(_1063_),
    .B(_1062_),
    .A_N(_1055_));
 sg13g2_xnor2_1 _5077_ (.Y(_1064_),
    .A(_1055_),
    .B(_1062_));
 sg13g2_a21oi_1 _5078_ (.A1(_0617_),
    .A2(_0627_),
    .Y(_1065_),
    .B1(_0599_));
 sg13g2_nor2_1 _5079_ (.A(_0628_),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_nand2b_1 _5080_ (.Y(_1067_),
    .B(_1064_),
    .A_N(_1066_));
 sg13g2_xor2_1 _5081_ (.B(_1066_),
    .A(_1064_),
    .X(_1068_));
 sg13g2_nor2b_1 _5082_ (.A(_1068_),
    .B_N(_1054_),
    .Y(_1069_));
 sg13g2_xnor2_1 _5083_ (.Y(_1070_),
    .A(_1054_),
    .B(_1068_));
 sg13g2_xnor2_1 _5084_ (.Y(_1071_),
    .A(_1053_),
    .B(_1070_));
 sg13g2_inv_1 _5085_ (.Y(_1072_),
    .A(_1071_));
 sg13g2_xor2_1 _5086_ (.B(\main.demo._t___stage___block_3_x[0] ),
    .A(\main.demo._t___stage___block_3_y[0] ),
    .X(_1073_));
 sg13g2_xnor2_1 _5087_ (.Y(_1074_),
    .A(\main.demo._t___stage___block_3_y[0] ),
    .B(\main.demo._t___stage___block_3_x[0] ));
 sg13g2_xnor2_1 _5088_ (.Y(_1075_),
    .A(_0545_),
    .B(_1071_));
 sg13g2_and3_1 _5089_ (.X(_1076_),
    .A(_0755_),
    .B(net436),
    .C(_1075_));
 sg13g2_nand3_1 _5090_ (.B(_0753_),
    .C(net439),
    .A(_0553_),
    .Y(_1077_));
 sg13g2_a22oi_1 _5091_ (.Y(_1078_),
    .B1(_1077_),
    .B2(_0755_),
    .A2(_1075_),
    .A1(net436));
 sg13g2_or2_2 _5092_ (.X(_1079_),
    .B(_1078_),
    .A(_1076_));
 sg13g2_inv_1 _5093_ (.Y(_1080_),
    .A(_1079_));
 sg13g2_nand2_1 _5094_ (.Y(_1081_),
    .A(\main.demo._q_speed[0] ),
    .B(_1080_));
 sg13g2_o21ai_1 _5095_ (.B1(_0743_),
    .Y(_1082_),
    .A1(_0744_),
    .A2(_0752_));
 sg13g2_a21oi_1 _5096_ (.A1(_0587_),
    .A2(_0735_),
    .Y(_1083_),
    .B1(_0733_));
 sg13g2_nand2b_1 _5097_ (.Y(_1084_),
    .B(_0626_),
    .A_N(_0637_));
 sg13g2_xnor2_1 _5098_ (.Y(_1085_),
    .A(_0626_),
    .B(_0637_));
 sg13g2_nand2b_1 _5099_ (.Y(_1086_),
    .B(_1085_),
    .A_N(_0649_));
 sg13g2_xnor2_1 _5100_ (.Y(_1087_),
    .A(_0649_),
    .B(_1085_));
 sg13g2_a21o_1 _5101_ (.A2(_0729_),
    .A1(_0629_),
    .B1(_0730_),
    .X(_1088_));
 sg13g2_and2_1 _5102_ (.A(_1087_),
    .B(_1088_),
    .X(_1089_));
 sg13g2_xor2_1 _5103_ (.B(_1088_),
    .A(_1087_),
    .X(_1090_));
 sg13g2_xnor2_1 _5104_ (.Y(_1091_),
    .A(_0628_),
    .B(_1090_));
 sg13g2_nor2_1 _5105_ (.A(_1083_),
    .B(_1091_),
    .Y(_1092_));
 sg13g2_xor2_1 _5106_ (.B(_1091_),
    .A(_1083_),
    .X(_1093_));
 sg13g2_xor2_1 _5107_ (.B(_1093_),
    .A(_1082_),
    .X(_1094_));
 sg13g2_nor2b_1 _5108_ (.A(_0545_),
    .B_N(_1094_),
    .Y(_1095_));
 sg13g2_xnor2_1 _5109_ (.Y(_1096_),
    .A(_0545_),
    .B(_1094_));
 sg13g2_xnor2_1 _5110_ (.Y(_1097_),
    .A(_0755_),
    .B(_1096_));
 sg13g2_a21oi_1 _5111_ (.A1(_1053_),
    .A2(_1070_),
    .Y(_1098_),
    .B1(_1069_));
 sg13g2_nand2_1 _5112_ (.Y(_1099_),
    .A(_1063_),
    .B(_1067_));
 sg13g2_o21ai_1 _5113_ (.B1(_1060_),
    .Y(_1100_),
    .A1(_0617_),
    .A2(_0690_));
 sg13g2_o21ai_1 _5114_ (.B1(_1056_),
    .Y(_1101_),
    .A1(_1057_),
    .A2(_1061_));
 sg13g2_nor2b_1 _5115_ (.A(_0633_),
    .B_N(_0694_),
    .Y(_1102_));
 sg13g2_xnor2_1 _5116_ (.Y(_1103_),
    .A(_0633_),
    .B(_0694_));
 sg13g2_xnor2_1 _5117_ (.Y(_1104_),
    .A(_0645_),
    .B(_0690_));
 sg13g2_nor2_1 _5118_ (.A(_0710_),
    .B(_1104_),
    .Y(_1105_));
 sg13g2_xor2_1 _5119_ (.B(_1104_),
    .A(_0710_),
    .X(_1106_));
 sg13g2_xnor2_1 _5120_ (.Y(_1107_),
    .A(_1103_),
    .B(_1106_));
 sg13g2_nor2b_1 _5121_ (.A(_1107_),
    .B_N(_1101_),
    .Y(_1108_));
 sg13g2_xor2_1 _5122_ (.B(_1107_),
    .A(_1101_),
    .X(_1109_));
 sg13g2_nor2b_1 _5123_ (.A(_1109_),
    .B_N(_1100_),
    .Y(_1110_));
 sg13g2_xnor2_1 _5124_ (.Y(_1111_),
    .A(_1100_),
    .B(_1109_));
 sg13g2_nand2_1 _5125_ (.Y(_1112_),
    .A(_1099_),
    .B(_1111_));
 sg13g2_nor2_1 _5126_ (.A(_1099_),
    .B(_1111_),
    .Y(_1113_));
 sg13g2_xor2_1 _5127_ (.B(_1111_),
    .A(_1099_),
    .X(_1114_));
 sg13g2_xnor2_1 _5128_ (.Y(_1115_),
    .A(_1098_),
    .B(_1114_));
 sg13g2_nand2b_1 _5129_ (.Y(_1116_),
    .B(_1115_),
    .A_N(net413));
 sg13g2_xor2_1 _5130_ (.B(_1115_),
    .A(net413),
    .X(_1117_));
 sg13g2_o21ai_1 _5131_ (.B1(_0756_),
    .Y(_1118_),
    .A1(_0757_),
    .A2(_1072_));
 sg13g2_or2_1 _5132_ (.X(_1119_),
    .B(_1118_),
    .A(_1117_));
 sg13g2_a21oi_1 _5133_ (.A1(_1117_),
    .A2(_1118_),
    .Y(_1120_),
    .B1(net439));
 sg13g2_a22oi_1 _5134_ (.Y(_1121_),
    .B1(_1119_),
    .B2(_1120_),
    .A2(_1097_),
    .A1(net439));
 sg13g2_or2_1 _5135_ (.X(_1122_),
    .B(_1121_),
    .A(_0015_));
 sg13g2_and2_1 _5136_ (.A(_0015_),
    .B(_1121_),
    .X(_1123_));
 sg13g2_xor2_1 _5137_ (.B(_1121_),
    .A(_0015_),
    .X(_1124_));
 sg13g2_xnor2_1 _5138_ (.Y(_1125_),
    .A(_1081_),
    .B(_1124_));
 sg13g2_nand2_1 _5139_ (.Y(_1126_),
    .A(_0987_),
    .B(_1125_));
 sg13g2_o21ai_1 _5140_ (.B1(_1122_),
    .Y(_1127_),
    .A1(_1081_),
    .A2(_1123_));
 sg13g2_a21oi_1 _5141_ (.A1(_0754_),
    .A2(_1096_),
    .Y(_1128_),
    .B1(_1095_));
 sg13g2_a21oi_2 _5142_ (.B1(_1092_),
    .Y(_1129_),
    .A2(_1093_),
    .A1(_1082_));
 sg13g2_a21o_1 _5143_ (.A2(_1090_),
    .A1(_0628_),
    .B1(_1089_),
    .X(_1130_));
 sg13g2_nand2_1 _5144_ (.Y(_1131_),
    .A(_1084_),
    .B(_1086_));
 sg13g2_nand2_1 _5145_ (.Y(_1132_),
    .A(_0688_),
    .B(_0696_));
 sg13g2_xnor2_1 _5146_ (.Y(_1133_),
    .A(_0688_),
    .B(_0696_));
 sg13g2_xor2_1 _5147_ (.B(_1133_),
    .A(_0712_),
    .X(_1134_));
 sg13g2_and2_1 _5148_ (.A(_1131_),
    .B(_1134_),
    .X(_1135_));
 sg13g2_xor2_1 _5149_ (.B(_1134_),
    .A(_1131_),
    .X(_1136_));
 sg13g2_xnor2_1 _5150_ (.Y(_1137_),
    .A(_0648_),
    .B(_1136_));
 sg13g2_nand2b_1 _5151_ (.Y(_1138_),
    .B(_1130_),
    .A_N(_1137_));
 sg13g2_xor2_1 _5152_ (.B(_1137_),
    .A(_1130_),
    .X(_1139_));
 sg13g2_xor2_1 _5153_ (.B(_1139_),
    .A(_1129_),
    .X(_1140_));
 sg13g2_nor2b_1 _5154_ (.A(net413),
    .B_N(_1140_),
    .Y(_1141_));
 sg13g2_xor2_1 _5155_ (.B(_1140_),
    .A(net413),
    .X(_1142_));
 sg13g2_nor2_1 _5156_ (.A(_1128_),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_a21oi_1 _5157_ (.A1(_1128_),
    .A2(_1142_),
    .Y(_1144_),
    .B1(net436));
 sg13g2_nand2b_1 _5158_ (.Y(_1145_),
    .B(_1144_),
    .A_N(_1143_));
 sg13g2_o21ai_1 _5159_ (.B1(_1116_),
    .Y(_1146_),
    .A1(_1117_),
    .A2(_1118_));
 sg13g2_o21ai_1 _5160_ (.B1(_1112_),
    .Y(_1147_),
    .A1(_1098_),
    .A2(_1113_));
 sg13g2_nor2_1 _5161_ (.A(_1108_),
    .B(_1110_),
    .Y(_1148_));
 sg13g2_a21oi_1 _5162_ (.A1(_0647_),
    .A2(_0770_),
    .Y(_1149_),
    .B1(_1105_));
 sg13g2_a21o_1 _5163_ (.A2(_1106_),
    .A1(_1103_),
    .B1(_1102_),
    .X(_1150_));
 sg13g2_nor2b_1 _5164_ (.A(_0693_),
    .B_N(_0769_),
    .Y(_1151_));
 sg13g2_xnor2_1 _5165_ (.Y(_1152_),
    .A(_0693_),
    .B(_0769_));
 sg13g2_nand3_1 _5166_ (.B(_0705_),
    .C(_0770_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .Y(_1153_));
 sg13g2_xor2_1 _5167_ (.B(_0775_),
    .A(_0770_),
    .X(_1154_));
 sg13g2_xor2_1 _5168_ (.B(_1154_),
    .A(_0774_),
    .X(_1155_));
 sg13g2_xor2_1 _5169_ (.B(_1155_),
    .A(_1152_),
    .X(_1156_));
 sg13g2_nand2_1 _5170_ (.Y(_1157_),
    .A(_1150_),
    .B(_1156_));
 sg13g2_xor2_1 _5171_ (.B(_1156_),
    .A(_1150_),
    .X(_1158_));
 sg13g2_inv_1 _5172_ (.Y(_1159_),
    .A(_1158_));
 sg13g2_xor2_1 _5173_ (.B(_1158_),
    .A(_1149_),
    .X(_1160_));
 sg13g2_nor2_1 _5174_ (.A(_1148_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_xor2_1 _5175_ (.B(_1160_),
    .A(_1148_),
    .X(_1162_));
 sg13g2_xnor2_1 _5176_ (.Y(_1163_),
    .A(_1147_),
    .B(_1162_));
 sg13g2_nor2b_1 _5177_ (.A(_1163_),
    .B_N(_0533_),
    .Y(_1164_));
 sg13g2_xnor2_1 _5178_ (.Y(_1165_),
    .A(_0533_),
    .B(_1163_));
 sg13g2_and2_1 _5179_ (.A(_1146_),
    .B(_1165_),
    .X(_1166_));
 sg13g2_o21ai_1 _5180_ (.B1(net436),
    .Y(_1167_),
    .A1(_1146_),
    .A2(_1165_));
 sg13g2_o21ai_1 _5181_ (.B1(_1145_),
    .Y(_1168_),
    .A1(_1166_),
    .A2(_1167_));
 sg13g2_xnor2_1 _5182_ (.Y(_1169_),
    .A(_2945_),
    .B(_1168_));
 sg13g2_xnor2_1 _5183_ (.Y(_1170_),
    .A(_1127_),
    .B(_1169_));
 sg13g2_o21ai_1 _5184_ (.B1(_1138_),
    .Y(_1171_),
    .A1(_1129_),
    .A2(_1139_));
 sg13g2_a21oi_1 _5185_ (.A1(_0648_),
    .A2(_1136_),
    .Y(_1172_),
    .B1(_1135_));
 sg13g2_o21ai_1 _5186_ (.B1(_1132_),
    .Y(_1173_),
    .A1(_0712_),
    .A2(_1133_));
 sg13g2_nor2_1 _5187_ (.A(_0763_),
    .B(_0771_),
    .Y(_1174_));
 sg13g2_xor2_1 _5188_ (.B(_0771_),
    .A(_0763_),
    .X(_1175_));
 sg13g2_xnor2_1 _5189_ (.Y(_1176_),
    .A(_0777_),
    .B(_1175_));
 sg13g2_nand2b_1 _5190_ (.Y(_1177_),
    .B(_1173_),
    .A_N(_1176_));
 sg13g2_xor2_1 _5191_ (.B(_1176_),
    .A(_1173_),
    .X(_1178_));
 sg13g2_xnor2_1 _5192_ (.Y(_1179_),
    .A(_0711_),
    .B(_1178_));
 sg13g2_nor2_1 _5193_ (.A(_1172_),
    .B(_1179_),
    .Y(_1180_));
 sg13g2_xor2_1 _5194_ (.B(_1179_),
    .A(_1172_),
    .X(_1181_));
 sg13g2_xnor2_1 _5195_ (.Y(_1182_),
    .A(_1171_),
    .B(_1181_));
 sg13g2_nand2b_1 _5196_ (.Y(_1183_),
    .B(_0533_),
    .A_N(_1182_));
 sg13g2_xnor2_1 _5197_ (.Y(_1184_),
    .A(_0533_),
    .B(_1182_));
 sg13g2_o21ai_1 _5198_ (.B1(_1184_),
    .Y(_1185_),
    .A1(_1141_),
    .A2(_1143_));
 sg13g2_a21oi_2 _5199_ (.B1(_1180_),
    .Y(_1186_),
    .A2(_1181_),
    .A1(_1171_));
 sg13g2_o21ai_1 _5200_ (.B1(_1177_),
    .Y(_1187_),
    .A1(_0711_),
    .A2(_1178_));
 sg13g2_a21oi_1 _5201_ (.A1(_0777_),
    .A2(_1175_),
    .Y(_1188_),
    .B1(_1174_));
 sg13g2_nor2_1 _5202_ (.A(_0799_),
    .B(_0809_),
    .Y(_1189_));
 sg13g2_xor2_1 _5203_ (.B(_0809_),
    .A(_0799_),
    .X(_1190_));
 sg13g2_xnor2_1 _5204_ (.Y(_1191_),
    .A(_0812_),
    .B(_1190_));
 sg13g2_xor2_1 _5205_ (.B(_1191_),
    .A(_1188_),
    .X(_1192_));
 sg13g2_nand2_1 _5206_ (.Y(_1193_),
    .A(_0776_),
    .B(_1192_));
 sg13g2_xnor2_1 _5207_ (.Y(_1194_),
    .A(_0776_),
    .B(_1192_));
 sg13g2_nand2b_1 _5208_ (.Y(_1195_),
    .B(_1187_),
    .A_N(_1194_));
 sg13g2_xor2_1 _5209_ (.B(_1194_),
    .A(_1187_),
    .X(_1196_));
 sg13g2_xor2_1 _5210_ (.B(_1196_),
    .A(_1186_),
    .X(_1197_));
 sg13g2_and2_1 _5211_ (.A(_0512_),
    .B(_1197_),
    .X(_1198_));
 sg13g2_xnor2_1 _5212_ (.Y(_1199_),
    .A(_0512_),
    .B(_1197_));
 sg13g2_nand3_1 _5213_ (.B(_1185_),
    .C(_1199_),
    .A(_1183_),
    .Y(_1200_));
 sg13g2_a21oi_1 _5214_ (.A1(_1183_),
    .A2(_1185_),
    .Y(_1201_),
    .B1(_1199_));
 sg13g2_a21o_1 _5215_ (.A2(_1185_),
    .A1(_1183_),
    .B1(_1199_),
    .X(_1202_));
 sg13g2_a21oi_1 _5216_ (.A1(_1200_),
    .A2(_1202_),
    .Y(_1203_),
    .B1(net436));
 sg13g2_a21oi_1 _5217_ (.A1(_1147_),
    .A2(_1162_),
    .Y(_1204_),
    .B1(_1161_));
 sg13g2_o21ai_1 _5218_ (.B1(_1157_),
    .Y(_1205_),
    .A1(_1149_),
    .A2(_1159_));
 sg13g2_o21ai_1 _5219_ (.B1(_1153_),
    .Y(_1206_),
    .A1(_0774_),
    .A2(_1154_));
 sg13g2_a21o_1 _5220_ (.A2(_1155_),
    .A1(_1152_),
    .B1(_1151_),
    .X(_1207_));
 sg13g2_xnor2_1 _5221_ (.Y(_1208_),
    .A(_0768_),
    .B(_0804_));
 sg13g2_nor2_1 _5222_ (.A(_0773_),
    .B(_0807_),
    .Y(_1209_));
 sg13g2_xor2_1 _5223_ (.B(_0807_),
    .A(_0773_),
    .X(_1210_));
 sg13g2_xnor2_1 _5224_ (.Y(_1211_),
    .A(_0708_),
    .B(_1210_));
 sg13g2_nor2b_1 _5225_ (.A(_1208_),
    .B_N(_1211_),
    .Y(_1212_));
 sg13g2_xnor2_1 _5226_ (.Y(_1213_),
    .A(_1208_),
    .B(_1211_));
 sg13g2_xor2_1 _5227_ (.B(_1213_),
    .A(_1207_),
    .X(_1214_));
 sg13g2_and2_1 _5228_ (.A(_1206_),
    .B(_1214_),
    .X(_1215_));
 sg13g2_xor2_1 _5229_ (.B(_1214_),
    .A(_1206_),
    .X(_1216_));
 sg13g2_nand2_1 _5230_ (.Y(_1217_),
    .A(_1205_),
    .B(_1216_));
 sg13g2_nor2_1 _5231_ (.A(_1205_),
    .B(_1216_),
    .Y(_1218_));
 sg13g2_xor2_1 _5232_ (.B(_1216_),
    .A(_1205_),
    .X(_1219_));
 sg13g2_xnor2_1 _5233_ (.Y(_1220_),
    .A(_1204_),
    .B(_1219_));
 sg13g2_nand2_1 _5234_ (.Y(_1221_),
    .A(_0512_),
    .B(_1220_));
 sg13g2_a21oi_1 _5235_ (.A1(_1146_),
    .A2(_1165_),
    .Y(_1222_),
    .B1(_1164_));
 sg13g2_xnor2_1 _5236_ (.Y(_1223_),
    .A(_0512_),
    .B(_1220_));
 sg13g2_or2_1 _5237_ (.X(_1224_),
    .B(_1223_),
    .A(_1222_));
 sg13g2_o21ai_1 _5238_ (.B1(_1221_),
    .Y(_1225_),
    .A1(_1222_),
    .A2(_1223_));
 sg13g2_o21ai_1 _5239_ (.B1(_1217_),
    .Y(_1226_),
    .A1(_1204_),
    .A2(_1218_));
 sg13g2_a21oi_1 _5240_ (.A1(_1207_),
    .A2(_1213_),
    .Y(_1227_),
    .B1(_1215_));
 sg13g2_a21oi_1 _5241_ (.A1(_0709_),
    .A2(_1210_),
    .Y(_1228_),
    .B1(_1209_));
 sg13g2_a21oi_1 _5242_ (.A1(_0768_),
    .A2(_0804_),
    .Y(_1229_),
    .B1(_1212_));
 sg13g2_inv_1 _5243_ (.Y(_1230_),
    .A(_1229_));
 sg13g2_xnor2_1 _5244_ (.Y(_1231_),
    .A(_0803_),
    .B(_0838_));
 sg13g2_xnor2_1 _5245_ (.Y(_1232_),
    .A(_0834_),
    .B(_0844_));
 sg13g2_nand2_1 _5246_ (.Y(_1233_),
    .A(_0840_),
    .B(_1232_));
 sg13g2_xor2_1 _5247_ (.B(_1232_),
    .A(_0840_),
    .X(_1234_));
 sg13g2_nand2b_1 _5248_ (.Y(_1235_),
    .B(_1234_),
    .A_N(_1231_));
 sg13g2_xnor2_1 _5249_ (.Y(_1236_),
    .A(_1231_),
    .B(_1234_));
 sg13g2_xnor2_1 _5250_ (.Y(_1237_),
    .A(_1229_),
    .B(_1236_));
 sg13g2_nor2b_1 _5251_ (.A(_1228_),
    .B_N(_1237_),
    .Y(_1238_));
 sg13g2_xnor2_1 _5252_ (.Y(_1239_),
    .A(_1228_),
    .B(_1237_));
 sg13g2_nor2b_1 _5253_ (.A(_1227_),
    .B_N(_1239_),
    .Y(_1240_));
 sg13g2_xnor2_1 _5254_ (.Y(_1241_),
    .A(_1227_),
    .B(_1239_));
 sg13g2_xnor2_1 _5255_ (.Y(_1242_),
    .A(_1226_),
    .B(_1241_));
 sg13g2_nand2_1 _5256_ (.Y(_1243_),
    .A(net412),
    .B(_1242_));
 sg13g2_nor2_1 _5257_ (.A(net412),
    .B(_1242_),
    .Y(_1244_));
 sg13g2_xor2_1 _5258_ (.B(_1242_),
    .A(net412),
    .X(_1245_));
 sg13g2_xnor2_1 _5259_ (.Y(_1246_),
    .A(_1225_),
    .B(_1245_));
 sg13g2_a21oi_2 _5260_ (.B1(_1203_),
    .Y(_1247_),
    .A2(_1246_),
    .A1(net436));
 sg13g2_nor2b_1 _5261_ (.A(_0012_),
    .B_N(_1247_),
    .Y(_1248_));
 sg13g2_or3_1 _5262_ (.A(_1141_),
    .B(_1143_),
    .C(_1184_),
    .X(_1249_));
 sg13g2_and2_1 _5263_ (.A(_1185_),
    .B(_1249_),
    .X(_1250_));
 sg13g2_a21oi_1 _5264_ (.A1(_1222_),
    .A2(_1223_),
    .Y(_1251_),
    .B1(net439));
 sg13g2_a22oi_1 _5265_ (.Y(_1252_),
    .B1(_1251_),
    .B2(_1224_),
    .A2(_1250_),
    .A1(net439));
 sg13g2_or2_1 _5266_ (.X(_1253_),
    .B(_1252_),
    .A(_0013_));
 sg13g2_a22oi_1 _5267_ (.Y(_1254_),
    .B1(_1169_),
    .B2(_1127_),
    .A2(_1168_),
    .A1(_2951_));
 sg13g2_xnor2_1 _5268_ (.Y(_1255_),
    .A(_0013_),
    .B(_1252_));
 sg13g2_o21ai_1 _5269_ (.B1(_1253_),
    .Y(_1256_),
    .A1(_1254_),
    .A2(_1255_));
 sg13g2_xnor2_1 _5270_ (.Y(_1257_),
    .A(_0012_),
    .B(_1247_));
 sg13g2_a21oi_1 _5271_ (.A1(_1256_),
    .A2(_1257_),
    .Y(_1258_),
    .B1(_1248_));
 sg13g2_o21ai_1 _5272_ (.B1(_1195_),
    .Y(_1259_),
    .A1(_1186_),
    .A2(_1196_));
 sg13g2_o21ai_1 _5273_ (.B1(_1193_),
    .Y(_1260_),
    .A1(_1188_),
    .A2(_1191_));
 sg13g2_a21oi_2 _5274_ (.B1(_1189_),
    .Y(_1261_),
    .A2(_1190_),
    .A1(_0812_));
 sg13g2_nand2_1 _5275_ (.Y(_1262_),
    .A(_0833_),
    .B(_0839_));
 sg13g2_xnor2_1 _5276_ (.Y(_1263_),
    .A(_0833_),
    .B(_0839_));
 sg13g2_xor2_1 _5277_ (.B(_1263_),
    .A(_0845_),
    .X(_1264_));
 sg13g2_nor2b_1 _5278_ (.A(_1261_),
    .B_N(_1264_),
    .Y(_1265_));
 sg13g2_xnor2_1 _5279_ (.Y(_1266_),
    .A(_1261_),
    .B(_1264_));
 sg13g2_xnor2_1 _5280_ (.Y(_1267_),
    .A(_0810_),
    .B(_1266_));
 sg13g2_nand2_1 _5281_ (.Y(_1268_),
    .A(_1260_),
    .B(_1267_));
 sg13g2_xor2_1 _5282_ (.B(_1267_),
    .A(_1260_),
    .X(_1269_));
 sg13g2_nand2_1 _5283_ (.Y(_1270_),
    .A(_1259_),
    .B(_1269_));
 sg13g2_xnor2_1 _5284_ (.Y(_1271_),
    .A(_1259_),
    .B(_1269_));
 sg13g2_nor2_1 _5285_ (.A(net412),
    .B(_1271_),
    .Y(_1272_));
 sg13g2_xor2_1 _5286_ (.B(_1271_),
    .A(net412),
    .X(_1273_));
 sg13g2_nor3_1 _5287_ (.A(_1198_),
    .B(_1201_),
    .C(_1273_),
    .Y(_1274_));
 sg13g2_o21ai_1 _5288_ (.B1(_1273_),
    .Y(_1275_),
    .A1(_1198_),
    .A2(_1201_));
 sg13g2_nor2_1 _5289_ (.A(net437),
    .B(_1274_),
    .Y(_1276_));
 sg13g2_a21oi_1 _5290_ (.A1(_1226_),
    .A2(_1241_),
    .Y(_1277_),
    .B1(_1240_));
 sg13g2_a21oi_2 _5291_ (.B1(_1238_),
    .Y(_1278_),
    .A2(_1236_),
    .A1(_1230_));
 sg13g2_o21ai_1 _5292_ (.B1(_1233_),
    .Y(_1279_),
    .A1(_0008_),
    .A2(_0834_));
 sg13g2_inv_1 _5293_ (.Y(_1280_),
    .A(_1279_));
 sg13g2_o21ai_1 _5294_ (.B1(_1235_),
    .Y(_1281_),
    .A1(_0803_),
    .A2(_0838_));
 sg13g2_nor2_1 _5295_ (.A(_0772_),
    .B(_0836_),
    .Y(_1282_));
 sg13g2_mux2_1 _5296_ (.A0(_0772_),
    .A1(_0866_),
    .S(_0836_),
    .X(_1283_));
 sg13g2_mux2_1 _5297_ (.A0(_0008_),
    .A1(_0841_),
    .S(_0894_),
    .X(_1284_));
 sg13g2_nand2_1 _5298_ (.Y(_1285_),
    .A(_0840_),
    .B(_1284_));
 sg13g2_nand2_1 _5299_ (.Y(_1286_),
    .A(_0840_),
    .B(_1285_));
 sg13g2_nor2_1 _5300_ (.A(_0806_),
    .B(_0841_),
    .Y(_1287_));
 sg13g2_o21ai_1 _5301_ (.B1(_1285_),
    .Y(_1288_),
    .A1(_0008_),
    .A2(_0894_));
 sg13g2_o21ai_1 _5302_ (.B1(_1286_),
    .Y(_1289_),
    .A1(_1287_),
    .A2(_1288_));
 sg13g2_xor2_1 _5303_ (.B(_1289_),
    .A(_1283_),
    .X(_1290_));
 sg13g2_nand2_1 _5304_ (.Y(_1291_),
    .A(_1281_),
    .B(_1290_));
 sg13g2_xnor2_1 _5305_ (.Y(_1292_),
    .A(_1281_),
    .B(_1290_));
 sg13g2_xnor2_1 _5306_ (.Y(_1293_),
    .A(_1280_),
    .B(_1292_));
 sg13g2_nor2_1 _5307_ (.A(_1278_),
    .B(_1293_),
    .Y(_1294_));
 sg13g2_xnor2_1 _5308_ (.Y(_1295_),
    .A(_1278_),
    .B(_1293_));
 sg13g2_nor2_1 _5309_ (.A(_1277_),
    .B(_1295_),
    .Y(_1296_));
 sg13g2_xor2_1 _5310_ (.B(_1295_),
    .A(_1277_),
    .X(_1297_));
 sg13g2_nand2_1 _5311_ (.Y(_1298_),
    .A(_0639_),
    .B(_1297_));
 sg13g2_xnor2_1 _5312_ (.Y(_1299_),
    .A(_0639_),
    .B(_1297_));
 sg13g2_a21oi_1 _5313_ (.A1(_1225_),
    .A2(_1243_),
    .Y(_1300_),
    .B1(_1244_));
 sg13g2_or2_1 _5314_ (.X(_1301_),
    .B(_1300_),
    .A(_1299_));
 sg13g2_a21oi_1 _5315_ (.A1(_1299_),
    .A2(_1300_),
    .Y(_1302_),
    .B1(net439));
 sg13g2_a22oi_1 _5316_ (.Y(_1303_),
    .B1(_1301_),
    .B2(_1302_),
    .A2(_1276_),
    .A1(_1275_));
 sg13g2_nor2_1 _5317_ (.A(_0007_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_xnor2_1 _5318_ (.Y(_1305_),
    .A(_0007_),
    .B(_1303_));
 sg13g2_nor2_1 _5319_ (.A(_1258_),
    .B(_1305_),
    .Y(_1306_));
 sg13g2_xor2_1 _5320_ (.B(_1305_),
    .A(_1258_),
    .X(_1307_));
 sg13g2_a21o_1 _5321_ (.A2(net392),
    .A1(_0920_),
    .B1(_0930_),
    .X(_1308_));
 sg13g2_nand3_1 _5322_ (.B(_0920_),
    .C(_1307_),
    .A(_2946_),
    .Y(_1309_));
 sg13g2_a21oi_1 _5323_ (.A1(_1308_),
    .A2(_1309_),
    .Y(_1310_),
    .B1(_2952_));
 sg13g2_nand3_1 _5324_ (.B(_1308_),
    .C(_1309_),
    .A(_2952_),
    .Y(_1311_));
 sg13g2_nand2b_2 _5325_ (.Y(_1312_),
    .B(_1311_),
    .A_N(_1310_));
 sg13g2_a21o_1 _5326_ (.A2(_1311_),
    .A1(_0920_),
    .B1(_1310_),
    .X(_1313_));
 sg13g2_nor2b_1 _5327_ (.A(_0945_),
    .B_N(net392),
    .Y(_1314_));
 sg13g2_xnor2_1 _5328_ (.Y(_1315_),
    .A(_0944_),
    .B(_1314_));
 sg13g2_xor2_1 _5329_ (.B(_1315_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ),
    .X(_1316_));
 sg13g2_xor2_1 _5330_ (.B(_1316_),
    .A(_1313_),
    .X(_1317_));
 sg13g2_nand2_1 _5331_ (.Y(_1318_),
    .A(net442),
    .B(_1317_));
 sg13g2_nor2_1 _5332_ (.A(_1170_),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_xnor2_1 _5333_ (.Y(_1320_),
    .A(_1170_),
    .B(_1318_));
 sg13g2_or2_1 _5334_ (.X(_1321_),
    .B(_1320_),
    .A(_1126_));
 sg13g2_nor2b_1 _5335_ (.A(_0018_),
    .B_N(_1315_),
    .Y(_1322_));
 sg13g2_a21o_1 _5336_ (.A2(_1316_),
    .A1(_1313_),
    .B1(_1322_),
    .X(_1323_));
 sg13g2_nand2_1 _5337_ (.Y(_1324_),
    .A(_0966_),
    .B(net392));
 sg13g2_xor2_1 _5338_ (.B(_1324_),
    .A(_0965_),
    .X(_1325_));
 sg13g2_xnor2_1 _5339_ (.Y(_1326_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[3] ),
    .B(_1325_));
 sg13g2_inv_1 _5340_ (.Y(_1327_),
    .A(_1326_));
 sg13g2_xnor2_1 _5341_ (.Y(_1328_),
    .A(_1323_),
    .B(_1327_));
 sg13g2_nor2_2 _5342_ (.A(_0936_),
    .B(net440),
    .Y(_1329_));
 sg13g2_xor2_1 _5343_ (.B(_1255_),
    .A(_1254_),
    .X(_1330_));
 sg13g2_xnor2_1 _5344_ (.Y(_1331_),
    .A(_1329_),
    .B(_1330_));
 sg13g2_nor3_1 _5345_ (.A(_0941_),
    .B(_1328_),
    .C(_1331_),
    .Y(_1332_));
 sg13g2_o21ai_1 _5346_ (.B1(_1331_),
    .Y(_1333_),
    .A1(_0941_),
    .A2(_1328_));
 sg13g2_nand2b_1 _5347_ (.Y(_1334_),
    .B(_1333_),
    .A_N(_1332_));
 sg13g2_nand3b_1 _5348_ (.B(_1333_),
    .C(_1319_),
    .Y(_1335_),
    .A_N(_1332_));
 sg13g2_xor2_1 _5349_ (.B(_1334_),
    .A(_1319_),
    .X(_1336_));
 sg13g2_or2_1 _5350_ (.X(_1337_),
    .B(_1336_),
    .A(_1321_));
 sg13g2_nor2_2 _5351_ (.A(net461),
    .B(net437),
    .Y(_1338_));
 sg13g2_nand2_2 _5352_ (.Y(_1339_),
    .A(net473),
    .B(net439));
 sg13g2_a21o_1 _5353_ (.A2(_1330_),
    .A1(_1329_),
    .B1(_1332_),
    .X(_1340_));
 sg13g2_a22oi_1 _5354_ (.Y(_1341_),
    .B1(_1327_),
    .B2(_1323_),
    .A2(_1325_),
    .A1(_2953_));
 sg13g2_nand2_1 _5355_ (.Y(_1342_),
    .A(_1010_),
    .B(net392));
 sg13g2_xor2_1 _5356_ (.B(_1342_),
    .A(_1009_),
    .X(_1343_));
 sg13g2_xnor2_1 _5357_ (.Y(_1344_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[4] ),
    .B(_1343_));
 sg13g2_xor2_1 _5358_ (.B(_1344_),
    .A(_1341_),
    .X(_1345_));
 sg13g2_xnor2_1 _5359_ (.Y(_1346_),
    .A(_0920_),
    .B(_1312_));
 sg13g2_nand2_1 _5360_ (.Y(_1347_),
    .A(_1329_),
    .B(_1346_));
 sg13g2_xnor2_1 _5361_ (.Y(_1348_),
    .A(_1256_),
    .B(_1257_));
 sg13g2_xor2_1 _5362_ (.B(_1348_),
    .A(_1347_),
    .X(_1349_));
 sg13g2_nand3_1 _5363_ (.B(_1345_),
    .C(_1349_),
    .A(net441),
    .Y(_1350_));
 sg13g2_a21o_1 _5364_ (.A2(_1345_),
    .A1(net441),
    .B1(_1349_),
    .X(_1351_));
 sg13g2_and3_1 _5365_ (.X(_1352_),
    .A(_1340_),
    .B(_1350_),
    .C(_1351_));
 sg13g2_a21oi_1 _5366_ (.A1(_1350_),
    .A2(_1351_),
    .Y(_1353_),
    .B1(_1340_));
 sg13g2_nor2_1 _5367_ (.A(_1352_),
    .B(_1353_),
    .Y(_1354_));
 sg13g2_xnor2_1 _5368_ (.Y(_1355_),
    .A(_1339_),
    .B(_1354_));
 sg13g2_nor2b_1 _5369_ (.A(_1335_),
    .B_N(_1355_),
    .Y(_1356_));
 sg13g2_xor2_1 _5370_ (.B(_1355_),
    .A(_1335_),
    .X(_1357_));
 sg13g2_nor2_1 _5371_ (.A(_1337_),
    .B(_1357_),
    .Y(_1358_));
 sg13g2_xor2_1 _5372_ (.B(_1320_),
    .A(_1126_),
    .X(_1359_));
 sg13g2_xnor2_1 _5373_ (.Y(_1360_),
    .A(_0987_),
    .B(_1125_));
 sg13g2_xor2_1 _5374_ (.B(_1079_),
    .A(\main.demo._q_speed[0] ),
    .X(_1361_));
 sg13g2_nor2_1 _5375_ (.A(_0941_),
    .B(_1361_),
    .Y(_1362_));
 sg13g2_nor2b_1 _5376_ (.A(_1360_),
    .B_N(_1362_),
    .Y(_1363_));
 sg13g2_nand2_1 _5377_ (.Y(_1364_),
    .A(_1359_),
    .B(_1363_));
 sg13g2_nor2_1 _5378_ (.A(_1336_),
    .B(_1364_),
    .Y(_1365_));
 sg13g2_nand2_1 _5379_ (.Y(_1366_),
    .A(_1337_),
    .B(_1357_));
 sg13g2_xnor2_1 _5380_ (.Y(_1367_),
    .A(_1337_),
    .B(_1357_));
 sg13g2_a21o_1 _5381_ (.A2(_1366_),
    .A1(_1365_),
    .B1(_1358_),
    .X(_1368_));
 sg13g2_nor3_2 _5382_ (.A(net460),
    .B(net437),
    .C(_1312_),
    .Y(_1369_));
 sg13g2_a21oi_1 _5383_ (.A1(_1338_),
    .A2(_1354_),
    .Y(_1370_),
    .B1(_1352_));
 sg13g2_o21ai_1 _5384_ (.B1(_1350_),
    .Y(_1371_),
    .A1(_1347_),
    .A2(_1348_));
 sg13g2_nand3_1 _5385_ (.B(_1317_),
    .C(_1329_),
    .A(_1307_),
    .Y(_1372_));
 sg13g2_a21o_1 _5386_ (.A2(_1329_),
    .A1(_1317_),
    .B1(net392),
    .X(_1373_));
 sg13g2_nand2_1 _5387_ (.Y(_1374_),
    .A(_1372_),
    .B(_1373_));
 sg13g2_xnor2_1 _5388_ (.Y(_1375_),
    .A(_0960_),
    .B(_1374_));
 sg13g2_nand2_1 _5389_ (.Y(_1376_),
    .A(_1371_),
    .B(_1375_));
 sg13g2_xnor2_1 _5390_ (.Y(_1377_),
    .A(_1371_),
    .B(_1375_));
 sg13g2_xnor2_1 _5391_ (.Y(_1378_),
    .A(_1016_),
    .B(_1377_));
 sg13g2_nor2_1 _5392_ (.A(_1370_),
    .B(_1378_),
    .Y(_1379_));
 sg13g2_xor2_1 _5393_ (.B(_1378_),
    .A(_1370_),
    .X(_1380_));
 sg13g2_xor2_1 _5394_ (.B(_1380_),
    .A(_1369_),
    .X(_1381_));
 sg13g2_and2_1 _5395_ (.A(_1356_),
    .B(_1381_),
    .X(_1382_));
 sg13g2_xor2_1 _5396_ (.B(_1381_),
    .A(_1356_),
    .X(_1383_));
 sg13g2_xnor2_1 _5397_ (.Y(_1384_),
    .A(_1368_),
    .B(_1383_));
 sg13g2_nand2b_1 _5398_ (.Y(_1385_),
    .B(_1343_),
    .A_N(_0016_));
 sg13g2_o21ai_1 _5399_ (.B1(_1385_),
    .Y(_1386_),
    .A1(_1341_),
    .A2(_1344_));
 sg13g2_nand2_2 _5400_ (.Y(_1387_),
    .A(net503),
    .B(net444));
 sg13g2_nand2b_1 _5401_ (.Y(_1388_),
    .B(_1009_),
    .A_N(_1010_));
 sg13g2_nand2_1 _5402_ (.Y(_1389_),
    .A(net392),
    .B(_1388_));
 sg13g2_xnor2_1 _5403_ (.Y(_1390_),
    .A(_1387_),
    .B(_1389_));
 sg13g2_xnor2_1 _5404_ (.Y(_1391_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[5] ),
    .B(_1390_));
 sg13g2_xor2_1 _5405_ (.B(_1391_),
    .A(_1386_),
    .X(_1392_));
 sg13g2_nor2_1 _5406_ (.A(net443),
    .B(_1392_),
    .Y(_1393_));
 sg13g2_xnor2_1 _5407_ (.Y(_1394_),
    .A(_1384_),
    .B(_1393_));
 sg13g2_nand2_1 _5408_ (.Y(_1395_),
    .A(net461),
    .B(_1032_));
 sg13g2_nor2_2 _5409_ (.A(_1394_),
    .B(_1395_),
    .Y(_1396_));
 sg13g2_nor2_1 _5410_ (.A(net443),
    .B(_1346_),
    .Y(_1397_));
 sg13g2_xnor2_1 _5411_ (.Y(_1398_),
    .A(_1360_),
    .B(_1362_));
 sg13g2_xnor2_1 _5412_ (.Y(_1399_),
    .A(_1397_),
    .B(_1398_));
 sg13g2_xnor2_1 _5413_ (.Y(_1400_),
    .A(_1359_),
    .B(_1363_));
 sg13g2_nor2_1 _5414_ (.A(net443),
    .B(_1317_),
    .Y(_1401_));
 sg13g2_xnor2_1 _5415_ (.Y(_1402_),
    .A(_1400_),
    .B(_1401_));
 sg13g2_nor2_1 _5416_ (.A(net434),
    .B(_1402_),
    .Y(_1403_));
 sg13g2_a21o_1 _5417_ (.A2(_1399_),
    .A1(net434),
    .B1(_1403_),
    .X(_1404_));
 sg13g2_a21oi_1 _5418_ (.A1(_0987_),
    .A2(_0988_),
    .Y(_1405_),
    .B1(_0995_));
 sg13g2_xnor2_1 _5419_ (.Y(_1406_),
    .A(_0986_),
    .B(_1405_));
 sg13g2_o21ai_1 _5420_ (.B1(_1026_),
    .Y(_1407_),
    .A1(_1002_),
    .A2(_1027_));
 sg13g2_nand2_1 _5421_ (.Y(_1408_),
    .A(_1021_),
    .B(_1023_));
 sg13g2_nand2_2 _5422_ (.Y(_1409_),
    .A(_0960_),
    .B(_1317_));
 sg13g2_nand2b_1 _5423_ (.Y(_1410_),
    .B(_1019_),
    .A_N(_1017_));
 sg13g2_nand2_1 _5424_ (.Y(_1411_),
    .A(_0935_),
    .B(_0973_));
 sg13g2_nor2_1 _5425_ (.A(_0021_),
    .B(_1390_),
    .Y(_1412_));
 sg13g2_a21oi_1 _5426_ (.A1(_1386_),
    .A2(_1391_),
    .Y(_1413_),
    .B1(_1412_));
 sg13g2_inv_1 _5427_ (.Y(_1414_),
    .A(_1413_));
 sg13g2_nand2_1 _5428_ (.Y(_1415_),
    .A(\main.demo._q_speed[8] ),
    .B(net444));
 sg13g2_nand3_1 _5429_ (.B(net444),
    .C(net392),
    .A(net503),
    .Y(_1416_));
 sg13g2_nand2_1 _5430_ (.Y(_1417_),
    .A(_1389_),
    .B(_1416_));
 sg13g2_xnor2_1 _5431_ (.Y(_1418_),
    .A(_1415_),
    .B(_1417_));
 sg13g2_xor2_1 _5432_ (.B(_1418_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ),
    .X(_1419_));
 sg13g2_xnor2_1 _5433_ (.Y(_1420_),
    .A(_1413_),
    .B(_1419_));
 sg13g2_nand2_2 _5434_ (.Y(_1421_),
    .A(net442),
    .B(_1420_));
 sg13g2_nor2_1 _5435_ (.A(_0913_),
    .B(_0915_),
    .Y(_1422_));
 sg13g2_a21oi_1 _5436_ (.A1(_0702_),
    .A2(_0909_),
    .Y(_1423_),
    .B1(_0911_));
 sg13g2_nand2b_2 _5437_ (.Y(_1424_),
    .B(_0701_),
    .A_N(_0534_));
 sg13g2_a21oi_1 _5438_ (.A1(_0892_),
    .A2(_0906_),
    .Y(_1425_),
    .B1(_0908_));
 sg13g2_a21o_1 _5439_ (.A2(_0903_),
    .A1(_0867_),
    .B1(_0905_),
    .X(_1426_));
 sg13g2_a21oi_1 _5440_ (.A1(_0895_),
    .A2(_0900_),
    .Y(_1427_),
    .B1(_0899_));
 sg13g2_nand3_1 _5441_ (.B(_0517_),
    .C(_0896_),
    .A(net484),
    .Y(_1428_));
 sg13g2_a21o_1 _5442_ (.A2(_0517_),
    .A1(net484),
    .B1(_0896_),
    .X(_1429_));
 sg13g2_nand2_2 _5443_ (.Y(_1430_),
    .A(_1428_),
    .B(_1429_));
 sg13g2_xnor2_1 _5444_ (.Y(_1431_),
    .A(_0895_),
    .B(_1430_));
 sg13g2_nor2_1 _5445_ (.A(_0863_),
    .B(_1431_),
    .Y(_1432_));
 sg13g2_nand2b_1 _5446_ (.Y(_1433_),
    .B(_1432_),
    .A_N(_0901_));
 sg13g2_xnor2_1 _5447_ (.Y(_1434_),
    .A(_0903_),
    .B(_1431_));
 sg13g2_xor2_1 _5448_ (.B(_1434_),
    .A(_1427_),
    .X(_1435_));
 sg13g2_nand2_1 _5449_ (.Y(_1436_),
    .A(_1426_),
    .B(_1435_));
 sg13g2_xnor2_1 _5450_ (.Y(_1437_),
    .A(_1426_),
    .B(_1435_));
 sg13g2_xor2_1 _5451_ (.B(_1437_),
    .A(_1425_),
    .X(_1438_));
 sg13g2_nand2_1 _5452_ (.Y(_1439_),
    .A(_1424_),
    .B(_1438_));
 sg13g2_xnor2_1 _5453_ (.Y(_1440_),
    .A(_1424_),
    .B(_1438_));
 sg13g2_xor2_1 _5454_ (.B(_1440_),
    .A(_1423_),
    .X(_1441_));
 sg13g2_xnor2_1 _5455_ (.Y(_1442_),
    .A(_0019_),
    .B(_1441_));
 sg13g2_nor2b_1 _5456_ (.A(_1422_),
    .B_N(_1442_),
    .Y(_1443_));
 sg13g2_xnor2_1 _5457_ (.Y(_1444_),
    .A(_1422_),
    .B(_1442_));
 sg13g2_inv_1 _5458_ (.Y(_1445_),
    .A(_1444_));
 sg13g2_xnor2_1 _5459_ (.Y(_1446_),
    .A(_1421_),
    .B(_1444_));
 sg13g2_nand2b_1 _5460_ (.Y(_1447_),
    .B(_1446_),
    .A_N(_1411_));
 sg13g2_xnor2_1 _5461_ (.Y(_1448_),
    .A(_1411_),
    .B(_1446_));
 sg13g2_nand2_1 _5462_ (.Y(_1449_),
    .A(_1410_),
    .B(_1448_));
 sg13g2_xnor2_1 _5463_ (.Y(_1450_),
    .A(_1410_),
    .B(_1448_));
 sg13g2_xor2_1 _5464_ (.B(_1450_),
    .A(_1409_),
    .X(_1451_));
 sg13g2_xnor2_1 _5465_ (.Y(_1452_),
    .A(_1408_),
    .B(_1451_));
 sg13g2_nor2b_1 _5466_ (.A(_1452_),
    .B_N(_1407_),
    .Y(_1453_));
 sg13g2_xor2_1 _5467_ (.B(_1452_),
    .A(_1407_),
    .X(_1454_));
 sg13g2_a22oi_1 _5468_ (.Y(_1455_),
    .B1(_1013_),
    .B2(_1008_),
    .A2(_1012_),
    .A1(_2956_));
 sg13g2_nor2_1 _5469_ (.A(_0967_),
    .B(_1388_),
    .Y(_1456_));
 sg13g2_nor2_1 _5470_ (.A(_0917_),
    .B(_1456_),
    .Y(_1457_));
 sg13g2_xnor2_1 _5471_ (.Y(_1458_),
    .A(_1387_),
    .B(_1457_));
 sg13g2_xnor2_1 _5472_ (.Y(_1459_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ),
    .B(_1458_));
 sg13g2_a21oi_1 _5473_ (.A1(_1455_),
    .A2(_1459_),
    .Y(_1460_),
    .B1(net443));
 sg13g2_o21ai_1 _5474_ (.B1(_1460_),
    .Y(_1461_),
    .A1(_1455_),
    .A2(_1459_));
 sg13g2_xor2_1 _5475_ (.B(_1461_),
    .A(_1454_),
    .X(_1462_));
 sg13g2_nand2_1 _5476_ (.Y(_1463_),
    .A(net446),
    .B(_0973_));
 sg13g2_xnor2_1 _5477_ (.Y(_1464_),
    .A(_0999_),
    .B(_1001_));
 sg13g2_xnor2_1 _5478_ (.Y(_1465_),
    .A(_1463_),
    .B(_1464_));
 sg13g2_nand2_1 _5479_ (.Y(_1466_),
    .A(net445),
    .B(_0934_));
 sg13g2_xnor2_1 _5480_ (.Y(_1467_),
    .A(_1406_),
    .B(_1466_));
 sg13g2_xnor2_1 _5481_ (.Y(_1468_),
    .A(_0996_),
    .B(_0998_));
 sg13g2_nand2_1 _5482_ (.Y(_1469_),
    .A(net445),
    .B(_0952_));
 sg13g2_xnor2_1 _5483_ (.Y(_1470_),
    .A(_1468_),
    .B(_1469_));
 sg13g2_a22oi_1 _5484_ (.Y(_1471_),
    .B1(_1470_),
    .B2(\main.demo._q_th[3] ),
    .A2(_1467_),
    .A1(\main.demo._q_th[2] ));
 sg13g2_nor2_1 _5485_ (.A(\main.demo._q_th[3] ),
    .B(_1470_),
    .Y(_1472_));
 sg13g2_nor2_1 _5486_ (.A(_1471_),
    .B(_1472_),
    .Y(_1473_));
 sg13g2_or2_1 _5487_ (.X(_1474_),
    .B(_1473_),
    .A(_1465_));
 sg13g2_o21ai_1 _5488_ (.B1(_1032_),
    .Y(_1475_),
    .A1(\main.demo._q_th[5] ),
    .A2(_1474_));
 sg13g2_nand2_1 _5489_ (.Y(_1476_),
    .A(\main.demo._q_th[5] ),
    .B(_1474_));
 sg13g2_xor2_1 _5490_ (.B(_1462_),
    .A(_0022_),
    .X(_1477_));
 sg13g2_and3_1 _5491_ (.X(_1478_),
    .A(_1475_),
    .B(_1476_),
    .C(_1477_));
 sg13g2_a21o_1 _5492_ (.A2(_1451_),
    .A1(_1408_),
    .B1(_1453_),
    .X(_1479_));
 sg13g2_nand2_1 _5493_ (.Y(_1480_),
    .A(_2955_),
    .B(_1458_));
 sg13g2_o21ai_1 _5494_ (.B1(_1480_),
    .Y(_1481_),
    .A1(_1455_),
    .A2(_1459_));
 sg13g2_xnor2_1 _5495_ (.Y(_1482_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ),
    .B(_1415_));
 sg13g2_a21oi_1 _5496_ (.A1(_1387_),
    .A2(_1456_),
    .Y(_1483_),
    .B1(_0917_));
 sg13g2_xnor2_1 _5497_ (.Y(_1484_),
    .A(_1482_),
    .B(_1483_));
 sg13g2_xnor2_1 _5498_ (.Y(_1485_),
    .A(_1481_),
    .B(_1484_));
 sg13g2_nand2_1 _5499_ (.Y(_1486_),
    .A(net445),
    .B(_1485_));
 sg13g2_o21ai_1 _5500_ (.B1(_1449_),
    .Y(_1487_),
    .A1(_1409_),
    .A2(_1450_));
 sg13g2_nand2_1 _5501_ (.Y(_1488_),
    .A(net441),
    .B(_1485_));
 sg13g2_nor2_1 _5502_ (.A(_0936_),
    .B(_1015_),
    .Y(_1489_));
 sg13g2_a21o_1 _5503_ (.A2(_1441_),
    .A1(_2954_),
    .B1(_1443_),
    .X(_1490_));
 sg13g2_o21ai_1 _5504_ (.B1(_1439_),
    .Y(_1491_),
    .A1(_1423_),
    .A2(_1440_));
 sg13g2_o21ai_1 _5505_ (.B1(_1436_),
    .Y(_1492_),
    .A1(_1425_),
    .A2(_1437_));
 sg13g2_o21ai_1 _5506_ (.B1(_1433_),
    .Y(_1493_),
    .A1(_1427_),
    .A2(_1434_));
 sg13g2_xor2_1 _5507_ (.B(_0550_),
    .A(\main.demo._q_speed[7] ),
    .X(_1494_));
 sg13g2_xnor2_1 _5508_ (.Y(_1495_),
    .A(_1432_),
    .B(_1494_));
 sg13g2_xor2_1 _5509_ (.B(net488),
    .A(net485),
    .X(_1496_));
 sg13g2_xnor2_1 _5510_ (.Y(_1497_),
    .A(_0009_),
    .B(_1496_));
 sg13g2_nand2_1 _5511_ (.Y(_1498_),
    .A(_0517_),
    .B(_1497_));
 sg13g2_o21ai_1 _5512_ (.B1(_1428_),
    .Y(_1499_),
    .A1(_0894_),
    .A2(_1430_));
 sg13g2_xnor2_1 _5513_ (.Y(_1500_),
    .A(_1498_),
    .B(_1499_));
 sg13g2_xnor2_1 _5514_ (.Y(_1501_),
    .A(_1495_),
    .B(_1500_));
 sg13g2_xnor2_1 _5515_ (.Y(_1502_),
    .A(_1493_),
    .B(_1501_));
 sg13g2_xnor2_1 _5516_ (.Y(_1503_),
    .A(_1492_),
    .B(_1502_));
 sg13g2_xnor2_1 _5517_ (.Y(_1504_),
    .A(_1491_),
    .B(_1503_));
 sg13g2_xnor2_1 _5518_ (.Y(_1505_),
    .A(_1490_),
    .B(_1504_));
 sg13g2_xnor2_1 _5519_ (.Y(_1506_),
    .A(_1489_),
    .B(_1505_));
 sg13g2_xnor2_1 _5520_ (.Y(_1507_),
    .A(_1488_),
    .B(_1506_));
 sg13g2_o21ai_1 _5521_ (.B1(_1447_),
    .Y(_1508_),
    .A1(_1421_),
    .A2(_1445_));
 sg13g2_a21oi_1 _5522_ (.A1(_0952_),
    .A2(_0960_),
    .Y(_1509_),
    .B1(_1508_));
 sg13g2_xnor2_1 _5523_ (.Y(_1510_),
    .A(_1507_),
    .B(_1509_));
 sg13g2_xnor2_1 _5524_ (.Y(_1511_),
    .A(_1487_),
    .B(_1510_));
 sg13g2_xnor2_1 _5525_ (.Y(_1512_),
    .A(_1486_),
    .B(_1511_));
 sg13g2_xor2_1 _5526_ (.B(_1512_),
    .A(_1479_),
    .X(_1513_));
 sg13g2_nand2_1 _5527_ (.Y(_1514_),
    .A(_2909_),
    .B(_1462_));
 sg13g2_o21ai_1 _5528_ (.B1(_1514_),
    .Y(_1515_),
    .A1(\main.demo._q_th[7] ),
    .A2(_1513_));
 sg13g2_a21oi_1 _5529_ (.A1(\main.demo._q_th[7] ),
    .A2(_1513_),
    .Y(_1516_),
    .B1(net461));
 sg13g2_o21ai_1 _5530_ (.B1(_1516_),
    .Y(_1517_),
    .A1(_1478_),
    .A2(_1515_));
 sg13g2_xnor2_1 _5531_ (.Y(_1518_),
    .A(_0992_),
    .B(_0994_));
 sg13g2_o21ai_1 _5532_ (.B1(net445),
    .Y(_1519_),
    .A1(_0921_),
    .A2(_0927_));
 sg13g2_a21oi_1 _5533_ (.A1(_0921_),
    .A2(_0927_),
    .Y(_1520_),
    .B1(_1519_));
 sg13g2_xnor2_1 _5534_ (.Y(_1521_),
    .A(_1518_),
    .B(_1520_));
 sg13g2_nand2b_1 _5535_ (.Y(_1522_),
    .B(net460),
    .A_N(_1521_));
 sg13g2_o21ai_1 _5536_ (.B1(_1522_),
    .Y(_1523_),
    .A1(net460),
    .A2(_1406_));
 sg13g2_a21oi_1 _5537_ (.A1(_1368_),
    .A2(_1383_),
    .Y(_1524_),
    .B1(_1382_));
 sg13g2_a21oi_1 _5538_ (.A1(_1369_),
    .A2(_1380_),
    .Y(_1525_),
    .B1(_1379_));
 sg13g2_nand2_1 _5539_ (.Y(_1526_),
    .A(_1317_),
    .B(_1338_));
 sg13g2_o21ai_1 _5540_ (.B1(_1376_),
    .Y(_1527_),
    .A1(_1016_),
    .A2(_1377_));
 sg13g2_o21ai_1 _5541_ (.B1(_1372_),
    .Y(_1528_),
    .A1(_0961_),
    .A2(_1374_));
 sg13g2_nor2b_1 _5542_ (.A(_1328_),
    .B_N(_1329_),
    .Y(_1529_));
 sg13g2_nor2_1 _5543_ (.A(_1304_),
    .B(_1306_),
    .Y(_1530_));
 sg13g2_nor2b_1 _5544_ (.A(_1272_),
    .B_N(_1275_),
    .Y(_1531_));
 sg13g2_a21oi_1 _5545_ (.A1(_0811_),
    .A2(_1266_),
    .Y(_1532_),
    .B1(_1265_));
 sg13g2_o21ai_1 _5546_ (.B1(_1262_),
    .Y(_1533_),
    .A1(_0845_),
    .A2(_1263_));
 sg13g2_or2_1 _5547_ (.X(_1534_),
    .B(_0863_),
    .A(_0842_));
 sg13g2_nand2_1 _5548_ (.Y(_1535_),
    .A(_0862_),
    .B(_0867_));
 sg13g2_xnor2_1 _5549_ (.Y(_1536_),
    .A(_0862_),
    .B(_0867_));
 sg13g2_xor2_1 _5550_ (.B(_1536_),
    .A(_1534_),
    .X(_1537_));
 sg13g2_and2_1 _5551_ (.A(_1533_),
    .B(_1537_),
    .X(_1538_));
 sg13g2_xor2_1 _5552_ (.B(_1537_),
    .A(_1533_),
    .X(_1539_));
 sg13g2_xnor2_1 _5553_ (.Y(_1540_),
    .A(_0842_),
    .B(_1539_));
 sg13g2_xnor2_1 _5554_ (.Y(_1541_),
    .A(_1532_),
    .B(_1540_));
 sg13g2_nand3_1 _5555_ (.B(_1270_),
    .C(_1541_),
    .A(_1268_),
    .Y(_1542_));
 sg13g2_a21o_1 _5556_ (.A2(_1270_),
    .A1(_1268_),
    .B1(_1541_),
    .X(_1543_));
 sg13g2_and2_1 _5557_ (.A(_1542_),
    .B(_1543_),
    .X(_1544_));
 sg13g2_xnor2_1 _5558_ (.Y(_1545_),
    .A(_0639_),
    .B(_1544_));
 sg13g2_nor2_1 _5559_ (.A(_1531_),
    .B(_1545_),
    .Y(_1546_));
 sg13g2_a21oi_1 _5560_ (.A1(_1531_),
    .A2(_1545_),
    .Y(_1547_),
    .B1(net437));
 sg13g2_nand2b_1 _5561_ (.Y(_1548_),
    .B(_1547_),
    .A_N(_1546_));
 sg13g2_nand2_1 _5562_ (.Y(_1549_),
    .A(_1298_),
    .B(_1301_));
 sg13g2_or2_1 _5563_ (.X(_1550_),
    .B(_1296_),
    .A(_1294_));
 sg13g2_o21ai_1 _5564_ (.B1(_1291_),
    .Y(_1551_),
    .A1(_1280_),
    .A2(_1292_));
 sg13g2_a21oi_1 _5565_ (.A1(_1283_),
    .A2(_1289_),
    .Y(_1552_),
    .B1(_1282_));
 sg13g2_xor2_1 _5566_ (.B(_0900_),
    .A(_0865_),
    .X(_1553_));
 sg13g2_xor2_1 _5567_ (.B(_1284_),
    .A(_0840_),
    .X(_1554_));
 sg13g2_xnor2_1 _5568_ (.Y(_1555_),
    .A(_1553_),
    .B(_1554_));
 sg13g2_nor2_1 _5569_ (.A(_1552_),
    .B(_1555_),
    .Y(_1556_));
 sg13g2_xor2_1 _5570_ (.B(_1555_),
    .A(_1552_),
    .X(_1557_));
 sg13g2_xnor2_1 _5571_ (.Y(_1558_),
    .A(_1288_),
    .B(_1557_));
 sg13g2_nor2b_1 _5572_ (.A(_1558_),
    .B_N(_1551_),
    .Y(_1559_));
 sg13g2_nand2b_1 _5573_ (.Y(_1560_),
    .B(_1558_),
    .A_N(_1551_));
 sg13g2_nor2b_1 _5574_ (.A(_1559_),
    .B_N(_1560_),
    .Y(_1561_));
 sg13g2_xnor2_1 _5575_ (.Y(_1562_),
    .A(_1550_),
    .B(_1561_));
 sg13g2_inv_1 _5576_ (.Y(_1563_),
    .A(_1562_));
 sg13g2_xnor2_1 _5577_ (.Y(_1564_),
    .A(_0702_),
    .B(_1562_));
 sg13g2_and2_1 _5578_ (.A(_1549_),
    .B(_1564_),
    .X(_1565_));
 sg13g2_o21ai_1 _5579_ (.B1(net436),
    .Y(_1566_),
    .A1(_1549_),
    .A2(_1564_));
 sg13g2_o21ai_1 _5580_ (.B1(_1548_),
    .Y(_1567_),
    .A1(_1565_),
    .A2(_1566_));
 sg13g2_nand2_1 _5581_ (.Y(_1568_),
    .A(_2954_),
    .B(_1567_));
 sg13g2_xnor2_1 _5582_ (.Y(_1569_),
    .A(_2954_),
    .B(_1567_));
 sg13g2_xor2_1 _5583_ (.B(_1569_),
    .A(_1530_),
    .X(_1570_));
 sg13g2_nand2_1 _5584_ (.Y(_1571_),
    .A(_1529_),
    .B(_1570_));
 sg13g2_xnor2_1 _5585_ (.Y(_1572_),
    .A(_1529_),
    .B(_1570_));
 sg13g2_xnor2_1 _5586_ (.Y(_1573_),
    .A(_1004_),
    .B(_1572_));
 sg13g2_nand2_1 _5587_ (.Y(_1574_),
    .A(_1528_),
    .B(_1573_));
 sg13g2_xnor2_1 _5588_ (.Y(_1575_),
    .A(_1528_),
    .B(_1573_));
 sg13g2_xor2_1 _5589_ (.B(_1575_),
    .A(_1421_),
    .X(_1576_));
 sg13g2_xnor2_1 _5590_ (.Y(_1577_),
    .A(_1527_),
    .B(_1576_));
 sg13g2_nor2_1 _5591_ (.A(_1526_),
    .B(_1577_),
    .Y(_1578_));
 sg13g2_xor2_1 _5592_ (.B(_1577_),
    .A(_1526_),
    .X(_1579_));
 sg13g2_nand2b_1 _5593_ (.Y(_1580_),
    .B(_1579_),
    .A_N(_1525_));
 sg13g2_nor2b_1 _5594_ (.A(_1579_),
    .B_N(_1525_),
    .Y(_1581_));
 sg13g2_xnor2_1 _5595_ (.Y(_1582_),
    .A(_1525_),
    .B(_1579_));
 sg13g2_xnor2_1 _5596_ (.Y(_1583_),
    .A(_1524_),
    .B(_1582_));
 sg13g2_nor2_1 _5597_ (.A(net443),
    .B(_1420_),
    .Y(_1584_));
 sg13g2_xnor2_1 _5598_ (.Y(_1585_),
    .A(_1583_),
    .B(_1584_));
 sg13g2_nor2_1 _5599_ (.A(net443),
    .B(_1345_),
    .Y(_1586_));
 sg13g2_xnor2_1 _5600_ (.Y(_1587_),
    .A(_1365_),
    .B(_1367_));
 sg13g2_xnor2_1 _5601_ (.Y(_1588_),
    .A(_1586_),
    .B(_1587_));
 sg13g2_nand2_1 _5602_ (.Y(_1589_),
    .A(\main.demo._q_th[2] ),
    .B(_1402_));
 sg13g2_nand2_1 _5603_ (.Y(_1590_),
    .A(net445),
    .B(_1328_));
 sg13g2_nand2_1 _5604_ (.Y(_1591_),
    .A(_1321_),
    .B(_1364_));
 sg13g2_xor2_1 _5605_ (.B(_1591_),
    .A(_1336_),
    .X(_1592_));
 sg13g2_xnor2_1 _5606_ (.Y(_1593_),
    .A(_1590_),
    .B(_1592_));
 sg13g2_o21ai_1 _5607_ (.B1(_2910_),
    .Y(_1594_),
    .A1(_1589_),
    .A2(_1593_));
 sg13g2_nand2_1 _5608_ (.Y(_1595_),
    .A(_1589_),
    .B(_1593_));
 sg13g2_nand2_1 _5609_ (.Y(_1596_),
    .A(_1594_),
    .B(_1595_));
 sg13g2_nand2_1 _5610_ (.Y(_1597_),
    .A(_1588_),
    .B(_1596_));
 sg13g2_a21o_1 _5611_ (.A2(_1597_),
    .A1(\main.demo._q_th[5] ),
    .B1(_1394_),
    .X(_1598_));
 sg13g2_o21ai_1 _5612_ (.B1(_1598_),
    .Y(_1599_),
    .A1(\main.demo._q_th[5] ),
    .A2(_1597_));
 sg13g2_xor2_1 _5613_ (.B(_1585_),
    .A(_0022_),
    .X(_1600_));
 sg13g2_o21ai_1 _5614_ (.B1(_1580_),
    .Y(_1601_),
    .A1(_1524_),
    .A2(_1581_));
 sg13g2_a21oi_1 _5615_ (.A1(_1527_),
    .A2(_1576_),
    .Y(_1602_),
    .B1(_1578_));
 sg13g2_o21ai_1 _5616_ (.B1(_1574_),
    .Y(_1603_),
    .A1(_1421_),
    .A2(_1575_));
 sg13g2_o21ai_1 _5617_ (.B1(_1571_),
    .Y(_1604_),
    .A1(_1005_),
    .A2(_1572_));
 sg13g2_nand2_1 _5618_ (.Y(_1605_),
    .A(_1329_),
    .B(_1345_));
 sg13g2_nor2_1 _5619_ (.A(_1328_),
    .B(_1339_),
    .Y(_1606_));
 sg13g2_o21ai_1 _5620_ (.B1(_1568_),
    .Y(_1607_),
    .A1(_1530_),
    .A2(_1569_));
 sg13g2_a21o_1 _5621_ (.A2(_1544_),
    .A1(_0639_),
    .B1(_1546_),
    .X(_1608_));
 sg13g2_o21ai_1 _5622_ (.B1(_1543_),
    .Y(_1609_),
    .A1(_1532_),
    .A2(_1540_));
 sg13g2_a21oi_1 _5623_ (.A1(_0842_),
    .A2(_1539_),
    .Y(_1610_),
    .B1(_1538_));
 sg13g2_xnor2_1 _5624_ (.Y(_1611_),
    .A(_0702_),
    .B(_1534_));
 sg13g2_xnor2_1 _5625_ (.Y(_1612_),
    .A(_0893_),
    .B(_1611_));
 sg13g2_xnor2_1 _5626_ (.Y(_1613_),
    .A(_0901_),
    .B(_1612_));
 sg13g2_o21ai_1 _5627_ (.B1(_1535_),
    .Y(_1614_),
    .A1(_1534_),
    .A2(_1536_));
 sg13g2_xnor2_1 _5628_ (.Y(_1615_),
    .A(_0843_),
    .B(_1614_));
 sg13g2_xnor2_1 _5629_ (.Y(_1616_),
    .A(_1613_),
    .B(_1615_));
 sg13g2_xnor2_1 _5630_ (.Y(_1617_),
    .A(_1610_),
    .B(_1616_));
 sg13g2_xnor2_1 _5631_ (.Y(_1618_),
    .A(_1609_),
    .B(_1617_));
 sg13g2_or2_1 _5632_ (.X(_1619_),
    .B(_1618_),
    .A(_1608_));
 sg13g2_a21oi_1 _5633_ (.A1(_1608_),
    .A2(_1618_),
    .Y(_1620_),
    .B1(net436));
 sg13g2_a21oi_1 _5634_ (.A1(_0702_),
    .A2(_1563_),
    .Y(_1621_),
    .B1(_1565_));
 sg13g2_a21oi_1 _5635_ (.A1(_1550_),
    .A2(_1560_),
    .Y(_1622_),
    .B1(_1559_));
 sg13g2_a21oi_1 _5636_ (.A1(_1288_),
    .A2(_1557_),
    .Y(_1623_),
    .B1(_1556_));
 sg13g2_a21oi_1 _5637_ (.A1(_0865_),
    .A2(_0900_),
    .Y(_1624_),
    .B1(_1554_));
 sg13g2_o21ai_1 _5638_ (.B1(_1554_),
    .Y(_1625_),
    .A1(_0865_),
    .A2(_0900_));
 sg13g2_nand2b_1 _5639_ (.Y(_1626_),
    .B(_1625_),
    .A_N(_1624_));
 sg13g2_xnor2_1 _5640_ (.Y(_1627_),
    .A(_0899_),
    .B(_1430_));
 sg13g2_xnor2_1 _5641_ (.Y(_1628_),
    .A(_1288_),
    .B(_1424_));
 sg13g2_xnor2_1 _5642_ (.Y(_1629_),
    .A(_1627_),
    .B(_1628_));
 sg13g2_xnor2_1 _5643_ (.Y(_1630_),
    .A(_1626_),
    .B(_1629_));
 sg13g2_xnor2_1 _5644_ (.Y(_1631_),
    .A(_1623_),
    .B(_1630_));
 sg13g2_xor2_1 _5645_ (.B(_1631_),
    .A(_1622_),
    .X(_1632_));
 sg13g2_or2_1 _5646_ (.X(_1633_),
    .B(_1632_),
    .A(_1621_));
 sg13g2_a21oi_1 _5647_ (.A1(_1621_),
    .A2(_1632_),
    .Y(_1634_),
    .B1(net439));
 sg13g2_a22oi_1 _5648_ (.Y(_1635_),
    .B1(_1633_),
    .B2(_1634_),
    .A2(_1620_),
    .A1(_1619_));
 sg13g2_xnor2_1 _5649_ (.Y(_1636_),
    .A(net503),
    .B(_1635_));
 sg13g2_xnor2_1 _5650_ (.Y(_1637_),
    .A(_1607_),
    .B(_1636_));
 sg13g2_xnor2_1 _5651_ (.Y(_1638_),
    .A(_1409_),
    .B(_1637_));
 sg13g2_xnor2_1 _5652_ (.Y(_1639_),
    .A(_1606_),
    .B(_1638_));
 sg13g2_xnor2_1 _5653_ (.Y(_1640_),
    .A(_1605_),
    .B(_1639_));
 sg13g2_xnor2_1 _5654_ (.Y(_1641_),
    .A(_1604_),
    .B(_1640_));
 sg13g2_xnor2_1 _5655_ (.Y(_1642_),
    .A(_1603_),
    .B(_1641_));
 sg13g2_a22oi_1 _5656_ (.Y(_1643_),
    .B1(_1419_),
    .B2(_1414_),
    .A2(_1418_),
    .A1(_2955_));
 sg13g2_nand2_1 _5657_ (.Y(_1644_),
    .A(\main.demo._q_speed[9] ),
    .B(net446));
 sg13g2_xnor2_1 _5658_ (.Y(_1645_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ),
    .B(_1644_));
 sg13g2_nand3_1 _5659_ (.B(net444),
    .C(net392),
    .A(\main.demo._q_speed[8] ),
    .Y(_1646_));
 sg13g2_nor2b_1 _5660_ (.A(_1417_),
    .B_N(_1646_),
    .Y(_1647_));
 sg13g2_xnor2_1 _5661_ (.Y(_1648_),
    .A(_1645_),
    .B(_1647_));
 sg13g2_xnor2_1 _5662_ (.Y(_1649_),
    .A(_1643_),
    .B(_1648_));
 sg13g2_o21ai_1 _5663_ (.B1(_1488_),
    .Y(_1650_),
    .A1(net443),
    .A2(_1649_));
 sg13g2_xnor2_1 _5664_ (.Y(_1651_),
    .A(_1642_),
    .B(_1650_));
 sg13g2_xnor2_1 _5665_ (.Y(_1652_),
    .A(_1602_),
    .B(_1651_));
 sg13g2_xnor2_1 _5666_ (.Y(_1653_),
    .A(_1601_),
    .B(_1652_));
 sg13g2_nor2_1 _5667_ (.A(\main.demo._q_th[7] ),
    .B(_1653_),
    .Y(_1654_));
 sg13g2_a221oi_1 _5668_ (.B2(_1600_),
    .C1(_1654_),
    .B1(_1599_),
    .A1(_2909_),
    .Y(_1655_),
    .A2(_1585_));
 sg13g2_nand2_1 _5669_ (.Y(_1656_),
    .A(\main.demo._q_th[7] ),
    .B(_1653_));
 sg13g2_nand3b_1 _5670_ (.B(_1656_),
    .C(net473),
    .Y(_1657_),
    .A_N(_1655_));
 sg13g2_or3_1 _5671_ (.A(net460),
    .B(net437),
    .C(_1361_),
    .X(_1658_));
 sg13g2_o21ai_1 _5672_ (.B1(_1658_),
    .Y(_1659_),
    .A1(net434),
    .A2(_1399_));
 sg13g2_inv_1 _5673_ (.Y(_1660_),
    .A(_1659_));
 sg13g2_a22oi_1 _5674_ (.Y(_1661_),
    .B1(net386),
    .B2(_1660_),
    .A2(_1523_),
    .A1(_1517_));
 sg13g2_nor2_2 _5675_ (.A(net473),
    .B(_1032_),
    .Y(_1662_));
 sg13g2_nor3_1 _5676_ (.A(net474),
    .B(_1032_),
    .C(_1521_),
    .Y(_1663_));
 sg13g2_nand4_1 _5677_ (.B(_1523_),
    .C(net386),
    .A(_1517_),
    .Y(_1664_),
    .D(_1660_));
 sg13g2_nor2b_1 _5678_ (.A(_1661_),
    .B_N(_1664_),
    .Y(_1665_));
 sg13g2_a221oi_1 _5679_ (.B2(net473),
    .C1(_1663_),
    .B1(_1665_),
    .A1(_1396_),
    .Y(_1666_),
    .A2(_1404_));
 sg13g2_inv_1 _5680_ (.Y(\main.demo._t___block_68_frag[0] ),
    .A(_1666_));
 sg13g2_or2_1 _5681_ (.X(_1667_),
    .B(_1467_),
    .A(net473));
 sg13g2_o21ai_1 _5682_ (.B1(_1667_),
    .Y(_1668_),
    .A1(net460),
    .A2(_1468_));
 sg13g2_nand2_1 _5683_ (.Y(_1669_),
    .A(_1517_),
    .B(_1668_));
 sg13g2_nand2_1 _5684_ (.Y(_1670_),
    .A(_1404_),
    .B(_1657_));
 sg13g2_nand4_1 _5685_ (.B(net387),
    .C(net386),
    .A(_1404_),
    .Y(_1671_),
    .D(_1668_));
 sg13g2_a22oi_1 _5686_ (.Y(_1672_),
    .B1(_1668_),
    .B2(net387),
    .A2(net386),
    .A1(_1404_));
 sg13g2_xor2_1 _5687_ (.B(_1670_),
    .A(_1669_),
    .X(_1673_));
 sg13g2_xnor2_1 _5688_ (.Y(_1674_),
    .A(_1664_),
    .B(_1673_));
 sg13g2_nor2_1 _5689_ (.A(net434),
    .B(_1593_),
    .Y(_1675_));
 sg13g2_a21oi_2 _5690_ (.B1(_1675_),
    .Y(_1676_),
    .A2(_1402_),
    .A1(net434));
 sg13g2_nor3_1 _5691_ (.A(net473),
    .B(_1032_),
    .C(_1669_),
    .Y(_1677_));
 sg13g2_a221oi_1 _5692_ (.B2(_1396_),
    .C1(_1677_),
    .B1(_1676_),
    .A1(net473),
    .Y(_1678_),
    .A2(_1674_));
 sg13g2_inv_1 _5693_ (.Y(\main.demo._t___block_68_frag[1] ),
    .A(_1678_));
 sg13g2_nand2b_1 _5694_ (.Y(_1679_),
    .B(net459),
    .A_N(_1470_));
 sg13g2_o21ai_1 _5695_ (.B1(_1679_),
    .Y(_1680_),
    .A1(net459),
    .A2(_1464_));
 sg13g2_and2_1 _5696_ (.A(net387),
    .B(_1680_),
    .X(_1681_));
 sg13g2_nand2_1 _5697_ (.Y(_1682_),
    .A(net386),
    .B(_1676_));
 sg13g2_nand4_1 _5698_ (.B(net386),
    .C(_1676_),
    .A(net387),
    .Y(_1683_),
    .D(_1680_));
 sg13g2_xnor2_1 _5699_ (.Y(_1684_),
    .A(_1681_),
    .B(_1682_));
 sg13g2_o21ai_1 _5700_ (.B1(_1671_),
    .Y(_1685_),
    .A1(_1664_),
    .A2(_1672_));
 sg13g2_nand2_1 _5701_ (.Y(_1686_),
    .A(_1684_),
    .B(_1685_));
 sg13g2_xnor2_1 _5702_ (.Y(_1687_),
    .A(_1684_),
    .B(_1685_));
 sg13g2_mux2_1 _5703_ (.A0(_1588_),
    .A1(_1593_),
    .S(net434),
    .X(_1688_));
 sg13g2_a22oi_1 _5704_ (.Y(_1689_),
    .B1(_1688_),
    .B2(_1396_),
    .A2(_1681_),
    .A1(_1662_));
 sg13g2_o21ai_1 _5705_ (.B1(_1689_),
    .Y(\main.demo._t___block_68_frag[2] ),
    .A1(net460),
    .A2(_1687_));
 sg13g2_nor2_1 _5706_ (.A(net459),
    .B(_1030_),
    .Y(_1690_));
 sg13g2_a21oi_1 _5707_ (.A1(net459),
    .A2(_1465_),
    .Y(_1691_),
    .B1(_1690_));
 sg13g2_nand2_1 _5708_ (.Y(_1692_),
    .A(net387),
    .B(_1691_));
 sg13g2_nand2_1 _5709_ (.Y(_1693_),
    .A(net386),
    .B(_1688_));
 sg13g2_and2_1 _5710_ (.A(_1692_),
    .B(_1693_),
    .X(_1694_));
 sg13g2_xnor2_1 _5711_ (.Y(_1695_),
    .A(_1692_),
    .B(_1693_));
 sg13g2_nand2_1 _5712_ (.Y(_1696_),
    .A(_1683_),
    .B(_1686_));
 sg13g2_xor2_1 _5713_ (.B(_1696_),
    .A(_1695_),
    .X(_1697_));
 sg13g2_nor3_1 _5714_ (.A(net474),
    .B(_1032_),
    .C(_1465_),
    .Y(_1698_));
 sg13g2_nor2_1 _5715_ (.A(_1396_),
    .B(_1698_),
    .Y(_1699_));
 sg13g2_o21ai_1 _5716_ (.B1(_1699_),
    .Y(\main.demo._t___block_68_frag[3] ),
    .A1(net459),
    .A2(_1697_));
 sg13g2_o21ai_1 _5717_ (.B1(_1683_),
    .Y(_1700_),
    .A1(_1692_),
    .A2(_1693_));
 sg13g2_a21oi_1 _5718_ (.A1(_1684_),
    .A2(_1685_),
    .Y(_1701_),
    .B1(_1700_));
 sg13g2_nor2_1 _5719_ (.A(_1339_),
    .B(_1588_),
    .Y(_1702_));
 sg13g2_a21oi_1 _5720_ (.A1(_1339_),
    .A2(_1394_),
    .Y(_1703_),
    .B1(_1702_));
 sg13g2_nand2_1 _5721_ (.Y(_1704_),
    .A(net386),
    .B(_1703_));
 sg13g2_nor2_1 _5722_ (.A(net459),
    .B(_1454_),
    .Y(_1705_));
 sg13g2_o21ai_1 _5723_ (.B1(net387),
    .Y(_1706_),
    .A1(_1662_),
    .A2(_1705_));
 sg13g2_xnor2_1 _5724_ (.Y(_1707_),
    .A(_1704_),
    .B(_1706_));
 sg13g2_o21ai_1 _5725_ (.B1(_1707_),
    .Y(_1708_),
    .A1(_1694_),
    .A2(_1701_));
 sg13g2_or3_1 _5726_ (.A(_1694_),
    .B(_1701_),
    .C(_1707_),
    .X(_1709_));
 sg13g2_and2_1 _5727_ (.A(net473),
    .B(_1709_),
    .X(_1710_));
 sg13g2_nor2_1 _5728_ (.A(net434),
    .B(_1585_),
    .Y(_1711_));
 sg13g2_a21oi_1 _5729_ (.A1(net434),
    .A2(_1394_),
    .Y(_1712_),
    .B1(_1711_));
 sg13g2_a221oi_1 _5730_ (.B2(_1396_),
    .C1(_1662_),
    .B1(_1712_),
    .A1(_1708_),
    .Y(_1713_),
    .A2(_1710_));
 sg13g2_inv_1 _5731_ (.Y(\main.demo._t___block_68_frag[4] ),
    .A(_1713_));
 sg13g2_nor2_1 _5732_ (.A(net474),
    .B(_1462_),
    .Y(_1714_));
 sg13g2_a21oi_1 _5733_ (.A1(net474),
    .A2(_1513_),
    .Y(_1715_),
    .B1(_1714_));
 sg13g2_nand2_1 _5734_ (.Y(_1716_),
    .A(net387),
    .B(_1715_));
 sg13g2_nand3_1 _5735_ (.B(_1662_),
    .C(_1715_),
    .A(net387),
    .Y(_1717_));
 sg13g2_o21ai_1 _5736_ (.B1(_1709_),
    .Y(_1718_),
    .A1(_1704_),
    .A2(_1706_));
 sg13g2_nand2_1 _5737_ (.Y(_1719_),
    .A(_1657_),
    .B(_1712_));
 sg13g2_xnor2_1 _5738_ (.Y(_1720_),
    .A(_1716_),
    .B(_1719_));
 sg13g2_xor2_1 _5739_ (.B(_1720_),
    .A(_1718_),
    .X(_1721_));
 sg13g2_o21ai_1 _5740_ (.B1(_1717_),
    .Y(\main.demo._t___block_68_frag[5] ),
    .A1(net460),
    .A2(_1721_));
 sg13g2_nor3_2 _5741_ (.A(\main.demo.zic._q_squ_env[5] ),
    .B(\main.demo.zic._q_squ_env[4] ),
    .C(\main.demo.zic._q_squ_env[3] ),
    .Y(_1722_));
 sg13g2_nor2_2 _5742_ (.A(\main.demo.zic._q_qpos[12] ),
    .B(_1722_),
    .Y(_1723_));
 sg13g2_or2_2 _5743_ (.X(_1724_),
    .B(_1722_),
    .A(\main.demo.zic._q_qpos[12] ));
 sg13g2_nor2b_1 _5744_ (.A(\main._w_demo_video_vs ),
    .B_N(\main.demo._q_prev_vs ),
    .Y(_1725_));
 sg13g2_nand2b_2 _5745_ (.Y(_1726_),
    .B(\main.demo._q_prev_vs ),
    .A_N(\main._w_demo_video_vs ));
 sg13g2_nand2_1 _5746_ (.Y(_1727_),
    .A(\main.demo._q_frame[1] ),
    .B(\main.demo._q_frame[0] ));
 sg13g2_nor2_2 _5747_ (.A(_1726_),
    .B(_1727_),
    .Y(_1728_));
 sg13g2_nand2_2 _5748_ (.Y(_1729_),
    .A(net640),
    .B(_1728_));
 sg13g2_nor2_1 _5749_ (.A(_2932_),
    .B(_1729_),
    .Y(_1730_));
 sg13g2_nor3_2 _5750_ (.A(_2930_),
    .B(_2932_),
    .C(_1729_),
    .Y(_1731_));
 sg13g2_and2_1 _5751_ (.A(_3237_),
    .B(_1731_),
    .X(_1732_));
 sg13g2_and2_1 _5752_ (.A(\main.demo._q_frame[7] ),
    .B(_1732_),
    .X(_1733_));
 sg13g2_and2_2 _5753_ (.A(net651),
    .B(_1733_),
    .X(_1734_));
 sg13g2_and2_1 _5754_ (.A(\main.demo._q_frame[9] ),
    .B(_1734_),
    .X(_1735_));
 sg13g2_xor2_1 _5755_ (.B(_1734_),
    .A(net639),
    .X(_1736_));
 sg13g2_nor2_2 _5756_ (.A(\main.demo._q_go ),
    .B(_1736_),
    .Y(_1737_));
 sg13g2_xnor2_1 _5757_ (.Y(_1738_),
    .A(\main.demo.zic._q_tpos[11] ),
    .B(_1724_));
 sg13g2_nand2_1 _5758_ (.Y(_1739_),
    .A(net539),
    .B(net535));
 sg13g2_xor2_1 _5759_ (.B(\main.demo.zic._q_tpos[10] ),
    .A(\main.demo.zic._q_tpos[11] ),
    .X(_1740_));
 sg13g2_xnor2_1 _5760_ (.Y(_1741_),
    .A(\main.demo.zic._q_tpos[9] ),
    .B(_1740_));
 sg13g2_xnor2_1 _5761_ (.Y(_1742_),
    .A(\main.demo.zic._q_tpos[8] ),
    .B(_1740_));
 sg13g2_inv_1 _5762_ (.Y(_1743_),
    .A(_1742_));
 sg13g2_xnor2_1 _5763_ (.Y(_1744_),
    .A(\main.demo.zic._q_tpos[7] ),
    .B(_1740_));
 sg13g2_or2_1 _5764_ (.X(_1745_),
    .B(_1744_),
    .A(_1724_));
 sg13g2_o21ai_1 _5765_ (.B1(\main.demo.zic._q_squ_env[5] ),
    .Y(_1746_),
    .A1(\main.demo.zic._q_squ_env[4] ),
    .A2(\main.demo.zic._q_squ_env[3] ));
 sg13g2_a22oi_1 _5766_ (.Y(_1747_),
    .B1(_1723_),
    .B2(_1746_),
    .A2(_2957_),
    .A1(\main.demo.zic._q_qpos[12] ));
 sg13g2_xnor2_1 _5767_ (.Y(_1748_),
    .A(\main.demo.zic._q_tpos[6] ),
    .B(_1740_));
 sg13g2_nor2_1 _5768_ (.A(_1747_),
    .B(_1748_),
    .Y(_1749_));
 sg13g2_xnor2_1 _5769_ (.Y(_1750_),
    .A(\main.demo.zic._q_tpos[5] ),
    .B(_1740_));
 sg13g2_xor2_1 _5770_ (.B(\main.demo.zic._q_squ_env[3] ),
    .A(\main.demo.zic._q_squ_env[4] ),
    .X(_1751_));
 sg13g2_nand2_1 _5771_ (.Y(_1752_),
    .A(\main.demo.zic._q_qpos[12] ),
    .B(_0023_));
 sg13g2_o21ai_1 _5772_ (.B1(_1752_),
    .Y(_1753_),
    .A1(\main.demo.zic._q_qpos[12] ),
    .A2(_1751_));
 sg13g2_nor2_1 _5773_ (.A(_1750_),
    .B(_1753_),
    .Y(_1754_));
 sg13g2_nor2_1 _5774_ (.A(\main.demo.zic._q_tpos[4] ),
    .B(_1740_),
    .Y(_1755_));
 sg13g2_nand2_1 _5775_ (.Y(_1756_),
    .A(\main.demo.zic._q_tpos[4] ),
    .B(_1740_));
 sg13g2_nand2_1 _5776_ (.Y(_1757_),
    .A(\main.demo.zic._q_squ_env[3] ),
    .B(_1756_));
 sg13g2_xnor2_1 _5777_ (.Y(_1758_),
    .A(_1750_),
    .B(_1753_));
 sg13g2_nor3_1 _5778_ (.A(_1755_),
    .B(_1757_),
    .C(_1758_),
    .Y(_1759_));
 sg13g2_nor2_1 _5779_ (.A(_1754_),
    .B(_1759_),
    .Y(_1760_));
 sg13g2_xor2_1 _5780_ (.B(_1748_),
    .A(_1747_),
    .X(_1761_));
 sg13g2_nor2b_1 _5781_ (.A(_1760_),
    .B_N(_1761_),
    .Y(_1762_));
 sg13g2_xnor2_1 _5782_ (.Y(_1763_),
    .A(_1724_),
    .B(_1744_));
 sg13g2_inv_1 _5783_ (.Y(_1764_),
    .A(_1763_));
 sg13g2_o21ai_1 _5784_ (.B1(_1764_),
    .Y(_1765_),
    .A1(_1749_),
    .A2(_1762_));
 sg13g2_xnor2_1 _5785_ (.Y(_1766_),
    .A(_1724_),
    .B(_1742_));
 sg13g2_a21oi_1 _5786_ (.A1(_1745_),
    .A2(_1765_),
    .Y(_1767_),
    .B1(_1766_));
 sg13g2_a21oi_1 _5787_ (.A1(_1723_),
    .A2(_1743_),
    .Y(_1768_),
    .B1(_1767_));
 sg13g2_a21o_1 _5788_ (.A2(_1741_),
    .A1(_1724_),
    .B1(_1768_),
    .X(_1769_));
 sg13g2_o21ai_1 _5789_ (.B1(_1769_),
    .Y(_1770_),
    .A1(_1724_),
    .A2(_1741_));
 sg13g2_a21oi_1 _5790_ (.A1(_1738_),
    .A2(_1770_),
    .Y(_1771_),
    .B1(_1737_));
 sg13g2_o21ai_1 _5791_ (.B1(_1771_),
    .Y(_1772_),
    .A1(\main.demo.zic._q_tpos[11] ),
    .A2(_1723_));
 sg13g2_nor2_1 _5792_ (.A(net311),
    .B(_1772_),
    .Y(_1773_));
 sg13g2_nor2_1 _5793_ (.A(_1738_),
    .B(_1770_),
    .Y(_1774_));
 sg13g2_nor2b_1 _5794_ (.A(_1774_),
    .B_N(_1771_),
    .Y(_1775_));
 sg13g2_xnor2_1 _5795_ (.Y(_1776_),
    .A(_1724_),
    .B(_1741_));
 sg13g2_xnor2_1 _5796_ (.Y(_1777_),
    .A(_1768_),
    .B(_1776_));
 sg13g2_nand3_1 _5797_ (.B(_1765_),
    .C(_1766_),
    .A(_1745_),
    .Y(_1778_));
 sg13g2_nor2b_1 _5798_ (.A(_1767_),
    .B_N(_1778_),
    .Y(_1779_));
 sg13g2_or3_1 _5799_ (.A(_1749_),
    .B(_1762_),
    .C(_1764_),
    .X(_1780_));
 sg13g2_nand2_1 _5800_ (.Y(_1781_),
    .A(_1765_),
    .B(_1780_));
 sg13g2_o21ai_1 _5801_ (.B1(_1758_),
    .Y(_1782_),
    .A1(_1755_),
    .A2(_1757_));
 sg13g2_nor2_1 _5802_ (.A(\main.demo.zic._q_clock_count[0] ),
    .B(_1759_),
    .Y(_1783_));
 sg13g2_nand2_1 _5803_ (.Y(_1784_),
    .A(_1782_),
    .B(_1783_));
 sg13g2_xor2_1 _5804_ (.B(_1761_),
    .A(_1760_),
    .X(_1785_));
 sg13g2_nor2_1 _5805_ (.A(\main.demo.zic._q_clock_count[1] ),
    .B(_1784_),
    .Y(_1786_));
 sg13g2_a21oi_1 _5806_ (.A1(\main.demo.zic._q_clock_count[1] ),
    .A2(_1784_),
    .Y(_1787_),
    .B1(_1785_));
 sg13g2_nor2_1 _5807_ (.A(_1786_),
    .B(_1787_),
    .Y(_1788_));
 sg13g2_o21ai_1 _5808_ (.B1(_1781_),
    .Y(_1789_),
    .A1(\main.demo.zic._q_clock_count[2] ),
    .A2(_1788_));
 sg13g2_nand2_1 _5809_ (.Y(_1790_),
    .A(\main.demo.zic._q_clock_count[2] ),
    .B(_1788_));
 sg13g2_a22oi_1 _5810_ (.Y(_1791_),
    .B1(_1789_),
    .B2(_1790_),
    .A2(_1779_),
    .A1(_0027_));
 sg13g2_inv_1 _5811_ (.Y(_1792_),
    .A(_1791_));
 sg13g2_o21ai_1 _5812_ (.B1(_1792_),
    .Y(_1793_),
    .A1(_0027_),
    .A2(_1779_));
 sg13g2_o21ai_1 _5813_ (.B1(_1793_),
    .Y(_1794_),
    .A1(\main.demo.zic._q_clock_count[4] ),
    .A2(_1777_));
 sg13g2_a21oi_1 _5814_ (.A1(\main.demo.zic._q_clock_count[4] ),
    .A2(_1777_),
    .Y(_1795_),
    .B1(_1737_));
 sg13g2_and2_1 _5815_ (.A(_1794_),
    .B(_1795_),
    .X(_1796_));
 sg13g2_o21ai_1 _5816_ (.B1(_1796_),
    .Y(_1797_),
    .A1(_0026_),
    .A2(_1775_));
 sg13g2_a22oi_1 _5817_ (.Y(_1798_),
    .B1(_1775_),
    .B2(_0026_),
    .A2(_1772_),
    .A1(net311));
 sg13g2_a21oi_1 _5818_ (.A1(_1797_),
    .A2(_1798_),
    .Y(\main._w_demo_audio1 ),
    .B1(net312));
 sg13g2_o21ai_1 _5819_ (.B1(net453),
    .Y(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ),
    .A1(net297),
    .A2(net338));
 sg13g2_a21oi_1 _5820_ (.A1(net338),
    .A2(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .Y(\main.demo._t___pip_58_1_3___block_87_atten_h[1] ),
    .B1(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ));
 sg13g2_xnor2_1 _5821_ (.Y(_1799_),
    .A(_2970_),
    .B(_3029_));
 sg13g2_nor2_1 _5822_ (.A(_2997_),
    .B(net405),
    .Y(_1800_));
 sg13g2_xnor2_1 _5823_ (.Y(_1801_),
    .A(_3007_),
    .B(_1800_));
 sg13g2_nor2_1 _5824_ (.A(_1799_),
    .B(_1801_),
    .Y(_1802_));
 sg13g2_xor2_1 _5825_ (.B(_1801_),
    .A(_1799_),
    .X(_1803_));
 sg13g2_xnor2_1 _5826_ (.Y(_1804_),
    .A(_2998_),
    .B(_1803_));
 sg13g2_nor3_1 _5827_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .B(_3053_),
    .C(_3058_),
    .Y(_1805_));
 sg13g2_a21o_1 _5828_ (.A2(_3058_),
    .A1(_3053_),
    .B1(_1805_),
    .X(_1806_));
 sg13g2_xor2_1 _5829_ (.B(_1806_),
    .A(_0051_),
    .X(_1807_));
 sg13g2_or2_1 _5830_ (.X(_1808_),
    .B(_3071_),
    .A(_3060_));
 sg13g2_o21ai_1 _5831_ (.B1(_1807_),
    .Y(_1809_),
    .A1(net405),
    .A2(_1808_));
 sg13g2_a21oi_1 _5832_ (.A1(_1807_),
    .A2(_1808_),
    .Y(_1810_),
    .B1(net405));
 sg13g2_a21o_2 _5833_ (.A2(_1807_),
    .A1(net405),
    .B1(_1810_),
    .X(_1811_));
 sg13g2_o21ai_1 _5834_ (.B1(_3090_),
    .Y(_1812_),
    .A1(_0046_),
    .A2(_3077_));
 sg13g2_xnor2_1 _5835_ (.Y(_1813_),
    .A(_3091_),
    .B(_1812_));
 sg13g2_nand2b_1 _5836_ (.Y(_1814_),
    .B(_1813_),
    .A_N(_1811_));
 sg13g2_nor2b_1 _5837_ (.A(_1813_),
    .B_N(_1811_),
    .Y(_1815_));
 sg13g2_xnor2_1 _5838_ (.Y(_1816_),
    .A(_3088_),
    .B(_3089_));
 sg13g2_nor2_1 _5839_ (.A(_1811_),
    .B(_1816_),
    .Y(_1817_));
 sg13g2_xor2_1 _5840_ (.B(_1816_),
    .A(_1811_),
    .X(_1818_));
 sg13g2_xnor2_1 _5841_ (.Y(_1819_),
    .A(_3085_),
    .B(_3087_));
 sg13g2_inv_1 _5842_ (.Y(_1820_),
    .A(_1819_));
 sg13g2_xnor2_1 _5843_ (.Y(_1821_),
    .A(_1811_),
    .B(_1819_));
 sg13g2_o21ai_1 _5844_ (.B1(_1811_),
    .Y(_1822_),
    .A1(_1807_),
    .A2(_1808_));
 sg13g2_xnor2_1 _5845_ (.Y(_1823_),
    .A(_3082_),
    .B(_3084_));
 sg13g2_nand2_1 _5846_ (.Y(_1824_),
    .A(_1822_),
    .B(_1823_));
 sg13g2_a21oi_1 _5847_ (.A1(_3100_),
    .A2(_3122_),
    .Y(_1825_),
    .B1(_3099_));
 sg13g2_xnor2_1 _5848_ (.Y(_1826_),
    .A(_1822_),
    .B(_1823_));
 sg13g2_o21ai_1 _5849_ (.B1(_1824_),
    .Y(_1827_),
    .A1(_1825_),
    .A2(_1826_));
 sg13g2_nand2_1 _5850_ (.Y(_1828_),
    .A(_1821_),
    .B(_1827_));
 sg13g2_o21ai_1 _5851_ (.B1(_1828_),
    .Y(_1829_),
    .A1(_1811_),
    .A2(_1820_));
 sg13g2_a21oi_1 _5852_ (.A1(_1818_),
    .A2(_1829_),
    .Y(_1830_),
    .B1(_1817_));
 sg13g2_a21oi_1 _5853_ (.A1(_1814_),
    .A2(_1830_),
    .Y(_1831_),
    .B1(_1815_));
 sg13g2_xnor2_1 _5854_ (.Y(_1832_),
    .A(_1809_),
    .B(_1831_));
 sg13g2_nor2_1 _5855_ (.A(_3123_),
    .B(_1832_),
    .Y(_1833_));
 sg13g2_xor2_1 _5856_ (.B(_1826_),
    .A(_1825_),
    .X(_1834_));
 sg13g2_xnor2_1 _5857_ (.Y(_1835_),
    .A(_1833_),
    .B(_1834_));
 sg13g2_nand2_1 _5858_ (.Y(_1836_),
    .A(_1804_),
    .B(_1835_));
 sg13g2_xnor2_1 _5859_ (.Y(_1837_),
    .A(_1804_),
    .B(_1835_));
 sg13g2_xor2_1 _5860_ (.B(_1837_),
    .A(_3125_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[1] ));
 sg13g2_o21ai_1 _5861_ (.B1(_1836_),
    .Y(_1838_),
    .A1(_3125_),
    .A2(_1837_));
 sg13g2_a21oi_1 _5862_ (.A1(_2999_),
    .A2(_1803_),
    .Y(_1839_),
    .B1(_1802_));
 sg13g2_xor2_1 _5863_ (.B(_3031_),
    .A(_3030_),
    .X(_1840_));
 sg13g2_inv_1 _5864_ (.Y(_1841_),
    .A(_1840_));
 sg13g2_nand2_1 _5865_ (.Y(_1842_),
    .A(_2997_),
    .B(_3007_));
 sg13g2_nand2_1 _5866_ (.Y(_1843_),
    .A(_3096_),
    .B(_1842_));
 sg13g2_xor2_1 _5867_ (.B(_1843_),
    .A(_1823_),
    .X(_1844_));
 sg13g2_xnor2_1 _5868_ (.Y(_1845_),
    .A(_1840_),
    .B(_1844_));
 sg13g2_nor2b_1 _5869_ (.A(_1839_),
    .B_N(_1845_),
    .Y(_1846_));
 sg13g2_xnor2_1 _5870_ (.Y(_1847_),
    .A(_1839_),
    .B(_1845_));
 sg13g2_nor2_1 _5871_ (.A(_3124_),
    .B(_1834_),
    .Y(_1848_));
 sg13g2_nor2_1 _5872_ (.A(_1832_),
    .B(_1848_),
    .Y(_1849_));
 sg13g2_xor2_1 _5873_ (.B(_1827_),
    .A(_1821_),
    .X(_1850_));
 sg13g2_xnor2_1 _5874_ (.Y(_1851_),
    .A(_1849_),
    .B(_1850_));
 sg13g2_nand2_1 _5875_ (.Y(_1852_),
    .A(_1847_),
    .B(_1851_));
 sg13g2_xnor2_1 _5876_ (.Y(_1853_),
    .A(_1847_),
    .B(_1851_));
 sg13g2_nand2b_1 _5877_ (.Y(_1854_),
    .B(_1838_),
    .A_N(_1853_));
 sg13g2_xnor2_1 _5878_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[2] ),
    .A(_1838_),
    .B(_1853_));
 sg13g2_a21oi_1 _5879_ (.A1(_1841_),
    .A2(_1844_),
    .Y(_1855_),
    .B1(_1846_));
 sg13g2_xor2_1 _5880_ (.B(_3034_),
    .A(_3033_),
    .X(_1856_));
 sg13g2_nor2_1 _5881_ (.A(_1823_),
    .B(_1842_),
    .Y(_1857_));
 sg13g2_nor2_1 _5882_ (.A(net404),
    .B(_1857_),
    .Y(_1858_));
 sg13g2_xnor2_1 _5883_ (.Y(_1859_),
    .A(_1819_),
    .B(_1858_));
 sg13g2_inv_1 _5884_ (.Y(_1860_),
    .A(_1859_));
 sg13g2_xnor2_1 _5885_ (.Y(_1861_),
    .A(_1856_),
    .B(_1859_));
 sg13g2_nand2b_1 _5886_ (.Y(_1862_),
    .B(_1861_),
    .A_N(_1855_));
 sg13g2_xnor2_1 _5887_ (.Y(_1863_),
    .A(_1855_),
    .B(_1861_));
 sg13g2_nand2b_1 _5888_ (.Y(_1864_),
    .B(_1848_),
    .A_N(_1850_));
 sg13g2_nor2b_1 _5889_ (.A(_1832_),
    .B_N(_1864_),
    .Y(_1865_));
 sg13g2_xor2_1 _5890_ (.B(_1829_),
    .A(_1818_),
    .X(_1866_));
 sg13g2_xnor2_1 _5891_ (.Y(_1867_),
    .A(_1865_),
    .B(_1866_));
 sg13g2_xnor2_1 _5892_ (.Y(_1868_),
    .A(_1863_),
    .B(_1867_));
 sg13g2_a21oi_1 _5893_ (.A1(_1852_),
    .A2(_1854_),
    .Y(_1869_),
    .B1(_1868_));
 sg13g2_nand3_1 _5894_ (.B(_1854_),
    .C(_1868_),
    .A(_1852_),
    .Y(_1870_));
 sg13g2_nor2b_1 _5895_ (.A(_1869_),
    .B_N(_1870_),
    .Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[3] ));
 sg13g2_a21o_1 _5896_ (.A2(_1867_),
    .A1(_1863_),
    .B1(_1869_),
    .X(_1871_));
 sg13g2_o21ai_1 _5897_ (.B1(_1862_),
    .Y(_1872_),
    .A1(_1856_),
    .A2(_1860_));
 sg13g2_nand2_1 _5898_ (.Y(_1873_),
    .A(_1820_),
    .B(_1857_));
 sg13g2_nor2b_1 _5899_ (.A(net404),
    .B_N(_1873_),
    .Y(_1874_));
 sg13g2_xnor2_1 _5900_ (.Y(_1875_),
    .A(_1816_),
    .B(_1874_));
 sg13g2_nor2_1 _5901_ (.A(_3066_),
    .B(_1875_),
    .Y(_1876_));
 sg13g2_xor2_1 _5902_ (.B(_1875_),
    .A(_3066_),
    .X(_1877_));
 sg13g2_xnor2_1 _5903_ (.Y(_1878_),
    .A(_1872_),
    .B(_1877_));
 sg13g2_or2_1 _5904_ (.X(_1879_),
    .B(_1866_),
    .A(_1864_));
 sg13g2_nand2b_1 _5905_ (.Y(_1880_),
    .B(_1879_),
    .A_N(_1832_));
 sg13g2_xnor2_1 _5906_ (.Y(_1881_),
    .A(_1811_),
    .B(_1813_));
 sg13g2_xnor2_1 _5907_ (.Y(_1882_),
    .A(_1830_),
    .B(_1881_));
 sg13g2_xnor2_1 _5908_ (.Y(_1883_),
    .A(_1880_),
    .B(_1882_));
 sg13g2_nor2_1 _5909_ (.A(_1878_),
    .B(_1883_),
    .Y(_1884_));
 sg13g2_xor2_1 _5910_ (.B(_1883_),
    .A(_1878_),
    .X(_1885_));
 sg13g2_xor2_1 _5911_ (.B(_1885_),
    .A(_1871_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_a21oi_1 _5912_ (.A1(_1871_),
    .A2(_1885_),
    .Y(_1886_),
    .B1(_1884_));
 sg13g2_or3_2 _5913_ (.A(_1832_),
    .B(_1879_),
    .C(_1882_),
    .X(_1887_));
 sg13g2_a21oi_1 _5914_ (.A1(_1872_),
    .A2(_1877_),
    .Y(_1888_),
    .B1(_1876_));
 sg13g2_nand2b_1 _5915_ (.Y(_1889_),
    .B(_1816_),
    .A_N(_1873_));
 sg13g2_nand2_1 _5916_ (.Y(_1890_),
    .A(_3096_),
    .B(_1889_));
 sg13g2_xor2_1 _5917_ (.B(_1890_),
    .A(_1813_),
    .X(_1891_));
 sg13g2_nand2_1 _5918_ (.Y(_1892_),
    .A(_3065_),
    .B(_1891_));
 sg13g2_xnor2_1 _5919_ (.Y(_1893_),
    .A(_3065_),
    .B(_1891_));
 sg13g2_xor2_1 _5920_ (.B(_1893_),
    .A(_1888_),
    .X(_1894_));
 sg13g2_inv_1 _5921_ (.Y(_1895_),
    .A(_1894_));
 sg13g2_xnor2_1 _5922_ (.Y(_1896_),
    .A(_1887_),
    .B(_1894_));
 sg13g2_xnor2_1 _5923_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[5] ),
    .A(_1886_),
    .B(_1896_));
 sg13g2_a21oi_1 _5924_ (.A1(_1887_),
    .A2(_1895_),
    .Y(_1897_),
    .B1(_1886_));
 sg13g2_nor3_2 _5925_ (.A(net404),
    .B(_1813_),
    .C(_1889_),
    .Y(_1898_));
 sg13g2_xnor2_1 _5926_ (.Y(_1899_),
    .A(_3064_),
    .B(_1898_));
 sg13g2_o21ai_1 _5927_ (.B1(_1892_),
    .Y(_1900_),
    .A1(_1888_),
    .A2(_1893_));
 sg13g2_nor2b_1 _5928_ (.A(_1899_),
    .B_N(_1900_),
    .Y(_1901_));
 sg13g2_xor2_1 _5929_ (.B(_1900_),
    .A(_1899_),
    .X(_1902_));
 sg13g2_nor2_1 _5930_ (.A(net391),
    .B(_1902_),
    .Y(_1903_));
 sg13g2_xor2_1 _5931_ (.B(_1902_),
    .A(net391),
    .X(_1904_));
 sg13g2_xor2_1 _5932_ (.B(_1904_),
    .A(_1897_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_a21oi_1 _5933_ (.A1(_1897_),
    .A2(_1904_),
    .Y(_1905_),
    .B1(_1903_));
 sg13g2_nand2_1 _5934_ (.Y(_1906_),
    .A(_3069_),
    .B(_1898_));
 sg13g2_xnor2_1 _5935_ (.Y(_1907_),
    .A(_3069_),
    .B(_1898_));
 sg13g2_a21oi_1 _5936_ (.A1(_3064_),
    .A2(_1898_),
    .Y(_1908_),
    .B1(_1901_));
 sg13g2_xnor2_1 _5937_ (.Y(_1909_),
    .A(_1907_),
    .B(_1908_));
 sg13g2_nor2_1 _5938_ (.A(net391),
    .B(_1909_),
    .Y(_1910_));
 sg13g2_xor2_1 _5939_ (.B(_1909_),
    .A(net391),
    .X(_1911_));
 sg13g2_nor2b_1 _5940_ (.A(_1905_),
    .B_N(_1911_),
    .Y(_1912_));
 sg13g2_xnor2_1 _5941_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[7] ),
    .A(_1905_),
    .B(_1911_));
 sg13g2_nor2b_1 _5942_ (.A(_3063_),
    .B_N(_1898_),
    .Y(_1913_));
 sg13g2_xnor2_1 _5943_ (.Y(_1914_),
    .A(_3063_),
    .B(_1898_));
 sg13g2_o21ai_1 _5944_ (.B1(_1906_),
    .Y(_1915_),
    .A1(_1907_),
    .A2(_1908_));
 sg13g2_xor2_1 _5945_ (.B(_1915_),
    .A(_1914_),
    .X(_1916_));
 sg13g2_inv_1 _5946_ (.Y(_1917_),
    .A(_1916_));
 sg13g2_xnor2_1 _5947_ (.Y(_1918_),
    .A(net391),
    .B(_1916_));
 sg13g2_o21ai_1 _5948_ (.B1(_1918_),
    .Y(_1919_),
    .A1(_1910_),
    .A2(_1912_));
 sg13g2_or3_1 _5949_ (.A(_1910_),
    .B(_1912_),
    .C(_1918_),
    .X(_1920_));
 sg13g2_and2_1 _5950_ (.A(_1919_),
    .B(_1920_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[8] ));
 sg13g2_o21ai_1 _5951_ (.B1(_1919_),
    .Y(_1921_),
    .A1(net391),
    .A2(_1917_));
 sg13g2_a21oi_1 _5952_ (.A1(_1914_),
    .A2(_1915_),
    .Y(_1922_),
    .B1(_1913_));
 sg13g2_xor2_1 _5953_ (.B(_1898_),
    .A(_3060_),
    .X(_1923_));
 sg13g2_xnor2_1 _5954_ (.Y(_1924_),
    .A(_1922_),
    .B(_1923_));
 sg13g2_xor2_1 _5955_ (.B(_1924_),
    .A(net391),
    .X(_1925_));
 sg13g2_xnor2_1 _5956_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[9] ),
    .A(_1921_),
    .B(_1925_));
 sg13g2_nand3_1 _5957_ (.B(_1921_),
    .C(_1924_),
    .A(net391),
    .Y(_1926_));
 sg13g2_nor3_1 _5958_ (.A(_3061_),
    .B(_1898_),
    .C(_1922_),
    .Y(_1927_));
 sg13g2_xnor2_1 _5959_ (.Y(_1928_),
    .A(_1807_),
    .B(_1927_));
 sg13g2_xnor2_1 _5960_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[10] ),
    .A(_1926_),
    .B(_1928_));
 sg13g2_xor2_1 _5961_ (.B(net656),
    .A(net498),
    .X(_1929_));
 sg13g2_nand2_1 _5962_ (.Y(_1930_),
    .A(_1832_),
    .B(_1929_));
 sg13g2_xor2_1 _5963_ (.B(_1929_),
    .A(_1832_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_a[1] ));
 sg13g2_a21oi_2 _5964_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ),
    .Y(_1931_),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ),
    .A1(net498));
 sg13g2_nand3_1 _5965_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ),
    .A(net498),
    .Y(_1932_));
 sg13g2_nand2b_1 _5966_ (.Y(_1933_),
    .B(_1932_),
    .A_N(_1931_));
 sg13g2_xnor2_1 _5967_ (.Y(_1934_),
    .A(net406),
    .B(_1933_));
 sg13g2_xnor2_1 _5968_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[2] ),
    .A(_1930_),
    .B(_1934_));
 sg13g2_nor2_1 _5969_ (.A(_2917_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ),
    .Y(_1935_));
 sg13g2_nor2b_2 _5970_ (.A(net499),
    .B_N(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ),
    .Y(_1936_));
 sg13g2_inv_1 _5971_ (.Y(_1937_),
    .A(_1936_));
 sg13g2_nor2_1 _5972_ (.A(_1935_),
    .B(_1936_),
    .Y(_1938_));
 sg13g2_xnor2_1 _5973_ (.Y(_1939_),
    .A(_1931_),
    .B(_1938_));
 sg13g2_nand2_1 _5974_ (.Y(_1940_),
    .A(_3096_),
    .B(_1939_));
 sg13g2_xnor2_1 _5975_ (.Y(_1941_),
    .A(net406),
    .B(_1939_));
 sg13g2_inv_1 _5976_ (.Y(_1942_),
    .A(_1941_));
 sg13g2_and2_1 _5977_ (.A(_1929_),
    .B(_1934_),
    .X(_1943_));
 sg13g2_nor2b_1 _5978_ (.A(_1832_),
    .B_N(_1943_),
    .Y(_1944_));
 sg13g2_a21oi_1 _5979_ (.A1(_3096_),
    .A2(_1933_),
    .Y(_1945_),
    .B1(_1943_));
 sg13g2_nor2_1 _5980_ (.A(_1944_),
    .B(_1945_),
    .Y(_1946_));
 sg13g2_nand2_1 _5981_ (.Y(_1947_),
    .A(_1941_),
    .B(_1944_));
 sg13g2_xnor2_1 _5982_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[3] ),
    .A(_1942_),
    .B(_1946_));
 sg13g2_xnor2_1 _5983_ (.Y(_1948_),
    .A(net498),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_o21ai_1 _5984_ (.B1(_1937_),
    .Y(_1949_),
    .A1(_1931_),
    .A2(_1935_));
 sg13g2_xnor2_1 _5985_ (.Y(_1950_),
    .A(_1948_),
    .B(_1949_));
 sg13g2_nor2_1 _5986_ (.A(net407),
    .B(_1950_),
    .Y(_1951_));
 sg13g2_xnor2_1 _5987_ (.Y(_1952_),
    .A(net407),
    .B(_1950_));
 sg13g2_o21ai_1 _5988_ (.B1(_1940_),
    .Y(_1953_),
    .A1(_1942_),
    .A2(_1945_));
 sg13g2_xnor2_1 _5989_ (.Y(_1954_),
    .A(_1952_),
    .B(_1953_));
 sg13g2_nor2_1 _5990_ (.A(_1947_),
    .B(_1954_),
    .Y(_1955_));
 sg13g2_xnor2_1 _5991_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[4] ),
    .A(_1947_),
    .B(_1954_));
 sg13g2_o21ai_1 _5992_ (.B1(_1949_),
    .Y(_1956_),
    .A1(_2917_),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_o21ai_1 _5993_ (.B1(_1956_),
    .Y(_1957_),
    .A1(net498),
    .A2(_2963_));
 sg13g2_nor2_1 _5994_ (.A(_1935_),
    .B(_1957_),
    .Y(_1958_));
 sg13g2_o21ai_1 _5995_ (.B1(_3096_),
    .Y(_1959_),
    .A1(_1936_),
    .A2(_1958_));
 sg13g2_nor3_1 _5996_ (.A(_3096_),
    .B(_1936_),
    .C(_1958_),
    .Y(_1960_));
 sg13g2_nor2_1 _5997_ (.A(_1951_),
    .B(_1953_),
    .Y(_1961_));
 sg13g2_a21oi_2 _5998_ (.B1(_1961_),
    .Y(_1962_),
    .A2(_1950_),
    .A1(net406));
 sg13g2_a21oi_1 _5999_ (.A1(_1959_),
    .A2(_1962_),
    .Y(_1963_),
    .B1(_1960_));
 sg13g2_or2_1 _6000_ (.X(\main.demo._d___pip_58_1_2___stage___block_3_a[5] ),
    .B(_1963_),
    .A(_1955_));
 sg13g2_or2_1 _6001_ (.X(_1964_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ),
    .A(net498));
 sg13g2_xor2_1 _6002_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ),
    .A(net498),
    .X(_1965_));
 sg13g2_xnor2_1 _6003_ (.Y(_1966_),
    .A(_1957_),
    .B(_1965_));
 sg13g2_inv_1 _6004_ (.Y(_1967_),
    .A(_1966_));
 sg13g2_nand2_1 _6005_ (.Y(_1968_),
    .A(net406),
    .B(_1967_));
 sg13g2_xnor2_1 _6006_ (.Y(_1969_),
    .A(net406),
    .B(_1966_));
 sg13g2_xnor2_1 _6007_ (.Y(_1970_),
    .A(_1962_),
    .B(_1969_));
 sg13g2_nand2_1 _6008_ (.Y(_1971_),
    .A(_1955_),
    .B(_1970_));
 sg13g2_xnor2_1 _6009_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[6] ),
    .A(_1955_),
    .B(_1970_));
 sg13g2_nand3b_1 _6010_ (.B(_1962_),
    .C(_1968_),
    .Y(_1972_),
    .A_N(_1960_));
 sg13g2_o21ai_1 _6011_ (.B1(_1972_),
    .Y(_1973_),
    .A1(net406),
    .A2(_1967_));
 sg13g2_nand4_1 _6012_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ),
    .A(net498),
    .Y(_1974_),
    .D(_1949_));
 sg13g2_o21ai_1 _6013_ (.B1(_1974_),
    .Y(_1975_),
    .A1(_1957_),
    .A2(_1964_));
 sg13g2_xnor2_1 _6014_ (.Y(_1976_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_a[7] ),
    .B(_1975_));
 sg13g2_xnor2_1 _6015_ (.Y(_1977_),
    .A(net406),
    .B(_1976_));
 sg13g2_xnor2_1 _6016_ (.Y(_1978_),
    .A(_1973_),
    .B(_1977_));
 sg13g2_xnor2_1 _6017_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[7] ),
    .A(_1971_),
    .B(_1978_));
 sg13g2_nor2_1 _6018_ (.A(net493),
    .B(_0067_),
    .Y(_1979_));
 sg13g2_xnor2_1 _6019_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_a[6] ),
    .A(net493),
    .B(net295));
 sg13g2_xor2_1 _6020_ (.B(_1979_),
    .A(net292),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[7] ));
 sg13g2_nor2_1 _6021_ (.A(net403),
    .B(_3201_),
    .Y(_1980_));
 sg13g2_xnor2_1 _6022_ (.Y(_1981_),
    .A(_3222_),
    .B(_1980_));
 sg13g2_xnor2_1 _6023_ (.Y(_1982_),
    .A(_3205_),
    .B(_1981_));
 sg13g2_nand2_1 _6024_ (.Y(_1983_),
    .A(_3202_),
    .B(_1982_));
 sg13g2_xor2_1 _6025_ (.B(_1982_),
    .A(_3202_),
    .X(_1984_));
 sg13g2_nor2b_1 _6026_ (.A(net390),
    .B_N(_3233_),
    .Y(_1985_));
 sg13g2_xnor2_1 _6027_ (.Y(_1986_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_xnor2_1 _6028_ (.Y(_1987_),
    .A(_1985_),
    .B(_1986_));
 sg13g2_and2_1 _6029_ (.A(_1984_),
    .B(_1987_),
    .X(_1988_));
 sg13g2_xor2_1 _6030_ (.B(_1987_),
    .A(_1984_),
    .X(_1989_));
 sg13g2_xor2_1 _6031_ (.B(_1989_),
    .A(_3234_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[1] ));
 sg13g2_a21oi_1 _6032_ (.A1(_3234_),
    .A2(_1989_),
    .Y(_1990_),
    .B1(_1988_));
 sg13g2_o21ai_1 _6033_ (.B1(_1983_),
    .Y(_1991_),
    .A1(_3206_),
    .A2(_1981_));
 sg13g2_nand2_1 _6034_ (.Y(_1992_),
    .A(_3201_),
    .B(_3222_));
 sg13g2_nand2_1 _6035_ (.Y(_1993_),
    .A(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .B(_1992_));
 sg13g2_xor2_1 _6036_ (.B(_1993_),
    .A(_0400_),
    .X(_1994_));
 sg13g2_nor2b_1 _6037_ (.A(_3212_),
    .B_N(_1994_),
    .Y(_1995_));
 sg13g2_xnor2_1 _6038_ (.Y(_1996_),
    .A(_3212_),
    .B(_1994_));
 sg13g2_xnor2_1 _6039_ (.Y(_1997_),
    .A(_1991_),
    .B(_1996_));
 sg13g2_inv_1 _6040_ (.Y(_1998_),
    .A(_1997_));
 sg13g2_nor2_1 _6041_ (.A(_3233_),
    .B(_1986_),
    .Y(_1999_));
 sg13g2_nor2_1 _6042_ (.A(net389),
    .B(_1999_),
    .Y(_2000_));
 sg13g2_xnor2_1 _6043_ (.Y(_2001_),
    .A(_0406_),
    .B(_0407_));
 sg13g2_xor2_1 _6044_ (.B(_2001_),
    .A(_2000_),
    .X(_2002_));
 sg13g2_xnor2_1 _6045_ (.Y(_2003_),
    .A(_1997_),
    .B(_2002_));
 sg13g2_nor2b_1 _6046_ (.A(_1990_),
    .B_N(_2003_),
    .Y(_2004_));
 sg13g2_xnor2_1 _6047_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[2] ),
    .A(_1990_),
    .B(_2003_));
 sg13g2_a21oi_2 _6048_ (.B1(_2004_),
    .Y(_2005_),
    .A2(_2002_),
    .A1(_1998_));
 sg13g2_a21o_1 _6049_ (.A2(_1996_),
    .A1(_1991_),
    .B1(_1995_),
    .X(_2006_));
 sg13g2_nor2_1 _6050_ (.A(_0400_),
    .B(_1992_),
    .Y(_2007_));
 sg13g2_nor2_1 _6051_ (.A(net402),
    .B(_2007_),
    .Y(_2008_));
 sg13g2_xnor2_1 _6052_ (.Y(_2009_),
    .A(_0394_),
    .B(_2008_));
 sg13g2_xnor2_1 _6053_ (.Y(_2010_),
    .A(_3228_),
    .B(_2009_));
 sg13g2_nand2_1 _6054_ (.Y(_2011_),
    .A(_2006_),
    .B(_2010_));
 sg13g2_xnor2_1 _6055_ (.Y(_2012_),
    .A(_2006_),
    .B(_2010_));
 sg13g2_nand2_1 _6056_ (.Y(_2013_),
    .A(_1999_),
    .B(_2001_));
 sg13g2_nand2_1 _6057_ (.Y(_2014_),
    .A(_0420_),
    .B(_2013_));
 sg13g2_xnor2_1 _6058_ (.Y(_2015_),
    .A(_0408_),
    .B(_0409_));
 sg13g2_xnor2_1 _6059_ (.Y(_2016_),
    .A(_2014_),
    .B(_2015_));
 sg13g2_nor2_1 _6060_ (.A(_2012_),
    .B(_2016_),
    .Y(_2017_));
 sg13g2_xor2_1 _6061_ (.B(_2016_),
    .A(_2012_),
    .X(_2018_));
 sg13g2_nor2b_1 _6062_ (.A(_2005_),
    .B_N(_2018_),
    .Y(_2019_));
 sg13g2_xnor2_1 _6063_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[3] ),
    .A(_2005_),
    .B(_2018_));
 sg13g2_nor2_1 _6064_ (.A(_2017_),
    .B(_2019_),
    .Y(_2020_));
 sg13g2_o21ai_1 _6065_ (.B1(_2011_),
    .Y(_2021_),
    .A1(_3229_),
    .A2(_2009_));
 sg13g2_nand2_1 _6066_ (.Y(_2022_),
    .A(_0394_),
    .B(_2007_));
 sg13g2_nand2_1 _6067_ (.Y(_2023_),
    .A(net396),
    .B(_2022_));
 sg13g2_xor2_1 _6068_ (.B(_2023_),
    .A(_0390_),
    .X(_2024_));
 sg13g2_nor2b_1 _6069_ (.A(_0333_),
    .B_N(_2024_),
    .Y(_2025_));
 sg13g2_xnor2_1 _6070_ (.Y(_2026_),
    .A(_0333_),
    .B(_2024_));
 sg13g2_xor2_1 _6071_ (.B(_2026_),
    .A(_2021_),
    .X(_2027_));
 sg13g2_xnor2_1 _6072_ (.Y(_2028_),
    .A(_2021_),
    .B(_2026_));
 sg13g2_nor2_1 _6073_ (.A(_2013_),
    .B(_2015_),
    .Y(_2029_));
 sg13g2_nor2_1 _6074_ (.A(net388),
    .B(_2029_),
    .Y(_2030_));
 sg13g2_xnor2_1 _6075_ (.Y(_2031_),
    .A(_0387_),
    .B(_0411_));
 sg13g2_xor2_1 _6076_ (.B(_2031_),
    .A(_2030_),
    .X(_2032_));
 sg13g2_xnor2_1 _6077_ (.Y(_2033_),
    .A(_2028_),
    .B(_2032_));
 sg13g2_nor2b_1 _6078_ (.A(_2020_),
    .B_N(_2033_),
    .Y(_2034_));
 sg13g2_xnor2_1 _6079_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[4] ),
    .A(_2020_),
    .B(_2033_));
 sg13g2_a21oi_1 _6080_ (.A1(_2027_),
    .A2(_2032_),
    .Y(_2035_),
    .B1(_2034_));
 sg13g2_a21o_1 _6081_ (.A2(_2026_),
    .A1(_2021_),
    .B1(_2025_),
    .X(_2036_));
 sg13g2_nor2_1 _6082_ (.A(_0390_),
    .B(_2022_),
    .Y(_2037_));
 sg13g2_nor2_1 _6083_ (.A(net402),
    .B(_2037_),
    .Y(_2038_));
 sg13g2_xnor2_1 _6084_ (.Y(_2039_),
    .A(_0382_),
    .B(_2038_));
 sg13g2_xnor2_1 _6085_ (.Y(_2040_),
    .A(_0337_),
    .B(_2039_));
 sg13g2_nand2_1 _6086_ (.Y(_2041_),
    .A(_2036_),
    .B(_2040_));
 sg13g2_xnor2_1 _6087_ (.Y(_2042_),
    .A(_2036_),
    .B(_2040_));
 sg13g2_nand2_1 _6088_ (.Y(_2043_),
    .A(_2029_),
    .B(_2031_));
 sg13g2_nand2_1 _6089_ (.Y(_2044_),
    .A(_0420_),
    .B(_2043_));
 sg13g2_xnor2_1 _6090_ (.Y(_2045_),
    .A(_0412_),
    .B(_0413_));
 sg13g2_xnor2_1 _6091_ (.Y(_2046_),
    .A(_2044_),
    .B(_2045_));
 sg13g2_nor2_1 _6092_ (.A(_2042_),
    .B(_2046_),
    .Y(_2047_));
 sg13g2_xor2_1 _6093_ (.B(_2046_),
    .A(_2042_),
    .X(_2048_));
 sg13g2_nor2b_1 _6094_ (.A(_2035_),
    .B_N(_2048_),
    .Y(_2049_));
 sg13g2_xnor2_1 _6095_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[5] ),
    .A(_2035_),
    .B(_2048_));
 sg13g2_nor2_1 _6096_ (.A(_2047_),
    .B(_2049_),
    .Y(_2050_));
 sg13g2_o21ai_1 _6097_ (.B1(_2041_),
    .Y(_2051_),
    .A1(_0338_),
    .A2(_2039_));
 sg13g2_nand2_1 _6098_ (.Y(_2052_),
    .A(_0382_),
    .B(_2037_));
 sg13g2_nand2_1 _6099_ (.Y(_2053_),
    .A(net396),
    .B(_2052_));
 sg13g2_xor2_1 _6100_ (.B(_2053_),
    .A(_0378_),
    .X(_2054_));
 sg13g2_nor2b_1 _6101_ (.A(_0344_),
    .B_N(_2054_),
    .Y(_2055_));
 sg13g2_xnor2_1 _6102_ (.Y(_2056_),
    .A(_0344_),
    .B(_2054_));
 sg13g2_xor2_1 _6103_ (.B(_2056_),
    .A(_2051_),
    .X(_2057_));
 sg13g2_xnor2_1 _6104_ (.Y(_2058_),
    .A(_2051_),
    .B(_2056_));
 sg13g2_nor2_1 _6105_ (.A(_2043_),
    .B(_2045_),
    .Y(_2059_));
 sg13g2_nor2_1 _6106_ (.A(net388),
    .B(_2059_),
    .Y(_2060_));
 sg13g2_xnor2_1 _6107_ (.Y(_2061_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_xor2_1 _6108_ (.B(_2061_),
    .A(_2060_),
    .X(_2062_));
 sg13g2_xnor2_1 _6109_ (.Y(_2063_),
    .A(_2058_),
    .B(_2062_));
 sg13g2_nor2b_1 _6110_ (.A(_2050_),
    .B_N(_2063_),
    .Y(_2064_));
 sg13g2_xnor2_1 _6111_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[6] ),
    .A(_2050_),
    .B(_2063_));
 sg13g2_a21oi_1 _6112_ (.A1(_2057_),
    .A2(_2062_),
    .Y(_2065_),
    .B1(_2064_));
 sg13g2_a21o_1 _6113_ (.A2(_2056_),
    .A1(_2051_),
    .B1(_2055_),
    .X(_2066_));
 sg13g2_nor2_1 _6114_ (.A(_0378_),
    .B(_2052_),
    .Y(_2067_));
 sg13g2_nor2_1 _6115_ (.A(net402),
    .B(_2067_),
    .Y(_2068_));
 sg13g2_xnor2_1 _6116_ (.Y(_2069_),
    .A(_0370_),
    .B(_2068_));
 sg13g2_xnor2_1 _6117_ (.Y(_2070_),
    .A(_0347_),
    .B(_2069_));
 sg13g2_nand2_1 _6118_ (.Y(_2071_),
    .A(_2066_),
    .B(_2070_));
 sg13g2_xnor2_1 _6119_ (.Y(_2072_),
    .A(_2066_),
    .B(_2070_));
 sg13g2_inv_1 _6120_ (.Y(_2073_),
    .A(_2072_));
 sg13g2_or3_1 _6121_ (.A(_0368_),
    .B(_0373_),
    .C(_0417_),
    .X(_2074_));
 sg13g2_and2_2 _6122_ (.A(_0418_),
    .B(_2074_),
    .X(_2075_));
 sg13g2_nand2_1 _6123_ (.Y(_2076_),
    .A(_2059_),
    .B(_2061_));
 sg13g2_nand2_1 _6124_ (.Y(_2077_),
    .A(_0420_),
    .B(_2076_));
 sg13g2_xor2_1 _6125_ (.B(_2077_),
    .A(_2075_),
    .X(_2078_));
 sg13g2_xnor2_1 _6126_ (.Y(_2079_),
    .A(_2072_),
    .B(_2078_));
 sg13g2_nor2b_1 _6127_ (.A(_2065_),
    .B_N(_2079_),
    .Y(_2080_));
 sg13g2_xnor2_1 _6128_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[7] ),
    .A(_2065_),
    .B(_2079_));
 sg13g2_or3_2 _6129_ (.A(net388),
    .B(_2075_),
    .C(_2076_),
    .X(_2081_));
 sg13g2_o21ai_1 _6130_ (.B1(_2071_),
    .Y(_2082_),
    .A1(_0348_),
    .A2(_2069_));
 sg13g2_a21o_1 _6131_ (.A2(_2067_),
    .A1(_0370_),
    .B1(net402),
    .X(_2083_));
 sg13g2_xor2_1 _6132_ (.B(_2083_),
    .A(_0365_),
    .X(_2084_));
 sg13g2_xor2_1 _6133_ (.B(_2084_),
    .A(_0353_),
    .X(_2085_));
 sg13g2_nand2_1 _6134_ (.Y(_2086_),
    .A(_2082_),
    .B(_2085_));
 sg13g2_xnor2_1 _6135_ (.Y(_2087_),
    .A(_2082_),
    .B(_2085_));
 sg13g2_nor2_1 _6136_ (.A(_2081_),
    .B(_2087_),
    .Y(_2088_));
 sg13g2_xor2_1 _6137_ (.B(_2087_),
    .A(_2081_),
    .X(_2089_));
 sg13g2_a21oi_2 _6138_ (.B1(_2080_),
    .Y(_2090_),
    .A2(_2078_),
    .A1(_2073_));
 sg13g2_nor2b_1 _6139_ (.A(_2090_),
    .B_N(_2089_),
    .Y(_2091_));
 sg13g2_xnor2_1 _6140_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[8] ),
    .A(_2089_),
    .B(_2090_));
 sg13g2_o21ai_1 _6141_ (.B1(_2086_),
    .Y(_2092_),
    .A1(_0353_),
    .A2(_2084_));
 sg13g2_nand4_1 _6142_ (.B(_0365_),
    .C(_0370_),
    .A(net396),
    .Y(_2093_),
    .D(_2067_));
 sg13g2_nand2_1 _6143_ (.Y(_2094_),
    .A(_2092_),
    .B(_2093_));
 sg13g2_nand3_1 _6144_ (.B(_2092_),
    .C(_2093_),
    .A(_0357_),
    .Y(_2095_));
 sg13g2_xnor2_1 _6145_ (.Y(_2096_),
    .A(_0357_),
    .B(_2094_));
 sg13g2_inv_1 _6146_ (.Y(_2097_),
    .A(_2096_));
 sg13g2_xnor2_1 _6147_ (.Y(_2098_),
    .A(_2081_),
    .B(_2096_));
 sg13g2_nor2_1 _6148_ (.A(_2088_),
    .B(_2091_),
    .Y(_2099_));
 sg13g2_xnor2_1 _6149_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[9] ),
    .A(_2098_),
    .B(_2099_));
 sg13g2_a21oi_1 _6150_ (.A1(_2081_),
    .A2(_2097_),
    .Y(_2100_),
    .B1(_2099_));
 sg13g2_xnor2_1 _6151_ (.Y(_2101_),
    .A(_0361_),
    .B(_2095_));
 sg13g2_xor2_1 _6152_ (.B(_2101_),
    .A(_2081_),
    .X(_2102_));
 sg13g2_xnor2_1 _6153_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[10] ),
    .A(_2100_),
    .B(_2102_));
 sg13g2_xnor2_1 _6154_ (.Y(_2103_),
    .A(_3196_),
    .B(_3205_));
 sg13g2_nand2_1 _6155_ (.Y(_2104_),
    .A(_1998_),
    .B(_2103_));
 sg13g2_xnor2_1 _6156_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[0] ),
    .A(_1997_),
    .B(_2103_));
 sg13g2_xnor2_1 _6157_ (.Y(_2105_),
    .A(_3215_),
    .B(_3217_));
 sg13g2_nor2_1 _6158_ (.A(net390),
    .B(_1997_),
    .Y(_2106_));
 sg13g2_xnor2_1 _6159_ (.Y(_2107_),
    .A(_2012_),
    .B(_2106_));
 sg13g2_xor2_1 _6160_ (.B(_2107_),
    .A(_2105_),
    .X(_2108_));
 sg13g2_nor2b_1 _6161_ (.A(_2104_),
    .B_N(_2108_),
    .Y(_2109_));
 sg13g2_xnor2_1 _6162_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[1] ),
    .A(_2104_),
    .B(_2108_));
 sg13g2_and2_1 _6163_ (.A(_1997_),
    .B(_2012_),
    .X(_2110_));
 sg13g2_nor2_1 _6164_ (.A(net389),
    .B(_2110_),
    .Y(_2111_));
 sg13g2_xnor2_1 _6165_ (.Y(_2112_),
    .A(_2027_),
    .B(_2111_));
 sg13g2_nand2b_1 _6166_ (.Y(_2113_),
    .B(_3233_),
    .A_N(_2112_));
 sg13g2_xnor2_1 _6167_ (.Y(_2114_),
    .A(_3233_),
    .B(_2112_));
 sg13g2_inv_1 _6168_ (.Y(_2115_),
    .A(_2114_));
 sg13g2_a21oi_1 _6169_ (.A1(_2105_),
    .A2(_2107_),
    .Y(_2116_),
    .B1(_2109_));
 sg13g2_xnor2_1 _6170_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[2] ),
    .A(_2114_),
    .B(_2116_));
 sg13g2_o21ai_1 _6171_ (.B1(_2113_),
    .Y(_2117_),
    .A1(_2115_),
    .A2(_2116_));
 sg13g2_and2_1 _6172_ (.A(_2028_),
    .B(_2110_),
    .X(_2118_));
 sg13g2_nor2_1 _6173_ (.A(net389),
    .B(_2118_),
    .Y(_2119_));
 sg13g2_xnor2_1 _6174_ (.Y(_2120_),
    .A(_2042_),
    .B(_2119_));
 sg13g2_xnor2_1 _6175_ (.Y(_2121_),
    .A(_1986_),
    .B(_2120_));
 sg13g2_nor2b_1 _6176_ (.A(_2121_),
    .B_N(_2117_),
    .Y(_2122_));
 sg13g2_xnor2_1 _6177_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[3] ),
    .A(_2117_),
    .B(_2121_));
 sg13g2_and2_1 _6178_ (.A(_2042_),
    .B(_2118_),
    .X(_2123_));
 sg13g2_nor2_1 _6179_ (.A(net388),
    .B(_2123_),
    .Y(_2124_));
 sg13g2_xnor2_1 _6180_ (.Y(_2125_),
    .A(_2057_),
    .B(_2124_));
 sg13g2_nor2_1 _6181_ (.A(_2001_),
    .B(_2125_),
    .Y(_2126_));
 sg13g2_nand2_1 _6182_ (.Y(_2127_),
    .A(_2001_),
    .B(_2125_));
 sg13g2_nand2b_1 _6183_ (.Y(_2128_),
    .B(_2127_),
    .A_N(_2126_));
 sg13g2_a21o_1 _6184_ (.A2(_2120_),
    .A1(_1986_),
    .B1(_2122_),
    .X(_2129_));
 sg13g2_xnor2_1 _6185_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[4] ),
    .A(_2128_),
    .B(_2129_));
 sg13g2_a21oi_1 _6186_ (.A1(_2127_),
    .A2(_2129_),
    .Y(_2130_),
    .B1(_2126_));
 sg13g2_and2_1 _6187_ (.A(_2058_),
    .B(_2123_),
    .X(_2131_));
 sg13g2_nor2_1 _6188_ (.A(net389),
    .B(_2131_),
    .Y(_2132_));
 sg13g2_xnor2_1 _6189_ (.Y(_2133_),
    .A(_2072_),
    .B(_2132_));
 sg13g2_nand2_1 _6190_ (.Y(_2134_),
    .A(_2015_),
    .B(_2133_));
 sg13g2_xnor2_1 _6191_ (.Y(_2135_),
    .A(_2015_),
    .B(_2133_));
 sg13g2_xor2_1 _6192_ (.B(_2135_),
    .A(_2130_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_o21ai_1 _6193_ (.B1(_2134_),
    .Y(_2136_),
    .A1(_2130_),
    .A2(_2135_));
 sg13g2_and2_1 _6194_ (.A(_2072_),
    .B(_2131_),
    .X(_2137_));
 sg13g2_nor2_1 _6195_ (.A(net388),
    .B(_2137_),
    .Y(_2138_));
 sg13g2_xor2_1 _6196_ (.B(_2138_),
    .A(_2087_),
    .X(_2139_));
 sg13g2_nor2_1 _6197_ (.A(_2031_),
    .B(_2139_),
    .Y(_2140_));
 sg13g2_xor2_1 _6198_ (.B(_2139_),
    .A(_2031_),
    .X(_2141_));
 sg13g2_xor2_1 _6199_ (.B(_2141_),
    .A(_2136_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[6] ));
 sg13g2_a21oi_1 _6200_ (.A1(_2136_),
    .A2(_2141_),
    .Y(_2142_),
    .B1(_2140_));
 sg13g2_and2_1 _6201_ (.A(_2087_),
    .B(_2137_),
    .X(_2143_));
 sg13g2_nor2_1 _6202_ (.A(net388),
    .B(_2143_),
    .Y(_2144_));
 sg13g2_xor2_1 _6203_ (.B(_2144_),
    .A(_2096_),
    .X(_2145_));
 sg13g2_xnor2_1 _6204_ (.Y(_2146_),
    .A(_2045_),
    .B(_2145_));
 sg13g2_nor2_1 _6205_ (.A(_2142_),
    .B(_2146_),
    .Y(_2147_));
 sg13g2_xor2_1 _6206_ (.B(_2146_),
    .A(_2142_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[7] ));
 sg13g2_nor2_1 _6207_ (.A(_0420_),
    .B(_2101_),
    .Y(_2148_));
 sg13g2_nor2b_1 _6208_ (.A(_2096_),
    .B_N(_2143_),
    .Y(_2149_));
 sg13g2_nor2_1 _6209_ (.A(_2101_),
    .B(_2149_),
    .Y(_2150_));
 sg13g2_nor2_1 _6210_ (.A(net388),
    .B(_2150_),
    .Y(_2151_));
 sg13g2_nor2_2 _6211_ (.A(_2148_),
    .B(_2151_),
    .Y(_2152_));
 sg13g2_a21oi_1 _6212_ (.A1(_2101_),
    .A2(_2149_),
    .Y(_2153_),
    .B1(_2152_));
 sg13g2_nor2_1 _6213_ (.A(_2061_),
    .B(_2153_),
    .Y(_2154_));
 sg13g2_xnor2_1 _6214_ (.Y(_2155_),
    .A(_2061_),
    .B(_2153_));
 sg13g2_a21oi_1 _6215_ (.A1(_2045_),
    .A2(_2145_),
    .Y(_2156_),
    .B1(_2147_));
 sg13g2_nor2_1 _6216_ (.A(_2155_),
    .B(_2156_),
    .Y(_2157_));
 sg13g2_xor2_1 _6217_ (.B(_2156_),
    .A(_2155_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[8] ));
 sg13g2_nand2_1 _6218_ (.Y(_2158_),
    .A(_2075_),
    .B(_2152_));
 sg13g2_nor2_1 _6219_ (.A(_2075_),
    .B(_2152_),
    .Y(_2159_));
 sg13g2_xor2_1 _6220_ (.B(_2152_),
    .A(_2075_),
    .X(_2160_));
 sg13g2_nor2_1 _6221_ (.A(_2154_),
    .B(_2157_),
    .Y(_2161_));
 sg13g2_xnor2_1 _6222_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[9] ),
    .A(_2160_),
    .B(_2161_));
 sg13g2_nor2_1 _6223_ (.A(_2148_),
    .B(_2150_),
    .Y(_2162_));
 sg13g2_o21ai_1 _6224_ (.B1(_2158_),
    .Y(_2163_),
    .A1(_2159_),
    .A2(_2161_));
 sg13g2_xnor2_1 _6225_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[10] ),
    .A(_2162_),
    .B(_2163_));
 sg13g2_xnor2_1 _6226_ (.Y(_2164_),
    .A(\main.demo._t___stage___block_3_y[2] ),
    .B(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_nor2b_1 _6227_ (.A(\main.demo._t___stage___block_3_y[2] ),
    .B_N(\main.demo._q_frame[0] ),
    .Y(_2165_));
 sg13g2_o21ai_1 _6228_ (.B1(_2164_),
    .Y(_2166_),
    .A1(\main.demo._q_frame[1] ),
    .A2(_2165_));
 sg13g2_o21ai_1 _6229_ (.B1(_2166_),
    .Y(_2167_),
    .A1(\main.demo._t___stage___block_3_y[2] ),
    .A2(_1727_));
 sg13g2_o21ai_1 _6230_ (.B1(_2167_),
    .Y(_2168_),
    .A1(net502),
    .A2(_2940_));
 sg13g2_xnor2_1 _6231_ (.Y(_2169_),
    .A(\main.demo._t___stage___block_3_y[1] ),
    .B(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_inv_1 _6232_ (.Y(_2170_),
    .A(_2169_));
 sg13g2_a22oi_1 _6233_ (.Y(_2171_),
    .B1(_2169_),
    .B2(net501),
    .A2(_2940_),
    .A1(net502));
 sg13g2_a22oi_1 _6234_ (.Y(_2172_),
    .B1(_2168_),
    .B2(_2171_),
    .A2(\main.demo._t___stage___block_3_y[0] ),
    .A1(_2930_));
 sg13g2_o21ai_1 _6235_ (.B1(_2172_),
    .Y(_2173_),
    .A1(net501),
    .A2(_2169_));
 sg13g2_a22oi_1 _6236_ (.Y(_2174_),
    .B1(net438),
    .B2(\main.demo._q_frame[5] ),
    .A2(_2938_),
    .A1(\main.demo._q_frame[4] ));
 sg13g2_nand4_1 _6237_ (.B(\main.demo._q_frame[6] ),
    .C(\main.demo._q_go ),
    .A(net546),
    .Y(_2175_),
    .D(\main.demo._q_frame[8] ));
 sg13g2_a221oi_1 _6238_ (.B2(_2174_),
    .C1(net652),
    .B1(_2173_),
    .A1(_2929_),
    .Y(_2176_),
    .A2(net440));
 sg13g2_inv_1 _6239_ (.Y(_2177_),
    .A(_2176_));
 sg13g2_nor2b_1 _6240_ (.A(\main.demo._t___stage___block_3_y[2] ),
    .B_N(\main.demo._d___pip_58_1_4___stage___block_3_cx[1] ),
    .Y(_2178_));
 sg13g2_o21ai_1 _6241_ (.B1(_2178_),
    .Y(_2179_),
    .A1(_2943_),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ));
 sg13g2_a22oi_1 _6242_ (.Y(_2180_),
    .B1(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ),
    .B2(_2164_),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[3] ),
    .A1(_2940_));
 sg13g2_a22oi_1 _6243_ (.Y(_2181_),
    .B1(_2179_),
    .B2(_2180_),
    .A2(_2966_),
    .A1(\main.demo._t___stage___block_3_y[1] ));
 sg13g2_o21ai_1 _6244_ (.B1(_2181_),
    .Y(_2182_),
    .A1(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ),
    .A2(_2169_));
 sg13g2_a22oi_1 _6245_ (.Y(_2183_),
    .B1(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ),
    .B2(_2169_),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ),
    .A1(_2938_));
 sg13g2_a22oi_1 _6246_ (.Y(_2184_),
    .B1(_2182_),
    .B2(_2183_),
    .A2(_2965_),
    .A1(\main.demo._t___stage___block_3_y[0] ));
 sg13g2_o21ai_1 _6247_ (.B1(_2184_),
    .Y(_2185_),
    .A1(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ),
    .A2(net438));
 sg13g2_a21oi_1 _6248_ (.A1(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ),
    .A2(net438),
    .Y(_2186_),
    .B1(\main.demo._d___pip_58_1_4___stage___block_3_cx[9] ));
 sg13g2_and2_2 _6249_ (.A(_2185_),
    .B(_2186_),
    .X(_2187_));
 sg13g2_nand2_1 _6250_ (.Y(_2188_),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[3] ));
 sg13g2_nand2_1 _6251_ (.Y(_2189_),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_l[0] ),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[4] ));
 sg13g2_nor2_1 _6252_ (.A(_2188_),
    .B(_2189_),
    .Y(_2190_));
 sg13g2_and2_1 _6253_ (.A(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[1] ),
    .X(_2191_));
 sg13g2_nand2_1 _6254_ (.Y(_2192_),
    .A(net479),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[1] ));
 sg13g2_nand2_1 _6255_ (.Y(_2193_),
    .A(net480),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[0] ));
 sg13g2_nor3_1 _6256_ (.A(_2964_),
    .B(_2192_),
    .C(_2193_),
    .Y(_2194_));
 sg13g2_nand2_2 _6257_ (.Y(_2195_),
    .A(net480),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[2] ));
 sg13g2_nor2_1 _6258_ (.A(_2188_),
    .B(_2195_),
    .Y(_2196_));
 sg13g2_nor2_1 _6259_ (.A(_2194_),
    .B(_2196_),
    .Y(_2197_));
 sg13g2_o21ai_1 _6260_ (.B1(_2197_),
    .Y(_2198_),
    .A1(_2192_),
    .A2(_2195_));
 sg13g2_xor2_1 _6261_ (.B(_2189_),
    .A(_2188_),
    .X(_2199_));
 sg13g2_a21oi_1 _6262_ (.A1(_2198_),
    .A2(_2199_),
    .Y(_2200_),
    .B1(_2190_));
 sg13g2_nand2_1 _6263_ (.Y(_2201_),
    .A(net479),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[5] ));
 sg13g2_nor2_1 _6264_ (.A(_2189_),
    .B(_2201_),
    .Y(_2202_));
 sg13g2_a22oi_1 _6265_ (.Y(_2203_),
    .B1(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .B2(net479),
    .A2(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .A1(net480));
 sg13g2_nor2_1 _6266_ (.A(_2202_),
    .B(_2203_),
    .Y(_2204_));
 sg13g2_xor2_1 _6267_ (.B(_2204_),
    .A(_2200_),
    .X(_2205_));
 sg13g2_nand2_1 _6268_ (.Y(_2206_),
    .A(net414),
    .B(_2205_));
 sg13g2_nand2_1 _6269_ (.Y(_2207_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ));
 sg13g2_nand2_1 _6270_ (.Y(_2208_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_and2_1 _6271_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ),
    .X(_2209_));
 sg13g2_nand2_1 _6272_ (.Y(_2210_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_nand2_1 _6273_ (.Y(_2211_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_or2_1 _6274_ (.X(_2212_),
    .B(_2211_),
    .A(_2210_));
 sg13g2_xnor2_1 _6275_ (.Y(_2213_),
    .A(_2209_),
    .B(_2211_));
 sg13g2_nand2b_1 _6276_ (.Y(_2214_),
    .B(_2213_),
    .A_N(_2207_));
 sg13g2_xnor2_1 _6277_ (.Y(_2215_),
    .A(_2207_),
    .B(_2213_));
 sg13g2_nand2_2 _6278_ (.Y(_2216_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[1] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_inv_1 _6279_ (.Y(_2217_),
    .A(_2216_));
 sg13g2_nand2_1 _6280_ (.Y(_2218_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ));
 sg13g2_a22oi_1 _6281_ (.Y(_2219_),
    .B1(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ),
    .B2(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .A2(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ),
    .A1(\main.demo._d___pip_58_1_4___block_68_frag[1] ));
 sg13g2_a21oi_1 _6282_ (.A1(_2209_),
    .A2(_2217_),
    .Y(_2220_),
    .B1(_2219_));
 sg13g2_nand2b_1 _6283_ (.Y(_2221_),
    .B(_2220_),
    .A_N(_2218_));
 sg13g2_o21ai_1 _6284_ (.B1(_2221_),
    .Y(_2222_),
    .A1(_2210_),
    .A2(_2216_));
 sg13g2_and2_1 _6285_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[0] ),
    .B(_2217_),
    .X(_2223_));
 sg13g2_nand2_1 _6286_ (.Y(_2224_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[0] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_and2_1 _6287_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ),
    .X(_2225_));
 sg13g2_nand2_1 _6288_ (.Y(_2226_),
    .A(_2216_),
    .B(_2224_));
 sg13g2_xnor2_1 _6289_ (.Y(_2227_),
    .A(_2216_),
    .B(_2224_));
 sg13g2_a22oi_1 _6290_ (.Y(_2228_),
    .B1(_2225_),
    .B2(_2226_),
    .A2(_2223_),
    .A1(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_xnor2_1 _6291_ (.Y(_2229_),
    .A(_2218_),
    .B(_2220_));
 sg13g2_nand2b_1 _6292_ (.Y(_2230_),
    .B(_2229_),
    .A_N(_2228_));
 sg13g2_xnor2_1 _6293_ (.Y(_2231_),
    .A(_2225_),
    .B(_2227_));
 sg13g2_nand2_1 _6294_ (.Y(_2232_),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ),
    .B(_2223_));
 sg13g2_nand3_1 _6295_ (.B(_2223_),
    .C(_2231_),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ),
    .Y(_2233_));
 sg13g2_xnor2_1 _6296_ (.Y(_2234_),
    .A(_2228_),
    .B(_2229_));
 sg13g2_nand2b_1 _6297_ (.Y(_2235_),
    .B(_2234_),
    .A_N(_2233_));
 sg13g2_xnor2_1 _6298_ (.Y(_2236_),
    .A(_2215_),
    .B(_2222_));
 sg13g2_a21oi_1 _6299_ (.A1(_2230_),
    .A2(_2235_),
    .Y(_2237_),
    .B1(_2236_));
 sg13g2_a21oi_1 _6300_ (.A1(_2215_),
    .A2(_2222_),
    .Y(_2238_),
    .B1(_2237_));
 sg13g2_and2_1 _6301_ (.A(_2212_),
    .B(_2214_),
    .X(_2239_));
 sg13g2_nand2_1 _6302_ (.Y(_2240_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ));
 sg13g2_nand2_1 _6303_ (.Y(_2241_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_nand2_1 _6304_ (.Y(_2242_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_xor2_1 _6305_ (.B(_2242_),
    .A(_2208_),
    .X(_2243_));
 sg13g2_nand2b_1 _6306_ (.Y(_2244_),
    .B(_2243_),
    .A_N(_2240_));
 sg13g2_xnor2_1 _6307_ (.Y(_2245_),
    .A(_2240_),
    .B(_2243_));
 sg13g2_nor2b_1 _6308_ (.A(_2239_),
    .B_N(_2245_),
    .Y(_2246_));
 sg13g2_xnor2_1 _6309_ (.Y(_2247_),
    .A(_2239_),
    .B(_2245_));
 sg13g2_nor2b_1 _6310_ (.A(_2238_),
    .B_N(_2247_),
    .Y(_2248_));
 sg13g2_xnor2_1 _6311_ (.Y(_2249_),
    .A(_2238_),
    .B(_2247_));
 sg13g2_o21ai_1 _6312_ (.B1(_2206_),
    .Y(_2250_),
    .A1(net414),
    .A2(_2249_));
 sg13g2_nand2_1 _6313_ (.Y(_2251_),
    .A(net440),
    .B(_2250_));
 sg13g2_nand2b_1 _6314_ (.Y(_2252_),
    .B(net438),
    .A_N(_2250_));
 sg13g2_a21oi_1 _6315_ (.A1(_2193_),
    .A2(_2195_),
    .Y(_2253_),
    .B1(_2192_));
 sg13g2_a22oi_1 _6316_ (.Y(_2254_),
    .B1(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .B2(net479),
    .A2(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .A1(net480));
 sg13g2_nor2_1 _6317_ (.A(_2196_),
    .B(_2254_),
    .Y(_2255_));
 sg13g2_xnor2_1 _6318_ (.Y(_2256_),
    .A(_2253_),
    .B(_2255_));
 sg13g2_nand2_1 _6319_ (.Y(_2257_),
    .A(_2187_),
    .B(_2256_));
 sg13g2_xnor2_1 _6320_ (.Y(_2258_),
    .A(_2233_),
    .B(_2234_));
 sg13g2_o21ai_1 _6321_ (.B1(_2257_),
    .Y(_2259_),
    .A1(net414),
    .A2(_2258_));
 sg13g2_nand3_1 _6322_ (.B(_2235_),
    .C(_2236_),
    .A(_2230_),
    .Y(_2260_));
 sg13g2_nor2_1 _6323_ (.A(_2187_),
    .B(_2237_),
    .Y(_2261_));
 sg13g2_xor2_1 _6324_ (.B(_2199_),
    .A(_2198_),
    .X(_2262_));
 sg13g2_a22oi_1 _6325_ (.Y(_2263_),
    .B1(_2262_),
    .B2(net414),
    .A2(_2261_),
    .A1(_2260_));
 sg13g2_xor2_1 _6326_ (.B(_2263_),
    .A(_0004_),
    .X(_2264_));
 sg13g2_a21oi_1 _6327_ (.A1(_2170_),
    .A2(_2259_),
    .Y(_2265_),
    .B1(_2264_));
 sg13g2_nor2_1 _6328_ (.A(_2170_),
    .B(_2259_),
    .Y(_2266_));
 sg13g2_a21oi_1 _6329_ (.A1(_2191_),
    .A2(_2193_),
    .Y(_2267_),
    .B1(_2195_));
 sg13g2_nand3_1 _6330_ (.B(_2193_),
    .C(_2195_),
    .A(_2191_),
    .Y(_2268_));
 sg13g2_xnor2_1 _6331_ (.Y(_2269_),
    .A(_2231_),
    .B(_2232_));
 sg13g2_nand3b_1 _6332_ (.B(_2268_),
    .C(_2187_),
    .Y(_2270_),
    .A_N(_2267_));
 sg13g2_o21ai_1 _6333_ (.B1(_2270_),
    .Y(_2271_),
    .A1(net414),
    .A2(_2269_));
 sg13g2_nand3b_1 _6334_ (.B(_2271_),
    .C(\main.demo._t___stage___block_3_x[1] ),
    .Y(_2272_),
    .A_N(_2266_));
 sg13g2_nand4_1 _6335_ (.B(_2252_),
    .C(_2265_),
    .A(_2251_),
    .Y(_2273_),
    .D(_2272_));
 sg13g2_nor2_1 _6336_ (.A(\main.demo._t___stage___block_3_x[0] ),
    .B(_2263_),
    .Y(_2274_));
 sg13g2_nand2_1 _6337_ (.Y(_2275_),
    .A(_2251_),
    .B(_2274_));
 sg13g2_nand3_1 _6338_ (.B(_2273_),
    .C(_2275_),
    .A(_2252_),
    .Y(_2276_));
 sg13g2_xor2_1 _6339_ (.B(_2271_),
    .A(_0005_),
    .X(_2277_));
 sg13g2_nor2_1 _6340_ (.A(_2266_),
    .B(_2277_),
    .Y(_2278_));
 sg13g2_nand4_1 _6341_ (.B(_2252_),
    .C(_2265_),
    .A(_2251_),
    .Y(_2279_),
    .D(_2278_));
 sg13g2_nand2_1 _6342_ (.Y(_2280_),
    .A(_2276_),
    .B(_2279_));
 sg13g2_nand2b_1 _6343_ (.Y(_2281_),
    .B(_2200_),
    .A_N(_2202_));
 sg13g2_nand2b_1 _6344_ (.Y(_2282_),
    .B(_2281_),
    .A_N(_2203_));
 sg13g2_o21ai_1 _6345_ (.B1(net414),
    .Y(_2283_),
    .A1(_2201_),
    .A2(_2282_));
 sg13g2_a21oi_1 _6346_ (.A1(_2201_),
    .A2(_2282_),
    .Y(_2284_),
    .B1(_2283_));
 sg13g2_o21ai_1 _6347_ (.B1(_2244_),
    .Y(_2285_),
    .A1(_2208_),
    .A2(_2242_));
 sg13g2_nand2_1 _6348_ (.Y(_2286_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_xor2_1 _6349_ (.B(_2286_),
    .A(_2241_),
    .X(_2287_));
 sg13g2_nand2_1 _6350_ (.Y(_2288_),
    .A(_2285_),
    .B(_2287_));
 sg13g2_xor2_1 _6351_ (.B(_2287_),
    .A(_2285_),
    .X(_2289_));
 sg13g2_nor3_1 _6352_ (.A(_2246_),
    .B(_2248_),
    .C(_2289_),
    .Y(_2290_));
 sg13g2_o21ai_1 _6353_ (.B1(_2289_),
    .Y(_2291_),
    .A1(_2246_),
    .A2(_2248_));
 sg13g2_nor2_1 _6354_ (.A(net414),
    .B(_2290_),
    .Y(_2292_));
 sg13g2_a21oi_1 _6355_ (.A1(_2291_),
    .A2(_2292_),
    .Y(_2293_),
    .B1(_2284_));
 sg13g2_nand2_1 _6356_ (.Y(_2294_),
    .A(_2280_),
    .B(_2293_));
 sg13g2_or2_1 _6357_ (.X(_2295_),
    .B(_2293_),
    .A(_2280_));
 sg13g2_nand3_1 _6358_ (.B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ),
    .C(_2242_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .Y(_2296_));
 sg13g2_nand2_1 _6359_ (.Y(_2297_),
    .A(_2288_),
    .B(_2291_));
 sg13g2_xnor2_1 _6360_ (.Y(_2298_),
    .A(_2296_),
    .B(_2297_));
 sg13g2_o21ai_1 _6361_ (.B1(_2283_),
    .Y(_2299_),
    .A1(net414),
    .A2(_2298_));
 sg13g2_nand2b_1 _6362_ (.Y(_2300_),
    .B(_2299_),
    .A_N(_2295_));
 sg13g2_a21o_1 _6363_ (.A2(_2300_),
    .A1(_2294_),
    .B1(_2176_),
    .X(\main.demo._d_prev_b[0] ));
 sg13g2_nor2_1 _6364_ (.A(net471),
    .B(\main.demo._w_vga_vga_y[5] ),
    .Y(_2301_));
 sg13g2_nor2_1 _6365_ (.A(_2931_),
    .B(\main.demo._w_vga_vga_y[6] ),
    .Y(_2302_));
 sg13g2_or2_1 _6366_ (.X(_2303_),
    .B(_2302_),
    .A(_2301_));
 sg13g2_a21oi_1 _6367_ (.A1(\main.demo._w_vga_vga_y[5] ),
    .A2(_2302_),
    .Y(_2304_),
    .B1(_2301_));
 sg13g2_nor2_1 _6368_ (.A(net469),
    .B(_2304_),
    .Y(_2305_));
 sg13g2_nor2_1 _6369_ (.A(net466),
    .B(net467),
    .Y(_2306_));
 sg13g2_nand2_1 _6370_ (.Y(_2307_),
    .A(_2305_),
    .B(_2306_));
 sg13g2_nand2_1 _6371_ (.Y(_2308_),
    .A(\main.demo._w_vga_vga_x[9] ),
    .B(_2307_));
 sg13g2_nand2_1 _6372_ (.Y(_2309_),
    .A(\main.demo._w_vga_vga_y[6] ),
    .B(\main.demo._w_vga_vga_y[5] ));
 sg13g2_inv_1 _6373_ (.Y(_2310_),
    .A(_2309_));
 sg13g2_nand2_1 _6374_ (.Y(_2311_),
    .A(net471),
    .B(_2309_));
 sg13g2_inv_1 _6375_ (.Y(_2312_),
    .A(_2311_));
 sg13g2_nor2_2 _6376_ (.A(\main.demo._w_vga_vga_y[6] ),
    .B(\main.demo._w_vga_vga_y[5] ),
    .Y(_2313_));
 sg13g2_nor2_1 _6377_ (.A(_2931_),
    .B(_2313_),
    .Y(_2314_));
 sg13g2_o21ai_1 _6378_ (.B1(\main.demo._w_vga_vga_x[5] ),
    .Y(_2315_),
    .A1(\main.demo._w_vga_vga_y[6] ),
    .A2(\main.demo._w_vga_vga_y[5] ));
 sg13g2_nor2_2 _6379_ (.A(_2310_),
    .B(_2315_),
    .Y(_2316_));
 sg13g2_nand2_1 _6380_ (.Y(_2317_),
    .A(net466),
    .B(net467));
 sg13g2_a22oi_1 _6381_ (.Y(_2318_),
    .B1(_2316_),
    .B2(_2317_),
    .A2(_2312_),
    .A1(net469));
 sg13g2_nor4_1 _6382_ (.A(net466),
    .B(net467),
    .C(_0055_),
    .D(_2302_),
    .Y(_2319_));
 sg13g2_a221oi_1 _6383_ (.B2(_2319_),
    .C1(\main.demo._w_vga_vga_x[9] ),
    .B1(_2309_),
    .A1(net466),
    .Y(_2320_),
    .A2(_2305_));
 sg13g2_o21ai_1 _6384_ (.B1(_2320_),
    .Y(_2321_),
    .A1(_2306_),
    .A2(_2318_));
 sg13g2_and2_1 _6385_ (.A(_2308_),
    .B(_2321_),
    .X(_2322_));
 sg13g2_nor2_1 _6386_ (.A(net467),
    .B(net469),
    .Y(_2323_));
 sg13g2_nand3_1 _6387_ (.B(_0053_),
    .C(_2323_),
    .A(\main.demo._w_vga_vga_x[9] ),
    .Y(_2324_));
 sg13g2_nand2b_1 _6388_ (.Y(_2325_),
    .B(_2303_),
    .A_N(_2324_));
 sg13g2_nand2_1 _6389_ (.Y(_2326_),
    .A(net469),
    .B(_2316_));
 sg13g2_a21oi_1 _6390_ (.A1(\main.demo._w_vga_vga_y[6] ),
    .A2(_0062_),
    .Y(_2327_),
    .B1(_2302_));
 sg13g2_o21ai_1 _6391_ (.B1(_2326_),
    .Y(_2328_),
    .A1(net469),
    .A2(_2327_));
 sg13g2_nor2b_1 _6392_ (.A(net468),
    .B_N(net470),
    .Y(_2329_));
 sg13g2_nor3_1 _6393_ (.A(net471),
    .B(_2310_),
    .C(_2313_),
    .Y(_2330_));
 sg13g2_a22oi_1 _6394_ (.Y(_2331_),
    .B1(_2329_),
    .B2(_2330_),
    .A2(_2328_),
    .A1(net468));
 sg13g2_a21oi_1 _6395_ (.A1(net471),
    .A2(\main.demo._w_vga_vga_y[5] ),
    .Y(_2332_),
    .B1(_2303_));
 sg13g2_nand2_1 _6396_ (.Y(_2333_),
    .A(net467),
    .B(_2332_));
 sg13g2_a21oi_1 _6397_ (.A1(_0056_),
    .A2(_2935_),
    .Y(_2334_),
    .B1(net468));
 sg13g2_a21oi_1 _6398_ (.A1(_2311_),
    .A2(_2334_),
    .Y(_2335_),
    .B1(net470));
 sg13g2_a221oi_1 _6399_ (.B2(_2335_),
    .C1(_2927_),
    .B1(_2333_),
    .A1(net470),
    .Y(_2336_),
    .A2(_2316_));
 sg13g2_a21o_1 _6400_ (.A2(_2331_),
    .A1(_2927_),
    .B1(_2336_),
    .X(_2337_));
 sg13g2_o21ai_1 _6401_ (.B1(_2325_),
    .Y(_2338_),
    .A1(\main.demo._w_vga_vga_x[9] ),
    .A2(_2337_));
 sg13g2_nor2_1 _6402_ (.A(net469),
    .B(net471),
    .Y(_2339_));
 sg13g2_a21oi_1 _6403_ (.A1(\main.demo._w_vga_vga_y[6] ),
    .A2(_2339_),
    .Y(_2340_),
    .B1(_2323_));
 sg13g2_nand3b_1 _6404_ (.B(_2326_),
    .C(_2340_),
    .Y(_2341_),
    .A_N(_2305_));
 sg13g2_nor2_1 _6405_ (.A(_2301_),
    .B(_2316_),
    .Y(_2342_));
 sg13g2_nand2_1 _6406_ (.Y(_2343_),
    .A(_2928_),
    .B(_2342_));
 sg13g2_nand3_1 _6407_ (.B(_2341_),
    .C(_2343_),
    .A(net466),
    .Y(_2344_));
 sg13g2_a21oi_1 _6408_ (.A1(net469),
    .A2(_2314_),
    .Y(_2345_),
    .B1(_2928_));
 sg13g2_nor3_1 _6409_ (.A(net470),
    .B(net471),
    .C(_2309_),
    .Y(_2346_));
 sg13g2_nor2_1 _6410_ (.A(_2316_),
    .B(_2346_),
    .Y(_2347_));
 sg13g2_nand2_1 _6411_ (.Y(_2348_),
    .A(_2345_),
    .B(_2347_));
 sg13g2_nor3_1 _6412_ (.A(_0055_),
    .B(net471),
    .C(_2313_),
    .Y(_2349_));
 sg13g2_o21ai_1 _6413_ (.B1(_2348_),
    .Y(_2350_),
    .A1(net467),
    .A2(_2349_));
 sg13g2_o21ai_1 _6414_ (.B1(_2344_),
    .Y(_2351_),
    .A1(net466),
    .A2(_2350_));
 sg13g2_o21ai_1 _6415_ (.B1(_2308_),
    .Y(_2352_),
    .A1(\main.demo._w_vga_vga_x[9] ),
    .A2(_2351_));
 sg13g2_o21ai_1 _6416_ (.B1(_2931_),
    .Y(_2353_),
    .A1(_2310_),
    .A2(_2313_));
 sg13g2_nand3_1 _6417_ (.B(_2311_),
    .C(_2353_),
    .A(net470),
    .Y(_2354_));
 sg13g2_nand2_1 _6418_ (.Y(_2355_),
    .A(net468),
    .B(_2314_));
 sg13g2_mux2_1 _6419_ (.A0(net467),
    .A1(_2355_),
    .S(_2354_),
    .X(_2356_));
 sg13g2_o21ai_1 _6420_ (.B1(_2345_),
    .Y(_2357_),
    .A1(net469),
    .A2(_2342_));
 sg13g2_o21ai_1 _6421_ (.B1(_2315_),
    .Y(_2358_),
    .A1(_2329_),
    .A2(_2334_));
 sg13g2_nand3_1 _6422_ (.B(_2357_),
    .C(_2358_),
    .A(net466),
    .Y(_2359_));
 sg13g2_o21ai_1 _6423_ (.B1(_2359_),
    .Y(_2360_),
    .A1(net466),
    .A2(_2356_));
 sg13g2_nand2b_1 _6424_ (.Y(_2361_),
    .B(_2360_),
    .A_N(\main.demo._w_vga_vga_x[9] ));
 sg13g2_o21ai_1 _6425_ (.B1(_2361_),
    .Y(_2362_),
    .A1(_2324_),
    .A2(_2342_));
 sg13g2_nand2b_1 _6426_ (.Y(_2363_),
    .B(_2352_),
    .A_N(_2362_));
 sg13g2_or2_2 _6427_ (.X(_2364_),
    .B(_2362_),
    .A(_2322_));
 sg13g2_xnor2_1 _6428_ (.Y(_2365_),
    .A(\main.demo._w_vga_vga_x[4] ),
    .B(_2364_));
 sg13g2_xnor2_1 _6429_ (.Y(_2366_),
    .A(\main.demo._w_vga_vga_x[3] ),
    .B(_2364_));
 sg13g2_xnor2_1 _6430_ (.Y(_2367_),
    .A(_2943_),
    .B(_2364_));
 sg13g2_xnor2_1 _6431_ (.Y(_2368_),
    .A(_2941_),
    .B(_2364_));
 sg13g2_nand2_1 _6432_ (.Y(_2369_),
    .A(_2940_),
    .B(_2368_));
 sg13g2_xnor2_1 _6433_ (.Y(_2370_),
    .A(_0004_),
    .B(_2364_));
 sg13g2_nor2_1 _6434_ (.A(_2938_),
    .B(_2370_),
    .Y(_2371_));
 sg13g2_nand2b_1 _6435_ (.Y(_2372_),
    .B(\main.demo._t___stage___block_3_y[1] ),
    .A_N(_2368_));
 sg13g2_xnor2_1 _6436_ (.Y(_2373_),
    .A(_0003_),
    .B(_2367_));
 sg13g2_a21oi_1 _6437_ (.A1(_2369_),
    .A2(_2371_),
    .Y(_2374_),
    .B1(_2373_));
 sg13g2_a22oi_1 _6438_ (.Y(_2375_),
    .B1(_2372_),
    .B2(_2374_),
    .A2(_2367_),
    .A1(_2942_));
 sg13g2_a21oi_1 _6439_ (.A1(\main.demo._w_vga_vga_y[3] ),
    .A2(_2366_),
    .Y(_2376_),
    .B1(_2375_));
 sg13g2_nor2_1 _6440_ (.A(\main.demo._w_vga_vga_y[4] ),
    .B(_2365_),
    .Y(_2377_));
 sg13g2_nor2_1 _6441_ (.A(\main.demo._w_vga_vga_y[3] ),
    .B(_2366_),
    .Y(_2378_));
 sg13g2_nor3_1 _6442_ (.A(_2376_),
    .B(_2377_),
    .C(_2378_),
    .Y(_2379_));
 sg13g2_a21oi_1 _6443_ (.A1(\main.demo._w_vga_vga_y[4] ),
    .A2(_2365_),
    .Y(_2380_),
    .B1(_2379_));
 sg13g2_xnor2_1 _6444_ (.Y(_2381_),
    .A(_2363_),
    .B(_2380_));
 sg13g2_a21o_1 _6445_ (.A2(_2338_),
    .A1(_2322_),
    .B1(_2381_),
    .X(_2382_));
 sg13g2_or3_1 _6446_ (.A(_2322_),
    .B(_2338_),
    .C(_2363_),
    .X(_2383_));
 sg13g2_and2_2 _6447_ (.A(\main.demo._q_go ),
    .B(_0960_),
    .X(_2384_));
 sg13g2_nand2_2 _6448_ (.Y(_2385_),
    .A(\main.demo._q_go ),
    .B(_0960_));
 sg13g2_nor2b_1 _6449_ (.A(\main.demo._w_vga_vga_y[7] ),
    .B_N(_0059_),
    .Y(_2386_));
 sg13g2_nor4_2 _6450_ (.A(\main.demo._w_vga_vga_y[10] ),
    .B(\main.demo._w_vga_vga_y[8] ),
    .C(_2385_),
    .Y(_2387_),
    .D(_2386_));
 sg13g2_a22oi_1 _6451_ (.Y(_2388_),
    .B1(_2941_),
    .B2(\main.demo._q_th[2] ),
    .A2(_2939_),
    .A1(\main.demo._q_th[1] ));
 sg13g2_a221oi_1 _6452_ (.B2(_2910_),
    .C1(_2388_),
    .B1(\main.demo._t___stage___block_3_x[2] ),
    .A1(_2911_),
    .Y(_2389_),
    .A2(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_a221oi_1 _6453_ (.B2(\main.demo._q_th[3] ),
    .C1(_2389_),
    .B1(_2943_),
    .A1(\main.demo._q_th[4] ),
    .Y(_2390_),
    .A2(_2933_));
 sg13g2_nand2b_1 _6454_ (.Y(_2391_),
    .B(\main.demo._w_vga_vga_x[4] ),
    .A_N(\main.demo._q_th[5] ));
 sg13g2_o21ai_1 _6455_ (.B1(_2391_),
    .Y(_2392_),
    .A1(\main.demo._q_th[4] ),
    .A2(_2933_));
 sg13g2_nor2b_1 _6456_ (.A(\main.demo._w_vga_vga_x[4] ),
    .B_N(\main.demo._q_th[5] ),
    .Y(_2393_));
 sg13g2_nor4_1 _6457_ (.A(\main.demo._q_th[8] ),
    .B(\main.demo._q_th[7] ),
    .C(\main.demo._q_th[6] ),
    .D(_2393_),
    .Y(_2394_));
 sg13g2_o21ai_1 _6458_ (.B1(_2394_),
    .Y(_2395_),
    .A1(_2390_),
    .A2(_2392_));
 sg13g2_nand4_1 _6459_ (.B(_2383_),
    .C(_2387_),
    .A(_2382_),
    .Y(_2396_),
    .D(_2395_));
 sg13g2_nand4_1 _6460_ (.B(_2295_),
    .C(_2299_),
    .A(_2177_),
    .Y(\main.demo._d_prev_b[1] ),
    .D(_2396_));
 sg13g2_or2_1 _6461_ (.X(_2397_),
    .B(_0231_),
    .A(net298));
 sg13g2_and2_1 _6462_ (.A(net319),
    .B(net317),
    .X(_2398_));
 sg13g2_nor3_1 _6463_ (.A(net298),
    .B(_3325_),
    .C(_2398_),
    .Y(_0069_));
 sg13g2_and2_1 _6464_ (.A(net321),
    .B(_2398_),
    .X(_2399_));
 sg13g2_nor2_1 _6465_ (.A(net321),
    .B(_2398_),
    .Y(_2400_));
 sg13g2_nor3_1 _6466_ (.A(_2397_),
    .B(_2399_),
    .C(_2400_),
    .Y(_0070_));
 sg13g2_and2_1 _6467_ (.A(net351),
    .B(_2399_),
    .X(_2401_));
 sg13g2_nand2_1 _6468_ (.Y(_2402_),
    .A(net351),
    .B(_2399_));
 sg13g2_nor2_1 _6469_ (.A(net351),
    .B(_2399_),
    .Y(_2403_));
 sg13g2_nor3_1 _6470_ (.A(_2397_),
    .B(_2401_),
    .C(_2403_),
    .Y(_0071_));
 sg13g2_xnor2_1 _6471_ (.Y(_2404_),
    .A(net331),
    .B(_2401_));
 sg13g2_nor2_1 _6472_ (.A(_2397_),
    .B(_2404_),
    .Y(_0072_));
 sg13g2_nand2_1 _6473_ (.Y(_2405_),
    .A(net307),
    .B(net331));
 sg13g2_nor2_2 _6474_ (.A(_2402_),
    .B(_2405_),
    .Y(_2406_));
 sg13g2_and3_1 _6475_ (.X(_2407_),
    .A(net356),
    .B(net382),
    .C(_2406_));
 sg13g2_a21oi_1 _6476_ (.A1(net325),
    .A2(_2406_),
    .Y(_2408_),
    .B1(net356));
 sg13g2_nor3_1 _6477_ (.A(_2397_),
    .B(_2407_),
    .C(_2408_),
    .Y(_0073_));
 sg13g2_nand2_1 _6478_ (.Y(_2409_),
    .A(net620),
    .B(\main.demo.vga._q_ycount[2] ));
 sg13g2_nand3_1 _6479_ (.B(net527),
    .C(net428),
    .A(net621),
    .Y(_2410_));
 sg13g2_inv_1 _6480_ (.Y(_2411_),
    .A(_2410_));
 sg13g2_nor2_2 _6481_ (.A(_2409_),
    .B(_2410_),
    .Y(_2412_));
 sg13g2_and3_1 _6482_ (.X(_2413_),
    .A(net334),
    .B(\main.demo.vga._q_ycount[4] ),
    .C(_2412_));
 sg13g2_nand2_1 _6483_ (.Y(_2414_),
    .A(_0236_),
    .B(_2413_));
 sg13g2_xor2_1 _6484_ (.B(_2414_),
    .A(net372),
    .X(_2415_));
 sg13g2_nand4_1 _6485_ (.B(net594),
    .C(net515),
    .A(net428),
    .Y(_2416_),
    .D(_0239_));
 sg13g2_a21oi_1 _6486_ (.A1(_2415_),
    .A2(_2416_),
    .Y(_0074_),
    .B1(net456));
 sg13g2_nor2_1 _6487_ (.A(\main.demo._q_speed[6] ),
    .B(_1726_),
    .Y(_2417_));
 sg13g2_o21ai_1 _6488_ (.B1(_2384_),
    .Y(_2418_),
    .A1(net607),
    .A2(_2417_));
 sg13g2_a21oi_1 _6489_ (.A1(net607),
    .A2(_2417_),
    .Y(_0075_),
    .B1(_2418_));
 sg13g2_nor2_1 _6490_ (.A(_1726_),
    .B(net425),
    .Y(_2419_));
 sg13g2_nand2_2 _6491_ (.Y(_2420_),
    .A(net435),
    .B(_2384_));
 sg13g2_nand2_1 _6492_ (.Y(_2421_),
    .A(net503),
    .B(\main.demo._q_speed[1] ));
 sg13g2_xnor2_1 _6493_ (.Y(_2422_),
    .A(net503),
    .B(\main.demo._q_speed[1] ));
 sg13g2_nor2_1 _6494_ (.A(\main.demo._q_speed[0] ),
    .B(\main.demo._q_speed[6] ),
    .Y(_2423_));
 sg13g2_xnor2_1 _6495_ (.Y(_2424_),
    .A(_2422_),
    .B(_2423_));
 sg13g2_nor2_1 _6496_ (.A(net435),
    .B(net425),
    .Y(_2425_));
 sg13g2_nor3_1 _6497_ (.A(net641),
    .B(net435),
    .C(net426),
    .Y(_2426_));
 sg13g2_xnor2_1 _6498_ (.Y(_2427_),
    .A(net645),
    .B(_1725_));
 sg13g2_a221oi_1 _6499_ (.B2(net426),
    .C1(_2426_),
    .B1(_2427_),
    .A1(net419),
    .Y(_0076_),
    .A2(_2424_));
 sg13g2_nand2_1 _6500_ (.Y(_2428_),
    .A(\main.demo._q_speed[2] ),
    .B(\main.demo._q_speed[8] ));
 sg13g2_xor2_1 _6501_ (.B(\main.demo._q_speed[8] ),
    .A(\main.demo._q_speed[2] ),
    .X(_2429_));
 sg13g2_o21ai_1 _6502_ (.B1(_2421_),
    .Y(_2430_),
    .A1(_2422_),
    .A2(_2423_));
 sg13g2_nand2_1 _6503_ (.Y(_2431_),
    .A(_2429_),
    .B(_2430_));
 sg13g2_or2_1 _6504_ (.X(_2432_),
    .B(_2430_),
    .A(_2429_));
 sg13g2_nand3_1 _6505_ (.B(_2431_),
    .C(_2432_),
    .A(_2384_),
    .Y(_2433_));
 sg13g2_a21oi_1 _6506_ (.A1(\main.demo._q_frame[0] ),
    .A2(net435),
    .Y(_2434_),
    .B1(net616));
 sg13g2_nor2_1 _6507_ (.A(_1728_),
    .B(_2434_),
    .Y(_2435_));
 sg13g2_a21oi_1 _6508_ (.A1(net426),
    .A2(_2435_),
    .Y(_2436_),
    .B1(net417));
 sg13g2_a22oi_1 _6509_ (.Y(_0077_),
    .B1(_2433_),
    .B2(_2436_),
    .A2(net417),
    .A1(_2945_));
 sg13g2_nand2_1 _6510_ (.Y(_2437_),
    .A(\main.demo._q_speed[3] ),
    .B(\main.demo._q_speed[9] ));
 sg13g2_xnor2_1 _6511_ (.Y(_2438_),
    .A(\main.demo._q_speed[3] ),
    .B(\main.demo._q_speed[9] ));
 sg13g2_nand3_1 _6512_ (.B(_2431_),
    .C(_2438_),
    .A(_2428_),
    .Y(_2439_));
 sg13g2_a21o_1 _6513_ (.A2(_2431_),
    .A1(_2428_),
    .B1(_2438_),
    .X(_2440_));
 sg13g2_nand3_1 _6514_ (.B(_2439_),
    .C(_2440_),
    .A(_2384_),
    .Y(_2441_));
 sg13g2_xor2_1 _6515_ (.B(_1728_),
    .A(net502),
    .X(_2442_));
 sg13g2_o21ai_1 _6516_ (.B1(_2420_),
    .Y(_2443_),
    .A1(_2384_),
    .A2(_2442_));
 sg13g2_a22oi_1 _6517_ (.Y(_0078_),
    .B1(_2441_),
    .B2(_2443_),
    .A2(net417),
    .A1(_2946_));
 sg13g2_xnor2_1 _6518_ (.Y(_2444_),
    .A(\main.demo._q_speed[10] ),
    .B(\main.demo._q_speed[4] ));
 sg13g2_a21oi_1 _6519_ (.A1(_2437_),
    .A2(_2440_),
    .Y(_2445_),
    .B1(_2444_));
 sg13g2_nand3_1 _6520_ (.B(_2440_),
    .C(_2444_),
    .A(_2437_),
    .Y(_2446_));
 sg13g2_nand2_1 _6521_ (.Y(_2447_),
    .A(net419),
    .B(_2446_));
 sg13g2_xnor2_1 _6522_ (.Y(_2448_),
    .A(net501),
    .B(_1729_));
 sg13g2_a22oi_1 _6523_ (.Y(_2449_),
    .B1(_2448_),
    .B2(net426),
    .A2(net417),
    .A1(net585));
 sg13g2_o21ai_1 _6524_ (.B1(net586),
    .Y(_0079_),
    .A1(_2445_),
    .A2(_2447_));
 sg13g2_a21oi_1 _6525_ (.A1(\main.demo._q_speed[10] ),
    .A2(\main.demo._q_speed[4] ),
    .Y(_2450_),
    .B1(_2445_));
 sg13g2_and2_1 _6526_ (.A(net658),
    .B(\main.demo._q_speed[5] ),
    .X(_2451_));
 sg13g2_nand2_1 _6527_ (.Y(_2452_),
    .A(\main.demo._q_speed[11] ),
    .B(\main.demo._q_speed[5] ));
 sg13g2_nor2_1 _6528_ (.A(net658),
    .B(\main.demo._q_speed[5] ),
    .Y(_2453_));
 sg13g2_nor3_1 _6529_ (.A(_2450_),
    .B(_2451_),
    .C(_2453_),
    .Y(_2454_));
 sg13g2_o21ai_1 _6530_ (.B1(_2450_),
    .Y(_2455_),
    .A1(_2451_),
    .A2(_2453_));
 sg13g2_nand2_1 _6531_ (.Y(_2456_),
    .A(net419),
    .B(_2455_));
 sg13g2_xnor2_1 _6532_ (.Y(_2457_),
    .A(_2930_),
    .B(_1730_));
 sg13g2_a22oi_1 _6533_ (.Y(_2458_),
    .B1(_2457_),
    .B2(net426),
    .A2(net417),
    .A1(net573));
 sg13g2_o21ai_1 _6534_ (.B1(_2458_),
    .Y(_0080_),
    .A1(_2454_),
    .A2(_2456_));
 sg13g2_and2_1 _6535_ (.A(\main.demo._q_speed[6] ),
    .B(\main.demo._q_speed[12] ),
    .X(_2459_));
 sg13g2_xor2_1 _6536_ (.B(\main.demo._q_speed[12] ),
    .A(\main.demo._q_speed[6] ),
    .X(_2460_));
 sg13g2_o21ai_1 _6537_ (.B1(_2452_),
    .Y(_2461_),
    .A1(_2450_),
    .A2(_2453_));
 sg13g2_xnor2_1 _6538_ (.Y(_2462_),
    .A(_2460_),
    .B(_2461_));
 sg13g2_xnor2_1 _6539_ (.Y(_2463_),
    .A(_2929_),
    .B(_1731_));
 sg13g2_a22oi_1 _6540_ (.Y(_2464_),
    .B1(_2463_),
    .B2(net426),
    .A2(net417),
    .A1(net622));
 sg13g2_o21ai_1 _6541_ (.B1(_2464_),
    .Y(_0081_),
    .A1(_2420_),
    .A2(_2462_));
 sg13g2_xor2_1 _6542_ (.B(\main.demo._q_speed[13] ),
    .A(net503),
    .X(_2465_));
 sg13g2_a21o_1 _6543_ (.A2(_2461_),
    .A1(_2460_),
    .B1(_2459_),
    .X(_2466_));
 sg13g2_and2_1 _6544_ (.A(_2465_),
    .B(_2466_),
    .X(_2467_));
 sg13g2_o21ai_1 _6545_ (.B1(net419),
    .Y(_2468_),
    .A1(_2465_),
    .A2(_2466_));
 sg13g2_mux2_1 _6546_ (.A0(\main.demo._q_frame[6] ),
    .A1(_3238_),
    .S(_1731_),
    .X(_2469_));
 sg13g2_a22oi_1 _6547_ (.Y(_2470_),
    .B1(_2469_),
    .B2(net426),
    .A2(net417),
    .A1(net503));
 sg13g2_o21ai_1 _6548_ (.B1(_2470_),
    .Y(_0082_),
    .A1(_2467_),
    .A2(_2468_));
 sg13g2_xnor2_1 _6549_ (.Y(_2471_),
    .A(\main.demo._q_speed[8] ),
    .B(\main.demo._q_speed[14] ));
 sg13g2_a21oi_1 _6550_ (.A1(net503),
    .A2(\main.demo._q_speed[13] ),
    .Y(_2472_),
    .B1(_2467_));
 sg13g2_nor2_1 _6551_ (.A(_2471_),
    .B(_2472_),
    .Y(_2473_));
 sg13g2_a21o_1 _6552_ (.A2(_2472_),
    .A1(_2471_),
    .B1(_2420_),
    .X(_2474_));
 sg13g2_xor2_1 _6553_ (.B(_1732_),
    .A(net500),
    .X(_2475_));
 sg13g2_a22oi_1 _6554_ (.Y(_2476_),
    .B1(_2475_),
    .B2(net425),
    .A2(net418),
    .A1(net627));
 sg13g2_o21ai_1 _6555_ (.B1(_2476_),
    .Y(_0083_),
    .A1(_2473_),
    .A2(_2474_));
 sg13g2_nand2_1 _6556_ (.Y(_2477_),
    .A(net574),
    .B(net417));
 sg13g2_a21oi_2 _6557_ (.B1(_2473_),
    .Y(_2478_),
    .A2(\main.demo._q_speed[14] ),
    .A1(\main.demo._q_speed[8] ));
 sg13g2_nor2_1 _6558_ (.A(\main.demo._q_speed[9] ),
    .B(\main.demo._q_speed[15] ),
    .Y(_2479_));
 sg13g2_nand2_1 _6559_ (.Y(_2480_),
    .A(\main.demo._q_speed[9] ),
    .B(net659));
 sg13g2_nor2b_1 _6560_ (.A(_2479_),
    .B_N(_2480_),
    .Y(_2481_));
 sg13g2_o21ai_1 _6561_ (.B1(_2384_),
    .Y(_2482_),
    .A1(_2478_),
    .A2(_2481_));
 sg13g2_a21oi_1 _6562_ (.A1(_2478_),
    .A2(_2481_),
    .Y(_2483_),
    .B1(_2482_));
 sg13g2_xor2_1 _6563_ (.B(_1733_),
    .A(net636),
    .X(_2484_));
 sg13g2_a21oi_1 _6564_ (.A1(net425),
    .A2(_2484_),
    .Y(_2485_),
    .B1(_2419_));
 sg13g2_o21ai_1 _6565_ (.B1(_2477_),
    .Y(_0084_),
    .A1(_2483_),
    .A2(_2485_));
 sg13g2_o21ai_1 _6566_ (.B1(_2480_),
    .Y(_2486_),
    .A1(_2478_),
    .A2(_2479_));
 sg13g2_and2_1 _6567_ (.A(net583),
    .B(_2486_),
    .X(_2487_));
 sg13g2_o21ai_1 _6568_ (.B1(net419),
    .Y(_2488_),
    .A1(net583),
    .A2(_2486_));
 sg13g2_a22oi_1 _6569_ (.Y(_2489_),
    .B1(net418),
    .B2(net583),
    .A2(net427),
    .A1(_1736_));
 sg13g2_o21ai_1 _6570_ (.B1(net584),
    .Y(_0085_),
    .A1(_2487_),
    .A2(_2488_));
 sg13g2_and2_1 _6571_ (.A(net604),
    .B(_2487_),
    .X(_2490_));
 sg13g2_o21ai_1 _6572_ (.B1(net419),
    .Y(_2491_),
    .A1(net604),
    .A2(_2487_));
 sg13g2_xor2_1 _6573_ (.B(_1735_),
    .A(net629),
    .X(_2492_));
 sg13g2_a22oi_1 _6574_ (.Y(_2493_),
    .B1(_2492_),
    .B2(net425),
    .A2(net418),
    .A1(net604));
 sg13g2_o21ai_1 _6575_ (.B1(net605),
    .Y(_0086_),
    .A1(_2490_),
    .A2(_2491_));
 sg13g2_and2_1 _6576_ (.A(net579),
    .B(_2490_),
    .X(_2494_));
 sg13g2_o21ai_1 _6577_ (.B1(_2419_),
    .Y(_2495_),
    .A1(net579),
    .A2(_2490_));
 sg13g2_a21oi_1 _6578_ (.A1(\main.demo._q_frame[10] ),
    .A2(_1735_),
    .Y(_2496_),
    .B1(net602));
 sg13g2_nand3_1 _6579_ (.B(\main.demo._q_frame[10] ),
    .C(_1735_),
    .A(\main.demo._q_frame[11] ),
    .Y(_2497_));
 sg13g2_nor2b_1 _6580_ (.A(net603),
    .B_N(_2497_),
    .Y(_2498_));
 sg13g2_a22oi_1 _6581_ (.Y(_2499_),
    .B1(_2498_),
    .B2(net427),
    .A2(net418),
    .A1(net579));
 sg13g2_o21ai_1 _6582_ (.B1(net580),
    .Y(_0087_),
    .A1(_2494_),
    .A2(_2495_));
 sg13g2_and2_1 _6583_ (.A(net595),
    .B(_2494_),
    .X(_2500_));
 sg13g2_o21ai_1 _6584_ (.B1(net419),
    .Y(_2501_),
    .A1(net595),
    .A2(_2494_));
 sg13g2_nand4_1 _6585_ (.B(\main.demo._q_frame[10] ),
    .C(\main.demo._q_frame[12] ),
    .A(net602),
    .Y(_2502_),
    .D(_1735_));
 sg13g2_xnor2_1 _6586_ (.Y(_2503_),
    .A(net649),
    .B(_2497_));
 sg13g2_a22oi_1 _6587_ (.Y(_2504_),
    .B1(_2503_),
    .B2(net427),
    .A2(net418),
    .A1(net595));
 sg13g2_o21ai_1 _6588_ (.B1(_2504_),
    .Y(_0088_),
    .A1(_2500_),
    .A2(_2501_));
 sg13g2_nand2_1 _6589_ (.Y(_2505_),
    .A(net598),
    .B(_2500_));
 sg13g2_nor2_1 _6590_ (.A(net598),
    .B(_2500_),
    .Y(_2506_));
 sg13g2_nand2_1 _6591_ (.Y(_2507_),
    .A(net419),
    .B(_2505_));
 sg13g2_nor2_1 _6592_ (.A(_2944_),
    .B(_2502_),
    .Y(_2508_));
 sg13g2_xnor2_1 _6593_ (.Y(_2509_),
    .A(net618),
    .B(_2502_));
 sg13g2_a22oi_1 _6594_ (.Y(_2510_),
    .B1(_2509_),
    .B2(net425),
    .A2(net418),
    .A1(net598));
 sg13g2_o21ai_1 _6595_ (.B1(net599),
    .Y(_0089_),
    .A1(_2506_),
    .A2(_2507_));
 sg13g2_or2_1 _6596_ (.X(_2511_),
    .B(_2505_),
    .A(net606));
 sg13g2_a21oi_1 _6597_ (.A1(net606),
    .A2(_2505_),
    .Y(_2512_),
    .B1(_2420_));
 sg13g2_xnor2_1 _6598_ (.Y(_2513_),
    .A(net562),
    .B(_2508_));
 sg13g2_nor3_1 _6599_ (.A(net606),
    .B(net435),
    .C(net425),
    .Y(_2514_));
 sg13g2_a221oi_1 _6600_ (.B2(net425),
    .C1(_2514_),
    .B1(net563),
    .A1(_2511_),
    .Y(_0090_),
    .A2(_2512_));
 sg13g2_nor2_1 _6601_ (.A(net458),
    .B(net646),
    .Y(_0091_));
 sg13g2_nor3_1 _6602_ (.A(net458),
    .B(_1728_),
    .C(net617),
    .Y(_0092_));
 sg13g2_and2_1 _6603_ (.A(net508),
    .B(_2442_),
    .X(_0093_));
 sg13g2_and2_1 _6604_ (.A(net508),
    .B(_2448_),
    .X(_0094_));
 sg13g2_and2_1 _6605_ (.A(net509),
    .B(_2457_),
    .X(_0095_));
 sg13g2_and2_1 _6606_ (.A(net509),
    .B(_2463_),
    .X(_0096_));
 sg13g2_and2_1 _6607_ (.A(net509),
    .B(_2469_),
    .X(_0097_));
 sg13g2_and2_1 _6608_ (.A(net509),
    .B(_2475_),
    .X(_0098_));
 sg13g2_and2_1 _6609_ (.A(net508),
    .B(net637),
    .X(_0099_));
 sg13g2_and2_1 _6610_ (.A(net509),
    .B(_1736_),
    .X(_0100_));
 sg13g2_and2_1 _6611_ (.A(net509),
    .B(_2492_),
    .X(_0101_));
 sg13g2_and2_1 _6612_ (.A(net508),
    .B(_2498_),
    .X(_0102_));
 sg13g2_and2_1 _6613_ (.A(net508),
    .B(net650),
    .X(_0103_));
 sg13g2_and2_1 _6614_ (.A(net508),
    .B(net619),
    .X(_0104_));
 sg13g2_nor2_1 _6615_ (.A(net458),
    .B(net563),
    .Y(_0105_));
 sg13g2_a21oi_2 _6616_ (.B1(_2503_),
    .Y(_2515_),
    .A2(_1734_),
    .A1(_0935_));
 sg13g2_o21ai_1 _6617_ (.B1(net509),
    .Y(_2516_),
    .A1(net308),
    .A2(_2515_));
 sg13g2_a21oi_1 _6618_ (.A1(_2913_),
    .A2(_2515_),
    .Y(_0106_),
    .B1(net309));
 sg13g2_mux2_1 _6619_ (.A0(net476),
    .A1(net547),
    .S(_1734_),
    .X(_2517_));
 sg13g2_and3_1 _6620_ (.X(_0107_),
    .A(net508),
    .B(\main.demo._q_go ),
    .C(_2517_));
 sg13g2_nand3_1 _6621_ (.B(\main.demo._q_go ),
    .C(_0961_),
    .A(net508),
    .Y(_2518_));
 sg13g2_a21oi_1 _6622_ (.A1(net441),
    .A2(_1734_),
    .Y(_2519_),
    .B1(_2518_));
 sg13g2_o21ai_1 _6623_ (.B1(_2519_),
    .Y(_0108_),
    .A1(net459),
    .A2(_1734_));
 sg13g2_nand4_1 _6624_ (.B(\main.demo._q_frame[4] ),
    .C(net501),
    .A(net500),
    .Y(_2520_),
    .D(_3237_));
 sg13g2_nand4_1 _6625_ (.B(\main.demo._q_frame[1] ),
    .C(\main.demo._q_frame[0] ),
    .A(net502),
    .Y(_2521_),
    .D(\main.demo._q_frame[8] ));
 sg13g2_o21ai_1 _6626_ (.B1(\main.demo._q_go ),
    .Y(_2522_),
    .A1(_2520_),
    .A2(_2521_));
 sg13g2_nand2_1 _6627_ (.Y(_2523_),
    .A(\main.demo._q_th[0] ),
    .B(_1726_));
 sg13g2_nand2_1 _6628_ (.Y(_2524_),
    .A(net287),
    .B(net435));
 sg13g2_a21oi_1 _6629_ (.A1(_2523_),
    .A2(_2524_),
    .Y(_0109_),
    .B1(net424));
 sg13g2_and3_1 _6630_ (.X(_2525_),
    .A(net304),
    .B(\main.demo._q_th[0] ),
    .C(net435));
 sg13g2_a21oi_1 _6631_ (.A1(\main.demo._q_th[0] ),
    .A2(net435),
    .Y(_2526_),
    .B1(net304));
 sg13g2_nor3_1 _6632_ (.A(net424),
    .B(_2525_),
    .C(net305),
    .Y(_0110_));
 sg13g2_and2_1 _6633_ (.A(net596),
    .B(_2525_),
    .X(_2527_));
 sg13g2_nor2_1 _6634_ (.A(net596),
    .B(_2525_),
    .Y(_2528_));
 sg13g2_nor3_1 _6635_ (.A(net424),
    .B(_2527_),
    .C(net597),
    .Y(_0111_));
 sg13g2_nor2_1 _6636_ (.A(net612),
    .B(_2527_),
    .Y(_2529_));
 sg13g2_and2_1 _6637_ (.A(net612),
    .B(_2527_),
    .X(_2530_));
 sg13g2_nor3_1 _6638_ (.A(net424),
    .B(_2529_),
    .C(_2530_),
    .Y(_0112_));
 sg13g2_nor2_1 _6639_ (.A(net379),
    .B(_2530_),
    .Y(_2531_));
 sg13g2_and2_1 _6640_ (.A(net379),
    .B(_2530_),
    .X(_2532_));
 sg13g2_nor3_1 _6641_ (.A(_2522_),
    .B(net380),
    .C(_2532_),
    .Y(_0113_));
 sg13g2_nor2_1 _6642_ (.A(net631),
    .B(_2532_),
    .Y(_2533_));
 sg13g2_and2_1 _6643_ (.A(\main.demo._q_th[5] ),
    .B(_2532_),
    .X(_2534_));
 sg13g2_nor3_1 _6644_ (.A(net424),
    .B(_2533_),
    .C(_2534_),
    .Y(_0114_));
 sg13g2_xnor2_1 _6645_ (.Y(_2535_),
    .A(net555),
    .B(_2534_));
 sg13g2_nor2_1 _6646_ (.A(net424),
    .B(_2535_),
    .Y(_0115_));
 sg13g2_nor2b_1 _6647_ (.A(net624),
    .B_N(_2534_),
    .Y(_2536_));
 sg13g2_xnor2_1 _6648_ (.Y(_2537_),
    .A(\main.demo._q_th[7] ),
    .B(_2536_));
 sg13g2_nor2_1 _6649_ (.A(net424),
    .B(net625),
    .Y(_0116_));
 sg13g2_nand3_1 _6650_ (.B(\main.demo._q_th[6] ),
    .C(_2534_),
    .A(\main.demo._q_th[7] ),
    .Y(_2538_));
 sg13g2_xor2_1 _6651_ (.B(_2538_),
    .A(net383),
    .X(_2539_));
 sg13g2_nor2_1 _6652_ (.A(net424),
    .B(net384),
    .Y(_0117_));
 sg13g2_mux4_1 _6653_ (.S0(net480),
    .A0(net537),
    .A1(net284),
    .A2(\main.demo._d_prev_b[5] ),
    .A3(\main.demo._d_prev_b[3] ),
    .S1(net479),
    .X(_2540_));
 sg13g2_and2_1 _6654_ (.A(net536),
    .B(net538),
    .X(_0118_));
 sg13g2_and2_1 _6655_ (.A(net536),
    .B(\main.demo._d_prev_b[1] ),
    .X(_0119_));
 sg13g2_mux4_1 _6656_ (.S0(net480),
    .A0(net283),
    .A1(net282),
    .A2(net284),
    .A3(net537),
    .S1(net479),
    .X(_2541_));
 sg13g2_and2_1 _6657_ (.A(net536),
    .B(_2541_),
    .X(_0120_));
 sg13g2_mux4_1 _6658_ (.S0(net480),
    .A0(net544),
    .A1(net278),
    .A2(net280),
    .A3(net281),
    .S1(net479),
    .X(_2542_));
 sg13g2_and2_1 _6659_ (.A(net536),
    .B(_2542_),
    .X(_0121_));
 sg13g2_and2_1 _6660_ (.A(net536),
    .B(\main.demo._d_prev_b[0] ),
    .X(_0122_));
 sg13g2_mux4_1 _6661_ (.S0(net480),
    .A0(net281),
    .A1(net280),
    .A2(net278),
    .A3(net544),
    .S1(net479),
    .X(_2543_));
 sg13g2_and2_1 _6662_ (.A(net536),
    .B(_2543_),
    .X(_0123_));
 sg13g2_nand2b_1 _6663_ (.Y(_2544_),
    .B(\main.demo.zic._q_rythm_count[12] ),
    .A_N(\main.demo.zic._q_rythm_count[11] ));
 sg13g2_nor4_2 _6664_ (.A(_2906_),
    .B(\main.demo.zic._q_rythm_count[9] ),
    .C(\main.demo.zic._q_rythm_count[8] ),
    .Y(_2545_),
    .D(_2544_));
 sg13g2_or4_1 _6665_ (.A(_2906_),
    .B(\main.demo.zic._q_rythm_count[9] ),
    .C(\main.demo.zic._q_rythm_count[8] ),
    .D(_2544_),
    .X(_2546_));
 sg13g2_nor3_1 _6666_ (.A(\main.demo.zic._q_clock_count[7] ),
    .B(\main.demo.zic._q_clock_count[6] ),
    .C(\main.demo.zic._q_clock_count[8] ),
    .Y(_2547_));
 sg13g2_nor2_1 _6667_ (.A(net609),
    .B(\main.demo.zic._q_clock_count[0] ),
    .Y(_2548_));
 sg13g2_nor4_1 _6668_ (.A(\main.demo.zic._q_clock_count[3] ),
    .B(\main.demo.zic._q_clock_count[2] ),
    .C(\main.demo.zic._q_clock_count[5] ),
    .D(\main.demo.zic._q_clock_count[4] ),
    .Y(_2549_));
 sg13g2_and3_2 _6669_ (.X(_2550_),
    .A(_2547_),
    .B(_2548_),
    .C(_2549_));
 sg13g2_nand3_1 _6670_ (.B(_2548_),
    .C(_2549_),
    .A(_2547_),
    .Y(_2551_));
 sg13g2_nor4_1 _6671_ (.A(\main.demo.zic._q_rythm_count[7] ),
    .B(\main.demo.zic._q_rythm_count[6] ),
    .C(\main.demo.zic._q_rythm_count[5] ),
    .D(\main.demo.zic._q_rythm_count[4] ),
    .Y(_2552_));
 sg13g2_nor4_1 _6672_ (.A(\main.demo.zic._q_rythm_count[3] ),
    .B(\main.demo.zic._q_rythm_count[2] ),
    .C(\main.demo.zic._q_rythm_count[1] ),
    .D(\main.demo.zic._q_rythm_count[0] ),
    .Y(_2553_));
 sg13g2_nand3_1 _6673_ (.B(_2552_),
    .C(_2553_),
    .A(net429),
    .Y(_2554_));
 sg13g2_and2_1 _6674_ (.A(net433),
    .B(_2554_),
    .X(_2555_));
 sg13g2_nand2_2 _6675_ (.Y(_2556_),
    .A(\main.demo.zic._q_idx[1] ),
    .B(\main.demo.zic._q_idx[0] ));
 sg13g2_and2_2 _6676_ (.A(\main.demo.zic._q_idx[3] ),
    .B(net464),
    .X(_2557_));
 sg13g2_nand2_2 _6677_ (.Y(_2558_),
    .A(net463),
    .B(net465));
 sg13g2_nor2_2 _6678_ (.A(_2556_),
    .B(_2558_),
    .Y(_2559_));
 sg13g2_nand2b_2 _6679_ (.Y(_2560_),
    .B(_2557_),
    .A_N(_2556_));
 sg13g2_nor2b_1 _6680_ (.A(\main.demo.zic._q_idx[5] ),
    .B_N(\main.demo.zic._q_idx[6] ),
    .Y(_2561_));
 sg13g2_nand2_2 _6681_ (.Y(_2562_),
    .A(net462),
    .B(_2561_));
 sg13g2_nor2_1 _6682_ (.A(_2560_),
    .B(_2562_),
    .Y(_2563_));
 sg13g2_nor2_2 _6683_ (.A(net433),
    .B(_2563_),
    .Y(_2564_));
 sg13g2_nand3_1 _6684_ (.B(net462),
    .C(_2559_),
    .A(\main.demo.zic._q_idx[5] ),
    .Y(_2565_));
 sg13g2_xor2_1 _6685_ (.B(_2565_),
    .A(_0033_),
    .X(_2566_));
 sg13g2_a22oi_1 _6686_ (.Y(_2567_),
    .B1(_2564_),
    .B2(_2566_),
    .A2(net433),
    .A1(net632));
 sg13g2_nor2_1 _6687_ (.A(_0032_),
    .B(_2560_),
    .Y(_2568_));
 sg13g2_xnor2_1 _6688_ (.Y(_2569_),
    .A(\main.demo.zic._q_idx[5] ),
    .B(_2568_));
 sg13g2_a22oi_1 _6689_ (.Y(_2570_),
    .B1(_2564_),
    .B2(_2569_),
    .A2(net433),
    .A1(net613));
 sg13g2_nand2b_1 _6690_ (.Y(_2571_),
    .B(_2567_),
    .A_N(_2570_));
 sg13g2_nand4_1 _6691_ (.B(\main.demo.zic._q_idx[1] ),
    .C(\main.demo.zic._q_idx[0] ),
    .A(net465),
    .Y(_2572_),
    .D(_2545_));
 sg13g2_or2_1 _6692_ (.X(_2573_),
    .B(_2556_),
    .A(_2546_));
 sg13g2_xnor2_1 _6693_ (.Y(_2574_),
    .A(_0032_),
    .B(_2559_));
 sg13g2_a22oi_1 _6694_ (.Y(_2575_),
    .B1(_2564_),
    .B2(_2574_),
    .A2(net433),
    .A1(net462));
 sg13g2_inv_1 _6695_ (.Y(_2576_),
    .A(_2575_));
 sg13g2_xor2_1 _6696_ (.B(_2573_),
    .A(net465),
    .X(_2577_));
 sg13g2_nor2_1 _6697_ (.A(net463),
    .B(_2577_),
    .Y(_2578_));
 sg13g2_a22oi_1 _6698_ (.Y(_2579_),
    .B1(_2572_),
    .B2(_2914_),
    .A2(_2559_),
    .A1(_2545_));
 sg13g2_xnor2_1 _6699_ (.Y(_2580_),
    .A(\main.demo.zic._q_idx[0] ),
    .B(net433));
 sg13g2_nand3_1 _6700_ (.B(\main.demo.zic._q_idx[1] ),
    .C(_2580_),
    .A(net463),
    .Y(_2581_));
 sg13g2_a22oi_1 _6701_ (.Y(_2582_),
    .B1(_2581_),
    .B2(_2577_),
    .A2(_2578_),
    .A1(_2575_));
 sg13g2_nor2_2 _6702_ (.A(_2914_),
    .B(net464),
    .Y(_2583_));
 sg13g2_nand2_1 _6703_ (.Y(_2584_),
    .A(_2575_),
    .B(_2583_));
 sg13g2_a21oi_1 _6704_ (.A1(_2556_),
    .A2(_2584_),
    .Y(_2585_),
    .B1(_2580_));
 sg13g2_nand3_1 _6705_ (.B(_2567_),
    .C(_2575_),
    .A(_2558_),
    .Y(_2586_));
 sg13g2_nand2_1 _6706_ (.Y(_2587_),
    .A(_2571_),
    .B(_2586_));
 sg13g2_nand2b_1 _6707_ (.Y(_2588_),
    .B(_2570_),
    .A_N(_2567_));
 sg13g2_a21oi_1 _6708_ (.A1(\main.demo.zic._q_idx[0] ),
    .A2(_2545_),
    .Y(_2589_),
    .B1(\main.demo.zic._q_idx[1] ));
 sg13g2_inv_1 _6709_ (.Y(_2590_),
    .A(_2589_));
 sg13g2_nand3_1 _6710_ (.B(_2588_),
    .C(_2590_),
    .A(_2572_),
    .Y(_2591_));
 sg13g2_nand2_1 _6711_ (.Y(_2592_),
    .A(_2573_),
    .B(_2590_));
 sg13g2_nor3_1 _6712_ (.A(net465),
    .B(_2580_),
    .C(_2592_),
    .Y(_2593_));
 sg13g2_nand2_1 _6713_ (.Y(_2594_),
    .A(_2579_),
    .B(_2593_));
 sg13g2_nor3_1 _6714_ (.A(_2585_),
    .B(_2587_),
    .C(_2591_),
    .Y(_2595_));
 sg13g2_nor4_1 _6715_ (.A(_2567_),
    .B(_2570_),
    .C(_2576_),
    .D(_2594_),
    .Y(_2596_));
 sg13g2_a21oi_1 _6716_ (.A1(_2571_),
    .A2(_2586_),
    .Y(_2597_),
    .B1(_2592_));
 sg13g2_nor4_1 _6717_ (.A(net433),
    .B(_2595_),
    .C(_2596_),
    .D(_2597_),
    .Y(_2598_));
 sg13g2_o21ai_1 _6718_ (.B1(_2598_),
    .Y(_2599_),
    .A1(_2571_),
    .A2(_2582_));
 sg13g2_nor3_1 _6719_ (.A(\main.demo.zic._q_drum_inc[0] ),
    .B(\main.demo.zic._q_drum_inc[1] ),
    .C(\main.demo.zic._q_drum_inc[2] ),
    .Y(_2600_));
 sg13g2_a21oi_1 _6720_ (.A1(_2960_),
    .A2(_2600_),
    .Y(_2601_),
    .B1(_2545_));
 sg13g2_a21oi_1 _6721_ (.A1(_2958_),
    .A2(_2601_),
    .Y(_2602_),
    .B1(net415));
 sg13g2_a22oi_1 _6722_ (.Y(_0124_),
    .B1(_2599_),
    .B2(_2602_),
    .A2(net415),
    .A1(_2958_));
 sg13g2_xnor2_1 _6723_ (.Y(_2603_),
    .A(\main.demo.zic._q_drum_inc[0] ),
    .B(net614));
 sg13g2_a21oi_1 _6724_ (.A1(_2601_),
    .A2(_2603_),
    .Y(_2604_),
    .B1(net415));
 sg13g2_a22oi_1 _6725_ (.Y(_0125_),
    .B1(_2599_),
    .B2(_2604_),
    .A2(net415),
    .A1(_2959_));
 sg13g2_o21ai_1 _6726_ (.B1(\main.demo.zic._q_drum_inc[2] ),
    .Y(_2605_),
    .A1(\main.demo.zic._q_drum_inc[0] ),
    .A2(net657));
 sg13g2_nand2b_1 _6727_ (.Y(_2606_),
    .B(_2605_),
    .A_N(_2600_));
 sg13g2_a21oi_1 _6728_ (.A1(_2601_),
    .A2(_2606_),
    .Y(_2607_),
    .B1(net415));
 sg13g2_a22oi_1 _6729_ (.Y(_0126_),
    .B1(_2599_),
    .B2(_2607_),
    .A2(net415),
    .A1(_2961_));
 sg13g2_nor3_1 _6730_ (.A(_2960_),
    .B(_2545_),
    .C(_2600_),
    .Y(_2608_));
 sg13g2_nor2_1 _6731_ (.A(net415),
    .B(_2608_),
    .Y(_2609_));
 sg13g2_a22oi_1 _6732_ (.Y(_0127_),
    .B1(_2599_),
    .B2(_2609_),
    .A2(net415),
    .A1(_2960_));
 sg13g2_and2_1 _6733_ (.A(net317),
    .B(net423),
    .X(_0128_));
 sg13g2_and2_1 _6734_ (.A(net319),
    .B(net423),
    .X(_0129_));
 sg13g2_and2_1 _6735_ (.A(net321),
    .B(net423),
    .X(_0130_));
 sg13g2_and2_1 _6736_ (.A(net351),
    .B(net422),
    .X(_0131_));
 sg13g2_and2_1 _6737_ (.A(net331),
    .B(net422),
    .X(_0132_));
 sg13g2_and2_1 _6738_ (.A(net307),
    .B(net423),
    .X(_0133_));
 sg13g2_and2_1 _6739_ (.A(net325),
    .B(net422),
    .X(_0134_));
 sg13g2_and2_1 _6740_ (.A(net356),
    .B(net422),
    .X(_0135_));
 sg13g2_and2_1 _6741_ (.A(net521),
    .B(net422),
    .X(_0136_));
 sg13g2_and2_1 _6742_ (.A(net520),
    .B(net422),
    .X(_0137_));
 sg13g2_and2_1 _6743_ (.A(net337),
    .B(net422),
    .X(_0138_));
 sg13g2_nor2_1 _6744_ (.A(net456),
    .B(net420),
    .Y(_0139_));
 sg13g2_nand4_1 _6745_ (.B(\main.demo.vga._q_ycount[4] ),
    .C(\main.demo.vga._d_vblank ),
    .A(_2907_),
    .Y(_2610_),
    .D(_0236_));
 sg13g2_nor3_1 _6746_ (.A(\main.demo.vga._q_ycount[0] ),
    .B(_2409_),
    .C(_2610_),
    .Y(_2611_));
 sg13g2_a21oi_1 _6747_ (.A1(net301),
    .A2(_2611_),
    .Y(_2612_),
    .B1(net291));
 sg13g2_nor4_1 _6748_ (.A(net301),
    .B(_2908_),
    .C(_2409_),
    .D(_2610_),
    .Y(_2613_));
 sg13g2_nor3_1 _6749_ (.A(net298),
    .B(net302),
    .C(_2613_),
    .Y(_0140_));
 sg13g2_nand4_1 _6750_ (.B(\main.demo.vga._q_xcount[9] ),
    .C(\main.demo.vga._q_xcount[8] ),
    .A(\main.demo.vga._q_xcount[6] ),
    .Y(_2614_),
    .D(\main.demo.vga._q_xcount[10] ));
 sg13g2_nor2_1 _6751_ (.A(_2402_),
    .B(_2614_),
    .Y(_2615_));
 sg13g2_a21oi_1 _6752_ (.A1(_3324_),
    .A2(_2615_),
    .Y(_2616_),
    .B1(net279));
 sg13g2_nor4_1 _6753_ (.A(\main.demo.vga._q_xcount[7] ),
    .B(_3327_),
    .C(_2405_),
    .D(_2614_),
    .Y(_2617_));
 sg13g2_nor3_1 _6754_ (.A(net298),
    .B(_2616_),
    .C(_2617_),
    .Y(_0141_));
 sg13g2_nor2_1 _6755_ (.A(net456),
    .B(_0235_),
    .Y(_0142_));
 sg13g2_nor2_1 _6756_ (.A(net458),
    .B(net317),
    .Y(_0143_));
 sg13g2_a21oi_1 _6757_ (.A1(net647),
    .A2(_2401_),
    .Y(_2618_),
    .B1(net307));
 sg13g2_nor2_1 _6758_ (.A(_2406_),
    .B(_2618_),
    .Y(_2619_));
 sg13g2_o21ai_1 _6759_ (.B1(net507),
    .Y(_2620_),
    .A1(net428),
    .A2(_2619_));
 sg13g2_inv_1 _6760_ (.Y(_0144_),
    .A(_2620_));
 sg13g2_xor2_1 _6761_ (.B(_2406_),
    .A(net325),
    .X(_2621_));
 sg13g2_o21ai_1 _6762_ (.B1(net507),
    .Y(_2622_),
    .A1(net428),
    .A2(_2621_));
 sg13g2_inv_1 _6763_ (.Y(_0145_),
    .A(_2622_));
 sg13g2_and2_1 _6764_ (.A(net521),
    .B(_2407_),
    .X(_2623_));
 sg13g2_xor2_1 _6765_ (.B(_2407_),
    .A(net521),
    .X(_2624_));
 sg13g2_o21ai_1 _6766_ (.B1(net510),
    .Y(_2625_),
    .A1(net428),
    .A2(_2624_));
 sg13g2_inv_1 _6767_ (.Y(_0146_),
    .A(_2625_));
 sg13g2_nand2_1 _6768_ (.Y(_2626_),
    .A(net520),
    .B(_2623_));
 sg13g2_o21ai_1 _6769_ (.B1(net506),
    .Y(_2627_),
    .A1(net520),
    .A2(_2623_));
 sg13g2_nor2b_1 _6770_ (.A(_2627_),
    .B_N(_2626_),
    .Y(_0147_));
 sg13g2_or2_1 _6771_ (.X(_2628_),
    .B(_2626_),
    .A(net337));
 sg13g2_a21oi_1 _6772_ (.A1(net337),
    .A2(_2626_),
    .Y(_2629_),
    .B1(net428));
 sg13g2_a21oi_1 _6773_ (.A1(_2628_),
    .A2(_2629_),
    .Y(_0148_),
    .B1(net456));
 sg13g2_nand2_1 _6774_ (.Y(_2630_),
    .A(net506),
    .B(_2416_));
 sg13g2_xnor2_1 _6775_ (.Y(_2631_),
    .A(net524),
    .B(net428));
 sg13g2_nor2_1 _6776_ (.A(_2630_),
    .B(_2631_),
    .Y(_0149_));
 sg13g2_a21oi_1 _6777_ (.A1(net524),
    .A2(net428),
    .Y(_2632_),
    .B1(net301));
 sg13g2_nor3_1 _6778_ (.A(net456),
    .B(_2411_),
    .C(_2632_),
    .Y(_0150_));
 sg13g2_xor2_1 _6779_ (.B(_2410_),
    .A(net600),
    .X(_2633_));
 sg13g2_a21oi_1 _6780_ (.A1(_2416_),
    .A2(_2633_),
    .Y(_0151_),
    .B1(net456));
 sg13g2_a21oi_1 _6781_ (.A1(\main.demo.vga._q_ycount[2] ),
    .A2(_2411_),
    .Y(_2634_),
    .B1(net364));
 sg13g2_nor3_1 _6782_ (.A(net456),
    .B(_2412_),
    .C(net365),
    .Y(_0152_));
 sg13g2_xnor2_1 _6783_ (.Y(_2635_),
    .A(net354),
    .B(_2412_));
 sg13g2_a21oi_1 _6784_ (.A1(_2416_),
    .A2(_2635_),
    .Y(_0153_),
    .B1(net456));
 sg13g2_a21oi_1 _6785_ (.A1(net354),
    .A2(_2412_),
    .Y(_2636_),
    .B1(net334));
 sg13g2_nor3_1 _6786_ (.A(_2413_),
    .B(_2630_),
    .C(_2636_),
    .Y(_0154_));
 sg13g2_and2_1 _6787_ (.A(net316),
    .B(_2413_),
    .X(_2637_));
 sg13g2_o21ai_1 _6788_ (.B1(net507),
    .Y(_2638_),
    .A1(net316),
    .A2(_2413_));
 sg13g2_nor2_1 _6789_ (.A(_2637_),
    .B(net572),
    .Y(_0155_));
 sg13g2_o21ai_1 _6790_ (.B1(net507),
    .Y(_2639_),
    .A1(net360),
    .A2(_2637_));
 sg13g2_a21oi_1 _6791_ (.A1(net360),
    .A2(_2637_),
    .Y(_0156_),
    .B1(_2639_));
 sg13g2_a21o_1 _6792_ (.A2(_2637_),
    .A1(net360),
    .B1(net320),
    .X(_2640_));
 sg13g2_and3_1 _6793_ (.X(_0157_),
    .A(net507),
    .B(_2414_),
    .C(_2640_));
 sg13g2_nor2_1 _6794_ (.A(net458),
    .B(_1737_),
    .Y(_0158_));
 sg13g2_or2_2 _6795_ (.X(_2641_),
    .B(_1737_),
    .A(net298));
 sg13g2_nor2_1 _6796_ (.A(_2967_),
    .B(net411),
    .Y(_0159_));
 sg13g2_and2_1 _6797_ (.A(net609),
    .B(\main.demo.zic._q_clock_count[0] ),
    .X(_2642_));
 sg13g2_nor3_1 _6798_ (.A(_2548_),
    .B(net411),
    .C(net610),
    .Y(_0160_));
 sg13g2_and2_1 _6799_ (.A(net530),
    .B(_2642_),
    .X(_2643_));
 sg13g2_nor2_1 _6800_ (.A(net530),
    .B(_2642_),
    .Y(_2644_));
 sg13g2_nor3_1 _6801_ (.A(net411),
    .B(_2643_),
    .C(net531),
    .Y(_0161_));
 sg13g2_and2_1 _6802_ (.A(net339),
    .B(_2643_),
    .X(_2645_));
 sg13g2_nor2_1 _6803_ (.A(net339),
    .B(_2643_),
    .Y(_2646_));
 sg13g2_nor3_1 _6804_ (.A(net411),
    .B(_2645_),
    .C(net340),
    .Y(_0162_));
 sg13g2_and2_1 _6805_ (.A(net540),
    .B(_2645_),
    .X(_2647_));
 sg13g2_nor2_1 _6806_ (.A(net540),
    .B(_2645_),
    .Y(_2648_));
 sg13g2_nor3_1 _6807_ (.A(net411),
    .B(_2647_),
    .C(_2648_),
    .Y(_0163_));
 sg13g2_and2_1 _6808_ (.A(net335),
    .B(_2647_),
    .X(_2649_));
 sg13g2_nor2_1 _6809_ (.A(net335),
    .B(_2647_),
    .Y(_2650_));
 sg13g2_nor3_1 _6810_ (.A(_2641_),
    .B(_2649_),
    .C(net336),
    .Y(_0164_));
 sg13g2_xnor2_1 _6811_ (.Y(_2651_),
    .A(net511),
    .B(_2649_));
 sg13g2_nor2_1 _6812_ (.A(net411),
    .B(_2651_),
    .Y(_0165_));
 sg13g2_nor2b_1 _6813_ (.A(net311),
    .B_N(_2649_),
    .Y(_2652_));
 sg13g2_xnor2_1 _6814_ (.Y(_2653_),
    .A(net367),
    .B(_2652_));
 sg13g2_nor2_1 _6815_ (.A(net411),
    .B(_2653_),
    .Y(_0166_));
 sg13g2_nand3_1 _6816_ (.B(\main.demo.zic._q_clock_count[6] ),
    .C(_2649_),
    .A(net367),
    .Y(_2654_));
 sg13g2_xor2_1 _6817_ (.B(_2654_),
    .A(net370),
    .X(_2655_));
 sg13g2_nor2_1 _6818_ (.A(net411),
    .B(net371),
    .Y(_0167_));
 sg13g2_nand2b_2 _6819_ (.Y(_2656_),
    .B(net433),
    .A_N(_2641_));
 sg13g2_nand2_1 _6820_ (.Y(_2657_),
    .A(\main.demo.zic._q_rythm_count[0] ),
    .B(_2551_));
 sg13g2_nand2_1 _6821_ (.Y(_2658_),
    .A(net289),
    .B(net429));
 sg13g2_a21oi_1 _6822_ (.A1(_2657_),
    .A2(_2658_),
    .Y(_0168_),
    .B1(net410));
 sg13g2_a21oi_1 _6823_ (.A1(\main.demo.zic._q_rythm_count[0] ),
    .A2(net429),
    .Y(_2659_),
    .B1(net326));
 sg13g2_and3_1 _6824_ (.X(_2660_),
    .A(net326),
    .B(\main.demo.zic._q_rythm_count[0] ),
    .C(net429));
 sg13g2_nor3_1 _6825_ (.A(net410),
    .B(net327),
    .C(_2660_),
    .Y(_0169_));
 sg13g2_and4_1 _6826_ (.A(net516),
    .B(net326),
    .C(\main.demo.zic._q_rythm_count[0] ),
    .D(net429),
    .X(_2661_));
 sg13g2_nor2_1 _6827_ (.A(net516),
    .B(_2660_),
    .Y(_2662_));
 sg13g2_and2_1 _6828_ (.A(net516),
    .B(_2660_),
    .X(_2663_));
 sg13g2_nor3_1 _6829_ (.A(net410),
    .B(net517),
    .C(_2663_),
    .Y(_0170_));
 sg13g2_nor2_1 _6830_ (.A(net518),
    .B(_2661_),
    .Y(_2664_));
 sg13g2_and2_1 _6831_ (.A(net518),
    .B(_2663_),
    .X(_2665_));
 sg13g2_nor3_1 _6832_ (.A(net410),
    .B(net519),
    .C(_2665_),
    .Y(_0171_));
 sg13g2_and3_1 _6833_ (.X(_2666_),
    .A(net344),
    .B(\main.demo.zic._q_rythm_count[3] ),
    .C(_2661_));
 sg13g2_nor2_1 _6834_ (.A(net344),
    .B(_2665_),
    .Y(_2667_));
 sg13g2_nor3_1 _6835_ (.A(net410),
    .B(_2666_),
    .C(net345),
    .Y(_0172_));
 sg13g2_nor2_1 _6836_ (.A(net512),
    .B(_2666_),
    .Y(_2668_));
 sg13g2_and3_1 _6837_ (.X(_2669_),
    .A(net512),
    .B(net344),
    .C(_2665_));
 sg13g2_nor3_1 _6838_ (.A(net409),
    .B(net513),
    .C(_2669_),
    .Y(_0173_));
 sg13g2_nor2_1 _6839_ (.A(net341),
    .B(_2669_),
    .Y(_2670_));
 sg13g2_and3_1 _6840_ (.X(_2671_),
    .A(net341),
    .B(\main.demo.zic._q_rythm_count[5] ),
    .C(_2666_));
 sg13g2_nor3_1 _6841_ (.A(net409),
    .B(net342),
    .C(_2671_),
    .Y(_0174_));
 sg13g2_and2_1 _6842_ (.A(net368),
    .B(_2671_),
    .X(_2672_));
 sg13g2_nor2_1 _6843_ (.A(net368),
    .B(_2671_),
    .Y(_2673_));
 sg13g2_nor3_1 _6844_ (.A(net409),
    .B(_2672_),
    .C(net369),
    .Y(_0175_));
 sg13g2_and2_1 _6845_ (.A(net526),
    .B(_2672_),
    .X(_2674_));
 sg13g2_nor2_1 _6846_ (.A(net526),
    .B(_2672_),
    .Y(_2675_));
 sg13g2_nor3_1 _6847_ (.A(net409),
    .B(_2674_),
    .C(_2675_),
    .Y(_0176_));
 sg13g2_nor2_1 _6848_ (.A(net543),
    .B(_2674_),
    .Y(_2676_));
 sg13g2_and2_1 _6849_ (.A(net543),
    .B(_2674_),
    .X(_2677_));
 sg13g2_nor3_1 _6850_ (.A(net409),
    .B(_2676_),
    .C(_2677_),
    .Y(_0177_));
 sg13g2_nor2_1 _6851_ (.A(net347),
    .B(_2677_),
    .Y(_2678_));
 sg13g2_and2_1 _6852_ (.A(net347),
    .B(_2677_),
    .X(_2679_));
 sg13g2_nor3_1 _6853_ (.A(net409),
    .B(net348),
    .C(_2679_),
    .Y(_0178_));
 sg13g2_nor2_1 _6854_ (.A(net357),
    .B(_2679_),
    .Y(_2680_));
 sg13g2_and2_1 _6855_ (.A(net357),
    .B(_2679_),
    .X(_2681_));
 sg13g2_nor3_1 _6856_ (.A(net409),
    .B(_2680_),
    .C(_2681_),
    .Y(_0179_));
 sg13g2_a21oi_1 _6857_ (.A1(net378),
    .A2(_2681_),
    .Y(_2682_),
    .B1(net409));
 sg13g2_o21ai_1 _6858_ (.B1(_2682_),
    .Y(_2683_),
    .A1(net378),
    .A2(_2681_));
 sg13g2_inv_1 _6859_ (.Y(_0180_),
    .A(_2683_));
 sg13g2_and2_1 _6860_ (.A(net504),
    .B(_2580_),
    .X(_0181_));
 sg13g2_nor2_1 _6861_ (.A(net454),
    .B(_2592_),
    .Y(_0182_));
 sg13g2_nor2_1 _6862_ (.A(net454),
    .B(_2577_),
    .Y(_0183_));
 sg13g2_and2_1 _6863_ (.A(net504),
    .B(_2579_),
    .X(_0184_));
 sg13g2_nor2_1 _6864_ (.A(net454),
    .B(_2575_),
    .Y(_0185_));
 sg13g2_and2_1 _6865_ (.A(net504),
    .B(_2570_),
    .X(_0186_));
 sg13g2_nor2_1 _6866_ (.A(net454),
    .B(net633),
    .Y(_0187_));
 sg13g2_nor2_1 _6867_ (.A(_2908_),
    .B(net420),
    .Y(_0188_));
 sg13g2_nor2b_1 _6868_ (.A(net420),
    .B_N(net301),
    .Y(_0189_));
 sg13g2_nor2b_1 _6869_ (.A(net420),
    .B_N(net600),
    .Y(_0190_));
 sg13g2_nor2b_1 _6870_ (.A(net420),
    .B_N(net364),
    .Y(_0191_));
 sg13g2_nor2b_1 _6871_ (.A(net420),
    .B_N(net354),
    .Y(_0192_));
 sg13g2_nor2_1 _6872_ (.A(_2907_),
    .B(net421),
    .Y(_0193_));
 sg13g2_nor2b_1 _6873_ (.A(net421),
    .B_N(net316),
    .Y(_0194_));
 sg13g2_and3_1 _6874_ (.X(_0195_),
    .A(\main.demo.vga._q_ycount[7] ),
    .B(net314),
    .C(_0240_));
 sg13g2_nor2b_1 _6875_ (.A(net420),
    .B_N(net320),
    .Y(_0196_));
 sg13g2_nor2b_1 _6876_ (.A(net420),
    .B_N(net372),
    .Y(_0197_));
 sg13g2_nand3b_1 _6877_ (.B(_2557_),
    .C(_2580_),
    .Y(_2684_),
    .A_N(\main.demo.zic._q_idx[1] ));
 sg13g2_nand2_1 _6878_ (.Y(_2685_),
    .A(_2594_),
    .B(_2684_));
 sg13g2_nand3_1 _6879_ (.B(_2588_),
    .C(_2685_),
    .A(_2575_),
    .Y(_2686_));
 sg13g2_nand3_1 _6880_ (.B(_2571_),
    .C(_2686_),
    .A(_2545_),
    .Y(_2687_));
 sg13g2_nand2_1 _6881_ (.Y(_2688_),
    .A(_2904_),
    .B(_2905_));
 sg13g2_nor2_1 _6882_ (.A(net385),
    .B(_2688_),
    .Y(_2689_));
 sg13g2_nor3_1 _6883_ (.A(\main.demo.zic._q_squ_env[3] ),
    .B(\main.demo.zic._q_squ_env[2] ),
    .C(_2688_),
    .Y(_2690_));
 sg13g2_nor2b_1 _6884_ (.A(\main.demo.zic._q_squ_env[4] ),
    .B_N(_2690_),
    .Y(_2691_));
 sg13g2_a21oi_1 _6885_ (.A1(_1722_),
    .A2(_2689_),
    .Y(_2692_),
    .B1(_2545_));
 sg13g2_a21oi_1 _6886_ (.A1(_2905_),
    .A2(_2692_),
    .Y(_2693_),
    .B1(net416));
 sg13g2_a221oi_1 _6887_ (.B2(_2693_),
    .C1(net455),
    .B1(_2687_),
    .A1(_2905_),
    .Y(_0198_),
    .A2(net416));
 sg13g2_xnor2_1 _6888_ (.Y(_2694_),
    .A(net522),
    .B(\main.demo.zic._q_squ_env[0] ));
 sg13g2_a21oi_1 _6889_ (.A1(_2692_),
    .A2(_2694_),
    .Y(_2695_),
    .B1(net416));
 sg13g2_a221oi_1 _6890_ (.B2(_2695_),
    .C1(net455),
    .B1(_2687_),
    .A1(_2904_),
    .Y(_0199_),
    .A2(net416));
 sg13g2_nor2b_2 _6891_ (.A(_2554_),
    .B_N(_2692_),
    .Y(_2696_));
 sg13g2_a21o_1 _6892_ (.A2(_2696_),
    .A1(_2688_),
    .B1(net416),
    .X(_2697_));
 sg13g2_a22oi_1 _6893_ (.Y(_2698_),
    .B1(_2697_),
    .B2(net385),
    .A2(_2696_),
    .A1(_2689_));
 sg13g2_a21oi_1 _6894_ (.A1(_2687_),
    .A2(_2698_),
    .Y(_0200_),
    .B1(net455));
 sg13g2_xor2_1 _6895_ (.B(_2689_),
    .A(\main.demo.zic._q_squ_env[3] ),
    .X(_2699_));
 sg13g2_a22oi_1 _6896_ (.Y(_2700_),
    .B1(_2696_),
    .B2(_2699_),
    .A2(net416),
    .A1(net630));
 sg13g2_a21oi_1 _6897_ (.A1(_2687_),
    .A2(_2700_),
    .Y(_0201_),
    .B1(net455));
 sg13g2_xnor2_1 _6898_ (.Y(_2701_),
    .A(net589),
    .B(_2690_));
 sg13g2_a22oi_1 _6899_ (.Y(_2702_),
    .B1(_2696_),
    .B2(net590),
    .A2(net416),
    .A1(\main.demo.zic._q_squ_env[4] ));
 sg13g2_a21oi_1 _6900_ (.A1(_2687_),
    .A2(net591),
    .Y(_0202_),
    .B1(net454));
 sg13g2_xnor2_1 _6901_ (.Y(_2703_),
    .A(_0024_),
    .B(_2691_));
 sg13g2_a22oi_1 _6902_ (.Y(_2704_),
    .B1(_2696_),
    .B2(_2703_),
    .A2(net416),
    .A1(net569));
 sg13g2_a21oi_1 _6903_ (.A1(_2687_),
    .A2(net570),
    .Y(_0203_),
    .B1(net454));
 sg13g2_nand2_1 _6904_ (.Y(_2705_),
    .A(_0032_),
    .B(\main.demo.zic._q_idx[4] ));
 sg13g2_nand2b_2 _6905_ (.Y(_2706_),
    .B(\main.demo.zic._q_idx[1] ),
    .A_N(\main.demo.zic._q_idx[0] ));
 sg13g2_nor2_2 _6906_ (.A(_2558_),
    .B(_2706_),
    .Y(_2707_));
 sg13g2_nor2_2 _6907_ (.A(\main.demo.zic._q_idx[1] ),
    .B(\main.demo.zic._q_idx[0] ),
    .Y(_2708_));
 sg13g2_nor2_2 _6908_ (.A(net463),
    .B(net464),
    .Y(_2709_));
 sg13g2_nand2_1 _6909_ (.Y(_2710_),
    .A(_2708_),
    .B(_2709_));
 sg13g2_nor2b_2 _6910_ (.A(\main.demo.zic._q_idx[1] ),
    .B_N(\main.demo.zic._q_idx[0] ),
    .Y(_2711_));
 sg13g2_nand2_1 _6911_ (.Y(_2712_),
    .A(_2583_),
    .B(_2711_));
 sg13g2_nand2_1 _6912_ (.Y(_2713_),
    .A(_2710_),
    .B(_2712_));
 sg13g2_o21ai_1 _6913_ (.B1(_2705_),
    .Y(_2714_),
    .A1(_2707_),
    .A2(_2713_));
 sg13g2_nor2_1 _6914_ (.A(_0032_),
    .B(\main.demo.zic._q_idx[4] ),
    .Y(_2715_));
 sg13g2_nand2_1 _6915_ (.Y(_2716_),
    .A(net464),
    .B(_2711_));
 sg13g2_nor2b_1 _6916_ (.A(net463),
    .B_N(net465),
    .Y(_2717_));
 sg13g2_nor2_1 _6917_ (.A(net463),
    .B(_2716_),
    .Y(_2718_));
 sg13g2_nand2b_1 _6918_ (.Y(_2719_),
    .B(_2718_),
    .A_N(_2715_));
 sg13g2_nand2_2 _6919_ (.Y(_2720_),
    .A(_2714_),
    .B(_2719_));
 sg13g2_nor2_1 _6920_ (.A(net463),
    .B(_2556_),
    .Y(_2721_));
 sg13g2_nor2b_1 _6921_ (.A(_2556_),
    .B_N(_2717_),
    .Y(_2722_));
 sg13g2_nor3_1 _6922_ (.A(_2914_),
    .B(net464),
    .C(_2556_),
    .Y(_2723_));
 sg13g2_nand2_1 _6923_ (.Y(_2724_),
    .A(_2557_),
    .B(_2711_));
 sg13g2_nor2_1 _6924_ (.A(_2722_),
    .B(_2723_),
    .Y(_2725_));
 sg13g2_a22oi_1 _6925_ (.Y(_2726_),
    .B1(_2724_),
    .B2(_2725_),
    .A2(\main.demo.zic._q_idx[4] ),
    .A1(_0032_));
 sg13g2_nand2_1 _6926_ (.Y(_2727_),
    .A(net464),
    .B(_2708_));
 sg13g2_nand2_1 _6927_ (.Y(_2728_),
    .A(_2708_),
    .B(_2717_));
 sg13g2_nor2_1 _6928_ (.A(_2715_),
    .B(_2728_),
    .Y(_2729_));
 sg13g2_nor2_1 _6929_ (.A(net464),
    .B(_2706_),
    .Y(_2730_));
 sg13g2_nor2b_1 _6930_ (.A(_2706_),
    .B_N(_2709_),
    .Y(_2731_));
 sg13g2_nor4_2 _6931_ (.A(_2720_),
    .B(_2726_),
    .C(_2729_),
    .Y(_2732_),
    .D(_2731_));
 sg13g2_nand2_1 _6932_ (.Y(_2733_),
    .A(\main.demo.zic._q_tpos[0] ),
    .B(_2732_));
 sg13g2_xnor2_1 _6933_ (.Y(_2734_),
    .A(net559),
    .B(_2732_));
 sg13g2_or2_1 _6934_ (.X(_2735_),
    .B(_2734_),
    .A(_2958_));
 sg13g2_xnor2_1 _6935_ (.Y(_2736_),
    .A(_2958_),
    .B(_2734_));
 sg13g2_o21ai_1 _6936_ (.B1(net505),
    .Y(_2737_),
    .A1(net559),
    .A2(net431));
 sg13g2_a21oi_1 _6937_ (.A1(net431),
    .A2(_2736_),
    .Y(_0204_),
    .B1(_2737_));
 sg13g2_nand2b_1 _6938_ (.Y(_2738_),
    .B(_2717_),
    .A_N(_2706_));
 sg13g2_a22oi_1 _6939_ (.Y(_2739_),
    .B1(_2560_),
    .B2(_2738_),
    .A2(net462),
    .A1(_0032_));
 sg13g2_nor2_2 _6940_ (.A(_2720_),
    .B(_2739_),
    .Y(_2740_));
 sg13g2_and3_1 _6941_ (.X(_2741_),
    .A(_2557_),
    .B(_2705_),
    .C(_2708_));
 sg13g2_nand2_1 _6942_ (.Y(_2742_),
    .A(_2583_),
    .B(_2708_));
 sg13g2_nand2b_1 _6943_ (.Y(_2743_),
    .B(_2709_),
    .A_N(_2556_));
 sg13g2_o21ai_1 _6944_ (.B1(_2743_),
    .Y(_2744_),
    .A1(_2715_),
    .A2(_2742_));
 sg13g2_nor4_2 _6945_ (.A(_2720_),
    .B(_2739_),
    .C(_2741_),
    .Y(_2745_),
    .D(_2744_));
 sg13g2_nand2_1 _6946_ (.Y(_2746_),
    .A(\main.demo.zic._q_tpos[1] ),
    .B(_2745_));
 sg13g2_xnor2_1 _6947_ (.Y(_2747_),
    .A(\main.demo.zic._q_tpos[1] ),
    .B(_2745_));
 sg13g2_xnor2_1 _6948_ (.Y(_2748_),
    .A(_2959_),
    .B(_2747_));
 sg13g2_a21oi_2 _6949_ (.B1(_2748_),
    .Y(_2749_),
    .A2(_2735_),
    .A1(_2733_));
 sg13g2_and3_1 _6950_ (.X(_2750_),
    .A(_2733_),
    .B(_2735_),
    .C(_2748_));
 sg13g2_o21ai_1 _6951_ (.B1(net431),
    .Y(_2751_),
    .A1(_2749_),
    .A2(_2750_));
 sg13g2_o21ai_1 _6952_ (.B1(_2751_),
    .Y(_2752_),
    .A1(net561),
    .A2(net431));
 sg13g2_nor2_1 _6953_ (.A(net454),
    .B(_2752_),
    .Y(_0205_));
 sg13g2_o21ai_1 _6954_ (.B1(_2746_),
    .Y(_2753_),
    .A1(_2959_),
    .A2(_2747_));
 sg13g2_and2_1 _6955_ (.A(\main.demo.zic._q_tpos[2] ),
    .B(_2740_),
    .X(_2754_));
 sg13g2_xor2_1 _6956_ (.B(_2740_),
    .A(\main.demo.zic._q_tpos[2] ),
    .X(_2755_));
 sg13g2_xnor2_1 _6957_ (.Y(_2756_),
    .A(\main.demo.zic._q_drum_inc[2] ),
    .B(_2755_));
 sg13g2_nand2b_1 _6958_ (.Y(_2757_),
    .B(_2753_),
    .A_N(_2756_));
 sg13g2_xnor2_1 _6959_ (.Y(_2758_),
    .A(_2753_),
    .B(_2756_));
 sg13g2_nand2_1 _6960_ (.Y(_2759_),
    .A(_2749_),
    .B(_2758_));
 sg13g2_xnor2_1 _6961_ (.Y(_2760_),
    .A(_2749_),
    .B(_2758_));
 sg13g2_o21ai_1 _6962_ (.B1(net505),
    .Y(_2761_),
    .A1(net552),
    .A2(net431));
 sg13g2_a21oi_1 _6963_ (.A1(net431),
    .A2(_2760_),
    .Y(_0206_),
    .B1(net553));
 sg13g2_a21oi_1 _6964_ (.A1(\main.demo.zic._q_drum_inc[2] ),
    .A2(_2755_),
    .Y(_2762_),
    .B1(_2754_));
 sg13g2_nor2b_1 _6965_ (.A(_2740_),
    .B_N(\main.demo.zic._q_tpos[3] ),
    .Y(_2763_));
 sg13g2_xnor2_1 _6966_ (.Y(_2764_),
    .A(\main.demo.zic._q_tpos[3] ),
    .B(_2740_));
 sg13g2_xnor2_1 _6967_ (.Y(_2765_),
    .A(\main.demo.zic._q_drum_inc[3] ),
    .B(_2764_));
 sg13g2_nor2_1 _6968_ (.A(_2762_),
    .B(_2765_),
    .Y(_2766_));
 sg13g2_xnor2_1 _6969_ (.Y(_2767_),
    .A(_2762_),
    .B(_2765_));
 sg13g2_and3_1 _6970_ (.X(_2768_),
    .A(_2757_),
    .B(_2759_),
    .C(_2767_));
 sg13g2_a21oi_1 _6971_ (.A1(_2757_),
    .A2(_2759_),
    .Y(_2769_),
    .B1(_2767_));
 sg13g2_o21ai_1 _6972_ (.B1(net431),
    .Y(_2770_),
    .A1(_2768_),
    .A2(_2769_));
 sg13g2_o21ai_1 _6973_ (.B1(_2770_),
    .Y(_2771_),
    .A1(net560),
    .A2(net431));
 sg13g2_nor2_1 _6974_ (.A(net455),
    .B(_2771_),
    .Y(_0207_));
 sg13g2_a21oi_1 _6975_ (.A1(\main.demo.zic._q_drum_inc[3] ),
    .A2(_2764_),
    .Y(_2772_),
    .B1(_2763_));
 sg13g2_nand2b_1 _6976_ (.Y(_2773_),
    .B(\main.demo.zic._q_tpos[4] ),
    .A_N(_2772_));
 sg13g2_xnor2_1 _6977_ (.Y(_2774_),
    .A(\main.demo.zic._q_tpos[4] ),
    .B(_2772_));
 sg13g2_or3_1 _6978_ (.A(_2766_),
    .B(_2769_),
    .C(_2774_),
    .X(_2775_));
 sg13g2_o21ai_1 _6979_ (.B1(_2774_),
    .Y(_2776_),
    .A1(_2766_),
    .A2(_2769_));
 sg13g2_a21oi_1 _6980_ (.A1(_2775_),
    .A2(_2776_),
    .Y(_2777_),
    .B1(_2551_));
 sg13g2_o21ai_1 _6981_ (.B1(net505),
    .Y(_2778_),
    .A1(net601),
    .A2(net432));
 sg13g2_nor2_1 _6982_ (.A(_2777_),
    .B(_2778_),
    .Y(_0208_));
 sg13g2_and2_1 _6983_ (.A(_2773_),
    .B(_2776_),
    .X(_2779_));
 sg13g2_nor3_1 _6984_ (.A(net376),
    .B(_2551_),
    .C(_2779_),
    .Y(_2780_));
 sg13g2_nand3_1 _6985_ (.B(net432),
    .C(_2779_),
    .A(net376),
    .Y(_2781_));
 sg13g2_o21ai_1 _6986_ (.B1(_2781_),
    .Y(_2782_),
    .A1(\main.demo.zic._q_tpos[5] ),
    .A2(net432));
 sg13g2_nor3_1 _6987_ (.A(net454),
    .B(_2780_),
    .C(net377),
    .Y(_0209_));
 sg13g2_o21ai_1 _6988_ (.B1(net505),
    .Y(_2783_),
    .A1(net578),
    .A2(_2780_));
 sg13g2_and2_1 _6989_ (.A(net578),
    .B(_2780_),
    .X(_2784_));
 sg13g2_nor2_1 _6990_ (.A(_2783_),
    .B(_2784_),
    .Y(_0210_));
 sg13g2_nor2_1 _6991_ (.A(net532),
    .B(_2784_),
    .Y(_2785_));
 sg13g2_and2_1 _6992_ (.A(net532),
    .B(_2784_),
    .X(_2786_));
 sg13g2_nor3_1 _6993_ (.A(net457),
    .B(net533),
    .C(_2786_),
    .Y(_0211_));
 sg13g2_o21ai_1 _6994_ (.B1(net506),
    .Y(_2787_),
    .A1(net358),
    .A2(_2786_));
 sg13g2_a21oi_1 _6995_ (.A1(net358),
    .A2(_2786_),
    .Y(_0212_),
    .B1(_2787_));
 sg13g2_a21oi_1 _6996_ (.A1(\main.demo.zic._q_tpos[8] ),
    .A2(_2786_),
    .Y(_2788_),
    .B1(net329));
 sg13g2_nand3_1 _6997_ (.B(net358),
    .C(_2786_),
    .A(net329),
    .Y(_2789_));
 sg13g2_inv_1 _6998_ (.Y(_2790_),
    .A(_2789_));
 sg13g2_nor3_1 _6999_ (.A(net457),
    .B(net330),
    .C(_2790_),
    .Y(_0213_));
 sg13g2_o21ai_1 _7000_ (.B1(net506),
    .Y(_2791_),
    .A1(_2903_),
    .A2(_2789_));
 sg13g2_a21oi_1 _7001_ (.A1(_2903_),
    .A2(_2789_),
    .Y(_0214_),
    .B1(_2791_));
 sg13g2_a21oi_1 _7002_ (.A1(net535),
    .A2(_2790_),
    .Y(_2792_),
    .B1(net539));
 sg13g2_o21ai_1 _7003_ (.B1(net506),
    .Y(_2793_),
    .A1(_1739_),
    .A2(_2789_));
 sg13g2_nor2_1 _7004_ (.A(_2792_),
    .B(_2793_),
    .Y(_0215_));
 sg13g2_nand2_1 _7005_ (.Y(_2794_),
    .A(\main.demo.zic._q_idx[5] ),
    .B(_0033_));
 sg13g2_nand3_1 _7006_ (.B(net462),
    .C(_0033_),
    .A(\main.demo.zic._q_idx[5] ),
    .Y(_2795_));
 sg13g2_nand2_1 _7007_ (.Y(_2796_),
    .A(_2738_),
    .B(_2743_));
 sg13g2_a21oi_1 _7008_ (.A1(\main.demo.zic._q_idx[0] ),
    .A2(_2583_),
    .Y(_2797_),
    .B1(_2796_));
 sg13g2_a21oi_1 _7009_ (.A1(_2710_),
    .A2(_2797_),
    .Y(_2798_),
    .B1(_2795_));
 sg13g2_nor2b_1 _7010_ (.A(_2561_),
    .B_N(_2794_),
    .Y(_2799_));
 sg13g2_nor2_1 _7011_ (.A(_2560_),
    .B(_2799_),
    .Y(_2800_));
 sg13g2_nand2b_1 _7012_ (.Y(_2801_),
    .B(_2742_),
    .A_N(_2722_));
 sg13g2_nor2_1 _7013_ (.A(_2730_),
    .B(_2801_),
    .Y(_2802_));
 sg13g2_nor2_1 _7014_ (.A(_2562_),
    .B(_2802_),
    .Y(_2803_));
 sg13g2_nor3_2 _7015_ (.A(_2798_),
    .B(_2800_),
    .C(_2803_),
    .Y(_2804_));
 sg13g2_nor2_1 _7016_ (.A(net462),
    .B(_2794_),
    .Y(_2805_));
 sg13g2_o21ai_1 _7017_ (.B1(_2805_),
    .Y(_2806_),
    .A1(_2713_),
    .A2(_2721_));
 sg13g2_or2_1 _7018_ (.X(_2807_),
    .B(_2710_),
    .A(_2562_));
 sg13g2_nand3_1 _7019_ (.B(_2806_),
    .C(_2807_),
    .A(_2804_),
    .Y(_2808_));
 sg13g2_a21oi_1 _7020_ (.A1(_2557_),
    .A2(_2708_),
    .Y(_2809_),
    .B1(_2718_));
 sg13g2_nor2b_2 _7021_ (.A(net462),
    .B_N(_2561_),
    .Y(_2810_));
 sg13g2_a21oi_1 _7022_ (.A1(_2718_),
    .A2(_2810_),
    .Y(_2811_),
    .B1(_2805_));
 sg13g2_nor2_1 _7023_ (.A(_2809_),
    .B(_2811_),
    .Y(_2812_));
 sg13g2_nand2_2 _7024_ (.Y(_2813_),
    .A(_2709_),
    .B(_2711_));
 sg13g2_nor2_1 _7025_ (.A(_2723_),
    .B(_2731_),
    .Y(_2814_));
 sg13g2_nand3_1 _7026_ (.B(_2813_),
    .C(_2814_),
    .A(_2727_),
    .Y(_2815_));
 sg13g2_o21ai_1 _7027_ (.B1(_2810_),
    .Y(_2816_),
    .A1(_2801_),
    .A2(_2815_));
 sg13g2_inv_1 _7028_ (.Y(_2817_),
    .A(_2816_));
 sg13g2_nor2_2 _7029_ (.A(_2727_),
    .B(_2795_),
    .Y(_2818_));
 sg13g2_nor2_1 _7030_ (.A(_2812_),
    .B(_2818_),
    .Y(_2819_));
 sg13g2_nand2_1 _7031_ (.Y(_2820_),
    .A(_2562_),
    .B(_2794_));
 sg13g2_nor2_1 _7032_ (.A(_2562_),
    .B(_2797_),
    .Y(_2821_));
 sg13g2_a21oi_2 _7033_ (.B1(_2821_),
    .Y(_2822_),
    .A2(_2820_),
    .A1(_2707_));
 sg13g2_nor2_1 _7034_ (.A(_2562_),
    .B(_2809_),
    .Y(_2823_));
 sg13g2_nor2_1 _7035_ (.A(_2716_),
    .B(_2795_),
    .Y(_2824_));
 sg13g2_nor2_1 _7036_ (.A(_2823_),
    .B(_2824_),
    .Y(_2825_));
 sg13g2_nand2_1 _7037_ (.Y(_2826_),
    .A(_2822_),
    .B(_2825_));
 sg13g2_nor4_2 _7038_ (.A(_2812_),
    .B(_2817_),
    .C(_2818_),
    .Y(_2827_),
    .D(_2826_));
 sg13g2_a21oi_1 _7039_ (.A1(_2802_),
    .A2(_2813_),
    .Y(_2828_),
    .B1(_2795_));
 sg13g2_a21oi_1 _7040_ (.A1(_2707_),
    .A2(_2810_),
    .Y(_2829_),
    .B1(_2828_));
 sg13g2_inv_1 _7041_ (.Y(_2830_),
    .A(_2829_));
 sg13g2_o21ai_1 _7042_ (.B1(_2810_),
    .Y(_2831_),
    .A1(_2713_),
    .A2(_2796_));
 sg13g2_nor2_1 _7043_ (.A(_2562_),
    .B(_2813_),
    .Y(_2832_));
 sg13g2_nand4_1 _7044_ (.B(_2742_),
    .C(_2813_),
    .A(_2738_),
    .Y(_2833_),
    .D(_2814_));
 sg13g2_o21ai_1 _7045_ (.B1(_2833_),
    .Y(_2834_),
    .A1(_2805_),
    .A2(_2832_));
 sg13g2_nand2_1 _7046_ (.Y(_2835_),
    .A(_2831_),
    .B(_2834_));
 sg13g2_o21ai_1 _7047_ (.B1(_2716_),
    .Y(_2836_),
    .A1(net464),
    .A2(_2706_));
 sg13g2_nor3_1 _7048_ (.A(_2914_),
    .B(net462),
    .C(_2799_),
    .Y(_2837_));
 sg13g2_nand2_1 _7049_ (.Y(_2838_),
    .A(_2836_),
    .B(_2837_));
 sg13g2_o21ai_1 _7050_ (.B1(_2838_),
    .Y(_2839_),
    .A1(\main.demo.zic._q_idx[5] ),
    .A2(\main.demo.zic._q_idx[6] ));
 sg13g2_a21oi_2 _7051_ (.B1(_2562_),
    .Y(_2840_),
    .A2(_2728_),
    .A1(_2724_));
 sg13g2_nor3_1 _7052_ (.A(_2835_),
    .B(_2839_),
    .C(_2840_),
    .Y(_2841_));
 sg13g2_nor2_1 _7053_ (.A(_2830_),
    .B(_2835_),
    .Y(_2842_));
 sg13g2_nand3_1 _7054_ (.B(_2829_),
    .C(_2841_),
    .A(_2827_),
    .Y(_2843_));
 sg13g2_nor3_1 _7055_ (.A(_2812_),
    .B(_2826_),
    .C(_2835_),
    .Y(_2844_));
 sg13g2_o21ai_1 _7056_ (.B1(_2844_),
    .Y(_2845_),
    .A1(_2808_),
    .A2(_2843_));
 sg13g2_a21oi_1 _7057_ (.A1(net429),
    .A2(_2845_),
    .Y(_2846_),
    .B1(net300));
 sg13g2_nand2_1 _7058_ (.Y(_2847_),
    .A(net300),
    .B(_2845_));
 sg13g2_o21ai_1 _7059_ (.B1(net504),
    .Y(_2848_),
    .A1(_2551_),
    .A2(_2847_));
 sg13g2_nor2_1 _7060_ (.A(_2846_),
    .B(_2848_),
    .Y(_0216_));
 sg13g2_a21oi_1 _7061_ (.A1(_2804_),
    .A2(_2827_),
    .Y(_2849_),
    .B1(_0028_));
 sg13g2_nand3_1 _7062_ (.B(_2804_),
    .C(_2827_),
    .A(_0028_),
    .Y(_2850_));
 sg13g2_nand2b_1 _7063_ (.Y(_2851_),
    .B(_2850_),
    .A_N(_2849_));
 sg13g2_nor2_1 _7064_ (.A(_2847_),
    .B(_2851_),
    .Y(_2852_));
 sg13g2_xnor2_1 _7065_ (.Y(_2853_),
    .A(_2847_),
    .B(_2851_));
 sg13g2_o21ai_1 _7066_ (.B1(net504),
    .Y(_2854_),
    .A1(net332),
    .A2(net430));
 sg13g2_a21oi_1 _7067_ (.A1(net429),
    .A2(_2853_),
    .Y(_0217_),
    .B1(_2854_));
 sg13g2_nor3_2 _7068_ (.A(_2818_),
    .B(_2830_),
    .C(_2840_),
    .Y(_2855_));
 sg13g2_nand2b_1 _7069_ (.Y(_2856_),
    .B(_2810_),
    .A_N(_2727_));
 sg13g2_nand4_1 _7070_ (.B(_2825_),
    .C(_2855_),
    .A(_2804_),
    .Y(_2857_),
    .D(_2856_));
 sg13g2_nand2_1 _7071_ (.Y(_2858_),
    .A(\main.demo.zic._q_qpos[2] ),
    .B(_2857_));
 sg13g2_xor2_1 _7072_ (.B(_2857_),
    .A(\main.demo.zic._q_qpos[2] ),
    .X(_2859_));
 sg13g2_or3_1 _7073_ (.A(_2849_),
    .B(_2852_),
    .C(_2859_),
    .X(_2860_));
 sg13g2_o21ai_1 _7074_ (.B1(_2859_),
    .Y(_2861_),
    .A1(_2849_),
    .A2(_2852_));
 sg13g2_a21oi_1 _7075_ (.A1(_2860_),
    .A2(_2861_),
    .Y(_2862_),
    .B1(_2551_));
 sg13g2_o21ai_1 _7076_ (.B1(net504),
    .Y(_2863_),
    .A1(net541),
    .A2(net429));
 sg13g2_nor2_1 _7077_ (.A(_2862_),
    .B(_2863_),
    .Y(_0218_));
 sg13g2_a21oi_1 _7078_ (.A1(_2822_),
    .A2(_2855_),
    .Y(_2864_),
    .B1(_0029_));
 sg13g2_nand3_1 _7079_ (.B(_2822_),
    .C(_2855_),
    .A(_0029_),
    .Y(_2865_));
 sg13g2_nand2b_1 _7080_ (.Y(_2866_),
    .B(_2865_),
    .A_N(_2864_));
 sg13g2_and3_1 _7081_ (.X(_2867_),
    .A(_2858_),
    .B(_2861_),
    .C(_2866_));
 sg13g2_a21oi_1 _7082_ (.A1(_2858_),
    .A2(_2861_),
    .Y(_2868_),
    .B1(_2866_));
 sg13g2_o21ai_1 _7083_ (.B1(_2550_),
    .Y(_2869_),
    .A1(_2867_),
    .A2(_2868_));
 sg13g2_o21ai_1 _7084_ (.B1(net507),
    .Y(_2870_),
    .A1(net352),
    .A2(net430));
 sg13g2_nor2b_1 _7085_ (.A(net353),
    .B_N(_2869_),
    .Y(_0219_));
 sg13g2_nand2_1 _7086_ (.Y(_2871_),
    .A(_2825_),
    .B(_2843_));
 sg13g2_nand2_1 _7087_ (.Y(_2872_),
    .A(\main.demo.zic._q_qpos[4] ),
    .B(_2871_));
 sg13g2_xor2_1 _7088_ (.B(_2871_),
    .A(\main.demo.zic._q_qpos[4] ),
    .X(_2873_));
 sg13g2_or3_1 _7089_ (.A(_2864_),
    .B(_2868_),
    .C(_2873_),
    .X(_2874_));
 sg13g2_o21ai_1 _7090_ (.B1(_2873_),
    .Y(_2875_),
    .A1(_2864_),
    .A2(_2868_));
 sg13g2_a21oi_1 _7091_ (.A1(_2874_),
    .A2(_2875_),
    .Y(_2876_),
    .B1(_2551_));
 sg13g2_o21ai_1 _7092_ (.B1(net505),
    .Y(_2877_),
    .A1(net549),
    .A2(net430));
 sg13g2_nor2_1 _7093_ (.A(_2876_),
    .B(net550),
    .Y(_0220_));
 sg13g2_nand2_1 _7094_ (.Y(_2878_),
    .A(_2819_),
    .B(_2842_));
 sg13g2_xnor2_1 _7095_ (.Y(_2879_),
    .A(_2962_),
    .B(_2878_));
 sg13g2_and3_1 _7096_ (.X(_2880_),
    .A(_2872_),
    .B(_2875_),
    .C(_2879_));
 sg13g2_a21oi_1 _7097_ (.A1(_2872_),
    .A2(_2875_),
    .Y(_2881_),
    .B1(_2879_));
 sg13g2_o21ai_1 _7098_ (.B1(net430),
    .Y(_2882_),
    .A1(_2880_),
    .A2(_2881_));
 sg13g2_o21ai_1 _7099_ (.B1(net507),
    .Y(_2883_),
    .A1(net349),
    .A2(net430));
 sg13g2_nor2b_1 _7100_ (.A(net350),
    .B_N(_2882_),
    .Y(_0221_));
 sg13g2_xor2_1 _7101_ (.B(_2816_),
    .A(net556),
    .X(_2884_));
 sg13g2_a21oi_1 _7102_ (.A1(_2962_),
    .A2(_2878_),
    .Y(_2885_),
    .B1(_2881_));
 sg13g2_nor2_1 _7103_ (.A(_2884_),
    .B(_2885_),
    .Y(_2886_));
 sg13g2_xnor2_1 _7104_ (.Y(_2887_),
    .A(_2884_),
    .B(_2885_));
 sg13g2_o21ai_1 _7105_ (.B1(net504),
    .Y(_2888_),
    .A1(net556),
    .A2(net430));
 sg13g2_a21oi_1 _7106_ (.A1(net430),
    .A2(_2887_),
    .Y(_0222_),
    .B1(_2888_));
 sg13g2_a21oi_1 _7107_ (.A1(\main.demo.zic._q_qpos[6] ),
    .A2(_2817_),
    .Y(_2889_),
    .B1(_2886_));
 sg13g2_nor3_2 _7108_ (.A(_0031_),
    .B(_2551_),
    .C(_2889_),
    .Y(_2890_));
 sg13g2_and3_1 _7109_ (.X(_2891_),
    .A(_0031_),
    .B(net432),
    .C(_2889_));
 sg13g2_o21ai_1 _7110_ (.B1(net504),
    .Y(_2892_),
    .A1(net362),
    .A2(net432));
 sg13g2_nor3_1 _7111_ (.A(_2890_),
    .B(_2891_),
    .C(_2892_),
    .Y(_0223_));
 sg13g2_and2_1 _7112_ (.A(net373),
    .B(_2890_),
    .X(_2893_));
 sg13g2_o21ai_1 _7113_ (.B1(net505),
    .Y(_2894_),
    .A1(net373),
    .A2(_2890_));
 sg13g2_nor2_1 _7114_ (.A(_2893_),
    .B(net374),
    .Y(_0224_));
 sg13g2_nand2_1 _7115_ (.Y(_2895_),
    .A(net528),
    .B(_2893_));
 sg13g2_o21ai_1 _7116_ (.B1(net506),
    .Y(_2896_),
    .A1(net528),
    .A2(_2893_));
 sg13g2_nor2b_1 _7117_ (.A(net529),
    .B_N(_2895_),
    .Y(_0225_));
 sg13g2_nand2b_1 _7118_ (.Y(_2897_),
    .B(_2895_),
    .A_N(net576));
 sg13g2_nand3_1 _7119_ (.B(net528),
    .C(_2893_),
    .A(net576),
    .Y(_2898_));
 sg13g2_and3_1 _7120_ (.X(_0226_),
    .A(net506),
    .B(_2897_),
    .C(_2898_));
 sg13g2_and2_1 _7121_ (.A(_2902_),
    .B(_2898_),
    .X(_2899_));
 sg13g2_nor2_1 _7122_ (.A(_2902_),
    .B(_2898_),
    .Y(_2900_));
 sg13g2_nor3_1 _7123_ (.A(net457),
    .B(net565),
    .C(_2900_),
    .Y(_0227_));
 sg13g2_o21ai_1 _7124_ (.B1(net505),
    .Y(_2901_),
    .A1(net582),
    .A2(_2900_));
 sg13g2_a21oi_1 _7125_ (.A1(net582),
    .A2(_2900_),
    .Y(_0228_),
    .B1(_2901_));
 sg13g2_xor2_1 _7126_ (.B(_0419_),
    .A(_0362_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[4] ));
 sg13g2_dfrbp_1 _7127_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net18),
    .D(net1),
    .Q_N(_0002_),
    .Q(rst_n_q));
 sg13g2_dfrbp_1 _7128_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net25),
    .D(net400),
    .Q_N(_3449_),
    .Q(_0067_));
 sg13g2_dfrbp_1 _7129_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net17),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .Q_N(_3448_),
    .Q(_0068_));
 sg13g2_dfrbp_1 _7130_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net227),
    .D(_0069_),
    .Q_N(_3447_),
    .Q(\main.demo.vga._q_xcount[1] ));
 sg13g2_dfrbp_1 _7131_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net226),
    .D(_0070_),
    .Q_N(_3446_),
    .Q(\main.demo.vga._q_xcount[2] ));
 sg13g2_dfrbp_1 _7132_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net225),
    .D(_0071_),
    .Q_N(_3445_),
    .Q(\main.demo.vga._q_xcount[3] ));
 sg13g2_dfrbp_1 _7133_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net224),
    .D(_0072_),
    .Q_N(_3444_),
    .Q(\main.demo.vga._q_xcount[4] ));
 sg13g2_dfrbp_1 _7134_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net223),
    .D(_0073_),
    .Q_N(_3443_),
    .Q(\main.demo.vga._q_xcount[7] ));
 sg13g2_dfrbp_1 _7135_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net26),
    .D(_0074_),
    .Q_N(_3450_),
    .Q(\main.demo.vga._d_vblank ));
 sg13g2_dfrbp_1 _7136_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net27),
    .D(net390),
    .Q_N(_3451_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ));
 sg13g2_dfrbp_1 _7137_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net28),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .Q_N(_3452_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ));
 sg13g2_dfrbp_1 _7138_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net29),
    .D(net403),
    .Q_N(_3453_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ));
 sg13g2_dfrbp_1 _7139_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net30),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[4] ),
    .Q_N(_3454_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_dfrbp_1 _7140_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net31),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[6] ),
    .Q_N(_3455_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ));
 sg13g2_dfrbp_1 _7141_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net63),
    .D(net293),
    .Q_N(_3456_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[7] ));
 sg13g2_dfrbp_1 _7142_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net222),
    .D(net313),
    .Q_N(_3442_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _7143_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net220),
    .D(net608),
    .Q_N(_3441_),
    .Q(\main.demo._q_speed[0] ));
 sg13g2_dfrbp_1 _7144_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net218),
    .D(net642),
    .Q_N(_0015_),
    .Q(\main.demo._q_speed[1] ));
 sg13g2_dfrbp_1 _7145_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net217),
    .D(_0077_),
    .Q_N(_0014_),
    .Q(\main.demo._q_speed[2] ));
 sg13g2_dfrbp_1 _7146_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net216),
    .D(_0078_),
    .Q_N(_0013_),
    .Q(\main.demo._q_speed[3] ));
 sg13g2_dfrbp_1 _7147_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net215),
    .D(net587),
    .Q_N(_0012_),
    .Q(\main.demo._q_speed[4] ));
 sg13g2_dfrbp_1 _7148_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net214),
    .D(_0080_),
    .Q_N(_0007_),
    .Q(\main.demo._q_speed[5] ));
 sg13g2_dfrbp_1 _7149_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net213),
    .D(net623),
    .Q_N(_0019_),
    .Q(\main.demo._q_speed[6] ));
 sg13g2_dfrbp_1 _7150_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net212),
    .D(_0082_),
    .Q_N(_3440_),
    .Q(\main.demo._q_speed[7] ));
 sg13g2_dfrbp_1 _7151_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net211),
    .D(_0083_),
    .Q_N(_3439_),
    .Q(\main.demo._q_speed[8] ));
 sg13g2_dfrbp_1 _7152_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net210),
    .D(net575),
    .Q_N(_3438_),
    .Q(\main.demo._q_speed[9] ));
 sg13g2_dfrbp_1 _7153_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net209),
    .D(_0085_),
    .Q_N(_3437_),
    .Q(\main.demo._q_speed[10] ));
 sg13g2_dfrbp_1 _7154_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net208),
    .D(_0086_),
    .Q_N(_3436_),
    .Q(\main.demo._q_speed[11] ));
 sg13g2_dfrbp_1 _7155_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net207),
    .D(net581),
    .Q_N(_3435_),
    .Q(\main.demo._q_speed[12] ));
 sg13g2_dfrbp_1 _7156_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net206),
    .D(_0088_),
    .Q_N(_3434_),
    .Q(\main.demo._q_speed[13] ));
 sg13g2_dfrbp_1 _7157_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net205),
    .D(_0089_),
    .Q_N(_3433_),
    .Q(\main.demo._q_speed[14] ));
 sg13g2_dfrbp_1 _7158_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net204),
    .D(_0090_),
    .Q_N(_3432_),
    .Q(\main.demo._q_speed[15] ));
 sg13g2_dfrbp_1 _7159_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net203),
    .D(_0091_),
    .Q_N(_3431_),
    .Q(\main.demo._q_frame[0] ));
 sg13g2_dfrbp_1 _7160_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net202),
    .D(_0092_),
    .Q_N(_3430_),
    .Q(\main.demo._q_frame[1] ));
 sg13g2_dfrbp_1 _7161_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net201),
    .D(_0093_),
    .Q_N(_3429_),
    .Q(\main.demo._q_frame[2] ));
 sg13g2_dfrbp_1 _7162_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net200),
    .D(_0094_),
    .Q_N(_3428_),
    .Q(\main.demo._q_frame[3] ));
 sg13g2_dfrbp_1 _7163_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net199),
    .D(_0095_),
    .Q_N(_3427_),
    .Q(\main.demo._q_frame[4] ));
 sg13g2_dfrbp_1 _7164_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net198),
    .D(_0096_),
    .Q_N(_3426_),
    .Q(\main.demo._q_frame[5] ));
 sg13g2_dfrbp_1 _7165_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net197),
    .D(_0097_),
    .Q_N(_3425_),
    .Q(\main.demo._q_frame[6] ));
 sg13g2_dfrbp_1 _7166_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net196),
    .D(_0098_),
    .Q_N(_3424_),
    .Q(\main.demo._q_frame[7] ));
 sg13g2_dfrbp_1 _7167_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net195),
    .D(_0099_),
    .Q_N(_3423_),
    .Q(\main.demo._q_frame[8] ));
 sg13g2_dfrbp_1 _7168_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net194),
    .D(_0100_),
    .Q_N(_3422_),
    .Q(\main.demo._q_frame[9] ));
 sg13g2_dfrbp_1 _7169_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net193),
    .D(_0101_),
    .Q_N(_3421_),
    .Q(\main.demo._q_frame[10] ));
 sg13g2_dfrbp_1 _7170_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net192),
    .D(_0102_),
    .Q_N(_3420_),
    .Q(\main.demo._q_frame[11] ));
 sg13g2_dfrbp_1 _7171_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net191),
    .D(_0103_),
    .Q_N(_3419_),
    .Q(\main.demo._q_frame[12] ));
 sg13g2_dfrbp_1 _7172_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net190),
    .D(_0104_),
    .Q_N(_3418_),
    .Q(\main.demo._q_frame[13] ));
 sg13g2_dfrbp_1 _7173_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net64),
    .D(_0105_),
    .Q_N(_3457_),
    .Q(\main.demo._q_frame[14] ));
 sg13g2_dfrbp_1 _7174_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net65),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[0] ),
    .Q_N(_3458_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ));
 sg13g2_dfrbp_1 _7175_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net66),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[1] ),
    .Q_N(_3459_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ));
 sg13g2_dfrbp_1 _7176_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net67),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[2] ),
    .Q_N(_3460_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ));
 sg13g2_dfrbp_1 _7177_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net68),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[3] ),
    .Q_N(_0038_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ));
 sg13g2_dfrbp_1 _7178_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net69),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[4] ),
    .Q_N(_0050_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ));
 sg13g2_dfrbp_1 _7179_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net70),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[5] ),
    .Q_N(_0049_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ));
 sg13g2_dfrbp_1 _7180_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net71),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[6] ),
    .Q_N(_0048_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ));
 sg13g2_dfrbp_1 _7181_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net72),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[7] ),
    .Q_N(_0047_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ));
 sg13g2_dfrbp_1 _7182_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net73),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[8] ),
    .Q_N(_0046_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ));
 sg13g2_dfrbp_1 _7183_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net74),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[9] ),
    .Q_N(_0045_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ));
 sg13g2_dfrbp_1 _7184_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net75),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[10] ),
    .Q_N(_0043_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[10] ));
 sg13g2_dfrbp_1 _7185_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net76),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[0] ),
    .Q_N(_3461_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_dfrbp_1 _7186_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net77),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[1] ),
    .Q_N(_3462_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ));
 sg13g2_dfrbp_1 _7187_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net78),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[2] ),
    .Q_N(_3463_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ));
 sg13g2_dfrbp_1 _7188_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net79),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[3] ),
    .Q_N(_3464_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ));
 sg13g2_dfrbp_1 _7189_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net80),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[4] ),
    .Q_N(_3465_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ));
 sg13g2_dfrbp_1 _7190_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net81),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[5] ),
    .Q_N(_3466_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_dfrbp_1 _7191_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net82),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[6] ),
    .Q_N(_3467_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ));
 sg13g2_dfrbp_1 _7192_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net83),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[7] ),
    .Q_N(_3468_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ));
 sg13g2_dfrbp_1 _7193_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net84),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[8] ),
    .Q_N(_3469_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ));
 sg13g2_dfrbp_1 _7194_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net85),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[9] ),
    .Q_N(_3470_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ));
 sg13g2_dfrbp_1 _7195_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net86),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[10] ),
    .Q_N(_3471_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ));
 sg13g2_dfrbp_1 _7196_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net87),
    .D(net592),
    .Q_N(_3472_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 _7197_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net88),
    .D(net286),
    .Q_N(_3473_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 _7198_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net89),
    .D(net486),
    .Q_N(_3474_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 _7199_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net90),
    .D(net545),
    .Q_N(_3475_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 _7200_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net91),
    .D(net296),
    .Q_N(_3476_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 _7201_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net92),
    .D(net318),
    .Q_N(_3477_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 _7202_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net93),
    .D(net294),
    .Q_N(_3478_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 _7203_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net94),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[0] ),
    .Q_N(_0011_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 _7204_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net95),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[1] ),
    .Q_N(_0008_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 _7205_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net96),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[2] ),
    .Q_N(_3479_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 _7206_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net97),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[3] ),
    .Q_N(_0010_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 _7207_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net98),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[4] ),
    .Q_N(_0009_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 _7208_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net99),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[5] ),
    .Q_N(_3480_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 _7209_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net100),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[6] ),
    .Q_N(_3481_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 _7210_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net101),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[7] ),
    .Q_N(_0036_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 _7211_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net102),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[8] ),
    .Q_N(_0006_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 _7212_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net103),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[9] ),
    .Q_N(_3482_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 _7213_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net104),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[10] ),
    .Q_N(_3483_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 _7214_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net105),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[0] ),
    .Q_N(_3484_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 _7215_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net106),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[1] ),
    .Q_N(_3485_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 _7216_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net107),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[2] ),
    .Q_N(_3486_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 _7217_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net108),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[3] ),
    .Q_N(_3487_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 _7218_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net109),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[4] ),
    .Q_N(_0041_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 _7219_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net110),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[5] ),
    .Q_N(_0040_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 _7220_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net111),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[6] ),
    .Q_N(_0039_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 _7221_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net112),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[7] ),
    .Q_N(_0037_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 _7222_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net113),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[8] ),
    .Q_N(_0044_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 _7223_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net114),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[9] ),
    .Q_N(_0042_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 _7224_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net115),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[10] ),
    .Q_N(_0051_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 _7225_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net116),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[0] ),
    .Q_N(_3488_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 _7226_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net117),
    .D(net324),
    .Q_N(_3489_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 _7227_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net118),
    .D(net568),
    .Q_N(_3490_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 _7228_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net119),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[3] ),
    .Q_N(_3491_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 _7229_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net120),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[4] ),
    .Q_N(_3492_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 _7230_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net121),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[5] ),
    .Q_N(_3493_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 _7231_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net122),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[6] ),
    .Q_N(_3494_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 _7232_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net123),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[7] ),
    .Q_N(_3495_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 _7233_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net124),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[8] ),
    .Q_N(_3496_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 _7234_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net125),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[9] ),
    .Q_N(_3497_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 _7235_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net126),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[10] ),
    .Q_N(_3498_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 _7236_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net127),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[1] ),
    .Q_N(_3499_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ));
 sg13g2_dfrbp_1 _7237_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net128),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[2] ),
    .Q_N(_0018_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ));
 sg13g2_dfrbp_1 _7238_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net129),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[3] ),
    .Q_N(_0017_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[3] ));
 sg13g2_dfrbp_1 _7239_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net130),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[4] ),
    .Q_N(_0016_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[4] ));
 sg13g2_dfrbp_1 _7240_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net131),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[5] ),
    .Q_N(_0021_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[5] ));
 sg13g2_dfrbp_1 _7241_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net132),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[6] ),
    .Q_N(_0020_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ));
 sg13g2_dfrbp_1 _7242_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net133),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[7] ),
    .Q_N(_3500_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ));
 sg13g2_dfrbp_1 _7243_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net134),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ),
    .Q_N(_3501_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_l[0] ));
 sg13g2_dfrbp_1 _7244_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net135),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .Q_N(_3502_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ));
 sg13g2_dfrbp_1 _7245_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net136),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .Q_N(_3503_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ));
 sg13g2_dfrbp_1 _7246_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net137),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_h[1] ),
    .Q_N(_3504_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_dfrbp_1 _7247_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net138),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ),
    .Q_N(_3505_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_dfrbp_1 _7248_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net139),
    .D(\main.demo._t___block_68_frag[0] ),
    .Q_N(_3506_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[0] ));
 sg13g2_dfrbp_1 _7249_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net140),
    .D(\main.demo._t___block_68_frag[1] ),
    .Q_N(_3507_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[1] ));
 sg13g2_dfrbp_1 _7250_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net141),
    .D(\main.demo._t___block_68_frag[2] ),
    .Q_N(_3508_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[2] ));
 sg13g2_dfrbp_1 _7251_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net142),
    .D(\main.demo._t___block_68_frag[3] ),
    .Q_N(_3509_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[3] ));
 sg13g2_dfrbp_1 _7252_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net155),
    .D(\main.demo._t___block_68_frag[4] ),
    .Q_N(_3510_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[4] ));
 sg13g2_dfrbp_1 _7253_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net189),
    .D(\main.demo._t___block_68_frag[5] ),
    .Q_N(_3417_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[5] ));
 sg13g2_dfrbp_1 _7254_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net188),
    .D(net310),
    .Q_N(_0000_),
    .Q(\main.demo._q_rot_en ));
 sg13g2_dfrbp_1 _7255_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net185),
    .D(net548),
    .Q_N(_0066_),
    .Q(\main.demo._q_effect[0] ));
 sg13g2_dfrbp_1 _7256_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net183),
    .D(_0108_),
    .Q_N(_3416_),
    .Q(\main.demo._q_effect[1] ));
 sg13g2_dfrbp_1 _7257_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net181),
    .D(net288),
    .Q_N(_0065_),
    .Q(\main.demo._q_th[0] ));
 sg13g2_dfrbp_1 _7258_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net179),
    .D(net306),
    .Q_N(_3415_),
    .Q(\main.demo._q_th[1] ));
 sg13g2_dfrbp_1 _7259_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net177),
    .D(_0111_),
    .Q_N(_3414_),
    .Q(\main.demo._q_th[2] ));
 sg13g2_dfrbp_1 _7260_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net175),
    .D(_0112_),
    .Q_N(_3413_),
    .Q(\main.demo._q_th[3] ));
 sg13g2_dfrbp_1 _7261_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net173),
    .D(net381),
    .Q_N(_3412_),
    .Q(\main.demo._q_th[4] ));
 sg13g2_dfrbp_1 _7262_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net171),
    .D(_0114_),
    .Q_N(_3411_),
    .Q(\main.demo._q_th[5] ));
 sg13g2_dfrbp_1 _7263_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net169),
    .D(_0115_),
    .Q_N(_0022_),
    .Q(\main.demo._q_th[6] ));
 sg13g2_dfrbp_1 _7264_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net167),
    .D(_0116_),
    .Q_N(_3410_),
    .Q(\main.demo._q_th[7] ));
 sg13g2_dfrbp_1 _7265_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net156),
    .D(_0117_),
    .Q_N(_3511_),
    .Q(\main.demo._q_th[8] ));
 sg13g2_dfrbp_1 _7266_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net157),
    .D(\main.demo._d_prev_b[0] ),
    .Q_N(_3512_),
    .Q(\main.demo._d_prev_b[2] ));
 sg13g2_dfrbp_1 _7267_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net158),
    .D(\main.demo._d_prev_b[1] ),
    .Q_N(_3513_),
    .Q(\main.demo._d_prev_b[3] ));
 sg13g2_dfrbp_1 _7268_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net159),
    .D(net281),
    .Q_N(_3514_),
    .Q(\main.demo._d_prev_b[4] ));
 sg13g2_dfrbp_1 _7269_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net160),
    .D(net283),
    .Q_N(_3515_),
    .Q(\main.demo._d_prev_b[5] ));
 sg13g2_dfrbp_1 _7270_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net161),
    .D(net280),
    .Q_N(_3516_),
    .Q(\main.demo._d_prev_b[6] ));
 sg13g2_dfrbp_1 _7271_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net162),
    .D(net282),
    .Q_N(_3517_),
    .Q(\main.demo._d_prev_b[7] ));
 sg13g2_dfrbp_1 _7272_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net163),
    .D(net278),
    .Q_N(_3518_),
    .Q(\main.demo._q_prev_b[6] ));
 sg13g2_dfrbp_1 _7273_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net164),
    .D(net284),
    .Q_N(_3519_),
    .Q(\main.demo._q_prev_b[7] ));
 sg13g2_dfrbp_1 _7274_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net187),
    .D(net291),
    .Q_N(_3520_),
    .Q(\main.demo._q_prev_vs ));
 sg13g2_dfrbp_1 _7275_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net165),
    .D(net279),
    .Q_N(_3409_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _7276_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net153),
    .D(_0118_),
    .Q_N(_3408_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _7277_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net152),
    .D(_0119_),
    .Q_N(_3407_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7278_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net151),
    .D(_0120_),
    .Q_N(_3406_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7279_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net150),
    .D(_0121_),
    .Q_N(_3405_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _7280_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net149),
    .D(_0122_),
    .Q_N(_3404_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7281_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net148),
    .D(_0123_),
    .Q_N(_3403_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7282_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net147),
    .D(_0124_),
    .Q_N(_3402_),
    .Q(\main.demo.zic._q_drum_inc[0] ));
 sg13g2_dfrbp_1 _7283_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net146),
    .D(net615),
    .Q_N(_3401_),
    .Q(\main.demo.zic._q_drum_inc[1] ));
 sg13g2_dfrbp_1 _7284_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net145),
    .D(_0126_),
    .Q_N(_3400_),
    .Q(\main.demo.zic._q_drum_inc[2] ));
 sg13g2_dfrbp_1 _7285_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net144),
    .D(_0127_),
    .Q_N(_3399_),
    .Q(\main.demo.zic._q_drum_inc[3] ));
 sg13g2_dfrbp_1 _7286_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net143),
    .D(_0128_),
    .Q_N(_0004_),
    .Q(\main.demo._t___stage___block_3_x[0] ));
 sg13g2_dfrbp_1 _7287_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net62),
    .D(_0129_),
    .Q_N(_0005_),
    .Q(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_dfrbp_1 _7288_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net61),
    .D(_0130_),
    .Q_N(_3398_),
    .Q(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_dfrbp_1 _7289_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net60),
    .D(_0131_),
    .Q_N(_0058_),
    .Q(\main.demo._w_vga_vga_x[3] ));
 sg13g2_dfrbp_1 _7290_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net59),
    .D(_0132_),
    .Q_N(_0057_),
    .Q(\main.demo._w_vga_vga_x[4] ));
 sg13g2_dfrbp_1 _7291_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net58),
    .D(_0133_),
    .Q_N(_0056_),
    .Q(\main.demo._w_vga_vga_x[5] ));
 sg13g2_dfrbp_1 _7292_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net57),
    .D(_0134_),
    .Q_N(_0055_),
    .Q(\main.demo._w_vga_vga_x[6] ));
 sg13g2_dfrbp_1 _7293_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net56),
    .D(_0135_),
    .Q_N(_0054_),
    .Q(\main.demo._w_vga_vga_x[7] ));
 sg13g2_dfrbp_1 _7294_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net55),
    .D(_0136_),
    .Q_N(_0053_),
    .Q(\main.demo._w_vga_vga_x[8] ));
 sg13g2_dfrbp_1 _7295_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net54),
    .D(_0137_),
    .Q_N(_0052_),
    .Q(\main.demo._w_vga_vga_x[9] ));
 sg13g2_dfrbp_1 _7296_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net53),
    .D(_0138_),
    .Q_N(_3397_),
    .Q(\main.demo._w_vga_vga_x[10] ));
 sg13g2_dfrbp_1 _7297_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net239),
    .D(_0139_),
    .Q_N(_3521_),
    .Q(\main.demo.vga._q_active_v ));
 sg13g2_dfrbp_1 _7298_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net52),
    .D(\main.demo.vga._d_active ),
    .Q_N(_3396_),
    .Q(\main.demo._w_vga_active ));
 sg13g2_dfrbp_1 _7299_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net51),
    .D(net303),
    .Q_N(_3395_),
    .Q(\main._w_demo_video_vs ));
 sg13g2_dfrbp_1 _7300_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net49),
    .D(net299),
    .Q_N(_3394_),
    .Q(\main._w_demo_video_hs ));
 sg13g2_dfrbp_1 _7301_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net47),
    .D(_0142_),
    .Q_N(_3393_),
    .Q(\main.demo.vga._q_active_h ));
 sg13g2_dfrbp_1 _7302_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net46),
    .D(_0143_),
    .Q_N(_3392_),
    .Q(\main.demo.vga._q_xcount[0] ));
 sg13g2_dfrbp_1 _7303_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net45),
    .D(_0144_),
    .Q_N(_3391_),
    .Q(\main.demo.vga._q_xcount[5] ));
 sg13g2_dfrbp_1 _7304_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net44),
    .D(_0145_),
    .Q_N(_3390_),
    .Q(\main.demo.vga._q_xcount[6] ));
 sg13g2_dfrbp_1 _7305_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net43),
    .D(_0146_),
    .Q_N(_3389_),
    .Q(\main.demo.vga._q_xcount[8] ));
 sg13g2_dfrbp_1 _7306_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net42),
    .D(_0147_),
    .Q_N(_3388_),
    .Q(\main.demo.vga._q_xcount[9] ));
 sg13g2_dfrbp_1 _7307_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net41),
    .D(_0148_),
    .Q_N(_3387_),
    .Q(\main.demo.vga._q_xcount[10] ));
 sg13g2_dfrbp_1 _7308_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net40),
    .D(_0149_),
    .Q_N(_3386_),
    .Q(\main.demo.vga._q_ycount[0] ));
 sg13g2_dfrbp_1 _7309_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net38),
    .D(net525),
    .Q_N(_3385_),
    .Q(\main.demo.vga._q_ycount[1] ));
 sg13g2_dfrbp_1 _7310_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net36),
    .D(_0151_),
    .Q_N(_3384_),
    .Q(\main.demo.vga._q_ycount[2] ));
 sg13g2_dfrbp_1 _7311_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net34),
    .D(net366),
    .Q_N(_3383_),
    .Q(\main.demo.vga._q_ycount[3] ));
 sg13g2_dfrbp_1 _7312_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net32),
    .D(_0153_),
    .Q_N(_3382_),
    .Q(\main.demo.vga._q_ycount[4] ));
 sg13g2_dfrbp_1 _7313_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net23),
    .D(net355),
    .Q_N(_3381_),
    .Q(\main.demo.vga._q_ycount[5] ));
 sg13g2_dfrbp_1 _7314_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net21),
    .D(_0155_),
    .Q_N(_3380_),
    .Q(\main.demo.vga._q_ycount[6] ));
 sg13g2_dfrbp_1 _7315_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net19),
    .D(net361),
    .Q_N(_3379_),
    .Q(\main.demo.vga._q_ycount[7] ));
 sg13g2_dfrbp_1 _7316_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net276),
    .D(_0157_),
    .Q_N(_3378_),
    .Q(\main.demo.vga._q_ycount[8] ));
 sg13g2_dfrbp_1 _7317_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net274),
    .D(_0158_),
    .Q_N(_3377_),
    .Q(\main.demo._q_go ));
 sg13g2_dfrbp_1 _7318_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net273),
    .D(_0159_),
    .Q_N(_0064_),
    .Q(\main.demo.zic._q_clock_count[0] ));
 sg13g2_dfrbp_1 _7319_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net272),
    .D(net611),
    .Q_N(_3376_),
    .Q(\main.demo.zic._q_clock_count[1] ));
 sg13g2_dfrbp_1 _7320_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net271),
    .D(_0161_),
    .Q_N(_3375_),
    .Q(\main.demo.zic._q_clock_count[2] ));
 sg13g2_dfrbp_1 _7321_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net270),
    .D(_0162_),
    .Q_N(_0027_),
    .Q(\main.demo.zic._q_clock_count[3] ));
 sg13g2_dfrbp_1 _7322_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net269),
    .D(_0163_),
    .Q_N(_3374_),
    .Q(\main.demo.zic._q_clock_count[4] ));
 sg13g2_dfrbp_1 _7323_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net268),
    .D(_0164_),
    .Q_N(_0026_),
    .Q(\main.demo.zic._q_clock_count[5] ));
 sg13g2_dfrbp_1 _7324_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net267),
    .D(_0165_),
    .Q_N(_0025_),
    .Q(\main.demo.zic._q_clock_count[6] ));
 sg13g2_dfrbp_1 _7325_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net266),
    .D(_0166_),
    .Q_N(_3373_),
    .Q(\main.demo.zic._q_clock_count[7] ));
 sg13g2_dfrbp_1 _7326_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net265),
    .D(_0167_),
    .Q_N(_3372_),
    .Q(\main.demo.zic._q_clock_count[8] ));
 sg13g2_dfrbp_1 _7327_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net264),
    .D(net290),
    .Q_N(_0063_),
    .Q(\main.demo.zic._q_rythm_count[0] ));
 sg13g2_dfrbp_1 _7328_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net262),
    .D(net328),
    .Q_N(_3371_),
    .Q(\main.demo.zic._q_rythm_count[1] ));
 sg13g2_dfrbp_1 _7329_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net260),
    .D(_0170_),
    .Q_N(_3370_),
    .Q(\main.demo.zic._q_rythm_count[2] ));
 sg13g2_dfrbp_1 _7330_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net258),
    .D(_0171_),
    .Q_N(_3369_),
    .Q(\main.demo.zic._q_rythm_count[3] ));
 sg13g2_dfrbp_1 _7331_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net256),
    .D(net346),
    .Q_N(_3368_),
    .Q(\main.demo.zic._q_rythm_count[4] ));
 sg13g2_dfrbp_1 _7332_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net254),
    .D(_0173_),
    .Q_N(_3367_),
    .Q(\main.demo.zic._q_rythm_count[5] ));
 sg13g2_dfrbp_1 _7333_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net252),
    .D(net343),
    .Q_N(_3366_),
    .Q(\main.demo.zic._q_rythm_count[6] ));
 sg13g2_dfrbp_1 _7334_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net250),
    .D(_0175_),
    .Q_N(_3365_),
    .Q(\main.demo.zic._q_rythm_count[7] ));
 sg13g2_dfrbp_1 _7335_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net248),
    .D(_0176_),
    .Q_N(_3364_),
    .Q(\main.demo.zic._q_rythm_count[8] ));
 sg13g2_dfrbp_1 _7336_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net246),
    .D(_0177_),
    .Q_N(_3363_),
    .Q(\main.demo.zic._q_rythm_count[9] ));
 sg13g2_dfrbp_1 _7337_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net244),
    .D(_0178_),
    .Q_N(_3362_),
    .Q(\main.demo.zic._q_rythm_count[10] ));
 sg13g2_dfrbp_1 _7338_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net242),
    .D(_0179_),
    .Q_N(_3361_),
    .Q(\main.demo.zic._q_rythm_count[11] ));
 sg13g2_dfrbp_1 _7339_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net240),
    .D(_0180_),
    .Q_N(_3360_),
    .Q(\main.demo.zic._q_rythm_count[12] ));
 sg13g2_dfrbp_1 _7340_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net238),
    .D(_0181_),
    .Q_N(_3359_),
    .Q(\main.demo.zic._q_idx[0] ));
 sg13g2_dfrbp_1 _7341_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net237),
    .D(_0182_),
    .Q_N(_3358_),
    .Q(\main.demo.zic._q_idx[1] ));
 sg13g2_dfrbp_1 _7342_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net236),
    .D(_0183_),
    .Q_N(_3357_),
    .Q(\main.demo.zic._q_idx[2] ));
 sg13g2_dfrbp_1 _7343_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net235),
    .D(_0184_),
    .Q_N(_3356_),
    .Q(\main.demo.zic._q_idx[3] ));
 sg13g2_dfrbp_1 _7344_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net234),
    .D(_0185_),
    .Q_N(_0032_),
    .Q(\main.demo.zic._q_idx[4] ));
 sg13g2_dfrbp_1 _7345_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net233),
    .D(_0186_),
    .Q_N(_0035_),
    .Q(\main.demo.zic._q_idx[5] ));
 sg13g2_dfrbp_1 _7346_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net232),
    .D(_0187_),
    .Q_N(_0033_),
    .Q(\main.demo.zic._q_idx[6] ));
 sg13g2_dfrbp_1 _7347_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net231),
    .D(_0188_),
    .Q_N(_3355_),
    .Q(\main.demo._t___stage___block_3_y[0] ));
 sg13g2_dfrbp_1 _7348_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net230),
    .D(_0189_),
    .Q_N(_3354_),
    .Q(\main.demo._t___stage___block_3_y[1] ));
 sg13g2_dfrbp_1 _7349_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net229),
    .D(_0190_),
    .Q_N(_0003_),
    .Q(\main.demo._t___stage___block_3_y[2] ));
 sg13g2_dfrbp_1 _7350_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net228),
    .D(_0191_),
    .Q_N(_0001_),
    .Q(\main.demo._w_vga_vga_y[3] ));
 sg13g2_dfrbp_1 _7351_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net221),
    .D(_0192_),
    .Q_N(_3353_),
    .Q(\main.demo._w_vga_vga_y[4] ));
 sg13g2_dfrbp_1 _7352_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net219),
    .D(_0193_),
    .Q_N(_0062_),
    .Q(\main.demo._w_vga_vga_y[5] ));
 sg13g2_dfrbp_1 _7353_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net186),
    .D(_0194_),
    .Q_N(_0061_),
    .Q(\main.demo._w_vga_vga_y[6] ));
 sg13g2_dfrbp_1 _7354_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net184),
    .D(net315),
    .Q_N(_0060_),
    .Q(\main.demo._w_vga_vga_y[7] ));
 sg13g2_dfrbp_1 _7355_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net182),
    .D(_0196_),
    .Q_N(_3352_),
    .Q(\main.demo._w_vga_vga_y[8] ));
 sg13g2_dfrbp_1 _7356_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net180),
    .D(_0197_),
    .Q_N(_0059_),
    .Q(\main.demo._w_vga_vga_y[10] ));
 sg13g2_dfrbp_1 _7357_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net178),
    .D(_0198_),
    .Q_N(_3351_),
    .Q(\main.demo.zic._q_squ_env[0] ));
 sg13g2_dfrbp_1 _7358_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net174),
    .D(net523),
    .Q_N(_3350_),
    .Q(\main.demo.zic._q_squ_env[1] ));
 sg13g2_dfrbp_1 _7359_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net170),
    .D(_0200_),
    .Q_N(_3349_),
    .Q(\main.demo.zic._q_squ_env[2] ));
 sg13g2_dfrbp_1 _7360_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net166),
    .D(_0201_),
    .Q_N(_3348_),
    .Q(\main.demo.zic._q_squ_env[3] ));
 sg13g2_dfrbp_1 _7361_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net50),
    .D(_0202_),
    .Q_N(_0023_),
    .Q(\main.demo.zic._q_squ_env[4] ));
 sg13g2_dfrbp_1 _7362_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net39),
    .D(_0203_),
    .Q_N(_0024_),
    .Q(\main.demo.zic._q_squ_env[5] ));
 sg13g2_dfrbp_1 _7363_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net35),
    .D(_0204_),
    .Q_N(_3347_),
    .Q(\main.demo.zic._q_tpos[0] ));
 sg13g2_dfrbp_1 _7364_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net24),
    .D(_0205_),
    .Q_N(_3346_),
    .Q(\main.demo.zic._q_tpos[1] ));
 sg13g2_dfrbp_1 _7365_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net20),
    .D(net554),
    .Q_N(_3345_),
    .Q(\main.demo.zic._q_tpos[2] ));
 sg13g2_dfrbp_1 _7366_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net275),
    .D(_0207_),
    .Q_N(_3344_),
    .Q(\main.demo.zic._q_tpos[3] ));
 sg13g2_dfrbp_1 _7367_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net261),
    .D(_0208_),
    .Q_N(_3343_),
    .Q(\main.demo.zic._q_tpos[4] ));
 sg13g2_dfrbp_1 _7368_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net257),
    .D(_0209_),
    .Q_N(_0034_),
    .Q(\main.demo.zic._q_tpos[5] ));
 sg13g2_dfrbp_1 _7369_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net253),
    .D(_0210_),
    .Q_N(_3342_),
    .Q(\main.demo.zic._q_tpos[6] ));
 sg13g2_dfrbp_1 _7370_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net249),
    .D(_0211_),
    .Q_N(_3341_),
    .Q(\main.demo.zic._q_tpos[7] ));
 sg13g2_dfrbp_1 _7371_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net245),
    .D(net359),
    .Q_N(_3340_),
    .Q(\main.demo.zic._q_tpos[8] ));
 sg13g2_dfrbp_1 _7372_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net241),
    .D(_0213_),
    .Q_N(_3339_),
    .Q(\main.demo.zic._q_tpos[9] ));
 sg13g2_dfrbp_1 _7373_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net176),
    .D(_0214_),
    .Q_N(_3338_),
    .Q(\main.demo.zic._q_tpos[10] ));
 sg13g2_dfrbp_1 _7374_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net168),
    .D(_0215_),
    .Q_N(_3337_),
    .Q(\main.demo.zic._q_tpos[11] ));
 sg13g2_dfrbp_1 _7375_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net48),
    .D(_0216_),
    .Q_N(_3336_),
    .Q(\main.demo.zic._q_qpos[0] ));
 sg13g2_dfrbp_1 _7376_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net33),
    .D(net333),
    .Q_N(_0028_),
    .Q(\main.demo.zic._q_qpos[1] ));
 sg13g2_dfrbp_1 _7377_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net16),
    .D(net542),
    .Q_N(_3335_),
    .Q(\main.demo.zic._q_qpos[2] ));
 sg13g2_dfrbp_1 _7378_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net259),
    .D(_0219_),
    .Q_N(_0029_),
    .Q(\main.demo.zic._q_qpos[3] ));
 sg13g2_dfrbp_1 _7379_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net251),
    .D(net551),
    .Q_N(_3334_),
    .Q(\main.demo.zic._q_qpos[4] ));
 sg13g2_dfrbp_1 _7380_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net243),
    .D(_0221_),
    .Q_N(_0030_),
    .Q(\main.demo.zic._q_qpos[5] ));
 sg13g2_dfrbp_1 _7381_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net172),
    .D(net557),
    .Q_N(_3333_),
    .Q(\main.demo.zic._q_qpos[6] ));
 sg13g2_dfrbp_1 _7382_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net37),
    .D(net363),
    .Q_N(_0031_),
    .Q(\main.demo.zic._q_qpos[7] ));
 sg13g2_dfrbp_1 _7383_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net263),
    .D(net375),
    .Q_N(_3332_),
    .Q(\main.demo.zic._q_qpos[8] ));
 sg13g2_dfrbp_1 _7384_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net247),
    .D(_0225_),
    .Q_N(_3331_),
    .Q(\main.demo.zic._q_qpos[9] ));
 sg13g2_dfrbp_1 _7385_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net154),
    .D(_0226_),
    .Q_N(_3330_),
    .Q(\main.demo.zic._q_qpos[10] ));
 sg13g2_dfrbp_1 _7386_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net255),
    .D(net566),
    .Q_N(_3329_),
    .Q(\main.demo.zic._q_qpos[11] ));
 sg13g2_dfrbp_1 _7387_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net22),
    .D(_0228_),
    .Q_N(_3328_),
    .Q(\main.demo.zic._q_qpos[12] ));
 sg13g2_tiehi _7129__17 (.L_HI(net17));
 sg13g2_tiehi _7127__18 (.L_HI(net18));
 sg13g2_tiehi _7315__19 (.L_HI(net19));
 sg13g2_tiehi _7365__20 (.L_HI(net20));
 sg13g2_tiehi _7314__21 (.L_HI(net21));
 sg13g2_tiehi _7387__22 (.L_HI(net22));
 sg13g2_tiehi _7313__23 (.L_HI(net23));
 sg13g2_tiehi _7364__24 (.L_HI(net24));
 sg13g2_tiehi _7128__25 (.L_HI(net25));
 sg13g2_tiehi _7135__26 (.L_HI(net26));
 sg13g2_tiehi _7136__27 (.L_HI(net27));
 sg13g2_tiehi _7137__28 (.L_HI(net28));
 sg13g2_tiehi _7138__29 (.L_HI(net29));
 sg13g2_tiehi _7139__30 (.L_HI(net30));
 sg13g2_tiehi _7140__31 (.L_HI(net31));
 sg13g2_tiehi _7312__32 (.L_HI(net32));
 sg13g2_tiehi _7376__33 (.L_HI(net33));
 sg13g2_tiehi _7311__34 (.L_HI(net34));
 sg13g2_tiehi _7363__35 (.L_HI(net35));
 sg13g2_tiehi _7310__36 (.L_HI(net36));
 sg13g2_tiehi _7382__37 (.L_HI(net37));
 sg13g2_tiehi _7309__38 (.L_HI(net38));
 sg13g2_tiehi _7362__39 (.L_HI(net39));
 sg13g2_tiehi _7308__40 (.L_HI(net40));
 sg13g2_tiehi _7307__41 (.L_HI(net41));
 sg13g2_tiehi _7306__42 (.L_HI(net42));
 sg13g2_tiehi _7305__43 (.L_HI(net43));
 sg13g2_tiehi _7304__44 (.L_HI(net44));
 sg13g2_tiehi _7303__45 (.L_HI(net45));
 sg13g2_tiehi _7302__46 (.L_HI(net46));
 sg13g2_tiehi _7301__47 (.L_HI(net47));
 sg13g2_tiehi _7375__48 (.L_HI(net48));
 sg13g2_tiehi _7300__49 (.L_HI(net49));
 sg13g2_tiehi _7361__50 (.L_HI(net50));
 sg13g2_tiehi _7299__51 (.L_HI(net51));
 sg13g2_tiehi _7298__52 (.L_HI(net52));
 sg13g2_tiehi _7296__53 (.L_HI(net53));
 sg13g2_tiehi _7295__54 (.L_HI(net54));
 sg13g2_tiehi _7294__55 (.L_HI(net55));
 sg13g2_tiehi _7293__56 (.L_HI(net56));
 sg13g2_tiehi _7292__57 (.L_HI(net57));
 sg13g2_tiehi _7291__58 (.L_HI(net58));
 sg13g2_tiehi _7290__59 (.L_HI(net59));
 sg13g2_tiehi _7289__60 (.L_HI(net60));
 sg13g2_tiehi _7288__61 (.L_HI(net61));
 sg13g2_tiehi _7287__62 (.L_HI(net62));
 sg13g2_tiehi _7141__63 (.L_HI(net63));
 sg13g2_tiehi _7173__64 (.L_HI(net64));
 sg13g2_tiehi _7174__65 (.L_HI(net65));
 sg13g2_tiehi _7175__66 (.L_HI(net66));
 sg13g2_tiehi _7176__67 (.L_HI(net67));
 sg13g2_tiehi _7177__68 (.L_HI(net68));
 sg13g2_tiehi _7178__69 (.L_HI(net69));
 sg13g2_tiehi _7179__70 (.L_HI(net70));
 sg13g2_tiehi _7180__71 (.L_HI(net71));
 sg13g2_tiehi _7181__72 (.L_HI(net72));
 sg13g2_tiehi _7182__73 (.L_HI(net73));
 sg13g2_tiehi _7183__74 (.L_HI(net74));
 sg13g2_tiehi _7184__75 (.L_HI(net75));
 sg13g2_tiehi _7185__76 (.L_HI(net76));
 sg13g2_tiehi _7186__77 (.L_HI(net77));
 sg13g2_tiehi _7187__78 (.L_HI(net78));
 sg13g2_tiehi _7188__79 (.L_HI(net79));
 sg13g2_tiehi _7189__80 (.L_HI(net80));
 sg13g2_tiehi _7190__81 (.L_HI(net81));
 sg13g2_tiehi _7191__82 (.L_HI(net82));
 sg13g2_tiehi _7192__83 (.L_HI(net83));
 sg13g2_tiehi _7193__84 (.L_HI(net84));
 sg13g2_tiehi _7194__85 (.L_HI(net85));
 sg13g2_tiehi _7195__86 (.L_HI(net86));
 sg13g2_tiehi _7196__87 (.L_HI(net87));
 sg13g2_tiehi _7197__88 (.L_HI(net88));
 sg13g2_tiehi _7198__89 (.L_HI(net89));
 sg13g2_tiehi _7199__90 (.L_HI(net90));
 sg13g2_tiehi _7200__91 (.L_HI(net91));
 sg13g2_tiehi _7201__92 (.L_HI(net92));
 sg13g2_tiehi _7202__93 (.L_HI(net93));
 sg13g2_tiehi _7203__94 (.L_HI(net94));
 sg13g2_tiehi _7204__95 (.L_HI(net95));
 sg13g2_tiehi _7205__96 (.L_HI(net96));
 sg13g2_tiehi _7206__97 (.L_HI(net97));
 sg13g2_tiehi _7207__98 (.L_HI(net98));
 sg13g2_tiehi _7208__99 (.L_HI(net99));
 sg13g2_tiehi _7209__100 (.L_HI(net100));
 sg13g2_tiehi _7210__101 (.L_HI(net101));
 sg13g2_tiehi _7211__102 (.L_HI(net102));
 sg13g2_tiehi _7212__103 (.L_HI(net103));
 sg13g2_tiehi _7213__104 (.L_HI(net104));
 sg13g2_tiehi _7214__105 (.L_HI(net105));
 sg13g2_tiehi _7215__106 (.L_HI(net106));
 sg13g2_tiehi _7216__107 (.L_HI(net107));
 sg13g2_tiehi _7217__108 (.L_HI(net108));
 sg13g2_tiehi _7218__109 (.L_HI(net109));
 sg13g2_tiehi _7219__110 (.L_HI(net110));
 sg13g2_tiehi _7220__111 (.L_HI(net111));
 sg13g2_tiehi _7221__112 (.L_HI(net112));
 sg13g2_tiehi _7222__113 (.L_HI(net113));
 sg13g2_tiehi _7223__114 (.L_HI(net114));
 sg13g2_tiehi _7224__115 (.L_HI(net115));
 sg13g2_tiehi _7225__116 (.L_HI(net116));
 sg13g2_tiehi _7226__117 (.L_HI(net117));
 sg13g2_tiehi _7227__118 (.L_HI(net118));
 sg13g2_tiehi _7228__119 (.L_HI(net119));
 sg13g2_tiehi _7229__120 (.L_HI(net120));
 sg13g2_tiehi _7230__121 (.L_HI(net121));
 sg13g2_tiehi _7231__122 (.L_HI(net122));
 sg13g2_tiehi _7232__123 (.L_HI(net123));
 sg13g2_tiehi _7233__124 (.L_HI(net124));
 sg13g2_tiehi _7234__125 (.L_HI(net125));
 sg13g2_tiehi _7235__126 (.L_HI(net126));
 sg13g2_tiehi _7236__127 (.L_HI(net127));
 sg13g2_tiehi _7237__128 (.L_HI(net128));
 sg13g2_tiehi _7238__129 (.L_HI(net129));
 sg13g2_tiehi _7239__130 (.L_HI(net130));
 sg13g2_tiehi _7240__131 (.L_HI(net131));
 sg13g2_tiehi _7241__132 (.L_HI(net132));
 sg13g2_tiehi _7242__133 (.L_HI(net133));
 sg13g2_tiehi _7243__134 (.L_HI(net134));
 sg13g2_tiehi _7244__135 (.L_HI(net135));
 sg13g2_tiehi _7245__136 (.L_HI(net136));
 sg13g2_tiehi _7246__137 (.L_HI(net137));
 sg13g2_tiehi _7247__138 (.L_HI(net138));
 sg13g2_tiehi _7248__139 (.L_HI(net139));
 sg13g2_tiehi _7249__140 (.L_HI(net140));
 sg13g2_tiehi _7250__141 (.L_HI(net141));
 sg13g2_tiehi _7251__142 (.L_HI(net142));
 sg13g2_tiehi _7286__143 (.L_HI(net143));
 sg13g2_tiehi _7285__144 (.L_HI(net144));
 sg13g2_tiehi _7284__145 (.L_HI(net145));
 sg13g2_tiehi _7283__146 (.L_HI(net146));
 sg13g2_tiehi _7282__147 (.L_HI(net147));
 sg13g2_tiehi _7281__148 (.L_HI(net148));
 sg13g2_tiehi _7280__149 (.L_HI(net149));
 sg13g2_tiehi _7279__150 (.L_HI(net150));
 sg13g2_tiehi _7278__151 (.L_HI(net151));
 sg13g2_tiehi _7277__152 (.L_HI(net152));
 sg13g2_tiehi _7276__153 (.L_HI(net153));
 sg13g2_tiehi _7385__154 (.L_HI(net154));
 sg13g2_tiehi _7252__155 (.L_HI(net155));
 sg13g2_tiehi _7265__156 (.L_HI(net156));
 sg13g2_tiehi _7266__157 (.L_HI(net157));
 sg13g2_tiehi _7267__158 (.L_HI(net158));
 sg13g2_tiehi _7268__159 (.L_HI(net159));
 sg13g2_tiehi _7269__160 (.L_HI(net160));
 sg13g2_tiehi _7270__161 (.L_HI(net161));
 sg13g2_tiehi _7271__162 (.L_HI(net162));
 sg13g2_tiehi _7272__163 (.L_HI(net163));
 sg13g2_tiehi _7273__164 (.L_HI(net164));
 sg13g2_tiehi _7275__165 (.L_HI(net165));
 sg13g2_tiehi _7360__166 (.L_HI(net166));
 sg13g2_tiehi _7264__167 (.L_HI(net167));
 sg13g2_tiehi _7374__168 (.L_HI(net168));
 sg13g2_tiehi _7263__169 (.L_HI(net169));
 sg13g2_tiehi _7359__170 (.L_HI(net170));
 sg13g2_tiehi _7262__171 (.L_HI(net171));
 sg13g2_tiehi _7381__172 (.L_HI(net172));
 sg13g2_tiehi _7261__173 (.L_HI(net173));
 sg13g2_tiehi _7358__174 (.L_HI(net174));
 sg13g2_tiehi _7260__175 (.L_HI(net175));
 sg13g2_tiehi _7373__176 (.L_HI(net176));
 sg13g2_tiehi _7259__177 (.L_HI(net177));
 sg13g2_tiehi _7357__178 (.L_HI(net178));
 sg13g2_tiehi _7258__179 (.L_HI(net179));
 sg13g2_tiehi _7356__180 (.L_HI(net180));
 sg13g2_tiehi _7257__181 (.L_HI(net181));
 sg13g2_tiehi _7355__182 (.L_HI(net182));
 sg13g2_tiehi _7256__183 (.L_HI(net183));
 sg13g2_tiehi _7354__184 (.L_HI(net184));
 sg13g2_tiehi _7255__185 (.L_HI(net185));
 sg13g2_tiehi _7353__186 (.L_HI(net186));
 sg13g2_tiehi _7274__187 (.L_HI(net187));
 sg13g2_tiehi _7254__188 (.L_HI(net188));
 sg13g2_tiehi _7253__189 (.L_HI(net189));
 sg13g2_tiehi _7172__190 (.L_HI(net190));
 sg13g2_tiehi _7171__191 (.L_HI(net191));
 sg13g2_tiehi _7170__192 (.L_HI(net192));
 sg13g2_tiehi _7169__193 (.L_HI(net193));
 sg13g2_tiehi _7168__194 (.L_HI(net194));
 sg13g2_tiehi _7167__195 (.L_HI(net195));
 sg13g2_tiehi _7166__196 (.L_HI(net196));
 sg13g2_tiehi _7165__197 (.L_HI(net197));
 sg13g2_tiehi _7164__198 (.L_HI(net198));
 sg13g2_tiehi _7163__199 (.L_HI(net199));
 sg13g2_tiehi _7162__200 (.L_HI(net200));
 sg13g2_tiehi _7161__201 (.L_HI(net201));
 sg13g2_tiehi _7160__202 (.L_HI(net202));
 sg13g2_tiehi _7159__203 (.L_HI(net203));
 sg13g2_tiehi _7158__204 (.L_HI(net204));
 sg13g2_tiehi _7157__205 (.L_HI(net205));
 sg13g2_tiehi _7156__206 (.L_HI(net206));
 sg13g2_tiehi _7155__207 (.L_HI(net207));
 sg13g2_tiehi _7154__208 (.L_HI(net208));
 sg13g2_tiehi _7153__209 (.L_HI(net209));
 sg13g2_tiehi _7152__210 (.L_HI(net210));
 sg13g2_tiehi _7151__211 (.L_HI(net211));
 sg13g2_tiehi _7150__212 (.L_HI(net212));
 sg13g2_tiehi _7149__213 (.L_HI(net213));
 sg13g2_tiehi _7148__214 (.L_HI(net214));
 sg13g2_tiehi _7147__215 (.L_HI(net215));
 sg13g2_tiehi _7146__216 (.L_HI(net216));
 sg13g2_tiehi _7145__217 (.L_HI(net217));
 sg13g2_tiehi _7144__218 (.L_HI(net218));
 sg13g2_tiehi _7352__219 (.L_HI(net219));
 sg13g2_tiehi _7143__220 (.L_HI(net220));
 sg13g2_tiehi _7351__221 (.L_HI(net221));
 sg13g2_tiehi _7142__222 (.L_HI(net222));
 sg13g2_tiehi _7134__223 (.L_HI(net223));
 sg13g2_tiehi _7133__224 (.L_HI(net224));
 sg13g2_tiehi _7132__225 (.L_HI(net225));
 sg13g2_tiehi _7131__226 (.L_HI(net226));
 sg13g2_tiehi _7130__227 (.L_HI(net227));
 sg13g2_tiehi _7350__228 (.L_HI(net228));
 sg13g2_tiehi _7349__229 (.L_HI(net229));
 sg13g2_tiehi _7348__230 (.L_HI(net230));
 sg13g2_tiehi _7347__231 (.L_HI(net231));
 sg13g2_tiehi _7346__232 (.L_HI(net232));
 sg13g2_tiehi _7345__233 (.L_HI(net233));
 sg13g2_tiehi _7344__234 (.L_HI(net234));
 sg13g2_tiehi _7343__235 (.L_HI(net235));
 sg13g2_tiehi _7342__236 (.L_HI(net236));
 sg13g2_tiehi _7341__237 (.L_HI(net237));
 sg13g2_tiehi _7340__238 (.L_HI(net238));
 sg13g2_tiehi _7297__239 (.L_HI(net239));
 sg13g2_tiehi _7339__240 (.L_HI(net240));
 sg13g2_tiehi _7372__241 (.L_HI(net241));
 sg13g2_tiehi _7338__242 (.L_HI(net242));
 sg13g2_tiehi _7380__243 (.L_HI(net243));
 sg13g2_tiehi _7337__244 (.L_HI(net244));
 sg13g2_tiehi _7371__245 (.L_HI(net245));
 sg13g2_tiehi _7336__246 (.L_HI(net246));
 sg13g2_tiehi _7384__247 (.L_HI(net247));
 sg13g2_tiehi _7335__248 (.L_HI(net248));
 sg13g2_tiehi _7370__249 (.L_HI(net249));
 sg13g2_tiehi _7334__250 (.L_HI(net250));
 sg13g2_tiehi _7379__251 (.L_HI(net251));
 sg13g2_tiehi _7333__252 (.L_HI(net252));
 sg13g2_tiehi _7369__253 (.L_HI(net253));
 sg13g2_tiehi _7332__254 (.L_HI(net254));
 sg13g2_tiehi _7386__255 (.L_HI(net255));
 sg13g2_tiehi _7331__256 (.L_HI(net256));
 sg13g2_tiehi _7368__257 (.L_HI(net257));
 sg13g2_tiehi _7330__258 (.L_HI(net258));
 sg13g2_tiehi _7378__259 (.L_HI(net259));
 sg13g2_tiehi _7329__260 (.L_HI(net260));
 sg13g2_tiehi _7367__261 (.L_HI(net261));
 sg13g2_tiehi _7328__262 (.L_HI(net262));
 sg13g2_tiehi _7383__263 (.L_HI(net263));
 sg13g2_tiehi _7327__264 (.L_HI(net264));
 sg13g2_tiehi _7326__265 (.L_HI(net265));
 sg13g2_tiehi _7325__266 (.L_HI(net266));
 sg13g2_tiehi _7324__267 (.L_HI(net267));
 sg13g2_tiehi _7323__268 (.L_HI(net268));
 sg13g2_tiehi _7322__269 (.L_HI(net269));
 sg13g2_tiehi _7321__270 (.L_HI(net270));
 sg13g2_tiehi _7320__271 (.L_HI(net271));
 sg13g2_tiehi _7319__272 (.L_HI(net272));
 sg13g2_tiehi _7318__273 (.L_HI(net273));
 sg13g2_tiehi _7317__274 (.L_HI(net274));
 sg13g2_tiehi _7366__275 (.L_HI(net275));
 sg13g2_tiehi _7316__276 (.L_HI(net276));
 sg13g2_tiehi tt_um_silice_277 (.L_HI(net277));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_silice_3 (.L_LO(net3));
 sg13g2_tielo tt_um_silice_4 (.L_LO(net4));
 sg13g2_tielo tt_um_silice_5 (.L_LO(net5));
 sg13g2_tielo tt_um_silice_6 (.L_LO(net6));
 sg13g2_tielo tt_um_silice_7 (.L_LO(net7));
 sg13g2_tielo tt_um_silice_8 (.L_LO(net8));
 sg13g2_tielo tt_um_silice_9 (.L_LO(net9));
 sg13g2_tielo tt_um_silice_10 (.L_LO(net10));
 sg13g2_tielo tt_um_silice_11 (.L_LO(net11));
 sg13g2_tielo tt_um_silice_12 (.L_LO(net12));
 sg13g2_tielo tt_um_silice_13 (.L_LO(net13));
 sg13g2_tielo tt_um_silice_14 (.L_LO(net14));
 sg13g2_tielo tt_um_silice_15 (.L_LO(net15));
 sg13g2_tiehi _7377__16 (.L_HI(net16));
 sg13g2_buf_2 _7664_ (.A(\main.demo._q_prev_vs ),
    .X(uo_out[3]));
 sg13g2_buf_2 fanout386 (.A(_1657_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_1517_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_1887_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_1307_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_0277_),
    .X(net393));
 sg13g2_buf_1 fanout394 (.A(_0277_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_3322_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(net399),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_1 fanout399 (.A(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ),
    .X(net400));
 sg13g2_buf_1 fanout401 (.A(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(net407),
    .X(net404));
 sg13g2_buf_1 fanout405 (.A(net407),
    .X(net405));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(net407));
 sg13g2_buf_2 fanout407 (.A(_3095_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_0704_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_2656_),
    .X(net409));
 sg13g2_buf_1 fanout410 (.A(_2656_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_2641_),
    .X(net411));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_0607_));
 sg13g2_buf_4 fanout413 (.X(net413),
    .A(_0505_));
 sg13g2_buf_2 fanout414 (.A(_2187_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_2555_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_2555_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_2425_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_2425_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_2419_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(net421),
    .X(net420));
 sg13g2_buf_1 fanout421 (.A(_0243_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_0234_),
    .X(net422));
 sg13g2_buf_1 fanout423 (.A(_0234_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_2522_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(net427),
    .X(net426));
 sg13g2_buf_1 fanout427 (.A(_2385_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_0231_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_2550_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_2550_),
    .X(net432));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(_2546_));
 sg13g2_buf_2 fanout434 (.A(_1338_),
    .X(net434));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(_1725_));
 sg13g2_buf_2 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_4 fanout437 (.X(net437),
    .A(net438));
 sg13g2_buf_2 fanout438 (.A(_1074_),
    .X(net438));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(net440));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(_1073_));
 sg13g2_buf_2 fanout441 (.A(_0940_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_0940_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_0919_),
    .X(net443));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(net446));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(net446));
 sg13g2_buf_1 fanout446 (.A(_0918_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_1 fanout448 (.A(_3238_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_2969_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net453),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(net453),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_2968_),
    .X(net453));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(net457));
 sg13g2_buf_2 fanout455 (.A(net457),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net457),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(net458),
    .X(net457));
 sg13g2_buf_4 fanout458 (.X(net458),
    .A(_2936_));
 sg13g2_buf_2 fanout459 (.A(net461),
    .X(net459));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(net461));
 sg13g2_buf_2 fanout461 (.A(_2912_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(\main.demo.zic._q_idx[4] ),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(\main.demo.zic._q_idx[3] ),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(net655),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(\main.demo._w_vga_vga_x[8] ),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(\main.demo._w_vga_vga_x[7] ),
    .X(net467));
 sg13g2_buf_1 fanout468 (.A(\main.demo._w_vga_vga_x[7] ),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(\main.demo._w_vga_vga_x[6] ),
    .X(net469));
 sg13g2_buf_1 fanout470 (.A(\main.demo._w_vga_vga_x[6] ),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(\main.demo._w_vga_vga_x[5] ),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(net475),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(\main.demo._q_effect[1] ),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(\main.demo._q_effect[0] ),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(\main.demo._q_effect[0] ),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(\main.demo._q_rot_en ),
    .X(net478));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_l[0] ));
 sg13g2_buf_2 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_1 fanout482 (.A(net338),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(net486),
    .X(net484));
 sg13g2_buf_1 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net322),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(net488));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ));
 sg13g2_buf_2 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(net492),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(net494),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net497),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net499),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[10] ));
 sg13g2_buf_2 fanout500 (.A(\main.demo._q_frame[7] ),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(\main.demo._q_frame[3] ),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(\main.demo._q_frame[2] ),
    .X(net502));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(\main.demo._q_speed[7] ));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(net505));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(net510));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(net510));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(net510));
 sg13g2_buf_2 fanout510 (.A(net571),
    .X(net510));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_silice_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload0 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload1 (.A(clknet_leaf_5_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_39_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_2_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_16_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_9_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_33_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_34_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_36_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_29_clk));
 sg13g2_inv_8 clkload12 (.A(clknet_leaf_31_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_32_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_23_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_24_clk));
 sg13g2_inv_8 clkload17 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_26_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\main.demo._d_prev_b[6] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold2 (.A(\main._w_demo_video_hs ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold3 (.A(\main.demo._d_prev_b[4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold4 (.A(\main.demo._d_prev_b[2] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold5 (.A(\main.demo._d_prev_b[5] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold6 (.A(\main.demo._d_prev_b[3] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold7 (.A(\main.demo._d_prev_b[7] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0064_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold9 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0065_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0109_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0063_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0168_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold14 (.A(\main._w_demo_video_vs ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0068_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold16 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[7] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold17 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0067_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold19 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0036_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0002_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0141_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold23 (.A(\main.demo.zic._q_qpos[0] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold24 (.A(\main.demo.vga._q_ycount[1] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold25 (.A(_2612_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0140_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold27 (.A(\main.demo._q_th[1] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold28 (.A(_2526_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0110_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold30 (.A(\main.demo.vga._q_xcount[5] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0000_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold32 (.A(_2516_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0106_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0025_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1773_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold36 (.A(\main._w_demo_audio1 ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold37 (.A(\main.demo.vga._q_active_v ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0195_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold39 (.A(\main.demo.vga._q_ycount[6] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold40 (.A(\main.demo.vga._q_xcount[0] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold41 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold42 (.A(\main.demo.vga._q_xcount[1] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold43 (.A(\main.demo.vga._q_ycount[8] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold44 (.A(\main.demo.vga._q_xcount[2] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold45 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0005_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold47 (.A(\main.demo._t___pip_58_1_0___stage___block_3_cx[1] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold48 (.A(\main.demo.vga._q_xcount[6] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold49 (.A(\main.demo.zic._q_rythm_count[1] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold50 (.A(_2659_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0169_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold52 (.A(\main.demo.zic._q_tpos[9] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold53 (.A(_2788_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold54 (.A(\main.demo.vga._q_xcount[4] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold55 (.A(\main.demo.zic._q_qpos[1] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0217_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold57 (.A(\main.demo.vga._q_ycount[5] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold58 (.A(\main.demo.zic._q_clock_count[5] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold59 (.A(_2650_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold60 (.A(\main.demo.vga._q_xcount[10] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0006_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold62 (.A(\main.demo.zic._q_clock_count[3] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold63 (.A(_2646_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold64 (.A(\main.demo.zic._q_rythm_count[6] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold65 (.A(_2670_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0174_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold67 (.A(\main.demo.zic._q_rythm_count[4] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold68 (.A(_2667_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0172_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold70 (.A(\main.demo.zic._q_rythm_count[10] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold71 (.A(_2678_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold72 (.A(\main.demo.zic._q_qpos[5] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold73 (.A(_2883_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold74 (.A(\main.demo.vga._q_xcount[3] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold75 (.A(\main.demo.zic._q_qpos[3] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold76 (.A(_2870_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold77 (.A(\main.demo.vga._q_ycount[4] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0154_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold79 (.A(\main.demo.vga._q_xcount[7] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold80 (.A(\main.demo.zic._q_rythm_count[11] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold81 (.A(\main.demo.zic._q_tpos[8] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0212_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold83 (.A(\main.demo.vga._q_ycount[7] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0156_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold85 (.A(\main.demo.zic._q_qpos[7] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0223_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold87 (.A(\main.demo.vga._q_ycount[3] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold88 (.A(_2634_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0152_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold90 (.A(\main.demo.zic._q_clock_count[7] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold91 (.A(\main.demo.zic._q_rythm_count[7] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold92 (.A(_2673_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold93 (.A(\main.demo.zic._q_clock_count[8] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold94 (.A(_2655_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold95 (.A(\main.demo.vga._d_vblank ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold96 (.A(\main.demo.zic._q_qpos[8] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold97 (.A(_2894_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0224_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0034_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold100 (.A(_2782_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold101 (.A(\main.demo.zic._q_rythm_count[12] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold102 (.A(\main.demo._q_th[4] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold103 (.A(_2531_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0113_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold105 (.A(\main.demo.vga._q_xcount[6] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold106 (.A(\main.demo._q_th[8] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold107 (.A(_2539_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold108 (.A(\main.demo.zic._q_squ_env[2] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold109 (.A(\main.demo.zic._q_clock_count[6] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold110 (.A(\main.demo.zic._q_rythm_count[5] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold111 (.A(_2668_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold112 (.A(\main.demo.vga._q_ycount[1] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0237_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold114 (.A(\main.demo.zic._q_rythm_count[2] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold115 (.A(_2662_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold116 (.A(\main.demo.zic._q_rythm_count[3] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold117 (.A(_2664_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold118 (.A(\main.demo.vga._q_xcount[9] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold119 (.A(\main.demo.vga._q_xcount[8] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold120 (.A(\main.demo.zic._q_squ_env[1] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0199_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold122 (.A(\main.demo.vga._q_ycount[0] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0150_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold124 (.A(\main.demo.zic._q_rythm_count[8] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold125 (.A(\main.demo.vga._q_ycount[0] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold126 (.A(\main.demo.zic._q_qpos[9] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold127 (.A(_2896_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold128 (.A(\main.demo.zic._q_clock_count[2] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold129 (.A(_2644_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold130 (.A(\main.demo.zic._q_tpos[7] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold131 (.A(_2785_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold132 (.A(\main.demo.zic._q_squ_env[0] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold133 (.A(\main.demo.zic._q_tpos[10] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold134 (.A(\main.demo._w_vga_active ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold135 (.A(\main.demo._q_prev_b[7] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold136 (.A(_2540_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold137 (.A(\main.demo.zic._q_tpos[11] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold138 (.A(\main.demo.zic._q_clock_count[4] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold139 (.A(\main.demo.zic._q_qpos[2] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0218_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold141 (.A(\main.demo.zic._q_rythm_count[9] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold142 (.A(\main.demo._q_prev_b[6] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold143 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold144 (.A(\main.demo._q_frame[7] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0066_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0107_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold147 (.A(\main.demo.zic._q_qpos[4] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold148 (.A(_2877_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0220_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold150 (.A(\main.demo.zic._q_tpos[2] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold151 (.A(_2761_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0206_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold153 (.A(\main.demo._q_th[6] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold154 (.A(\main.demo.zic._q_qpos[6] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0222_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold156 (.A(\main.demo.zic._q_drum_inc[2] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold157 (.A(\main.demo.zic._q_tpos[0] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold158 (.A(\main.demo.zic._q_tpos[3] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold159 (.A(\main.demo.zic._q_tpos[1] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold160 (.A(\main.demo._q_frame[14] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold161 (.A(_2513_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold162 (.A(\main.demo.zic._q_qpos[11] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold163 (.A(_2899_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0227_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold165 (.A(\main.demo._t___stage___block_3_y[2] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold166 (.A(\main.demo._t___pip_58_1_0___stage___block_3_cx[2] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold167 (.A(\main.demo.zic._q_squ_env[5] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold168 (.A(_2704_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold169 (.A(rst_n_q),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold170 (.A(_2638_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold171 (.A(\main.demo._q_speed[5] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold172 (.A(\main.demo._q_speed[9] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0084_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold174 (.A(\main.demo.zic._q_qpos[10] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold175 (.A(\main.demo.zic._q_drum_inc[3] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold176 (.A(\main.demo.zic._q_tpos[6] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold177 (.A(\main.demo._q_speed[12] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold178 (.A(_2499_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0087_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold180 (.A(\main.demo.zic._q_qpos[12] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold181 (.A(\main.demo._q_speed[10] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold182 (.A(_2489_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold183 (.A(\main.demo._q_speed[4] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold184 (.A(_2449_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0079_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0003_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0023_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold188 (.A(_2701_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold189 (.A(_2702_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold190 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold191 (.A(\main.demo.vga._q_ycount[6] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0236_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold193 (.A(\main.demo._q_speed[13] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold194 (.A(\main.demo._q_th[2] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold195 (.A(_2528_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold196 (.A(\main.demo._q_speed[14] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold197 (.A(_2510_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold198 (.A(\main.demo.vga._q_ycount[2] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold199 (.A(\main.demo.zic._q_tpos[4] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold200 (.A(\main.demo._q_frame[11] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold201 (.A(_2496_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold202 (.A(\main.demo._q_speed[11] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold203 (.A(_2493_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold204 (.A(\main.demo._q_speed[15] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold205 (.A(\main.demo._q_speed[0] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0075_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold207 (.A(\main.demo.zic._q_clock_count[1] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold208 (.A(_2642_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0160_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold210 (.A(\main.demo._q_th[3] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0035_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold212 (.A(\main.demo.zic._q_drum_inc[1] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0125_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold214 (.A(\main.demo._q_frame[1] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold215 (.A(_2434_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold216 (.A(\main.demo._q_frame[13] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold217 (.A(_2509_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold218 (.A(\main.demo.vga._q_ycount[3] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold219 (.A(\main.demo.vga._q_ycount[1] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold220 (.A(\main.demo._q_speed[6] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0081_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0022_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold223 (.A(_2537_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0001_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold225 (.A(\main.demo._q_speed[8] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold226 (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold227 (.A(\main.demo._q_frame[10] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold228 (.A(\main.demo.zic._q_squ_env[3] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold229 (.A(\main.demo._q_th[5] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold230 (.A(\main.demo.zic._q_idx[6] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold231 (.A(_2567_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold232 (.A(\main.demo._q_speed[3] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold233 (.A(\main.demo.zic._q_drum_inc[0] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold234 (.A(\main.demo._q_frame[8] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold235 (.A(_2484_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0001_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold237 (.A(\main.demo._q_frame[9] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold238 (.A(\main.demo._q_frame[2] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold239 (.A(\main.demo._q_speed[1] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0076_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold241 (.A(\main.demo._t___stage___block_3_y[1] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold242 (.A(\main.demo._t___stage___block_3_y[0] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold243 (.A(\main.demo._q_frame[0] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold244 (.A(_2427_),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold245 (.A(\main.demo.vga._q_xcount[4] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0004_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold247 (.A(\main.demo._q_frame[12] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold248 (.A(_2503_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold249 (.A(\main.demo._q_frame[8] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold250 (.A(_2175_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold251 (.A(\main.demo._q_frame[5] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold252 (.A(\main.demo._q_speed[2] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold253 (.A(\main.demo.zic._q_idx[2] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold254 (.A(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold255 (.A(\main.demo.zic._q_drum_inc[1] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold256 (.A(\main.demo._q_speed[11] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold257 (.A(\main.demo._q_speed[15] ),
    .X(net659));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_8 FILLER_22_404 ();
 sg13g2_decap_8 FILLER_22_411 ();
 sg13g2_decap_8 FILLER_22_418 ();
 sg13g2_decap_8 FILLER_22_425 ();
 sg13g2_decap_8 FILLER_22_432 ();
 sg13g2_decap_8 FILLER_22_439 ();
 sg13g2_decap_8 FILLER_22_446 ();
 sg13g2_decap_8 FILLER_22_453 ();
 sg13g2_decap_8 FILLER_22_460 ();
 sg13g2_decap_8 FILLER_22_467 ();
 sg13g2_decap_8 FILLER_22_474 ();
 sg13g2_decap_8 FILLER_22_481 ();
 sg13g2_decap_8 FILLER_22_488 ();
 sg13g2_decap_8 FILLER_22_495 ();
 sg13g2_decap_8 FILLER_22_502 ();
 sg13g2_decap_8 FILLER_22_509 ();
 sg13g2_decap_8 FILLER_22_516 ();
 sg13g2_decap_8 FILLER_22_523 ();
 sg13g2_decap_8 FILLER_22_530 ();
 sg13g2_decap_8 FILLER_22_537 ();
 sg13g2_decap_8 FILLER_22_544 ();
 sg13g2_decap_8 FILLER_22_551 ();
 sg13g2_decap_8 FILLER_22_558 ();
 sg13g2_decap_8 FILLER_22_565 ();
 sg13g2_decap_8 FILLER_22_572 ();
 sg13g2_decap_8 FILLER_22_579 ();
 sg13g2_decap_8 FILLER_22_586 ();
 sg13g2_decap_8 FILLER_22_593 ();
 sg13g2_decap_8 FILLER_22_600 ();
 sg13g2_decap_8 FILLER_22_607 ();
 sg13g2_decap_8 FILLER_22_614 ();
 sg13g2_decap_8 FILLER_22_621 ();
 sg13g2_decap_8 FILLER_22_628 ();
 sg13g2_decap_8 FILLER_22_635 ();
 sg13g2_decap_8 FILLER_22_642 ();
 sg13g2_decap_8 FILLER_22_649 ();
 sg13g2_decap_8 FILLER_22_656 ();
 sg13g2_decap_8 FILLER_22_663 ();
 sg13g2_decap_8 FILLER_22_670 ();
 sg13g2_decap_8 FILLER_22_677 ();
 sg13g2_decap_8 FILLER_22_684 ();
 sg13g2_decap_8 FILLER_22_691 ();
 sg13g2_decap_8 FILLER_22_698 ();
 sg13g2_decap_8 FILLER_22_705 ();
 sg13g2_decap_8 FILLER_22_712 ();
 sg13g2_decap_8 FILLER_22_719 ();
 sg13g2_decap_8 FILLER_22_726 ();
 sg13g2_decap_8 FILLER_22_733 ();
 sg13g2_decap_8 FILLER_22_740 ();
 sg13g2_decap_8 FILLER_22_747 ();
 sg13g2_decap_8 FILLER_22_754 ();
 sg13g2_decap_8 FILLER_22_761 ();
 sg13g2_decap_8 FILLER_22_768 ();
 sg13g2_decap_8 FILLER_22_775 ();
 sg13g2_decap_8 FILLER_22_782 ();
 sg13g2_decap_8 FILLER_22_789 ();
 sg13g2_decap_8 FILLER_22_796 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_decap_8 FILLER_22_810 ();
 sg13g2_decap_8 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_decap_8 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_838 ();
 sg13g2_decap_8 FILLER_22_845 ();
 sg13g2_decap_8 FILLER_22_852 ();
 sg13g2_fill_2 FILLER_22_859 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_4 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_286 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_307 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_4 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_339 ();
 sg13g2_decap_4 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_348 ();
 sg13g2_decap_4 FILLER_23_401 ();
 sg13g2_fill_2 FILLER_23_410 ();
 sg13g2_fill_1 FILLER_23_412 ();
 sg13g2_fill_1 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_23_472 ();
 sg13g2_decap_8 FILLER_23_479 ();
 sg13g2_decap_8 FILLER_23_486 ();
 sg13g2_decap_8 FILLER_23_493 ();
 sg13g2_decap_8 FILLER_23_500 ();
 sg13g2_decap_8 FILLER_23_507 ();
 sg13g2_decap_8 FILLER_23_514 ();
 sg13g2_decap_8 FILLER_23_521 ();
 sg13g2_decap_8 FILLER_23_528 ();
 sg13g2_decap_8 FILLER_23_535 ();
 sg13g2_decap_8 FILLER_23_542 ();
 sg13g2_decap_8 FILLER_23_549 ();
 sg13g2_decap_8 FILLER_23_556 ();
 sg13g2_decap_8 FILLER_23_563 ();
 sg13g2_decap_8 FILLER_23_570 ();
 sg13g2_decap_8 FILLER_23_577 ();
 sg13g2_decap_8 FILLER_23_584 ();
 sg13g2_decap_8 FILLER_23_591 ();
 sg13g2_decap_8 FILLER_23_598 ();
 sg13g2_decap_8 FILLER_23_605 ();
 sg13g2_decap_8 FILLER_23_612 ();
 sg13g2_decap_8 FILLER_23_619 ();
 sg13g2_decap_8 FILLER_23_626 ();
 sg13g2_decap_8 FILLER_23_633 ();
 sg13g2_decap_4 FILLER_23_640 ();
 sg13g2_fill_2 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_650 ();
 sg13g2_fill_2 FILLER_23_657 ();
 sg13g2_fill_1 FILLER_23_659 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_fill_2 FILLER_23_679 ();
 sg13g2_fill_1 FILLER_23_681 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_fill_1 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_724 ();
 sg13g2_decap_8 FILLER_23_731 ();
 sg13g2_decap_8 FILLER_23_738 ();
 sg13g2_decap_8 FILLER_23_745 ();
 sg13g2_decap_8 FILLER_23_752 ();
 sg13g2_decap_8 FILLER_23_759 ();
 sg13g2_decap_8 FILLER_23_766 ();
 sg13g2_decap_8 FILLER_23_773 ();
 sg13g2_decap_8 FILLER_23_780 ();
 sg13g2_decap_8 FILLER_23_787 ();
 sg13g2_decap_8 FILLER_23_794 ();
 sg13g2_decap_8 FILLER_23_801 ();
 sg13g2_decap_8 FILLER_23_808 ();
 sg13g2_decap_8 FILLER_23_815 ();
 sg13g2_decap_8 FILLER_23_822 ();
 sg13g2_decap_8 FILLER_23_829 ();
 sg13g2_decap_8 FILLER_23_836 ();
 sg13g2_decap_8 FILLER_23_843 ();
 sg13g2_decap_8 FILLER_23_850 ();
 sg13g2_decap_4 FILLER_23_857 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_4 FILLER_24_324 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_4 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_389 ();
 sg13g2_fill_1 FILLER_24_391 ();
 sg13g2_decap_4 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_24_419 ();
 sg13g2_decap_8 FILLER_24_445 ();
 sg13g2_fill_1 FILLER_24_452 ();
 sg13g2_fill_2 FILLER_24_474 ();
 sg13g2_fill_1 FILLER_24_476 ();
 sg13g2_fill_1 FILLER_24_482 ();
 sg13g2_decap_8 FILLER_24_491 ();
 sg13g2_decap_4 FILLER_24_498 ();
 sg13g2_decap_8 FILLER_24_507 ();
 sg13g2_decap_8 FILLER_24_514 ();
 sg13g2_decap_8 FILLER_24_521 ();
 sg13g2_decap_8 FILLER_24_528 ();
 sg13g2_decap_8 FILLER_24_545 ();
 sg13g2_decap_8 FILLER_24_552 ();
 sg13g2_decap_8 FILLER_24_559 ();
 sg13g2_decap_8 FILLER_24_566 ();
 sg13g2_decap_8 FILLER_24_573 ();
 sg13g2_decap_8 FILLER_24_580 ();
 sg13g2_decap_8 FILLER_24_587 ();
 sg13g2_decap_8 FILLER_24_594 ();
 sg13g2_decap_8 FILLER_24_601 ();
 sg13g2_decap_8 FILLER_24_608 ();
 sg13g2_decap_8 FILLER_24_615 ();
 sg13g2_decap_8 FILLER_24_622 ();
 sg13g2_decap_8 FILLER_24_629 ();
 sg13g2_decap_4 FILLER_24_636 ();
 sg13g2_fill_2 FILLER_24_640 ();
 sg13g2_fill_1 FILLER_24_673 ();
 sg13g2_decap_8 FILLER_24_692 ();
 sg13g2_decap_4 FILLER_24_699 ();
 sg13g2_fill_1 FILLER_24_703 ();
 sg13g2_decap_8 FILLER_24_726 ();
 sg13g2_fill_2 FILLER_24_737 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_fill_2 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_785 ();
 sg13g2_decap_8 FILLER_24_792 ();
 sg13g2_decap_8 FILLER_24_799 ();
 sg13g2_decap_8 FILLER_24_806 ();
 sg13g2_decap_8 FILLER_24_813 ();
 sg13g2_decap_8 FILLER_24_820 ();
 sg13g2_decap_8 FILLER_24_827 ();
 sg13g2_decap_8 FILLER_24_834 ();
 sg13g2_decap_8 FILLER_24_841 ();
 sg13g2_decap_8 FILLER_24_848 ();
 sg13g2_decap_8 FILLER_24_855 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_388 ();
 sg13g2_fill_2 FILLER_25_395 ();
 sg13g2_fill_1 FILLER_25_414 ();
 sg13g2_fill_2 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_437 ();
 sg13g2_fill_2 FILLER_25_444 ();
 sg13g2_fill_1 FILLER_25_446 ();
 sg13g2_fill_2 FILLER_25_452 ();
 sg13g2_fill_1 FILLER_25_482 ();
 sg13g2_decap_8 FILLER_25_496 ();
 sg13g2_decap_4 FILLER_25_525 ();
 sg13g2_fill_2 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_559 ();
 sg13g2_decap_8 FILLER_25_566 ();
 sg13g2_decap_8 FILLER_25_573 ();
 sg13g2_decap_8 FILLER_25_580 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_decap_8 FILLER_25_594 ();
 sg13g2_decap_8 FILLER_25_601 ();
 sg13g2_decap_8 FILLER_25_608 ();
 sg13g2_decap_8 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_622 ();
 sg13g2_decap_4 FILLER_25_629 ();
 sg13g2_fill_2 FILLER_25_641 ();
 sg13g2_fill_1 FILLER_25_643 ();
 sg13g2_fill_1 FILLER_25_671 ();
 sg13g2_decap_8 FILLER_25_699 ();
 sg13g2_decap_4 FILLER_25_706 ();
 sg13g2_fill_2 FILLER_25_726 ();
 sg13g2_decap_4 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_803 ();
 sg13g2_decap_8 FILLER_25_810 ();
 sg13g2_decap_8 FILLER_25_817 ();
 sg13g2_decap_8 FILLER_25_824 ();
 sg13g2_decap_8 FILLER_25_831 ();
 sg13g2_decap_8 FILLER_25_838 ();
 sg13g2_decap_8 FILLER_25_845 ();
 sg13g2_decap_8 FILLER_25_852 ();
 sg13g2_fill_2 FILLER_25_859 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_4 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_fill_2 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_275 ();
 sg13g2_fill_2 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_fill_2 FILLER_26_309 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_decap_4 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_decap_4 FILLER_26_354 ();
 sg13g2_fill_2 FILLER_26_358 ();
 sg13g2_fill_2 FILLER_26_389 ();
 sg13g2_fill_2 FILLER_26_409 ();
 sg13g2_fill_1 FILLER_26_411 ();
 sg13g2_fill_2 FILLER_26_418 ();
 sg13g2_fill_1 FILLER_26_434 ();
 sg13g2_fill_1 FILLER_26_446 ();
 sg13g2_fill_1 FILLER_26_464 ();
 sg13g2_fill_2 FILLER_26_486 ();
 sg13g2_decap_8 FILLER_26_493 ();
 sg13g2_decap_4 FILLER_26_500 ();
 sg13g2_decap_4 FILLER_26_517 ();
 sg13g2_decap_4 FILLER_26_526 ();
 sg13g2_fill_1 FILLER_26_530 ();
 sg13g2_fill_1 FILLER_26_543 ();
 sg13g2_fill_1 FILLER_26_557 ();
 sg13g2_fill_2 FILLER_26_563 ();
 sg13g2_fill_1 FILLER_26_575 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_fill_1 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_652 ();
 sg13g2_decap_8 FILLER_26_659 ();
 sg13g2_decap_8 FILLER_26_666 ();
 sg13g2_decap_4 FILLER_26_673 ();
 sg13g2_fill_1 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_696 ();
 sg13g2_fill_1 FILLER_26_703 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_4 FILLER_26_733 ();
 sg13g2_fill_1 FILLER_26_737 ();
 sg13g2_decap_8 FILLER_26_751 ();
 sg13g2_fill_1 FILLER_26_758 ();
 sg13g2_decap_8 FILLER_26_772 ();
 sg13g2_decap_8 FILLER_26_779 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_decap_4 FILLER_27_383 ();
 sg13g2_fill_1 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_392 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_fill_2 FILLER_27_403 ();
 sg13g2_fill_1 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_8 FILLER_27_436 ();
 sg13g2_decap_8 FILLER_27_443 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_4 FILLER_27_496 ();
 sg13g2_decap_8 FILLER_27_533 ();
 sg13g2_decap_4 FILLER_27_540 ();
 sg13g2_fill_1 FILLER_27_544 ();
 sg13g2_fill_1 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_594 ();
 sg13g2_decap_8 FILLER_27_601 ();
 sg13g2_decap_8 FILLER_27_608 ();
 sg13g2_decap_8 FILLER_27_615 ();
 sg13g2_decap_4 FILLER_27_622 ();
 sg13g2_fill_2 FILLER_27_626 ();
 sg13g2_fill_1 FILLER_27_641 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_fill_2 FILLER_27_680 ();
 sg13g2_decap_8 FILLER_27_724 ();
 sg13g2_fill_1 FILLER_27_731 ();
 sg13g2_decap_8 FILLER_27_752 ();
 sg13g2_decap_8 FILLER_27_759 ();
 sg13g2_fill_2 FILLER_27_766 ();
 sg13g2_decap_8 FILLER_27_785 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_4 FILLER_27_856 ();
 sg13g2_fill_2 FILLER_27_860 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_4 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_382 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_fill_2 FILLER_28_409 ();
 sg13g2_fill_1 FILLER_28_433 ();
 sg13g2_decap_8 FILLER_28_445 ();
 sg13g2_fill_2 FILLER_28_452 ();
 sg13g2_fill_1 FILLER_28_454 ();
 sg13g2_fill_2 FILLER_28_460 ();
 sg13g2_fill_1 FILLER_28_462 ();
 sg13g2_decap_8 FILLER_28_471 ();
 sg13g2_fill_2 FILLER_28_478 ();
 sg13g2_fill_1 FILLER_28_480 ();
 sg13g2_fill_2 FILLER_28_505 ();
 sg13g2_fill_1 FILLER_28_507 ();
 sg13g2_decap_4 FILLER_28_527 ();
 sg13g2_fill_2 FILLER_28_531 ();
 sg13g2_fill_2 FILLER_28_550 ();
 sg13g2_fill_1 FILLER_28_552 ();
 sg13g2_decap_8 FILLER_28_561 ();
 sg13g2_decap_4 FILLER_28_568 ();
 sg13g2_fill_1 FILLER_28_572 ();
 sg13g2_fill_2 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_594 ();
 sg13g2_decap_8 FILLER_28_601 ();
 sg13g2_decap_8 FILLER_28_608 ();
 sg13g2_decap_8 FILLER_28_615 ();
 sg13g2_decap_8 FILLER_28_622 ();
 sg13g2_fill_2 FILLER_28_629 ();
 sg13g2_fill_1 FILLER_28_652 ();
 sg13g2_fill_2 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_fill_2 FILLER_28_679 ();
 sg13g2_fill_1 FILLER_28_681 ();
 sg13g2_fill_2 FILLER_28_704 ();
 sg13g2_fill_1 FILLER_28_706 ();
 sg13g2_fill_2 FILLER_28_728 ();
 sg13g2_fill_1 FILLER_28_746 ();
 sg13g2_fill_1 FILLER_28_763 ();
 sg13g2_decap_4 FILLER_28_783 ();
 sg13g2_fill_2 FILLER_28_808 ();
 sg13g2_decap_8 FILLER_28_831 ();
 sg13g2_decap_8 FILLER_28_838 ();
 sg13g2_decap_8 FILLER_28_845 ();
 sg13g2_decap_8 FILLER_28_852 ();
 sg13g2_fill_2 FILLER_28_859 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_4 FILLER_29_245 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_261 ();
 sg13g2_fill_2 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_fill_2 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_decap_4 FILLER_29_312 ();
 sg13g2_fill_2 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_fill_2 FILLER_29_371 ();
 sg13g2_decap_4 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_393 ();
 sg13g2_decap_4 FILLER_29_400 ();
 sg13g2_fill_1 FILLER_29_404 ();
 sg13g2_fill_2 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_431 ();
 sg13g2_fill_1 FILLER_29_433 ();
 sg13g2_decap_8 FILLER_29_442 ();
 sg13g2_fill_1 FILLER_29_449 ();
 sg13g2_fill_1 FILLER_29_482 ();
 sg13g2_decap_8 FILLER_29_492 ();
 sg13g2_decap_4 FILLER_29_499 ();
 sg13g2_fill_1 FILLER_29_503 ();
 sg13g2_decap_4 FILLER_29_524 ();
 sg13g2_fill_1 FILLER_29_528 ();
 sg13g2_fill_1 FILLER_29_540 ();
 sg13g2_fill_2 FILLER_29_554 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_fill_1 FILLER_29_574 ();
 sg13g2_fill_1 FILLER_29_587 ();
 sg13g2_decap_8 FILLER_29_606 ();
 sg13g2_fill_2 FILLER_29_613 ();
 sg13g2_fill_1 FILLER_29_615 ();
 sg13g2_decap_8 FILLER_29_620 ();
 sg13g2_decap_4 FILLER_29_627 ();
 sg13g2_fill_1 FILLER_29_636 ();
 sg13g2_decap_8 FILLER_29_643 ();
 sg13g2_decap_4 FILLER_29_674 ();
 sg13g2_decap_8 FILLER_29_690 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_decap_8 FILLER_29_726 ();
 sg13g2_fill_1 FILLER_29_733 ();
 sg13g2_fill_1 FILLER_29_743 ();
 sg13g2_fill_2 FILLER_29_757 ();
 sg13g2_fill_1 FILLER_29_759 ();
 sg13g2_fill_2 FILLER_29_766 ();
 sg13g2_decap_8 FILLER_29_774 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_fill_2 FILLER_29_788 ();
 sg13g2_fill_1 FILLER_29_790 ();
 sg13g2_fill_2 FILLER_29_815 ();
 sg13g2_fill_1 FILLER_29_817 ();
 sg13g2_fill_2 FILLER_29_825 ();
 sg13g2_fill_1 FILLER_29_827 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_4 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_decap_4 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_405 ();
 sg13g2_fill_1 FILLER_30_412 ();
 sg13g2_decap_8 FILLER_30_439 ();
 sg13g2_decap_4 FILLER_30_446 ();
 sg13g2_decap_8 FILLER_30_471 ();
 sg13g2_fill_1 FILLER_30_478 ();
 sg13g2_decap_8 FILLER_30_496 ();
 sg13g2_decap_4 FILLER_30_503 ();
 sg13g2_fill_1 FILLER_30_507 ();
 sg13g2_fill_1 FILLER_30_512 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_4 FILLER_30_547 ();
 sg13g2_fill_2 FILLER_30_551 ();
 sg13g2_decap_8 FILLER_30_557 ();
 sg13g2_fill_1 FILLER_30_564 ();
 sg13g2_decap_4 FILLER_30_601 ();
 sg13g2_fill_1 FILLER_30_640 ();
 sg13g2_decap_4 FILLER_30_653 ();
 sg13g2_decap_8 FILLER_30_673 ();
 sg13g2_fill_1 FILLER_30_680 ();
 sg13g2_fill_2 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_fill_2 FILLER_30_700 ();
 sg13g2_decap_4 FILLER_30_723 ();
 sg13g2_decap_8 FILLER_30_747 ();
 sg13g2_decap_8 FILLER_30_754 ();
 sg13g2_fill_2 FILLER_30_761 ();
 sg13g2_fill_1 FILLER_30_763 ();
 sg13g2_fill_2 FILLER_30_769 ();
 sg13g2_decap_4 FILLER_30_790 ();
 sg13g2_fill_1 FILLER_30_794 ();
 sg13g2_fill_1 FILLER_30_822 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_fill_2 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_298 ();
 sg13g2_decap_8 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_decap_8 FILLER_31_360 ();
 sg13g2_decap_4 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_decap_4 FILLER_31_380 ();
 sg13g2_fill_2 FILLER_31_384 ();
 sg13g2_fill_2 FILLER_31_429 ();
 sg13g2_decap_4 FILLER_31_444 ();
 sg13g2_fill_2 FILLER_31_469 ();
 sg13g2_decap_4 FILLER_31_500 ();
 sg13g2_fill_2 FILLER_31_514 ();
 sg13g2_fill_1 FILLER_31_516 ();
 sg13g2_fill_1 FILLER_31_541 ();
 sg13g2_decap_8 FILLER_31_550 ();
 sg13g2_fill_2 FILLER_31_557 ();
 sg13g2_fill_2 FILLER_31_564 ();
 sg13g2_decap_8 FILLER_31_573 ();
 sg13g2_decap_4 FILLER_31_580 ();
 sg13g2_fill_2 FILLER_31_589 ();
 sg13g2_decap_4 FILLER_31_601 ();
 sg13g2_fill_2 FILLER_31_605 ();
 sg13g2_decap_8 FILLER_31_611 ();
 sg13g2_decap_8 FILLER_31_618 ();
 sg13g2_fill_1 FILLER_31_625 ();
 sg13g2_fill_1 FILLER_31_652 ();
 sg13g2_fill_1 FILLER_31_667 ();
 sg13g2_decap_4 FILLER_31_700 ();
 sg13g2_fill_2 FILLER_31_704 ();
 sg13g2_decap_8 FILLER_31_723 ();
 sg13g2_decap_8 FILLER_31_730 ();
 sg13g2_fill_1 FILLER_31_737 ();
 sg13g2_fill_2 FILLER_31_755 ();
 sg13g2_fill_1 FILLER_31_757 ();
 sg13g2_fill_2 FILLER_31_783 ();
 sg13g2_fill_1 FILLER_31_785 ();
 sg13g2_decap_8 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_806 ();
 sg13g2_decap_8 FILLER_31_813 ();
 sg13g2_decap_4 FILLER_31_820 ();
 sg13g2_fill_2 FILLER_31_824 ();
 sg13g2_decap_8 FILLER_31_842 ();
 sg13g2_decap_8 FILLER_31_849 ();
 sg13g2_decap_4 FILLER_31_856 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_4 FILLER_32_252 ();
 sg13g2_decap_4 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_299 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_decap_4 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_390 ();
 sg13g2_fill_2 FILLER_32_398 ();
 sg13g2_decap_8 FILLER_32_408 ();
 sg13g2_decap_4 FILLER_32_415 ();
 sg13g2_fill_1 FILLER_32_419 ();
 sg13g2_fill_2 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_438 ();
 sg13g2_decap_8 FILLER_32_458 ();
 sg13g2_decap_4 FILLER_32_465 ();
 sg13g2_fill_1 FILLER_32_469 ();
 sg13g2_decap_4 FILLER_32_497 ();
 sg13g2_fill_1 FILLER_32_501 ();
 sg13g2_decap_4 FILLER_32_548 ();
 sg13g2_decap_8 FILLER_32_572 ();
 sg13g2_decap_4 FILLER_32_579 ();
 sg13g2_decap_8 FILLER_32_587 ();
 sg13g2_fill_2 FILLER_32_594 ();
 sg13g2_decap_4 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_647 ();
 sg13g2_decap_8 FILLER_32_654 ();
 sg13g2_decap_8 FILLER_32_661 ();
 sg13g2_decap_8 FILLER_32_668 ();
 sg13g2_decap_8 FILLER_32_675 ();
 sg13g2_fill_1 FILLER_32_682 ();
 sg13g2_decap_8 FILLER_32_692 ();
 sg13g2_decap_4 FILLER_32_699 ();
 sg13g2_fill_1 FILLER_32_703 ();
 sg13g2_fill_2 FILLER_32_725 ();
 sg13g2_fill_1 FILLER_32_743 ();
 sg13g2_decap_4 FILLER_32_760 ();
 sg13g2_fill_2 FILLER_32_764 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_fill_2 FILLER_32_777 ();
 sg13g2_fill_1 FILLER_32_779 ();
 sg13g2_decap_8 FILLER_32_807 ();
 sg13g2_fill_2 FILLER_32_814 ();
 sg13g2_fill_1 FILLER_32_816 ();
 sg13g2_decap_4 FILLER_32_843 ();
 sg13g2_fill_2 FILLER_32_847 ();
 sg13g2_decap_4 FILLER_32_857 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_297 ();
 sg13g2_decap_4 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_decap_4 FILLER_33_362 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_fill_2 FILLER_33_416 ();
 sg13g2_decap_4 FILLER_33_426 ();
 sg13g2_decap_8 FILLER_33_443 ();
 sg13g2_decap_4 FILLER_33_450 ();
 sg13g2_fill_1 FILLER_33_454 ();
 sg13g2_fill_2 FILLER_33_464 ();
 sg13g2_decap_4 FILLER_33_486 ();
 sg13g2_fill_2 FILLER_33_490 ();
 sg13g2_fill_2 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_507 ();
 sg13g2_decap_4 FILLER_33_514 ();
 sg13g2_decap_8 FILLER_33_538 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_fill_1 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_565 ();
 sg13g2_decap_8 FILLER_33_624 ();
 sg13g2_decap_4 FILLER_33_647 ();
 sg13g2_fill_2 FILLER_33_651 ();
 sg13g2_fill_1 FILLER_33_674 ();
 sg13g2_fill_2 FILLER_33_683 ();
 sg13g2_decap_8 FILLER_33_698 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_fill_2 FILLER_33_728 ();
 sg13g2_fill_1 FILLER_33_730 ();
 sg13g2_decap_4 FILLER_33_745 ();
 sg13g2_fill_1 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_fill_2 FILLER_33_800 ();
 sg13g2_fill_1 FILLER_33_802 ();
 sg13g2_fill_2 FILLER_33_817 ();
 sg13g2_fill_2 FILLER_33_839 ();
 sg13g2_fill_1 FILLER_33_841 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_fill_2 FILLER_34_259 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_decap_4 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_decap_4 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_decap_4 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_331 ();
 sg13g2_fill_2 FILLER_34_337 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_348 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_370 ();
 sg13g2_fill_1 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_4 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_418 ();
 sg13g2_fill_1 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_34_432 ();
 sg13g2_fill_2 FILLER_34_444 ();
 sg13g2_fill_1 FILLER_34_446 ();
 sg13g2_decap_8 FILLER_34_468 ();
 sg13g2_fill_2 FILLER_34_475 ();
 sg13g2_fill_1 FILLER_34_477 ();
 sg13g2_fill_1 FILLER_34_483 ();
 sg13g2_fill_2 FILLER_34_509 ();
 sg13g2_fill_1 FILLER_34_511 ();
 sg13g2_fill_2 FILLER_34_520 ();
 sg13g2_fill_1 FILLER_34_522 ();
 sg13g2_decap_8 FILLER_34_528 ();
 sg13g2_fill_2 FILLER_34_535 ();
 sg13g2_decap_8 FILLER_34_581 ();
 sg13g2_decap_4 FILLER_34_588 ();
 sg13g2_fill_2 FILLER_34_592 ();
 sg13g2_decap_8 FILLER_34_612 ();
 sg13g2_decap_8 FILLER_34_619 ();
 sg13g2_fill_2 FILLER_34_681 ();
 sg13g2_decap_4 FILLER_34_696 ();
 sg13g2_fill_1 FILLER_34_700 ();
 sg13g2_decap_4 FILLER_34_714 ();
 sg13g2_fill_1 FILLER_34_718 ();
 sg13g2_fill_2 FILLER_34_726 ();
 sg13g2_fill_1 FILLER_34_728 ();
 sg13g2_decap_4 FILLER_34_753 ();
 sg13g2_decap_8 FILLER_34_762 ();
 sg13g2_fill_2 FILLER_34_769 ();
 sg13g2_fill_2 FILLER_34_775 ();
 sg13g2_fill_1 FILLER_34_777 ();
 sg13g2_fill_2 FILLER_34_798 ();
 sg13g2_decap_4 FILLER_34_818 ();
 sg13g2_fill_1 FILLER_34_822 ();
 sg13g2_fill_1 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_855 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_248 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_fill_1 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_295 ();
 sg13g2_decap_4 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_318 ();
 sg13g2_decap_4 FILLER_35_325 ();
 sg13g2_fill_1 FILLER_35_342 ();
 sg13g2_fill_2 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_353 ();
 sg13g2_decap_4 FILLER_35_388 ();
 sg13g2_fill_1 FILLER_35_392 ();
 sg13g2_fill_2 FILLER_35_408 ();
 sg13g2_decap_4 FILLER_35_436 ();
 sg13g2_fill_2 FILLER_35_440 ();
 sg13g2_decap_8 FILLER_35_446 ();
 sg13g2_decap_8 FILLER_35_457 ();
 sg13g2_decap_4 FILLER_35_464 ();
 sg13g2_fill_2 FILLER_35_481 ();
 sg13g2_decap_8 FILLER_35_491 ();
 sg13g2_fill_2 FILLER_35_498 ();
 sg13g2_fill_1 FILLER_35_504 ();
 sg13g2_decap_4 FILLER_35_510 ();
 sg13g2_decap_4 FILLER_35_531 ();
 sg13g2_fill_1 FILLER_35_535 ();
 sg13g2_fill_2 FILLER_35_541 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_4 FILLER_35_560 ();
 sg13g2_fill_1 FILLER_35_564 ();
 sg13g2_fill_2 FILLER_35_570 ();
 sg13g2_fill_2 FILLER_35_580 ();
 sg13g2_decap_8 FILLER_35_615 ();
 sg13g2_decap_4 FILLER_35_622 ();
 sg13g2_fill_2 FILLER_35_651 ();
 sg13g2_fill_1 FILLER_35_653 ();
 sg13g2_fill_2 FILLER_35_659 ();
 sg13g2_decap_4 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_674 ();
 sg13g2_fill_1 FILLER_35_681 ();
 sg13g2_decap_8 FILLER_35_699 ();
 sg13g2_decap_8 FILLER_35_706 ();
 sg13g2_fill_1 FILLER_35_738 ();
 sg13g2_fill_1 FILLER_35_757 ();
 sg13g2_fill_2 FILLER_35_763 ();
 sg13g2_fill_1 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_793 ();
 sg13g2_decap_4 FILLER_35_800 ();
 sg13g2_fill_1 FILLER_35_826 ();
 sg13g2_fill_2 FILLER_35_831 ();
 sg13g2_fill_2 FILLER_35_839 ();
 sg13g2_fill_1 FILLER_35_841 ();
 sg13g2_fill_2 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_245 ();
 sg13g2_decap_4 FILLER_36_251 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_decap_4 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_decap_4 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_fill_2 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_404 ();
 sg13g2_fill_2 FILLER_36_409 ();
 sg13g2_decap_8 FILLER_36_424 ();
 sg13g2_decap_4 FILLER_36_457 ();
 sg13g2_fill_2 FILLER_36_461 ();
 sg13g2_decap_4 FILLER_36_487 ();
 sg13g2_fill_2 FILLER_36_499 ();
 sg13g2_decap_8 FILLER_36_514 ();
 sg13g2_fill_2 FILLER_36_529 ();
 sg13g2_fill_1 FILLER_36_531 ();
 sg13g2_decap_8 FILLER_36_536 ();
 sg13g2_decap_4 FILLER_36_543 ();
 sg13g2_fill_1 FILLER_36_547 ();
 sg13g2_fill_2 FILLER_36_558 ();
 sg13g2_fill_1 FILLER_36_560 ();
 sg13g2_decap_4 FILLER_36_585 ();
 sg13g2_fill_2 FILLER_36_589 ();
 sg13g2_fill_1 FILLER_36_619 ();
 sg13g2_decap_8 FILLER_36_645 ();
 sg13g2_decap_4 FILLER_36_652 ();
 sg13g2_fill_1 FILLER_36_656 ();
 sg13g2_fill_1 FILLER_36_674 ();
 sg13g2_fill_2 FILLER_36_686 ();
 sg13g2_fill_1 FILLER_36_688 ();
 sg13g2_fill_1 FILLER_36_697 ();
 sg13g2_decap_8 FILLER_36_719 ();
 sg13g2_fill_1 FILLER_36_726 ();
 sg13g2_decap_8 FILLER_36_736 ();
 sg13g2_decap_4 FILLER_36_743 ();
 sg13g2_fill_2 FILLER_36_747 ();
 sg13g2_decap_8 FILLER_36_765 ();
 sg13g2_decap_4 FILLER_36_772 ();
 sg13g2_decap_4 FILLER_36_784 ();
 sg13g2_fill_2 FILLER_36_794 ();
 sg13g2_fill_1 FILLER_36_796 ();
 sg13g2_decap_4 FILLER_36_818 ();
 sg13g2_fill_2 FILLER_36_822 ();
 sg13g2_fill_1 FILLER_36_828 ();
 sg13g2_fill_1 FILLER_36_841 ();
 sg13g2_decap_8 FILLER_36_855 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_fill_2 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_281 ();
 sg13g2_decap_8 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_decap_4 FILLER_37_324 ();
 sg13g2_fill_2 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_334 ();
 sg13g2_decap_8 FILLER_37_341 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_418 ();
 sg13g2_fill_1 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_4 FILLER_37_462 ();
 sg13g2_fill_2 FILLER_37_466 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_fill_1 FILLER_37_488 ();
 sg13g2_fill_2 FILLER_37_497 ();
 sg13g2_decap_4 FILLER_37_506 ();
 sg13g2_decap_4 FILLER_37_518 ();
 sg13g2_fill_2 FILLER_37_548 ();
 sg13g2_fill_2 FILLER_37_558 ();
 sg13g2_fill_1 FILLER_37_560 ();
 sg13g2_fill_1 FILLER_37_580 ();
 sg13g2_fill_1 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_614 ();
 sg13g2_fill_1 FILLER_37_631 ();
 sg13g2_decap_4 FILLER_37_650 ();
 sg13g2_fill_1 FILLER_37_654 ();
 sg13g2_decap_8 FILLER_37_667 ();
 sg13g2_decap_4 FILLER_37_674 ();
 sg13g2_fill_1 FILLER_37_678 ();
 sg13g2_decap_8 FILLER_37_698 ();
 sg13g2_decap_4 FILLER_37_705 ();
 sg13g2_decap_4 FILLER_37_714 ();
 sg13g2_fill_2 FILLER_37_726 ();
 sg13g2_fill_1 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_741 ();
 sg13g2_fill_2 FILLER_37_760 ();
 sg13g2_decap_8 FILLER_37_790 ();
 sg13g2_fill_2 FILLER_37_813 ();
 sg13g2_fill_1 FILLER_37_815 ();
 sg13g2_fill_1 FILLER_37_837 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_245 ();
 sg13g2_decap_4 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_decap_4 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_300 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_fill_2 FILLER_38_328 ();
 sg13g2_decap_4 FILLER_38_346 ();
 sg13g2_decap_8 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_fill_2 FILLER_38_384 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_fill_1 FILLER_38_405 ();
 sg13g2_decap_4 FILLER_38_409 ();
 sg13g2_fill_1 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_419 ();
 sg13g2_fill_2 FILLER_38_426 ();
 sg13g2_decap_4 FILLER_38_436 ();
 sg13g2_fill_1 FILLER_38_444 ();
 sg13g2_fill_1 FILLER_38_477 ();
 sg13g2_fill_2 FILLER_38_512 ();
 sg13g2_fill_1 FILLER_38_514 ();
 sg13g2_decap_8 FILLER_38_519 ();
 sg13g2_fill_1 FILLER_38_526 ();
 sg13g2_decap_8 FILLER_38_536 ();
 sg13g2_decap_4 FILLER_38_543 ();
 sg13g2_fill_1 FILLER_38_547 ();
 sg13g2_fill_1 FILLER_38_560 ();
 sg13g2_decap_8 FILLER_38_569 ();
 sg13g2_fill_1 FILLER_38_576 ();
 sg13g2_fill_2 FILLER_38_582 ();
 sg13g2_decap_4 FILLER_38_589 ();
 sg13g2_fill_2 FILLER_38_593 ();
 sg13g2_decap_8 FILLER_38_615 ();
 sg13g2_decap_8 FILLER_38_622 ();
 sg13g2_fill_2 FILLER_38_629 ();
 sg13g2_fill_2 FILLER_38_648 ();
 sg13g2_fill_1 FILLER_38_650 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_fill_2 FILLER_38_670 ();
 sg13g2_fill_1 FILLER_38_672 ();
 sg13g2_fill_2 FILLER_38_683 ();
 sg13g2_fill_1 FILLER_38_685 ();
 sg13g2_fill_2 FILLER_38_690 ();
 sg13g2_fill_2 FILLER_38_701 ();
 sg13g2_fill_1 FILLER_38_726 ();
 sg13g2_fill_1 FILLER_38_747 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_4 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_793 ();
 sg13g2_fill_1 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_829 ();
 sg13g2_decap_4 FILLER_38_836 ();
 sg13g2_fill_1 FILLER_38_840 ();
 sg13g2_fill_2 FILLER_38_859 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_fill_2 FILLER_39_217 ();
 sg13g2_fill_1 FILLER_39_219 ();
 sg13g2_fill_1 FILLER_39_247 ();
 sg13g2_fill_2 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_270 ();
 sg13g2_fill_2 FILLER_39_275 ();
 sg13g2_fill_1 FILLER_39_277 ();
 sg13g2_fill_1 FILLER_39_291 ();
 sg13g2_fill_1 FILLER_39_319 ();
 sg13g2_fill_2 FILLER_39_335 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_decap_8 FILLER_39_346 ();
 sg13g2_fill_1 FILLER_39_361 ();
 sg13g2_fill_2 FILLER_39_395 ();
 sg13g2_fill_1 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_39_431 ();
 sg13g2_decap_8 FILLER_39_438 ();
 sg13g2_decap_8 FILLER_39_445 ();
 sg13g2_decap_4 FILLER_39_452 ();
 sg13g2_decap_4 FILLER_39_460 ();
 sg13g2_fill_1 FILLER_39_464 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_decap_8 FILLER_39_477 ();
 sg13g2_fill_2 FILLER_39_484 ();
 sg13g2_fill_1 FILLER_39_486 ();
 sg13g2_decap_4 FILLER_39_576 ();
 sg13g2_fill_1 FILLER_39_580 ();
 sg13g2_decap_4 FILLER_39_586 ();
 sg13g2_fill_1 FILLER_39_590 ();
 sg13g2_fill_1 FILLER_39_623 ();
 sg13g2_decap_4 FILLER_39_647 ();
 sg13g2_fill_1 FILLER_39_651 ();
 sg13g2_decap_4 FILLER_39_663 ();
 sg13g2_fill_1 FILLER_39_667 ();
 sg13g2_fill_1 FILLER_39_689 ();
 sg13g2_fill_1 FILLER_39_708 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_4 FILLER_39_728 ();
 sg13g2_decap_8 FILLER_39_737 ();
 sg13g2_fill_2 FILLER_39_744 ();
 sg13g2_fill_2 FILLER_39_764 ();
 sg13g2_fill_1 FILLER_39_766 ();
 sg13g2_decap_8 FILLER_39_783 ();
 sg13g2_decap_4 FILLER_39_790 ();
 sg13g2_decap_8 FILLER_39_802 ();
 sg13g2_decap_4 FILLER_39_809 ();
 sg13g2_fill_2 FILLER_39_813 ();
 sg13g2_fill_1 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_decap_4 FILLER_39_840 ();
 sg13g2_fill_1 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_853 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_fill_2 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_83 ();
 sg13g2_decap_8 FILLER_40_90 ();
 sg13g2_decap_8 FILLER_40_97 ();
 sg13g2_decap_8 FILLER_40_104 ();
 sg13g2_decap_8 FILLER_40_111 ();
 sg13g2_decap_8 FILLER_40_118 ();
 sg13g2_decap_8 FILLER_40_125 ();
 sg13g2_decap_8 FILLER_40_132 ();
 sg13g2_decap_8 FILLER_40_139 ();
 sg13g2_decap_8 FILLER_40_146 ();
 sg13g2_decap_8 FILLER_40_153 ();
 sg13g2_decap_8 FILLER_40_160 ();
 sg13g2_decap_8 FILLER_40_167 ();
 sg13g2_decap_8 FILLER_40_174 ();
 sg13g2_decap_8 FILLER_40_181 ();
 sg13g2_decap_8 FILLER_40_188 ();
 sg13g2_decap_8 FILLER_40_195 ();
 sg13g2_fill_1 FILLER_40_202 ();
 sg13g2_decap_8 FILLER_40_211 ();
 sg13g2_decap_8 FILLER_40_218 ();
 sg13g2_decap_4 FILLER_40_242 ();
 sg13g2_fill_1 FILLER_40_254 ();
 sg13g2_fill_2 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_262 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_2 FILLER_40_313 ();
 sg13g2_fill_1 FILLER_40_323 ();
 sg13g2_fill_2 FILLER_40_333 ();
 sg13g2_fill_1 FILLER_40_335 ();
 sg13g2_decap_8 FILLER_40_354 ();
 sg13g2_decap_8 FILLER_40_373 ();
 sg13g2_fill_2 FILLER_40_380 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_fill_1 FILLER_40_395 ();
 sg13g2_fill_2 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_406 ();
 sg13g2_fill_2 FILLER_40_415 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_501 ();
 sg13g2_decap_8 FILLER_40_508 ();
 sg13g2_decap_4 FILLER_40_515 ();
 sg13g2_fill_1 FILLER_40_519 ();
 sg13g2_fill_1 FILLER_40_537 ();
 sg13g2_fill_2 FILLER_40_551 ();
 sg13g2_decap_4 FILLER_40_571 ();
 sg13g2_fill_1 FILLER_40_575 ();
 sg13g2_decap_8 FILLER_40_662 ();
 sg13g2_fill_2 FILLER_40_669 ();
 sg13g2_decap_8 FILLER_40_676 ();
 sg13g2_decap_8 FILLER_40_683 ();
 sg13g2_fill_2 FILLER_40_690 ();
 sg13g2_decap_8 FILLER_40_697 ();
 sg13g2_decap_4 FILLER_40_704 ();
 sg13g2_fill_1 FILLER_40_708 ();
 sg13g2_fill_1 FILLER_40_721 ();
 sg13g2_fill_2 FILLER_40_734 ();
 sg13g2_fill_1 FILLER_40_736 ();
 sg13g2_fill_1 FILLER_40_742 ();
 sg13g2_fill_1 FILLER_40_752 ();
 sg13g2_fill_2 FILLER_40_764 ();
 sg13g2_fill_1 FILLER_40_766 ();
 sg13g2_decap_4 FILLER_40_789 ();
 sg13g2_fill_1 FILLER_40_793 ();
 sg13g2_fill_2 FILLER_40_834 ();
 sg13g2_fill_1 FILLER_40_836 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_4 FILLER_41_63 ();
 sg13g2_fill_2 FILLER_41_67 ();
 sg13g2_fill_2 FILLER_41_94 ();
 sg13g2_fill_2 FILLER_41_100 ();
 sg13g2_decap_8 FILLER_41_111 ();
 sg13g2_decap_8 FILLER_41_118 ();
 sg13g2_decap_8 FILLER_41_125 ();
 sg13g2_decap_8 FILLER_41_132 ();
 sg13g2_decap_8 FILLER_41_139 ();
 sg13g2_decap_8 FILLER_41_146 ();
 sg13g2_decap_8 FILLER_41_153 ();
 sg13g2_decap_8 FILLER_41_160 ();
 sg13g2_decap_8 FILLER_41_167 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_decap_4 FILLER_41_209 ();
 sg13g2_decap_8 FILLER_41_229 ();
 sg13g2_decap_4 FILLER_41_241 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_254 ();
 sg13g2_fill_1 FILLER_41_261 ();
 sg13g2_decap_8 FILLER_41_270 ();
 sg13g2_decap_8 FILLER_41_277 ();
 sg13g2_decap_4 FILLER_41_284 ();
 sg13g2_fill_1 FILLER_41_288 ();
 sg13g2_decap_8 FILLER_41_293 ();
 sg13g2_decap_4 FILLER_41_300 ();
 sg13g2_fill_1 FILLER_41_304 ();
 sg13g2_fill_2 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_331 ();
 sg13g2_fill_2 FILLER_41_363 ();
 sg13g2_fill_1 FILLER_41_365 ();
 sg13g2_decap_8 FILLER_41_370 ();
 sg13g2_fill_1 FILLER_41_385 ();
 sg13g2_fill_2 FILLER_41_409 ();
 sg13g2_fill_1 FILLER_41_411 ();
 sg13g2_fill_2 FILLER_41_424 ();
 sg13g2_decap_8 FILLER_41_431 ();
 sg13g2_decap_4 FILLER_41_438 ();
 sg13g2_fill_1 FILLER_41_442 ();
 sg13g2_decap_8 FILLER_41_456 ();
 sg13g2_decap_8 FILLER_41_463 ();
 sg13g2_decap_8 FILLER_41_478 ();
 sg13g2_fill_2 FILLER_41_542 ();
 sg13g2_fill_1 FILLER_41_544 ();
 sg13g2_decap_4 FILLER_41_561 ();
 sg13g2_fill_1 FILLER_41_565 ();
 sg13g2_decap_4 FILLER_41_578 ();
 sg13g2_fill_1 FILLER_41_582 ();
 sg13g2_decap_8 FILLER_41_598 ();
 sg13g2_decap_4 FILLER_41_620 ();
 sg13g2_fill_2 FILLER_41_642 ();
 sg13g2_fill_1 FILLER_41_644 ();
 sg13g2_decap_4 FILLER_41_672 ();
 sg13g2_fill_1 FILLER_41_676 ();
 sg13g2_fill_2 FILLER_41_685 ();
 sg13g2_fill_1 FILLER_41_687 ();
 sg13g2_fill_1 FILLER_41_708 ();
 sg13g2_fill_2 FILLER_41_725 ();
 sg13g2_fill_1 FILLER_41_727 ();
 sg13g2_decap_4 FILLER_41_733 ();
 sg13g2_fill_1 FILLER_41_737 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_4 FILLER_41_784 ();
 sg13g2_fill_1 FILLER_41_796 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_4 FILLER_41_812 ();
 sg13g2_fill_1 FILLER_41_816 ();
 sg13g2_fill_2 FILLER_41_825 ();
 sg13g2_fill_1 FILLER_41_827 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_fill_2 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_89 ();
 sg13g2_decap_8 FILLER_42_117 ();
 sg13g2_decap_8 FILLER_42_124 ();
 sg13g2_decap_8 FILLER_42_131 ();
 sg13g2_decap_8 FILLER_42_138 ();
 sg13g2_decap_8 FILLER_42_145 ();
 sg13g2_decap_8 FILLER_42_152 ();
 sg13g2_decap_8 FILLER_42_159 ();
 sg13g2_decap_8 FILLER_42_166 ();
 sg13g2_decap_8 FILLER_42_173 ();
 sg13g2_decap_4 FILLER_42_180 ();
 sg13g2_fill_1 FILLER_42_184 ();
 sg13g2_fill_1 FILLER_42_198 ();
 sg13g2_decap_4 FILLER_42_222 ();
 sg13g2_decap_8 FILLER_42_241 ();
 sg13g2_fill_2 FILLER_42_260 ();
 sg13g2_decap_4 FILLER_42_270 ();
 sg13g2_fill_2 FILLER_42_274 ();
 sg13g2_fill_2 FILLER_42_281 ();
 sg13g2_decap_4 FILLER_42_297 ();
 sg13g2_decap_8 FILLER_42_306 ();
 sg13g2_fill_2 FILLER_42_313 ();
 sg13g2_fill_1 FILLER_42_315 ();
 sg13g2_fill_2 FILLER_42_321 ();
 sg13g2_fill_1 FILLER_42_323 ();
 sg13g2_decap_8 FILLER_42_328 ();
 sg13g2_decap_4 FILLER_42_335 ();
 sg13g2_fill_1 FILLER_42_339 ();
 sg13g2_fill_1 FILLER_42_348 ();
 sg13g2_decap_4 FILLER_42_353 ();
 sg13g2_fill_2 FILLER_42_357 ();
 sg13g2_fill_2 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_2 FILLER_42_433 ();
 sg13g2_decap_4 FILLER_42_487 ();
 sg13g2_fill_2 FILLER_42_491 ();
 sg13g2_decap_8 FILLER_42_506 ();
 sg13g2_fill_1 FILLER_42_513 ();
 sg13g2_fill_2 FILLER_42_533 ();
 sg13g2_fill_2 FILLER_42_554 ();
 sg13g2_fill_1 FILLER_42_556 ();
 sg13g2_fill_2 FILLER_42_566 ();
 sg13g2_decap_4 FILLER_42_600 ();
 sg13g2_fill_2 FILLER_42_604 ();
 sg13g2_fill_1 FILLER_42_634 ();
 sg13g2_fill_2 FILLER_42_641 ();
 sg13g2_decap_8 FILLER_42_663 ();
 sg13g2_decap_4 FILLER_42_670 ();
 sg13g2_decap_4 FILLER_42_687 ();
 sg13g2_fill_1 FILLER_42_691 ();
 sg13g2_decap_8 FILLER_42_702 ();
 sg13g2_fill_2 FILLER_42_709 ();
 sg13g2_fill_2 FILLER_42_741 ();
 sg13g2_fill_1 FILLER_42_759 ();
 sg13g2_decap_8 FILLER_42_768 ();
 sg13g2_fill_1 FILLER_42_775 ();
 sg13g2_fill_1 FILLER_42_793 ();
 sg13g2_decap_8 FILLER_42_820 ();
 sg13g2_fill_1 FILLER_42_827 ();
 sg13g2_fill_1 FILLER_42_833 ();
 sg13g2_decap_8 FILLER_42_842 ();
 sg13g2_fill_1 FILLER_42_849 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_fill_2 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_142 ();
 sg13g2_decap_8 FILLER_43_149 ();
 sg13g2_decap_8 FILLER_43_156 ();
 sg13g2_decap_8 FILLER_43_163 ();
 sg13g2_decap_8 FILLER_43_170 ();
 sg13g2_decap_8 FILLER_43_177 ();
 sg13g2_decap_8 FILLER_43_184 ();
 sg13g2_decap_4 FILLER_43_191 ();
 sg13g2_decap_4 FILLER_43_199 ();
 sg13g2_fill_2 FILLER_43_208 ();
 sg13g2_fill_2 FILLER_43_215 ();
 sg13g2_fill_1 FILLER_43_217 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_fill_2 FILLER_43_252 ();
 sg13g2_fill_1 FILLER_43_273 ();
 sg13g2_decap_4 FILLER_43_305 ();
 sg13g2_fill_2 FILLER_43_309 ();
 sg13g2_fill_2 FILLER_43_319 ();
 sg13g2_decap_8 FILLER_43_344 ();
 sg13g2_decap_4 FILLER_43_351 ();
 sg13g2_fill_1 FILLER_43_355 ();
 sg13g2_decap_4 FILLER_43_368 ();
 sg13g2_fill_2 FILLER_43_372 ();
 sg13g2_decap_8 FILLER_43_379 ();
 sg13g2_fill_1 FILLER_43_386 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_decap_8 FILLER_43_409 ();
 sg13g2_fill_2 FILLER_43_416 ();
 sg13g2_decap_8 FILLER_43_433 ();
 sg13g2_decap_8 FILLER_43_440 ();
 sg13g2_fill_1 FILLER_43_447 ();
 sg13g2_decap_8 FILLER_43_452 ();
 sg13g2_decap_4 FILLER_43_459 ();
 sg13g2_fill_1 FILLER_43_463 ();
 sg13g2_decap_8 FILLER_43_480 ();
 sg13g2_fill_1 FILLER_43_487 ();
 sg13g2_decap_8 FILLER_43_501 ();
 sg13g2_decap_4 FILLER_43_508 ();
 sg13g2_fill_2 FILLER_43_512 ();
 sg13g2_fill_1 FILLER_43_540 ();
 sg13g2_fill_1 FILLER_43_545 ();
 sg13g2_fill_1 FILLER_43_556 ();
 sg13g2_fill_1 FILLER_43_563 ();
 sg13g2_fill_2 FILLER_43_576 ();
 sg13g2_fill_1 FILLER_43_578 ();
 sg13g2_fill_1 FILLER_43_592 ();
 sg13g2_decap_4 FILLER_43_601 ();
 sg13g2_fill_2 FILLER_43_623 ();
 sg13g2_fill_1 FILLER_43_625 ();
 sg13g2_fill_2 FILLER_43_632 ();
 sg13g2_decap_4 FILLER_43_651 ();
 sg13g2_fill_1 FILLER_43_655 ();
 sg13g2_fill_2 FILLER_43_669 ();
 sg13g2_fill_1 FILLER_43_671 ();
 sg13g2_fill_2 FILLER_43_685 ();
 sg13g2_fill_2 FILLER_43_707 ();
 sg13g2_fill_1 FILLER_43_709 ();
 sg13g2_decap_8 FILLER_43_730 ();
 sg13g2_decap_8 FILLER_43_737 ();
 sg13g2_decap_8 FILLER_43_760 ();
 sg13g2_decap_8 FILLER_43_767 ();
 sg13g2_fill_2 FILLER_43_778 ();
 sg13g2_fill_1 FILLER_43_792 ();
 sg13g2_decap_4 FILLER_43_796 ();
 sg13g2_fill_1 FILLER_43_800 ();
 sg13g2_decap_8 FILLER_43_809 ();
 sg13g2_fill_1 FILLER_43_816 ();
 sg13g2_fill_1 FILLER_43_823 ();
 sg13g2_fill_2 FILLER_43_834 ();
 sg13g2_decap_4 FILLER_43_856 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_9 ();
 sg13g2_fill_2 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_146 ();
 sg13g2_decap_8 FILLER_44_153 ();
 sg13g2_decap_8 FILLER_44_160 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_decap_8 FILLER_44_174 ();
 sg13g2_decap_4 FILLER_44_181 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_fill_2 FILLER_44_196 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_decap_4 FILLER_44_245 ();
 sg13g2_fill_2 FILLER_44_249 ();
 sg13g2_decap_4 FILLER_44_254 ();
 sg13g2_fill_1 FILLER_44_258 ();
 sg13g2_decap_8 FILLER_44_264 ();
 sg13g2_decap_8 FILLER_44_271 ();
 sg13g2_fill_2 FILLER_44_278 ();
 sg13g2_fill_2 FILLER_44_297 ();
 sg13g2_fill_1 FILLER_44_299 ();
 sg13g2_decap_4 FILLER_44_328 ();
 sg13g2_fill_1 FILLER_44_352 ();
 sg13g2_fill_2 FILLER_44_380 ();
 sg13g2_decap_4 FILLER_44_433 ();
 sg13g2_decap_4 FILLER_44_463 ();
 sg13g2_fill_1 FILLER_44_467 ();
 sg13g2_decap_4 FILLER_44_509 ();
 sg13g2_fill_1 FILLER_44_521 ();
 sg13g2_fill_2 FILLER_44_526 ();
 sg13g2_fill_1 FILLER_44_528 ();
 sg13g2_decap_4 FILLER_44_596 ();
 sg13g2_fill_2 FILLER_44_600 ();
 sg13g2_decap_8 FILLER_44_610 ();
 sg13g2_decap_8 FILLER_44_617 ();
 sg13g2_fill_2 FILLER_44_624 ();
 sg13g2_fill_1 FILLER_44_626 ();
 sg13g2_fill_1 FILLER_44_640 ();
 sg13g2_decap_8 FILLER_44_653 ();
 sg13g2_decap_4 FILLER_44_660 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_fill_1 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_697 ();
 sg13g2_fill_1 FILLER_44_704 ();
 sg13g2_decap_4 FILLER_44_723 ();
 sg13g2_fill_2 FILLER_44_727 ();
 sg13g2_decap_4 FILLER_44_741 ();
 sg13g2_fill_1 FILLER_44_794 ();
 sg13g2_decap_4 FILLER_44_811 ();
 sg13g2_fill_2 FILLER_44_815 ();
 sg13g2_fill_2 FILLER_44_838 ();
 sg13g2_fill_1 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_853 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_4 ();
 sg13g2_fill_1 FILLER_45_42 ();
 sg13g2_fill_2 FILLER_45_134 ();
 sg13g2_fill_1 FILLER_45_136 ();
 sg13g2_decap_8 FILLER_45_150 ();
 sg13g2_decap_8 FILLER_45_157 ();
 sg13g2_decap_8 FILLER_45_164 ();
 sg13g2_decap_4 FILLER_45_171 ();
 sg13g2_decap_4 FILLER_45_201 ();
 sg13g2_fill_2 FILLER_45_218 ();
 sg13g2_decap_8 FILLER_45_240 ();
 sg13g2_fill_2 FILLER_45_272 ();
 sg13g2_decap_4 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_319 ();
 sg13g2_decap_4 FILLER_45_326 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_fill_1 FILLER_45_365 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_4 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_400 ();
 sg13g2_decap_8 FILLER_45_407 ();
 sg13g2_fill_2 FILLER_45_414 ();
 sg13g2_decap_8 FILLER_45_443 ();
 sg13g2_decap_8 FILLER_45_450 ();
 sg13g2_decap_8 FILLER_45_457 ();
 sg13g2_fill_2 FILLER_45_464 ();
 sg13g2_fill_1 FILLER_45_466 ();
 sg13g2_fill_2 FILLER_45_494 ();
 sg13g2_fill_2 FILLER_45_501 ();
 sg13g2_fill_1 FILLER_45_503 ();
 sg13g2_fill_1 FILLER_45_514 ();
 sg13g2_fill_2 FILLER_45_535 ();
 sg13g2_fill_1 FILLER_45_537 ();
 sg13g2_fill_2 FILLER_45_563 ();
 sg13g2_fill_1 FILLER_45_565 ();
 sg13g2_fill_2 FILLER_45_592 ();
 sg13g2_fill_1 FILLER_45_594 ();
 sg13g2_decap_8 FILLER_45_621 ();
 sg13g2_fill_2 FILLER_45_628 ();
 sg13g2_fill_1 FILLER_45_630 ();
 sg13g2_decap_8 FILLER_45_642 ();
 sg13g2_decap_4 FILLER_45_666 ();
 sg13g2_fill_2 FILLER_45_670 ();
 sg13g2_decap_8 FILLER_45_676 ();
 sg13g2_fill_2 FILLER_45_683 ();
 sg13g2_decap_4 FILLER_45_703 ();
 sg13g2_fill_2 FILLER_45_720 ();
 sg13g2_fill_1 FILLER_45_722 ();
 sg13g2_fill_2 FILLER_45_740 ();
 sg13g2_fill_1 FILLER_45_750 ();
 sg13g2_decap_4 FILLER_45_759 ();
 sg13g2_fill_2 FILLER_45_763 ();
 sg13g2_fill_1 FILLER_45_769 ();
 sg13g2_decap_8 FILLER_45_786 ();
 sg13g2_fill_2 FILLER_45_793 ();
 sg13g2_fill_1 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_806 ();
 sg13g2_decap_4 FILLER_45_813 ();
 sg13g2_fill_1 FILLER_45_817 ();
 sg13g2_fill_1 FILLER_45_823 ();
 sg13g2_decap_8 FILLER_45_832 ();
 sg13g2_fill_2 FILLER_45_839 ();
 sg13g2_fill_1 FILLER_45_841 ();
 sg13g2_fill_2 FILLER_45_846 ();
 sg13g2_decap_4 FILLER_45_856 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_16 ();
 sg13g2_fill_2 FILLER_46_21 ();
 sg13g2_fill_1 FILLER_46_55 ();
 sg13g2_fill_2 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_157 ();
 sg13g2_decap_8 FILLER_46_164 ();
 sg13g2_decap_8 FILLER_46_171 ();
 sg13g2_fill_1 FILLER_46_178 ();
 sg13g2_decap_4 FILLER_46_231 ();
 sg13g2_fill_1 FILLER_46_235 ();
 sg13g2_decap_8 FILLER_46_272 ();
 sg13g2_decap_4 FILLER_46_279 ();
 sg13g2_decap_8 FILLER_46_288 ();
 sg13g2_decap_8 FILLER_46_295 ();
 sg13g2_fill_2 FILLER_46_302 ();
 sg13g2_decap_4 FILLER_46_319 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_372 ();
 sg13g2_fill_2 FILLER_46_379 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_2 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_46_414 ();
 sg13g2_fill_2 FILLER_46_421 ();
 sg13g2_fill_2 FILLER_46_475 ();
 sg13g2_decap_8 FILLER_46_502 ();
 sg13g2_decap_8 FILLER_46_521 ();
 sg13g2_fill_1 FILLER_46_528 ();
 sg13g2_fill_2 FILLER_46_537 ();
 sg13g2_fill_1 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_565 ();
 sg13g2_decap_8 FILLER_46_592 ();
 sg13g2_decap_8 FILLER_46_599 ();
 sg13g2_decap_4 FILLER_46_614 ();
 sg13g2_fill_2 FILLER_46_618 ();
 sg13g2_fill_2 FILLER_46_646 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_4 FILLER_46_679 ();
 sg13g2_fill_1 FILLER_46_683 ();
 sg13g2_decap_8 FILLER_46_703 ();
 sg13g2_fill_1 FILLER_46_710 ();
 sg13g2_decap_8 FILLER_46_719 ();
 sg13g2_decap_4 FILLER_46_726 ();
 sg13g2_fill_2 FILLER_46_730 ();
 sg13g2_fill_1 FILLER_46_747 ();
 sg13g2_fill_1 FILLER_46_753 ();
 sg13g2_fill_2 FILLER_46_771 ();
 sg13g2_decap_8 FILLER_46_778 ();
 sg13g2_fill_1 FILLER_46_785 ();
 sg13g2_fill_2 FILLER_46_823 ();
 sg13g2_fill_1 FILLER_46_825 ();
 sg13g2_decap_4 FILLER_46_839 ();
 sg13g2_fill_2 FILLER_46_859 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_16 ();
 sg13g2_fill_2 FILLER_47_77 ();
 sg13g2_fill_1 FILLER_47_79 ();
 sg13g2_fill_2 FILLER_47_111 ();
 sg13g2_fill_2 FILLER_47_131 ();
 sg13g2_fill_1 FILLER_47_133 ();
 sg13g2_fill_2 FILLER_47_148 ();
 sg13g2_decap_8 FILLER_47_195 ();
 sg13g2_fill_2 FILLER_47_202 ();
 sg13g2_fill_1 FILLER_47_204 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_fill_2 FILLER_47_238 ();
 sg13g2_fill_2 FILLER_47_244 ();
 sg13g2_fill_1 FILLER_47_246 ();
 sg13g2_decap_8 FILLER_47_251 ();
 sg13g2_fill_1 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_264 ();
 sg13g2_fill_2 FILLER_47_369 ();
 sg13g2_fill_1 FILLER_47_371 ();
 sg13g2_fill_2 FILLER_47_389 ();
 sg13g2_fill_2 FILLER_47_396 ();
 sg13g2_fill_1 FILLER_47_398 ();
 sg13g2_fill_2 FILLER_47_433 ();
 sg13g2_decap_4 FILLER_47_439 ();
 sg13g2_fill_1 FILLER_47_443 ();
 sg13g2_fill_2 FILLER_47_452 ();
 sg13g2_fill_1 FILLER_47_462 ();
 sg13g2_decap_4 FILLER_47_480 ();
 sg13g2_fill_1 FILLER_47_484 ();
 sg13g2_decap_4 FILLER_47_493 ();
 sg13g2_fill_2 FILLER_47_497 ();
 sg13g2_fill_1 FILLER_47_515 ();
 sg13g2_fill_2 FILLER_47_537 ();
 sg13g2_fill_2 FILLER_47_544 ();
 sg13g2_decap_8 FILLER_47_558 ();
 sg13g2_decap_8 FILLER_47_565 ();
 sg13g2_fill_2 FILLER_47_572 ();
 sg13g2_decap_8 FILLER_47_578 ();
 sg13g2_decap_8 FILLER_47_585 ();
 sg13g2_fill_2 FILLER_47_592 ();
 sg13g2_decap_8 FILLER_47_639 ();
 sg13g2_decap_4 FILLER_47_646 ();
 sg13g2_decap_4 FILLER_47_658 ();
 sg13g2_fill_2 FILLER_47_680 ();
 sg13g2_fill_2 FILLER_47_699 ();
 sg13g2_fill_1 FILLER_47_701 ();
 sg13g2_decap_8 FILLER_47_720 ();
 sg13g2_fill_1 FILLER_47_727 ();
 sg13g2_decap_4 FILLER_47_747 ();
 sg13g2_decap_8 FILLER_47_754 ();
 sg13g2_fill_1 FILLER_47_761 ();
 sg13g2_decap_4 FILLER_47_771 ();
 sg13g2_fill_1 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_decap_4 FILLER_47_814 ();
 sg13g2_fill_1 FILLER_47_818 ();
 sg13g2_fill_2 FILLER_47_836 ();
 sg13g2_fill_1 FILLER_47_838 ();
 sg13g2_fill_2 FILLER_47_859 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_4 ();
 sg13g2_fill_1 FILLER_48_53 ();
 sg13g2_fill_2 FILLER_48_71 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_210 ();
 sg13g2_fill_2 FILLER_48_219 ();
 sg13g2_fill_1 FILLER_48_221 ();
 sg13g2_fill_2 FILLER_48_274 ();
 sg13g2_fill_1 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_286 ();
 sg13g2_decap_8 FILLER_48_293 ();
 sg13g2_fill_2 FILLER_48_300 ();
 sg13g2_decap_8 FILLER_48_306 ();
 sg13g2_decap_8 FILLER_48_313 ();
 sg13g2_decap_8 FILLER_48_320 ();
 sg13g2_fill_1 FILLER_48_327 ();
 sg13g2_decap_8 FILLER_48_332 ();
 sg13g2_decap_8 FILLER_48_339 ();
 sg13g2_decap_8 FILLER_48_346 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_fill_1 FILLER_48_364 ();
 sg13g2_decap_4 FILLER_48_417 ();
 sg13g2_fill_2 FILLER_48_421 ();
 sg13g2_fill_1 FILLER_48_462 ();
 sg13g2_fill_2 FILLER_48_489 ();
 sg13g2_fill_1 FILLER_48_491 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_fill_2 FILLER_48_504 ();
 sg13g2_fill_1 FILLER_48_506 ();
 sg13g2_fill_2 FILLER_48_510 ();
 sg13g2_decap_4 FILLER_48_520 ();
 sg13g2_fill_1 FILLER_48_524 ();
 sg13g2_fill_2 FILLER_48_533 ();
 sg13g2_decap_8 FILLER_48_551 ();
 sg13g2_decap_4 FILLER_48_558 ();
 sg13g2_fill_1 FILLER_48_562 ();
 sg13g2_fill_2 FILLER_48_619 ();
 sg13g2_fill_1 FILLER_48_621 ();
 sg13g2_decap_4 FILLER_48_648 ();
 sg13g2_decap_8 FILLER_48_669 ();
 sg13g2_decap_8 FILLER_48_676 ();
 sg13g2_fill_1 FILLER_48_683 ();
 sg13g2_decap_8 FILLER_48_701 ();
 sg13g2_fill_2 FILLER_48_708 ();
 sg13g2_fill_1 FILLER_48_710 ();
 sg13g2_decap_8 FILLER_48_724 ();
 sg13g2_fill_2 FILLER_48_731 ();
 sg13g2_decap_4 FILLER_48_751 ();
 sg13g2_fill_1 FILLER_48_755 ();
 sg13g2_decap_8 FILLER_48_779 ();
 sg13g2_decap_8 FILLER_48_786 ();
 sg13g2_fill_2 FILLER_48_793 ();
 sg13g2_fill_1 FILLER_48_795 ();
 sg13g2_decap_4 FILLER_48_813 ();
 sg13g2_fill_1 FILLER_48_817 ();
 sg13g2_fill_2 FILLER_48_826 ();
 sg13g2_decap_4 FILLER_48_833 ();
 sg13g2_decap_4 FILLER_48_858 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_28 ();
 sg13g2_fill_1 FILLER_49_30 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_fill_1 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_86 ();
 sg13g2_fill_1 FILLER_49_88 ();
 sg13g2_fill_2 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_178 ();
 sg13g2_decap_8 FILLER_49_185 ();
 sg13g2_decap_8 FILLER_49_192 ();
 sg13g2_decap_8 FILLER_49_199 ();
 sg13g2_decap_8 FILLER_49_206 ();
 sg13g2_fill_2 FILLER_49_213 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_1 FILLER_49_258 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_fill_1 FILLER_49_430 ();
 sg13g2_fill_2 FILLER_49_457 ();
 sg13g2_fill_2 FILLER_49_485 ();
 sg13g2_fill_1 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_514 ();
 sg13g2_decap_8 FILLER_49_521 ();
 sg13g2_decap_4 FILLER_49_528 ();
 sg13g2_fill_2 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_586 ();
 sg13g2_fill_2 FILLER_49_593 ();
 sg13g2_decap_8 FILLER_49_633 ();
 sg13g2_decap_8 FILLER_49_640 ();
 sg13g2_fill_2 FILLER_49_647 ();
 sg13g2_fill_1 FILLER_49_649 ();
 sg13g2_fill_1 FILLER_49_663 ();
 sg13g2_decap_4 FILLER_49_668 ();
 sg13g2_fill_2 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_682 ();
 sg13g2_decap_4 FILLER_49_689 ();
 sg13g2_fill_2 FILLER_49_693 ();
 sg13g2_decap_4 FILLER_49_705 ();
 sg13g2_fill_1 FILLER_49_730 ();
 sg13g2_fill_2 FILLER_49_761 ();
 sg13g2_fill_1 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_778 ();
 sg13g2_decap_8 FILLER_49_785 ();
 sg13g2_fill_2 FILLER_49_792 ();
 sg13g2_fill_1 FILLER_49_840 ();
 sg13g2_fill_2 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_11 ();
 sg13g2_fill_2 FILLER_50_43 ();
 sg13g2_fill_2 FILLER_50_62 ();
 sg13g2_fill_1 FILLER_50_64 ();
 sg13g2_fill_2 FILLER_50_88 ();
 sg13g2_fill_2 FILLER_50_120 ();
 sg13g2_fill_1 FILLER_50_122 ();
 sg13g2_decap_4 FILLER_50_128 ();
 sg13g2_decap_8 FILLER_50_151 ();
 sg13g2_fill_2 FILLER_50_158 ();
 sg13g2_fill_1 FILLER_50_160 ();
 sg13g2_decap_8 FILLER_50_178 ();
 sg13g2_fill_1 FILLER_50_185 ();
 sg13g2_fill_1 FILLER_50_190 ();
 sg13g2_decap_8 FILLER_50_199 ();
 sg13g2_fill_1 FILLER_50_206 ();
 sg13g2_decap_8 FILLER_50_248 ();
 sg13g2_fill_1 FILLER_50_255 ();
 sg13g2_decap_8 FILLER_50_265 ();
 sg13g2_fill_2 FILLER_50_272 ();
 sg13g2_decap_4 FILLER_50_287 ();
 sg13g2_fill_1 FILLER_50_291 ();
 sg13g2_fill_1 FILLER_50_301 ();
 sg13g2_decap_4 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_326 ();
 sg13g2_decap_4 FILLER_50_331 ();
 sg13g2_fill_1 FILLER_50_335 ();
 sg13g2_decap_4 FILLER_50_341 ();
 sg13g2_fill_2 FILLER_50_349 ();
 sg13g2_fill_1 FILLER_50_351 ();
 sg13g2_decap_8 FILLER_50_382 ();
 sg13g2_decap_4 FILLER_50_389 ();
 sg13g2_fill_1 FILLER_50_402 ();
 sg13g2_fill_2 FILLER_50_412 ();
 sg13g2_fill_1 FILLER_50_414 ();
 sg13g2_decap_8 FILLER_50_423 ();
 sg13g2_decap_4 FILLER_50_430 ();
 sg13g2_fill_1 FILLER_50_441 ();
 sg13g2_decap_8 FILLER_50_446 ();
 sg13g2_fill_2 FILLER_50_453 ();
 sg13g2_fill_2 FILLER_50_467 ();
 sg13g2_fill_1 FILLER_50_469 ();
 sg13g2_decap_4 FILLER_50_474 ();
 sg13g2_fill_2 FILLER_50_478 ();
 sg13g2_decap_8 FILLER_50_484 ();
 sg13g2_decap_8 FILLER_50_491 ();
 sg13g2_decap_8 FILLER_50_524 ();
 sg13g2_fill_1 FILLER_50_531 ();
 sg13g2_decap_8 FILLER_50_558 ();
 sg13g2_decap_4 FILLER_50_565 ();
 sg13g2_fill_1 FILLER_50_569 ();
 sg13g2_decap_8 FILLER_50_574 ();
 sg13g2_fill_1 FILLER_50_581 ();
 sg13g2_decap_8 FILLER_50_615 ();
 sg13g2_fill_1 FILLER_50_622 ();
 sg13g2_decap_8 FILLER_50_639 ();
 sg13g2_fill_1 FILLER_50_646 ();
 sg13g2_fill_1 FILLER_50_691 ();
 sg13g2_fill_1 FILLER_50_714 ();
 sg13g2_fill_2 FILLER_50_720 ();
 sg13g2_decap_8 FILLER_50_727 ();
 sg13g2_decap_4 FILLER_50_734 ();
 sg13g2_fill_2 FILLER_50_738 ();
 sg13g2_decap_8 FILLER_50_756 ();
 sg13g2_fill_2 FILLER_50_789 ();
 sg13g2_fill_1 FILLER_50_816 ();
 sg13g2_fill_2 FILLER_50_822 ();
 sg13g2_decap_4 FILLER_50_831 ();
 sg13g2_fill_2 FILLER_50_835 ();
 sg13g2_fill_2 FILLER_50_842 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_13 ();
 sg13g2_decap_4 FILLER_51_20 ();
 sg13g2_decap_4 FILLER_51_55 ();
 sg13g2_fill_1 FILLER_51_87 ();
 sg13g2_fill_2 FILLER_51_92 ();
 sg13g2_fill_2 FILLER_51_103 ();
 sg13g2_fill_1 FILLER_51_105 ();
 sg13g2_fill_2 FILLER_51_126 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_decap_4 FILLER_51_156 ();
 sg13g2_fill_1 FILLER_51_160 ();
 sg13g2_fill_2 FILLER_51_178 ();
 sg13g2_fill_2 FILLER_51_206 ();
 sg13g2_fill_1 FILLER_51_208 ();
 sg13g2_fill_2 FILLER_51_230 ();
 sg13g2_decap_4 FILLER_51_245 ();
 sg13g2_fill_2 FILLER_51_292 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_fill_2 FILLER_51_360 ();
 sg13g2_fill_1 FILLER_51_362 ();
 sg13g2_fill_1 FILLER_51_399 ();
 sg13g2_fill_2 FILLER_51_411 ();
 sg13g2_fill_1 FILLER_51_413 ();
 sg13g2_fill_1 FILLER_51_422 ();
 sg13g2_fill_1 FILLER_51_445 ();
 sg13g2_fill_1 FILLER_51_468 ();
 sg13g2_decap_8 FILLER_51_495 ();
 sg13g2_fill_1 FILLER_51_502 ();
 sg13g2_decap_8 FILLER_51_535 ();
 sg13g2_decap_4 FILLER_51_551 ();
 sg13g2_fill_1 FILLER_51_602 ();
 sg13g2_decap_4 FILLER_51_619 ();
 sg13g2_decap_8 FILLER_51_640 ();
 sg13g2_fill_2 FILLER_51_652 ();
 sg13g2_fill_2 FILLER_51_666 ();
 sg13g2_fill_1 FILLER_51_668 ();
 sg13g2_fill_1 FILLER_51_676 ();
 sg13g2_fill_1 FILLER_51_687 ();
 sg13g2_fill_2 FILLER_51_703 ();
 sg13g2_decap_8 FILLER_51_734 ();
 sg13g2_decap_4 FILLER_51_741 ();
 sg13g2_fill_1 FILLER_51_745 ();
 sg13g2_fill_2 FILLER_51_762 ();
 sg13g2_fill_2 FILLER_51_772 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_decap_8 FILLER_51_786 ();
 sg13g2_decap_4 FILLER_51_793 ();
 sg13g2_fill_1 FILLER_51_797 ();
 sg13g2_fill_2 FILLER_51_803 ();
 sg13g2_fill_2 FILLER_51_818 ();
 sg13g2_fill_1 FILLER_51_836 ();
 sg13g2_decap_8 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_27 ();
 sg13g2_fill_2 FILLER_52_51 ();
 sg13g2_fill_1 FILLER_52_82 ();
 sg13g2_decap_8 FILLER_52_87 ();
 sg13g2_fill_1 FILLER_52_94 ();
 sg13g2_fill_2 FILLER_52_108 ();
 sg13g2_fill_1 FILLER_52_114 ();
 sg13g2_fill_2 FILLER_52_128 ();
 sg13g2_fill_1 FILLER_52_135 ();
 sg13g2_decap_4 FILLER_52_169 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_fill_2 FILLER_52_206 ();
 sg13g2_decap_4 FILLER_52_230 ();
 sg13g2_fill_1 FILLER_52_234 ();
 sg13g2_fill_2 FILLER_52_238 ();
 sg13g2_fill_1 FILLER_52_240 ();
 sg13g2_fill_1 FILLER_52_251 ();
 sg13g2_fill_2 FILLER_52_260 ();
 sg13g2_fill_2 FILLER_52_271 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_decap_4 FILLER_52_285 ();
 sg13g2_fill_1 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_300 ();
 sg13g2_decap_4 FILLER_52_305 ();
 sg13g2_fill_1 FILLER_52_314 ();
 sg13g2_fill_1 FILLER_52_324 ();
 sg13g2_decap_4 FILLER_52_338 ();
 sg13g2_decap_8 FILLER_52_347 ();
 sg13g2_fill_2 FILLER_52_354 ();
 sg13g2_fill_2 FILLER_52_369 ();
 sg13g2_fill_2 FILLER_52_389 ();
 sg13g2_fill_1 FILLER_52_391 ();
 sg13g2_fill_2 FILLER_52_397 ();
 sg13g2_fill_1 FILLER_52_399 ();
 sg13g2_decap_4 FILLER_52_408 ();
 sg13g2_fill_2 FILLER_52_412 ();
 sg13g2_fill_2 FILLER_52_422 ();
 sg13g2_fill_1 FILLER_52_424 ();
 sg13g2_fill_2 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_52_442 ();
 sg13g2_fill_2 FILLER_52_449 ();
 sg13g2_fill_2 FILLER_52_464 ();
 sg13g2_decap_4 FILLER_52_496 ();
 sg13g2_fill_1 FILLER_52_529 ();
 sg13g2_fill_1 FILLER_52_534 ();
 sg13g2_decap_8 FILLER_52_561 ();
 sg13g2_decap_4 FILLER_52_568 ();
 sg13g2_fill_2 FILLER_52_582 ();
 sg13g2_fill_1 FILLER_52_584 ();
 sg13g2_fill_2 FILLER_52_596 ();
 sg13g2_fill_2 FILLER_52_603 ();
 sg13g2_fill_1 FILLER_52_605 ();
 sg13g2_fill_1 FILLER_52_615 ();
 sg13g2_fill_2 FILLER_52_624 ();
 sg13g2_decap_4 FILLER_52_634 ();
 sg13g2_fill_2 FILLER_52_638 ();
 sg13g2_fill_1 FILLER_52_660 ();
 sg13g2_fill_1 FILLER_52_666 ();
 sg13g2_decap_4 FILLER_52_675 ();
 sg13g2_decap_4 FILLER_52_685 ();
 sg13g2_decap_8 FILLER_52_697 ();
 sg13g2_decap_4 FILLER_52_704 ();
 sg13g2_fill_2 FILLER_52_721 ();
 sg13g2_fill_1 FILLER_52_723 ();
 sg13g2_decap_4 FILLER_52_732 ();
 sg13g2_decap_8 FILLER_52_744 ();
 sg13g2_fill_1 FILLER_52_751 ();
 sg13g2_decap_8 FILLER_52_776 ();
 sg13g2_fill_2 FILLER_52_783 ();
 sg13g2_decap_4 FILLER_52_806 ();
 sg13g2_fill_2 FILLER_52_810 ();
 sg13g2_decap_8 FILLER_52_816 ();
 sg13g2_decap_4 FILLER_52_823 ();
 sg13g2_decap_8 FILLER_52_835 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_8 FILLER_52_854 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_16 ();
 sg13g2_decap_8 FILLER_53_23 ();
 sg13g2_decap_4 FILLER_53_30 ();
 sg13g2_fill_1 FILLER_53_45 ();
 sg13g2_decap_8 FILLER_53_55 ();
 sg13g2_fill_2 FILLER_53_74 ();
 sg13g2_fill_1 FILLER_53_76 ();
 sg13g2_fill_2 FILLER_53_102 ();
 sg13g2_fill_1 FILLER_53_117 ();
 sg13g2_fill_1 FILLER_53_123 ();
 sg13g2_decap_8 FILLER_53_132 ();
 sg13g2_fill_2 FILLER_53_139 ();
 sg13g2_decap_4 FILLER_53_149 ();
 sg13g2_fill_2 FILLER_53_179 ();
 sg13g2_fill_1 FILLER_53_181 ();
 sg13g2_decap_8 FILLER_53_208 ();
 sg13g2_decap_4 FILLER_53_215 ();
 sg13g2_fill_2 FILLER_53_219 ();
 sg13g2_fill_2 FILLER_53_225 ();
 sg13g2_fill_1 FILLER_53_227 ();
 sg13g2_fill_1 FILLER_53_232 ();
 sg13g2_decap_8 FILLER_53_241 ();
 sg13g2_decap_8 FILLER_53_248 ();
 sg13g2_fill_1 FILLER_53_255 ();
 sg13g2_decap_8 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_fill_2 FILLER_53_280 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_decap_4 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_305 ();
 sg13g2_decap_8 FILLER_53_345 ();
 sg13g2_decap_8 FILLER_53_352 ();
 sg13g2_fill_1 FILLER_53_359 ();
 sg13g2_fill_2 FILLER_53_416 ();
 sg13g2_fill_1 FILLER_53_418 ();
 sg13g2_fill_1 FILLER_53_424 ();
 sg13g2_fill_1 FILLER_53_436 ();
 sg13g2_fill_1 FILLER_53_441 ();
 sg13g2_decap_8 FILLER_53_446 ();
 sg13g2_fill_2 FILLER_53_453 ();
 sg13g2_fill_1 FILLER_53_455 ();
 sg13g2_fill_2 FILLER_53_478 ();
 sg13g2_fill_1 FILLER_53_531 ();
 sg13g2_fill_2 FILLER_53_547 ();
 sg13g2_fill_1 FILLER_53_549 ();
 sg13g2_fill_2 FILLER_53_556 ();
 sg13g2_fill_1 FILLER_53_558 ();
 sg13g2_fill_2 FILLER_53_594 ();
 sg13g2_fill_2 FILLER_53_604 ();
 sg13g2_fill_1 FILLER_53_606 ();
 sg13g2_fill_2 FILLER_53_612 ();
 sg13g2_fill_2 FILLER_53_622 ();
 sg13g2_decap_8 FILLER_53_629 ();
 sg13g2_fill_1 FILLER_53_640 ();
 sg13g2_decap_4 FILLER_53_650 ();
 sg13g2_fill_2 FILLER_53_654 ();
 sg13g2_fill_2 FILLER_53_677 ();
 sg13g2_fill_1 FILLER_53_679 ();
 sg13g2_decap_8 FILLER_53_688 ();
 sg13g2_fill_2 FILLER_53_695 ();
 sg13g2_decap_8 FILLER_53_709 ();
 sg13g2_fill_1 FILLER_53_716 ();
 sg13g2_decap_8 FILLER_53_730 ();
 sg13g2_fill_2 FILLER_53_737 ();
 sg13g2_fill_1 FILLER_53_739 ();
 sg13g2_fill_1 FILLER_53_745 ();
 sg13g2_fill_2 FILLER_53_810 ();
 sg13g2_decap_8 FILLER_53_836 ();
 sg13g2_decap_8 FILLER_53_843 ();
 sg13g2_decap_8 FILLER_53_850 ();
 sg13g2_decap_4 FILLER_53_857 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_fill_1 FILLER_54_26 ();
 sg13g2_decap_4 FILLER_54_48 ();
 sg13g2_fill_1 FILLER_54_52 ();
 sg13g2_decap_8 FILLER_54_64 ();
 sg13g2_fill_1 FILLER_54_71 ();
 sg13g2_fill_2 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_85 ();
 sg13g2_fill_1 FILLER_54_87 ();
 sg13g2_decap_4 FILLER_54_104 ();
 sg13g2_fill_2 FILLER_54_108 ();
 sg13g2_fill_2 FILLER_54_122 ();
 sg13g2_decap_4 FILLER_54_133 ();
 sg13g2_fill_1 FILLER_54_137 ();
 sg13g2_fill_1 FILLER_54_164 ();
 sg13g2_fill_2 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_fill_1 FILLER_54_210 ();
 sg13g2_decap_8 FILLER_54_232 ();
 sg13g2_decap_8 FILLER_54_239 ();
 sg13g2_decap_4 FILLER_54_246 ();
 sg13g2_fill_1 FILLER_54_250 ();
 sg13g2_decap_4 FILLER_54_264 ();
 sg13g2_fill_1 FILLER_54_281 ();
 sg13g2_decap_8 FILLER_54_303 ();
 sg13g2_fill_2 FILLER_54_310 ();
 sg13g2_fill_2 FILLER_54_322 ();
 sg13g2_fill_1 FILLER_54_324 ();
 sg13g2_fill_1 FILLER_54_341 ();
 sg13g2_decap_8 FILLER_54_355 ();
 sg13g2_fill_1 FILLER_54_362 ();
 sg13g2_fill_2 FILLER_54_389 ();
 sg13g2_fill_1 FILLER_54_457 ();
 sg13g2_fill_1 FILLER_54_490 ();
 sg13g2_decap_4 FILLER_54_496 ();
 sg13g2_fill_2 FILLER_54_508 ();
 sg13g2_fill_1 FILLER_54_510 ();
 sg13g2_fill_2 FILLER_54_542 ();
 sg13g2_decap_4 FILLER_54_580 ();
 sg13g2_fill_1 FILLER_54_584 ();
 sg13g2_fill_1 FILLER_54_590 ();
 sg13g2_decap_4 FILLER_54_596 ();
 sg13g2_fill_2 FILLER_54_618 ();
 sg13g2_fill_2 FILLER_54_643 ();
 sg13g2_decap_8 FILLER_54_658 ();
 sg13g2_fill_2 FILLER_54_665 ();
 sg13g2_fill_1 FILLER_54_667 ();
 sg13g2_fill_2 FILLER_54_676 ();
 sg13g2_decap_8 FILLER_54_690 ();
 sg13g2_fill_2 FILLER_54_697 ();
 sg13g2_fill_1 FILLER_54_699 ();
 sg13g2_fill_2 FILLER_54_712 ();
 sg13g2_fill_1 FILLER_54_714 ();
 sg13g2_fill_1 FILLER_54_723 ();
 sg13g2_decap_8 FILLER_54_729 ();
 sg13g2_decap_8 FILLER_54_736 ();
 sg13g2_decap_4 FILLER_54_743 ();
 sg13g2_fill_2 FILLER_54_747 ();
 sg13g2_decap_4 FILLER_54_754 ();
 sg13g2_fill_2 FILLER_54_766 ();
 sg13g2_fill_2 FILLER_54_776 ();
 sg13g2_fill_1 FILLER_54_790 ();
 sg13g2_fill_2 FILLER_54_795 ();
 sg13g2_fill_1 FILLER_54_797 ();
 sg13g2_decap_8 FILLER_54_805 ();
 sg13g2_decap_8 FILLER_54_812 ();
 sg13g2_decap_8 FILLER_54_819 ();
 sg13g2_decap_8 FILLER_54_826 ();
 sg13g2_decap_8 FILLER_54_833 ();
 sg13g2_decap_8 FILLER_54_840 ();
 sg13g2_decap_8 FILLER_54_847 ();
 sg13g2_decap_8 FILLER_54_854 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_19 ();
 sg13g2_decap_4 FILLER_55_50 ();
 sg13g2_fill_2 FILLER_55_54 ();
 sg13g2_fill_2 FILLER_55_76 ();
 sg13g2_fill_1 FILLER_55_78 ();
 sg13g2_fill_2 FILLER_55_92 ();
 sg13g2_fill_2 FILLER_55_99 ();
 sg13g2_fill_1 FILLER_55_129 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_decap_8 FILLER_55_201 ();
 sg13g2_fill_2 FILLER_55_208 ();
 sg13g2_decap_4 FILLER_55_241 ();
 sg13g2_fill_2 FILLER_55_257 ();
 sg13g2_decap_8 FILLER_55_274 ();
 sg13g2_fill_1 FILLER_55_281 ();
 sg13g2_fill_2 FILLER_55_294 ();
 sg13g2_fill_2 FILLER_55_303 ();
 sg13g2_fill_2 FILLER_55_325 ();
 sg13g2_fill_1 FILLER_55_327 ();
 sg13g2_decap_8 FILLER_55_347 ();
 sg13g2_fill_1 FILLER_55_354 ();
 sg13g2_decap_4 FILLER_55_397 ();
 sg13g2_fill_1 FILLER_55_401 ();
 sg13g2_decap_8 FILLER_55_406 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_fill_2 FILLER_55_420 ();
 sg13g2_fill_1 FILLER_55_422 ();
 sg13g2_fill_2 FILLER_55_456 ();
 sg13g2_fill_2 FILLER_55_463 ();
 sg13g2_fill_1 FILLER_55_474 ();
 sg13g2_decap_8 FILLER_55_479 ();
 sg13g2_decap_8 FILLER_55_486 ();
 sg13g2_fill_2 FILLER_55_509 ();
 sg13g2_fill_1 FILLER_55_511 ();
 sg13g2_fill_2 FILLER_55_518 ();
 sg13g2_fill_1 FILLER_55_525 ();
 sg13g2_decap_4 FILLER_55_572 ();
 sg13g2_decap_8 FILLER_55_603 ();
 sg13g2_decap_4 FILLER_55_622 ();
 sg13g2_decap_8 FILLER_55_634 ();
 sg13g2_decap_8 FILLER_55_641 ();
 sg13g2_decap_4 FILLER_55_656 ();
 sg13g2_decap_8 FILLER_55_665 ();
 sg13g2_decap_4 FILLER_55_700 ();
 sg13g2_fill_2 FILLER_55_704 ();
 sg13g2_fill_1 FILLER_55_715 ();
 sg13g2_decap_8 FILLER_55_792 ();
 sg13g2_decap_8 FILLER_55_799 ();
 sg13g2_decap_8 FILLER_55_806 ();
 sg13g2_decap_8 FILLER_55_813 ();
 sg13g2_decap_8 FILLER_55_820 ();
 sg13g2_decap_8 FILLER_55_827 ();
 sg13g2_decap_8 FILLER_55_834 ();
 sg13g2_decap_8 FILLER_55_841 ();
 sg13g2_decap_8 FILLER_55_848 ();
 sg13g2_decap_8 FILLER_55_855 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_50 ();
 sg13g2_fill_2 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_58 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_4 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_105 ();
 sg13g2_fill_1 FILLER_56_107 ();
 sg13g2_fill_2 FILLER_56_114 ();
 sg13g2_fill_1 FILLER_56_116 ();
 sg13g2_decap_8 FILLER_56_125 ();
 sg13g2_decap_8 FILLER_56_132 ();
 sg13g2_decap_4 FILLER_56_139 ();
 sg13g2_fill_1 FILLER_56_143 ();
 sg13g2_fill_2 FILLER_56_170 ();
 sg13g2_fill_2 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_188 ();
 sg13g2_fill_1 FILLER_56_238 ();
 sg13g2_decap_4 FILLER_56_255 ();
 sg13g2_fill_2 FILLER_56_259 ();
 sg13g2_fill_2 FILLER_56_274 ();
 sg13g2_fill_1 FILLER_56_276 ();
 sg13g2_decap_4 FILLER_56_283 ();
 sg13g2_fill_1 FILLER_56_287 ();
 sg13g2_fill_2 FILLER_56_296 ();
 sg13g2_fill_2 FILLER_56_368 ();
 sg13g2_fill_1 FILLER_56_370 ();
 sg13g2_fill_1 FILLER_56_385 ();
 sg13g2_fill_2 FILLER_56_394 ();
 sg13g2_fill_1 FILLER_56_427 ();
 sg13g2_fill_1 FILLER_56_465 ();
 sg13g2_decap_8 FILLER_56_492 ();
 sg13g2_fill_1 FILLER_56_509 ();
 sg13g2_fill_1 FILLER_56_573 ();
 sg13g2_fill_2 FILLER_56_580 ();
 sg13g2_fill_1 FILLER_56_586 ();
 sg13g2_fill_1 FILLER_56_593 ();
 sg13g2_decap_4 FILLER_56_642 ();
 sg13g2_fill_2 FILLER_56_676 ();
 sg13g2_fill_2 FILLER_56_689 ();
 sg13g2_decap_4 FILLER_56_699 ();
 sg13g2_decap_4 FILLER_56_738 ();
 sg13g2_fill_1 FILLER_56_742 ();
 sg13g2_decap_8 FILLER_56_756 ();
 sg13g2_decap_8 FILLER_56_763 ();
 sg13g2_decap_8 FILLER_56_770 ();
 sg13g2_fill_2 FILLER_56_777 ();
 sg13g2_decap_8 FILLER_56_783 ();
 sg13g2_decap_8 FILLER_56_790 ();
 sg13g2_decap_8 FILLER_56_797 ();
 sg13g2_decap_8 FILLER_56_804 ();
 sg13g2_decap_8 FILLER_56_811 ();
 sg13g2_decap_8 FILLER_56_818 ();
 sg13g2_decap_8 FILLER_56_825 ();
 sg13g2_decap_8 FILLER_56_832 ();
 sg13g2_decap_8 FILLER_56_839 ();
 sg13g2_decap_8 FILLER_56_846 ();
 sg13g2_decap_8 FILLER_56_853 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_12 ();
 sg13g2_fill_1 FILLER_57_16 ();
 sg13g2_fill_2 FILLER_57_21 ();
 sg13g2_fill_2 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_47 ();
 sg13g2_fill_2 FILLER_57_54 ();
 sg13g2_decap_8 FILLER_57_60 ();
 sg13g2_fill_2 FILLER_57_67 ();
 sg13g2_fill_1 FILLER_57_69 ();
 sg13g2_decap_4 FILLER_57_74 ();
 sg13g2_fill_2 FILLER_57_78 ();
 sg13g2_fill_1 FILLER_57_86 ();
 sg13g2_fill_2 FILLER_57_94 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_4 FILLER_57_126 ();
 sg13g2_fill_2 FILLER_57_130 ();
 sg13g2_fill_2 FILLER_57_153 ();
 sg13g2_fill_1 FILLER_57_172 ();
 sg13g2_decap_4 FILLER_57_199 ();
 sg13g2_fill_2 FILLER_57_245 ();
 sg13g2_decap_8 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_302 ();
 sg13g2_decap_4 FILLER_57_309 ();
 sg13g2_decap_4 FILLER_57_323 ();
 sg13g2_decap_4 FILLER_57_344 ();
 sg13g2_fill_1 FILLER_57_348 ();
 sg13g2_fill_1 FILLER_57_353 ();
 sg13g2_fill_2 FILLER_57_363 ();
 sg13g2_fill_1 FILLER_57_379 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_decap_4 FILLER_57_407 ();
 sg13g2_fill_2 FILLER_57_425 ();
 sg13g2_fill_1 FILLER_57_427 ();
 sg13g2_decap_4 FILLER_57_434 ();
 sg13g2_decap_4 FILLER_57_449 ();
 sg13g2_fill_1 FILLER_57_453 ();
 sg13g2_fill_2 FILLER_57_462 ();
 sg13g2_decap_8 FILLER_57_469 ();
 sg13g2_decap_8 FILLER_57_480 ();
 sg13g2_fill_2 FILLER_57_525 ();
 sg13g2_fill_1 FILLER_57_541 ();
 sg13g2_fill_1 FILLER_57_551 ();
 sg13g2_decap_8 FILLER_57_577 ();
 sg13g2_fill_2 FILLER_57_603 ();
 sg13g2_fill_1 FILLER_57_605 ();
 sg13g2_decap_4 FILLER_57_612 ();
 sg13g2_decap_4 FILLER_57_632 ();
 sg13g2_fill_2 FILLER_57_644 ();
 sg13g2_fill_1 FILLER_57_646 ();
 sg13g2_decap_8 FILLER_57_659 ();
 sg13g2_fill_1 FILLER_57_666 ();
 sg13g2_decap_8 FILLER_57_677 ();
 sg13g2_fill_2 FILLER_57_684 ();
 sg13g2_fill_1 FILLER_57_686 ();
 sg13g2_decap_8 FILLER_57_699 ();
 sg13g2_decap_8 FILLER_57_706 ();
 sg13g2_fill_2 FILLER_57_713 ();
 sg13g2_fill_2 FILLER_57_718 ();
 sg13g2_fill_2 FILLER_57_728 ();
 sg13g2_fill_1 FILLER_57_751 ();
 sg13g2_decap_4 FILLER_57_760 ();
 sg13g2_fill_1 FILLER_57_764 ();
 sg13g2_decap_8 FILLER_57_773 ();
 sg13g2_decap_8 FILLER_57_780 ();
 sg13g2_decap_8 FILLER_57_787 ();
 sg13g2_decap_8 FILLER_57_794 ();
 sg13g2_decap_8 FILLER_57_801 ();
 sg13g2_decap_8 FILLER_57_808 ();
 sg13g2_decap_8 FILLER_57_815 ();
 sg13g2_decap_8 FILLER_57_822 ();
 sg13g2_decap_8 FILLER_57_829 ();
 sg13g2_decap_8 FILLER_57_836 ();
 sg13g2_decap_8 FILLER_57_843 ();
 sg13g2_decap_8 FILLER_57_850 ();
 sg13g2_decap_4 FILLER_57_857 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_fill_2 FILLER_58_26 ();
 sg13g2_fill_2 FILLER_58_51 ();
 sg13g2_fill_1 FILLER_58_53 ();
 sg13g2_decap_4 FILLER_58_101 ();
 sg13g2_fill_1 FILLER_58_105 ();
 sg13g2_decap_4 FILLER_58_204 ();
 sg13g2_fill_1 FILLER_58_208 ();
 sg13g2_decap_8 FILLER_58_222 ();
 sg13g2_fill_1 FILLER_58_229 ();
 sg13g2_decap_8 FILLER_58_235 ();
 sg13g2_decap_4 FILLER_58_242 ();
 sg13g2_fill_1 FILLER_58_246 ();
 sg13g2_decap_8 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_265 ();
 sg13g2_fill_1 FILLER_58_267 ();
 sg13g2_decap_4 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_280 ();
 sg13g2_fill_1 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_305 ();
 sg13g2_fill_1 FILLER_58_312 ();
 sg13g2_decap_8 FILLER_58_318 ();
 sg13g2_fill_2 FILLER_58_325 ();
 sg13g2_fill_2 FILLER_58_337 ();
 sg13g2_fill_2 FILLER_58_349 ();
 sg13g2_decap_4 FILLER_58_387 ();
 sg13g2_fill_2 FILLER_58_391 ();
 sg13g2_decap_4 FILLER_58_398 ();
 sg13g2_fill_1 FILLER_58_402 ();
 sg13g2_decap_4 FILLER_58_407 ();
 sg13g2_decap_4 FILLER_58_419 ();
 sg13g2_fill_2 FILLER_58_434 ();
 sg13g2_fill_1 FILLER_58_436 ();
 sg13g2_fill_1 FILLER_58_454 ();
 sg13g2_decap_8 FILLER_58_463 ();
 sg13g2_fill_2 FILLER_58_470 ();
 sg13g2_fill_1 FILLER_58_472 ();
 sg13g2_decap_4 FILLER_58_477 ();
 sg13g2_fill_2 FILLER_58_481 ();
 sg13g2_fill_2 FILLER_58_494 ();
 sg13g2_fill_1 FILLER_58_501 ();
 sg13g2_fill_2 FILLER_58_508 ();
 sg13g2_fill_2 FILLER_58_523 ();
 sg13g2_fill_1 FILLER_58_555 ();
 sg13g2_fill_2 FILLER_58_572 ();
 sg13g2_fill_1 FILLER_58_574 ();
 sg13g2_fill_2 FILLER_58_584 ();
 sg13g2_fill_1 FILLER_58_586 ();
 sg13g2_decap_8 FILLER_58_595 ();
 sg13g2_decap_8 FILLER_58_602 ();
 sg13g2_decap_4 FILLER_58_609 ();
 sg13g2_fill_2 FILLER_58_613 ();
 sg13g2_fill_2 FILLER_58_631 ();
 sg13g2_fill_1 FILLER_58_633 ();
 sg13g2_decap_8 FILLER_58_642 ();
 sg13g2_fill_1 FILLER_58_649 ();
 sg13g2_decap_4 FILLER_58_677 ();
 sg13g2_fill_1 FILLER_58_681 ();
 sg13g2_decap_4 FILLER_58_701 ();
 sg13g2_fill_1 FILLER_58_705 ();
 sg13g2_decap_8 FILLER_58_712 ();
 sg13g2_decap_4 FILLER_58_719 ();
 sg13g2_fill_1 FILLER_58_723 ();
 sg13g2_decap_8 FILLER_58_741 ();
 sg13g2_fill_2 FILLER_58_748 ();
 sg13g2_fill_2 FILLER_58_758 ();
 sg13g2_fill_1 FILLER_58_760 ();
 sg13g2_decap_8 FILLER_58_786 ();
 sg13g2_decap_8 FILLER_58_793 ();
 sg13g2_decap_8 FILLER_58_800 ();
 sg13g2_decap_8 FILLER_58_807 ();
 sg13g2_decap_8 FILLER_58_814 ();
 sg13g2_decap_8 FILLER_58_821 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_19 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_decap_4 FILLER_59_72 ();
 sg13g2_fill_1 FILLER_59_76 ();
 sg13g2_fill_2 FILLER_59_89 ();
 sg13g2_decap_4 FILLER_59_96 ();
 sg13g2_fill_2 FILLER_59_100 ();
 sg13g2_decap_4 FILLER_59_124 ();
 sg13g2_fill_2 FILLER_59_262 ();
 sg13g2_fill_1 FILLER_59_280 ();
 sg13g2_fill_1 FILLER_59_293 ();
 sg13g2_fill_1 FILLER_59_298 ();
 sg13g2_fill_2 FILLER_59_311 ();
 sg13g2_fill_1 FILLER_59_334 ();
 sg13g2_fill_1 FILLER_59_418 ();
 sg13g2_fill_2 FILLER_59_460 ();
 sg13g2_fill_1 FILLER_59_462 ();
 sg13g2_fill_2 FILLER_59_505 ();
 sg13g2_fill_1 FILLER_59_507 ();
 sg13g2_fill_1 FILLER_59_518 ();
 sg13g2_fill_2 FILLER_59_528 ();
 sg13g2_fill_1 FILLER_59_530 ();
 sg13g2_fill_1 FILLER_59_536 ();
 sg13g2_fill_2 FILLER_59_566 ();
 sg13g2_fill_2 FILLER_59_601 ();
 sg13g2_fill_1 FILLER_59_621 ();
 sg13g2_fill_2 FILLER_59_626 ();
 sg13g2_fill_1 FILLER_59_628 ();
 sg13g2_fill_2 FILLER_59_657 ();
 sg13g2_decap_8 FILLER_59_662 ();
 sg13g2_fill_1 FILLER_59_669 ();
 sg13g2_decap_4 FILLER_59_673 ();
 sg13g2_fill_1 FILLER_59_677 ();
 sg13g2_fill_2 FILLER_59_689 ();
 sg13g2_fill_1 FILLER_59_691 ();
 sg13g2_decap_8 FILLER_59_700 ();
 sg13g2_fill_1 FILLER_59_707 ();
 sg13g2_decap_4 FILLER_59_720 ();
 sg13g2_decap_8 FILLER_59_745 ();
 sg13g2_decap_8 FILLER_59_752 ();
 sg13g2_fill_1 FILLER_59_759 ();
 sg13g2_fill_1 FILLER_59_765 ();
 sg13g2_decap_8 FILLER_59_774 ();
 sg13g2_decap_8 FILLER_59_781 ();
 sg13g2_decap_8 FILLER_59_788 ();
 sg13g2_decap_8 FILLER_59_795 ();
 sg13g2_decap_8 FILLER_59_802 ();
 sg13g2_decap_8 FILLER_59_809 ();
 sg13g2_decap_8 FILLER_59_816 ();
 sg13g2_decap_8 FILLER_59_823 ();
 sg13g2_decap_8 FILLER_59_830 ();
 sg13g2_decap_8 FILLER_59_837 ();
 sg13g2_decap_8 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_851 ();
 sg13g2_decap_4 FILLER_59_858 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_176 ();
 sg13g2_fill_2 FILLER_60_236 ();
 sg13g2_fill_1 FILLER_60_264 ();
 sg13g2_decap_4 FILLER_60_288 ();
 sg13g2_fill_1 FILLER_60_292 ();
 sg13g2_fill_2 FILLER_60_301 ();
 sg13g2_fill_1 FILLER_60_303 ();
 sg13g2_decap_8 FILLER_60_308 ();
 sg13g2_decap_8 FILLER_60_315 ();
 sg13g2_fill_2 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_324 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_332 ();
 sg13g2_decap_4 FILLER_60_359 ();
 sg13g2_decap_8 FILLER_60_390 ();
 sg13g2_decap_4 FILLER_60_414 ();
 sg13g2_fill_2 FILLER_60_418 ();
 sg13g2_fill_2 FILLER_60_447 ();
 sg13g2_fill_2 FILLER_60_480 ();
 sg13g2_fill_1 FILLER_60_482 ();
 sg13g2_fill_2 FILLER_60_518 ();
 sg13g2_decap_4 FILLER_60_565 ();
 sg13g2_fill_1 FILLER_60_569 ();
 sg13g2_fill_2 FILLER_60_574 ();
 sg13g2_fill_1 FILLER_60_576 ();
 sg13g2_decap_4 FILLER_60_581 ();
 sg13g2_fill_1 FILLER_60_585 ();
 sg13g2_decap_4 FILLER_60_594 ();
 sg13g2_fill_2 FILLER_60_598 ();
 sg13g2_decap_4 FILLER_60_612 ();
 sg13g2_fill_1 FILLER_60_636 ();
 sg13g2_decap_4 FILLER_60_641 ();
 sg13g2_fill_2 FILLER_60_645 ();
 sg13g2_fill_1 FILLER_60_674 ();
 sg13g2_fill_2 FILLER_60_701 ();
 sg13g2_decap_4 FILLER_60_719 ();
 sg13g2_decap_4 FILLER_60_749 ();
 sg13g2_fill_2 FILLER_60_753 ();
 sg13g2_decap_8 FILLER_60_775 ();
 sg13g2_decap_8 FILLER_60_782 ();
 sg13g2_decap_8 FILLER_60_789 ();
 sg13g2_decap_8 FILLER_60_796 ();
 sg13g2_decap_8 FILLER_60_803 ();
 sg13g2_decap_8 FILLER_60_810 ();
 sg13g2_decap_8 FILLER_60_817 ();
 sg13g2_decap_8 FILLER_60_824 ();
 sg13g2_decap_8 FILLER_60_831 ();
 sg13g2_decap_8 FILLER_60_838 ();
 sg13g2_decap_8 FILLER_60_845 ();
 sg13g2_decap_8 FILLER_60_852 ();
 sg13g2_fill_2 FILLER_60_859 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_fill_1 FILLER_61_26 ();
 sg13g2_fill_2 FILLER_61_44 ();
 sg13g2_fill_1 FILLER_61_46 ();
 sg13g2_fill_2 FILLER_61_51 ();
 sg13g2_fill_1 FILLER_61_53 ();
 sg13g2_decap_4 FILLER_61_58 ();
 sg13g2_decap_8 FILLER_61_66 ();
 sg13g2_decap_4 FILLER_61_73 ();
 sg13g2_fill_2 FILLER_61_96 ();
 sg13g2_fill_1 FILLER_61_98 ();
 sg13g2_fill_1 FILLER_61_104 ();
 sg13g2_fill_2 FILLER_61_114 ();
 sg13g2_fill_1 FILLER_61_125 ();
 sg13g2_fill_2 FILLER_61_135 ();
 sg13g2_fill_1 FILLER_61_157 ();
 sg13g2_fill_1 FILLER_61_174 ();
 sg13g2_fill_1 FILLER_61_203 ();
 sg13g2_fill_2 FILLER_61_209 ();
 sg13g2_fill_1 FILLER_61_236 ();
 sg13g2_decap_8 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_278 ();
 sg13g2_fill_2 FILLER_61_285 ();
 sg13g2_decap_4 FILLER_61_292 ();
 sg13g2_fill_1 FILLER_61_296 ();
 sg13g2_fill_2 FILLER_61_306 ();
 sg13g2_fill_1 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_fill_1 FILLER_61_329 ();
 sg13g2_decap_4 FILLER_61_338 ();
 sg13g2_fill_2 FILLER_61_342 ();
 sg13g2_fill_1 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_364 ();
 sg13g2_fill_2 FILLER_61_373 ();
 sg13g2_fill_2 FILLER_61_401 ();
 sg13g2_fill_1 FILLER_61_403 ();
 sg13g2_fill_1 FILLER_61_465 ();
 sg13g2_fill_2 FILLER_61_516 ();
 sg13g2_fill_1 FILLER_61_526 ();
 sg13g2_fill_1 FILLER_61_573 ();
 sg13g2_fill_1 FILLER_61_593 ();
 sg13g2_fill_2 FILLER_61_610 ();
 sg13g2_fill_2 FILLER_61_626 ();
 sg13g2_decap_4 FILLER_61_656 ();
 sg13g2_decap_8 FILLER_61_668 ();
 sg13g2_fill_2 FILLER_61_675 ();
 sg13g2_fill_1 FILLER_61_677 ();
 sg13g2_decap_8 FILLER_61_683 ();
 sg13g2_decap_4 FILLER_61_690 ();
 sg13g2_fill_2 FILLER_61_698 ();
 sg13g2_fill_1 FILLER_61_700 ();
 sg13g2_decap_4 FILLER_61_725 ();
 sg13g2_fill_2 FILLER_61_729 ();
 sg13g2_fill_1 FILLER_61_736 ();
 sg13g2_fill_2 FILLER_61_755 ();
 sg13g2_decap_8 FILLER_61_782 ();
 sg13g2_decap_8 FILLER_61_789 ();
 sg13g2_decap_8 FILLER_61_796 ();
 sg13g2_decap_8 FILLER_61_803 ();
 sg13g2_decap_8 FILLER_61_810 ();
 sg13g2_decap_8 FILLER_61_817 ();
 sg13g2_decap_8 FILLER_61_824 ();
 sg13g2_decap_8 FILLER_61_831 ();
 sg13g2_decap_8 FILLER_61_838 ();
 sg13g2_decap_8 FILLER_61_845 ();
 sg13g2_decap_8 FILLER_61_852 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_30 ();
 sg13g2_fill_1 FILLER_62_32 ();
 sg13g2_fill_2 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_54 ();
 sg13g2_decap_4 FILLER_62_61 ();
 sg13g2_fill_1 FILLER_62_65 ();
 sg13g2_fill_1 FILLER_62_90 ();
 sg13g2_fill_2 FILLER_62_130 ();
 sg13g2_fill_1 FILLER_62_132 ();
 sg13g2_fill_1 FILLER_62_167 ();
 sg13g2_fill_2 FILLER_62_204 ();
 sg13g2_fill_1 FILLER_62_206 ();
 sg13g2_fill_1 FILLER_62_234 ();
 sg13g2_fill_1 FILLER_62_244 ();
 sg13g2_fill_2 FILLER_62_288 ();
 sg13g2_fill_1 FILLER_62_290 ();
 sg13g2_fill_2 FILLER_62_347 ();
 sg13g2_fill_1 FILLER_62_349 ();
 sg13g2_decap_8 FILLER_62_355 ();
 sg13g2_fill_2 FILLER_62_362 ();
 sg13g2_fill_1 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_377 ();
 sg13g2_fill_1 FILLER_62_384 ();
 sg13g2_decap_8 FILLER_62_389 ();
 sg13g2_fill_2 FILLER_62_414 ();
 sg13g2_fill_1 FILLER_62_416 ();
 sg13g2_fill_1 FILLER_62_426 ();
 sg13g2_decap_4 FILLER_62_431 ();
 sg13g2_fill_2 FILLER_62_435 ();
 sg13g2_fill_1 FILLER_62_460 ();
 sg13g2_fill_2 FILLER_62_471 ();
 sg13g2_fill_2 FILLER_62_481 ();
 sg13g2_fill_1 FILLER_62_483 ();
 sg13g2_fill_1 FILLER_62_506 ();
 sg13g2_fill_1 FILLER_62_521 ();
 sg13g2_fill_2 FILLER_62_536 ();
 sg13g2_decap_8 FILLER_62_581 ();
 sg13g2_fill_2 FILLER_62_588 ();
 sg13g2_decap_8 FILLER_62_611 ();
 sg13g2_decap_8 FILLER_62_618 ();
 sg13g2_decap_4 FILLER_62_625 ();
 sg13g2_decap_8 FILLER_62_642 ();
 sg13g2_fill_2 FILLER_62_649 ();
 sg13g2_fill_1 FILLER_62_651 ();
 sg13g2_decap_4 FILLER_62_664 ();
 sg13g2_fill_1 FILLER_62_668 ();
 sg13g2_fill_2 FILLER_62_693 ();
 sg13g2_fill_1 FILLER_62_695 ();
 sg13g2_decap_8 FILLER_62_720 ();
 sg13g2_fill_2 FILLER_62_727 ();
 sg13g2_fill_1 FILLER_62_729 ();
 sg13g2_decap_8 FILLER_62_778 ();
 sg13g2_decap_8 FILLER_62_785 ();
 sg13g2_decap_8 FILLER_62_792 ();
 sg13g2_decap_8 FILLER_62_799 ();
 sg13g2_decap_8 FILLER_62_806 ();
 sg13g2_decap_8 FILLER_62_813 ();
 sg13g2_decap_8 FILLER_62_820 ();
 sg13g2_decap_8 FILLER_62_827 ();
 sg13g2_decap_8 FILLER_62_834 ();
 sg13g2_decap_8 FILLER_62_841 ();
 sg13g2_decap_8 FILLER_62_848 ();
 sg13g2_decap_8 FILLER_62_855 ();
 sg13g2_fill_1 FILLER_63_38 ();
 sg13g2_fill_2 FILLER_63_44 ();
 sg13g2_fill_1 FILLER_63_46 ();
 sg13g2_fill_2 FILLER_63_57 ();
 sg13g2_fill_2 FILLER_63_77 ();
 sg13g2_decap_4 FILLER_63_84 ();
 sg13g2_fill_1 FILLER_63_88 ();
 sg13g2_fill_2 FILLER_63_121 ();
 sg13g2_fill_2 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_152 ();
 sg13g2_fill_2 FILLER_63_188 ();
 sg13g2_fill_1 FILLER_63_190 ();
 sg13g2_fill_2 FILLER_63_230 ();
 sg13g2_decap_4 FILLER_63_267 ();
 sg13g2_fill_2 FILLER_63_271 ();
 sg13g2_decap_8 FILLER_63_277 ();
 sg13g2_fill_2 FILLER_63_284 ();
 sg13g2_fill_1 FILLER_63_300 ();
 sg13g2_fill_2 FILLER_63_334 ();
 sg13g2_fill_1 FILLER_63_336 ();
 sg13g2_decap_4 FILLER_63_342 ();
 sg13g2_fill_1 FILLER_63_346 ();
 sg13g2_decap_4 FILLER_63_352 ();
 sg13g2_fill_1 FILLER_63_361 ();
 sg13g2_fill_2 FILLER_63_376 ();
 sg13g2_fill_1 FILLER_63_415 ();
 sg13g2_fill_2 FILLER_63_449 ();
 sg13g2_fill_2 FILLER_63_481 ();
 sg13g2_fill_1 FILLER_63_483 ();
 sg13g2_fill_1 FILLER_63_488 ();
 sg13g2_fill_1 FILLER_63_509 ();
 sg13g2_fill_2 FILLER_63_560 ();
 sg13g2_fill_1 FILLER_63_569 ();
 sg13g2_fill_2 FILLER_63_589 ();
 sg13g2_fill_1 FILLER_63_596 ();
 sg13g2_decap_8 FILLER_63_605 ();
 sg13g2_fill_2 FILLER_63_624 ();
 sg13g2_fill_1 FILLER_63_626 ();
 sg13g2_decap_8 FILLER_63_644 ();
 sg13g2_decap_4 FILLER_63_651 ();
 sg13g2_fill_1 FILLER_63_655 ();
 sg13g2_fill_1 FILLER_63_674 ();
 sg13g2_decap_4 FILLER_63_688 ();
 sg13g2_decap_4 FILLER_63_701 ();
 sg13g2_fill_1 FILLER_63_705 ();
 sg13g2_decap_4 FILLER_63_711 ();
 sg13g2_fill_2 FILLER_63_715 ();
 sg13g2_decap_4 FILLER_63_730 ();
 sg13g2_decap_8 FILLER_63_739 ();
 sg13g2_fill_1 FILLER_63_746 ();
 sg13g2_fill_1 FILLER_63_760 ();
 sg13g2_fill_2 FILLER_63_769 ();
 sg13g2_decap_8 FILLER_63_776 ();
 sg13g2_decap_8 FILLER_63_783 ();
 sg13g2_decap_8 FILLER_63_790 ();
 sg13g2_decap_8 FILLER_63_797 ();
 sg13g2_decap_8 FILLER_63_804 ();
 sg13g2_decap_8 FILLER_63_811 ();
 sg13g2_decap_8 FILLER_63_818 ();
 sg13g2_decap_8 FILLER_63_825 ();
 sg13g2_decap_8 FILLER_63_832 ();
 sg13g2_decap_8 FILLER_63_839 ();
 sg13g2_decap_8 FILLER_63_846 ();
 sg13g2_decap_8 FILLER_63_853 ();
 sg13g2_fill_2 FILLER_63_860 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_43 ();
 sg13g2_fill_1 FILLER_64_57 ();
 sg13g2_fill_2 FILLER_64_79 ();
 sg13g2_fill_1 FILLER_64_81 ();
 sg13g2_fill_2 FILLER_64_103 ();
 sg13g2_fill_1 FILLER_64_105 ();
 sg13g2_fill_1 FILLER_64_111 ();
 sg13g2_fill_2 FILLER_64_146 ();
 sg13g2_fill_2 FILLER_64_174 ();
 sg13g2_fill_1 FILLER_64_176 ();
 sg13g2_fill_2 FILLER_64_184 ();
 sg13g2_fill_1 FILLER_64_186 ();
 sg13g2_fill_2 FILLER_64_256 ();
 sg13g2_fill_1 FILLER_64_258 ();
 sg13g2_fill_1 FILLER_64_285 ();
 sg13g2_fill_2 FILLER_64_294 ();
 sg13g2_fill_1 FILLER_64_301 ();
 sg13g2_fill_2 FILLER_64_323 ();
 sg13g2_fill_1 FILLER_64_340 ();
 sg13g2_decap_8 FILLER_64_356 ();
 sg13g2_fill_1 FILLER_64_363 ();
 sg13g2_fill_2 FILLER_64_378 ();
 sg13g2_decap_8 FILLER_64_449 ();
 sg13g2_decap_4 FILLER_64_456 ();
 sg13g2_fill_1 FILLER_64_460 ();
 sg13g2_fill_1 FILLER_64_465 ();
 sg13g2_fill_2 FILLER_64_516 ();
 sg13g2_fill_2 FILLER_64_562 ();
 sg13g2_decap_4 FILLER_64_601 ();
 sg13g2_fill_2 FILLER_64_605 ();
 sg13g2_decap_8 FILLER_64_619 ();
 sg13g2_fill_1 FILLER_64_626 ();
 sg13g2_decap_4 FILLER_64_649 ();
 sg13g2_fill_2 FILLER_64_673 ();
 sg13g2_decap_8 FILLER_64_688 ();
 sg13g2_fill_2 FILLER_64_695 ();
 sg13g2_fill_1 FILLER_64_697 ();
 sg13g2_fill_2 FILLER_64_726 ();
 sg13g2_decap_4 FILLER_64_756 ();
 sg13g2_fill_2 FILLER_64_760 ();
 sg13g2_decap_8 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_782 ();
 sg13g2_decap_8 FILLER_64_789 ();
 sg13g2_decap_8 FILLER_64_796 ();
 sg13g2_decap_8 FILLER_64_803 ();
 sg13g2_decap_8 FILLER_64_810 ();
 sg13g2_decap_8 FILLER_64_817 ();
 sg13g2_decap_8 FILLER_64_824 ();
 sg13g2_decap_8 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_87 ();
 sg13g2_decap_4 FILLER_65_118 ();
 sg13g2_fill_1 FILLER_65_131 ();
 sg13g2_fill_2 FILLER_65_182 ();
 sg13g2_fill_1 FILLER_65_200 ();
 sg13g2_fill_2 FILLER_65_247 ();
 sg13g2_fill_1 FILLER_65_249 ();
 sg13g2_decap_8 FILLER_65_280 ();
 sg13g2_decap_4 FILLER_65_287 ();
 sg13g2_fill_1 FILLER_65_301 ();
 sg13g2_fill_2 FILLER_65_312 ();
 sg13g2_decap_4 FILLER_65_323 ();
 sg13g2_fill_2 FILLER_65_327 ();
 sg13g2_fill_1 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_349 ();
 sg13g2_decap_8 FILLER_65_356 ();
 sg13g2_fill_1 FILLER_65_373 ();
 sg13g2_fill_2 FILLER_65_391 ();
 sg13g2_fill_1 FILLER_65_393 ();
 sg13g2_fill_1 FILLER_65_402 ();
 sg13g2_decap_8 FILLER_65_463 ();
 sg13g2_decap_4 FILLER_65_470 ();
 sg13g2_decap_4 FILLER_65_478 ();
 sg13g2_fill_2 FILLER_65_482 ();
 sg13g2_fill_2 FILLER_65_560 ();
 sg13g2_fill_1 FILLER_65_562 ();
 sg13g2_fill_1 FILLER_65_627 ();
 sg13g2_decap_8 FILLER_65_674 ();
 sg13g2_decap_8 FILLER_65_681 ();
 sg13g2_fill_1 FILLER_65_688 ();
 sg13g2_decap_4 FILLER_65_695 ();
 sg13g2_fill_1 FILLER_65_699 ();
 sg13g2_decap_8 FILLER_65_704 ();
 sg13g2_decap_4 FILLER_65_711 ();
 sg13g2_decap_8 FILLER_65_723 ();
 sg13g2_fill_2 FILLER_65_730 ();
 sg13g2_fill_1 FILLER_65_732 ();
 sg13g2_fill_1 FILLER_65_737 ();
 sg13g2_decap_4 FILLER_65_753 ();
 sg13g2_fill_1 FILLER_65_757 ();
 sg13g2_fill_2 FILLER_65_763 ();
 sg13g2_fill_1 FILLER_65_765 ();
 sg13g2_decap_8 FILLER_65_784 ();
 sg13g2_decap_8 FILLER_65_791 ();
 sg13g2_decap_8 FILLER_65_798 ();
 sg13g2_decap_8 FILLER_65_805 ();
 sg13g2_decap_8 FILLER_65_812 ();
 sg13g2_decap_8 FILLER_65_819 ();
 sg13g2_decap_8 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_833 ();
 sg13g2_decap_8 FILLER_65_840 ();
 sg13g2_decap_8 FILLER_65_847 ();
 sg13g2_decap_8 FILLER_65_854 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_59 ();
 sg13g2_fill_2 FILLER_66_65 ();
 sg13g2_fill_1 FILLER_66_67 ();
 sg13g2_fill_2 FILLER_66_115 ();
 sg13g2_fill_1 FILLER_66_129 ();
 sg13g2_decap_4 FILLER_66_156 ();
 sg13g2_fill_2 FILLER_66_160 ();
 sg13g2_decap_8 FILLER_66_265 ();
 sg13g2_decap_4 FILLER_66_280 ();
 sg13g2_fill_1 FILLER_66_292 ();
 sg13g2_fill_2 FILLER_66_308 ();
 sg13g2_fill_1 FILLER_66_326 ();
 sg13g2_fill_1 FILLER_66_337 ();
 sg13g2_fill_2 FILLER_66_390 ();
 sg13g2_fill_1 FILLER_66_392 ();
 sg13g2_fill_2 FILLER_66_460 ();
 sg13g2_fill_1 FILLER_66_462 ();
 sg13g2_fill_2 FILLER_66_511 ();
 sg13g2_fill_2 FILLER_66_536 ();
 sg13g2_fill_1 FILLER_66_538 ();
 sg13g2_fill_2 FILLER_66_588 ();
 sg13g2_fill_1 FILLER_66_590 ();
 sg13g2_decap_8 FILLER_66_621 ();
 sg13g2_decap_4 FILLER_66_628 ();
 sg13g2_fill_2 FILLER_66_640 ();
 sg13g2_fill_2 FILLER_66_648 ();
 sg13g2_fill_1 FILLER_66_650 ();
 sg13g2_fill_2 FILLER_66_659 ();
 sg13g2_decap_4 FILLER_66_679 ();
 sg13g2_fill_2 FILLER_66_691 ();
 sg13g2_fill_1 FILLER_66_693 ();
 sg13g2_fill_1 FILLER_66_701 ();
 sg13g2_fill_2 FILLER_66_715 ();
 sg13g2_fill_1 FILLER_66_717 ();
 sg13g2_decap_8 FILLER_66_748 ();
 sg13g2_fill_2 FILLER_66_755 ();
 sg13g2_fill_1 FILLER_66_757 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_fill_1 FILLER_67_26 ();
 sg13g2_fill_2 FILLER_67_138 ();
 sg13g2_decap_8 FILLER_67_144 ();
 sg13g2_fill_1 FILLER_67_151 ();
 sg13g2_decap_4 FILLER_67_155 ();
 sg13g2_fill_1 FILLER_67_159 ();
 sg13g2_fill_2 FILLER_67_165 ();
 sg13g2_fill_1 FILLER_67_189 ();
 sg13g2_fill_2 FILLER_67_220 ();
 sg13g2_fill_2 FILLER_67_231 ();
 sg13g2_fill_1 FILLER_67_233 ();
 sg13g2_decap_8 FILLER_67_286 ();
 sg13g2_fill_2 FILLER_67_304 ();
 sg13g2_fill_1 FILLER_67_306 ();
 sg13g2_decap_8 FILLER_67_334 ();
 sg13g2_decap_8 FILLER_67_341 ();
 sg13g2_fill_2 FILLER_67_348 ();
 sg13g2_fill_1 FILLER_67_350 ();
 sg13g2_decap_4 FILLER_67_355 ();
 sg13g2_fill_1 FILLER_67_367 ();
 sg13g2_fill_1 FILLER_67_390 ();
 sg13g2_fill_2 FILLER_67_412 ();
 sg13g2_fill_1 FILLER_67_414 ();
 sg13g2_fill_2 FILLER_67_425 ();
 sg13g2_fill_1 FILLER_67_432 ();
 sg13g2_fill_1 FILLER_67_460 ();
 sg13g2_fill_1 FILLER_67_492 ();
 sg13g2_fill_1 FILLER_67_569 ();
 sg13g2_decap_8 FILLER_67_578 ();
 sg13g2_decap_8 FILLER_67_585 ();
 sg13g2_decap_4 FILLER_67_592 ();
 sg13g2_fill_2 FILLER_67_596 ();
 sg13g2_fill_2 FILLER_67_614 ();
 sg13g2_decap_4 FILLER_67_633 ();
 sg13g2_fill_1 FILLER_67_637 ();
 sg13g2_decap_8 FILLER_67_652 ();
 sg13g2_decap_8 FILLER_67_659 ();
 sg13g2_fill_2 FILLER_67_666 ();
 sg13g2_fill_2 FILLER_67_678 ();
 sg13g2_fill_1 FILLER_67_680 ();
 sg13g2_decap_4 FILLER_67_689 ();
 sg13g2_decap_8 FILLER_67_712 ();
 sg13g2_decap_8 FILLER_67_740 ();
 sg13g2_decap_8 FILLER_67_747 ();
 sg13g2_decap_8 FILLER_67_754 ();
 sg13g2_fill_1 FILLER_67_761 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_decap_8 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_784 ();
 sg13g2_decap_8 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_798 ();
 sg13g2_decap_8 FILLER_67_805 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_854 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_9 ();
 sg13g2_fill_2 FILLER_68_38 ();
 sg13g2_fill_1 FILLER_68_40 ();
 sg13g2_decap_8 FILLER_68_54 ();
 sg13g2_fill_2 FILLER_68_61 ();
 sg13g2_fill_1 FILLER_68_63 ();
 sg13g2_fill_2 FILLER_68_78 ();
 sg13g2_fill_2 FILLER_68_102 ();
 sg13g2_fill_2 FILLER_68_113 ();
 sg13g2_fill_1 FILLER_68_125 ();
 sg13g2_fill_1 FILLER_68_152 ();
 sg13g2_decap_4 FILLER_68_162 ();
 sg13g2_fill_1 FILLER_68_176 ();
 sg13g2_fill_1 FILLER_68_200 ();
 sg13g2_fill_1 FILLER_68_216 ();
 sg13g2_fill_1 FILLER_68_226 ();
 sg13g2_fill_2 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_247 ();
 sg13g2_fill_2 FILLER_68_265 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_decap_4 FILLER_68_302 ();
 sg13g2_fill_1 FILLER_68_306 ();
 sg13g2_decap_4 FILLER_68_311 ();
 sg13g2_fill_2 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_403 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_fill_1 FILLER_68_439 ();
 sg13g2_fill_2 FILLER_68_470 ();
 sg13g2_fill_1 FILLER_68_472 ();
 sg13g2_decap_4 FILLER_68_491 ();
 sg13g2_decap_4 FILLER_68_541 ();
 sg13g2_fill_1 FILLER_68_545 ();
 sg13g2_fill_2 FILLER_68_563 ();
 sg13g2_fill_1 FILLER_68_565 ();
 sg13g2_decap_8 FILLER_68_592 ();
 sg13g2_decap_4 FILLER_68_599 ();
 sg13g2_fill_1 FILLER_68_603 ();
 sg13g2_decap_4 FILLER_68_612 ();
 sg13g2_fill_1 FILLER_68_616 ();
 sg13g2_fill_2 FILLER_68_625 ();
 sg13g2_fill_1 FILLER_68_627 ();
 sg13g2_fill_2 FILLER_68_648 ();
 sg13g2_decap_8 FILLER_68_668 ();
 sg13g2_fill_2 FILLER_68_690 ();
 sg13g2_fill_1 FILLER_68_692 ();
 sg13g2_fill_2 FILLER_68_715 ();
 sg13g2_fill_1 FILLER_68_717 ();
 sg13g2_fill_2 FILLER_68_729 ();
 sg13g2_fill_1 FILLER_68_731 ();
 sg13g2_decap_8 FILLER_68_749 ();
 sg13g2_decap_8 FILLER_68_756 ();
 sg13g2_decap_8 FILLER_68_763 ();
 sg13g2_decap_8 FILLER_68_770 ();
 sg13g2_decap_8 FILLER_68_777 ();
 sg13g2_decap_8 FILLER_68_784 ();
 sg13g2_decap_8 FILLER_68_791 ();
 sg13g2_decap_8 FILLER_68_798 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_decap_8 FILLER_68_812 ();
 sg13g2_decap_8 FILLER_68_819 ();
 sg13g2_decap_8 FILLER_68_826 ();
 sg13g2_decap_8 FILLER_68_833 ();
 sg13g2_decap_8 FILLER_68_840 ();
 sg13g2_decap_8 FILLER_68_847 ();
 sg13g2_decap_8 FILLER_68_854 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_94 ();
 sg13g2_fill_1 FILLER_69_121 ();
 sg13g2_fill_2 FILLER_69_185 ();
 sg13g2_fill_1 FILLER_69_187 ();
 sg13g2_fill_2 FILLER_69_267 ();
 sg13g2_decap_8 FILLER_69_274 ();
 sg13g2_fill_2 FILLER_69_281 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_fill_2 FILLER_69_294 ();
 sg13g2_decap_4 FILLER_69_327 ();
 sg13g2_fill_1 FILLER_69_331 ();
 sg13g2_decap_4 FILLER_69_336 ();
 sg13g2_fill_1 FILLER_69_345 ();
 sg13g2_decap_4 FILLER_69_350 ();
 sg13g2_fill_1 FILLER_69_354 ();
 sg13g2_decap_8 FILLER_69_368 ();
 sg13g2_fill_2 FILLER_69_375 ();
 sg13g2_fill_1 FILLER_69_377 ();
 sg13g2_fill_2 FILLER_69_382 ();
 sg13g2_fill_1 FILLER_69_398 ();
 sg13g2_fill_2 FILLER_69_418 ();
 sg13g2_fill_1 FILLER_69_420 ();
 sg13g2_fill_1 FILLER_69_460 ();
 sg13g2_decap_8 FILLER_69_527 ();
 sg13g2_fill_2 FILLER_69_534 ();
 sg13g2_decap_8 FILLER_69_567 ();
 sg13g2_fill_2 FILLER_69_574 ();
 sg13g2_decap_8 FILLER_69_580 ();
 sg13g2_decap_4 FILLER_69_587 ();
 sg13g2_decap_8 FILLER_69_594 ();
 sg13g2_decap_4 FILLER_69_601 ();
 sg13g2_decap_4 FILLER_69_609 ();
 sg13g2_decap_8 FILLER_69_651 ();
 sg13g2_decap_4 FILLER_69_658 ();
 sg13g2_fill_2 FILLER_69_662 ();
 sg13g2_fill_1 FILLER_69_672 ();
 sg13g2_decap_8 FILLER_69_707 ();
 sg13g2_fill_2 FILLER_69_718 ();
 sg13g2_decap_8 FILLER_69_739 ();
 sg13g2_decap_8 FILLER_69_746 ();
 sg13g2_decap_8 FILLER_69_753 ();
 sg13g2_decap_8 FILLER_69_760 ();
 sg13g2_decap_8 FILLER_69_767 ();
 sg13g2_decap_8 FILLER_69_774 ();
 sg13g2_decap_8 FILLER_69_781 ();
 sg13g2_decap_8 FILLER_69_788 ();
 sg13g2_decap_8 FILLER_69_795 ();
 sg13g2_decap_8 FILLER_69_802 ();
 sg13g2_decap_8 FILLER_69_809 ();
 sg13g2_decap_8 FILLER_69_816 ();
 sg13g2_decap_8 FILLER_69_823 ();
 sg13g2_decap_8 FILLER_69_830 ();
 sg13g2_decap_8 FILLER_69_837 ();
 sg13g2_decap_8 FILLER_69_844 ();
 sg13g2_decap_8 FILLER_69_851 ();
 sg13g2_decap_4 FILLER_69_858 ();
 sg13g2_fill_2 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_37 ();
 sg13g2_fill_1 FILLER_70_49 ();
 sg13g2_decap_4 FILLER_70_60 ();
 sg13g2_decap_4 FILLER_70_68 ();
 sg13g2_fill_1 FILLER_70_72 ();
 sg13g2_fill_1 FILLER_70_97 ();
 sg13g2_fill_2 FILLER_70_117 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_190 ();
 sg13g2_fill_2 FILLER_70_202 ();
 sg13g2_fill_1 FILLER_70_226 ();
 sg13g2_fill_2 FILLER_70_235 ();
 sg13g2_fill_2 FILLER_70_260 ();
 sg13g2_decap_4 FILLER_70_278 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_fill_2 FILLER_70_292 ();
 sg13g2_fill_2 FILLER_70_308 ();
 sg13g2_decap_4 FILLER_70_341 ();
 sg13g2_fill_2 FILLER_70_397 ();
 sg13g2_fill_2 FILLER_70_430 ();
 sg13g2_fill_1 FILLER_70_436 ();
 sg13g2_fill_1 FILLER_70_464 ();
 sg13g2_fill_1 FILLER_70_512 ();
 sg13g2_fill_2 FILLER_70_518 ();
 sg13g2_fill_2 FILLER_70_529 ();
 sg13g2_fill_1 FILLER_70_531 ();
 sg13g2_fill_1 FILLER_70_535 ();
 sg13g2_fill_1 FILLER_70_562 ();
 sg13g2_decap_8 FILLER_70_615 ();
 sg13g2_fill_2 FILLER_70_633 ();
 sg13g2_fill_1 FILLER_70_639 ();
 sg13g2_decap_8 FILLER_70_644 ();
 sg13g2_decap_4 FILLER_70_688 ();
 sg13g2_fill_1 FILLER_70_697 ();
 sg13g2_fill_2 FILLER_70_712 ();
 sg13g2_decap_8 FILLER_70_727 ();
 sg13g2_decap_8 FILLER_70_734 ();
 sg13g2_decap_8 FILLER_70_741 ();
 sg13g2_decap_8 FILLER_70_748 ();
 sg13g2_decap_8 FILLER_70_755 ();
 sg13g2_decap_8 FILLER_70_762 ();
 sg13g2_decap_8 FILLER_70_769 ();
 sg13g2_decap_8 FILLER_70_776 ();
 sg13g2_decap_8 FILLER_70_783 ();
 sg13g2_decap_8 FILLER_70_790 ();
 sg13g2_decap_8 FILLER_70_797 ();
 sg13g2_decap_8 FILLER_70_804 ();
 sg13g2_decap_8 FILLER_70_811 ();
 sg13g2_decap_8 FILLER_70_818 ();
 sg13g2_decap_8 FILLER_70_825 ();
 sg13g2_decap_8 FILLER_70_832 ();
 sg13g2_decap_8 FILLER_70_839 ();
 sg13g2_decap_8 FILLER_70_846 ();
 sg13g2_decap_8 FILLER_70_853 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_59 ();
 sg13g2_fill_2 FILLER_71_92 ();
 sg13g2_fill_2 FILLER_71_120 ();
 sg13g2_fill_1 FILLER_71_136 ();
 sg13g2_fill_2 FILLER_71_146 ();
 sg13g2_fill_1 FILLER_71_148 ();
 sg13g2_fill_2 FILLER_71_162 ();
 sg13g2_decap_4 FILLER_71_195 ();
 sg13g2_fill_1 FILLER_71_199 ();
 sg13g2_fill_1 FILLER_71_236 ();
 sg13g2_fill_1 FILLER_71_273 ();
 sg13g2_fill_2 FILLER_71_300 ();
 sg13g2_fill_1 FILLER_71_302 ();
 sg13g2_fill_2 FILLER_71_334 ();
 sg13g2_fill_1 FILLER_71_336 ();
 sg13g2_fill_2 FILLER_71_367 ();
 sg13g2_fill_1 FILLER_71_369 ();
 sg13g2_fill_2 FILLER_71_414 ();
 sg13g2_decap_4 FILLER_71_474 ();
 sg13g2_fill_2 FILLER_71_486 ();
 sg13g2_fill_1 FILLER_71_488 ();
 sg13g2_decap_4 FILLER_71_537 ();
 sg13g2_fill_2 FILLER_71_558 ();
 sg13g2_fill_2 FILLER_71_572 ();
 sg13g2_decap_8 FILLER_71_578 ();
 sg13g2_decap_4 FILLER_71_585 ();
 sg13g2_fill_1 FILLER_71_589 ();
 sg13g2_fill_1 FILLER_71_596 ();
 sg13g2_decap_8 FILLER_71_601 ();
 sg13g2_fill_2 FILLER_71_608 ();
 sg13g2_fill_1 FILLER_71_613 ();
 sg13g2_fill_2 FILLER_71_629 ();
 sg13g2_fill_2 FILLER_71_652 ();
 sg13g2_fill_1 FILLER_71_660 ();
 sg13g2_fill_1 FILLER_71_683 ();
 sg13g2_decap_4 FILLER_71_707 ();
 sg13g2_decap_8 FILLER_71_719 ();
 sg13g2_decap_8 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_733 ();
 sg13g2_decap_8 FILLER_71_740 ();
 sg13g2_decap_8 FILLER_71_747 ();
 sg13g2_decap_8 FILLER_71_754 ();
 sg13g2_decap_8 FILLER_71_761 ();
 sg13g2_decap_8 FILLER_71_768 ();
 sg13g2_decap_8 FILLER_71_775 ();
 sg13g2_decap_8 FILLER_71_782 ();
 sg13g2_decap_8 FILLER_71_789 ();
 sg13g2_decap_8 FILLER_71_796 ();
 sg13g2_decap_8 FILLER_71_803 ();
 sg13g2_decap_8 FILLER_71_810 ();
 sg13g2_decap_8 FILLER_71_817 ();
 sg13g2_decap_8 FILLER_71_824 ();
 sg13g2_decap_8 FILLER_71_831 ();
 sg13g2_decap_8 FILLER_71_838 ();
 sg13g2_decap_8 FILLER_71_845 ();
 sg13g2_decap_8 FILLER_71_852 ();
 sg13g2_fill_2 FILLER_71_859 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_9 ();
 sg13g2_fill_2 FILLER_72_36 ();
 sg13g2_fill_2 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_97 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_fill_1 FILLER_72_148 ();
 sg13g2_decap_4 FILLER_72_158 ();
 sg13g2_decap_4 FILLER_72_174 ();
 sg13g2_fill_1 FILLER_72_178 ();
 sg13g2_decap_4 FILLER_72_192 ();
 sg13g2_fill_1 FILLER_72_196 ();
 sg13g2_fill_1 FILLER_72_213 ();
 sg13g2_decap_4 FILLER_72_222 ();
 sg13g2_fill_1 FILLER_72_248 ();
 sg13g2_fill_2 FILLER_72_284 ();
 sg13g2_fill_2 FILLER_72_303 ();
 sg13g2_fill_1 FILLER_72_305 ();
 sg13g2_fill_2 FILLER_72_365 ();
 sg13g2_fill_1 FILLER_72_367 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_decap_8 FILLER_72_384 ();
 sg13g2_fill_1 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_decap_8 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_72_415 ();
 sg13g2_decap_8 FILLER_72_422 ();
 sg13g2_fill_2 FILLER_72_429 ();
 sg13g2_fill_1 FILLER_72_431 ();
 sg13g2_decap_4 FILLER_72_436 ();
 sg13g2_fill_1 FILLER_72_440 ();
 sg13g2_decap_8 FILLER_72_459 ();
 sg13g2_decap_8 FILLER_72_466 ();
 sg13g2_fill_1 FILLER_72_473 ();
 sg13g2_decap_8 FILLER_72_478 ();
 sg13g2_decap_4 FILLER_72_485 ();
 sg13g2_fill_2 FILLER_72_489 ();
 sg13g2_fill_2 FILLER_72_509 ();
 sg13g2_fill_1 FILLER_72_511 ();
 sg13g2_decap_8 FILLER_72_533 ();
 sg13g2_decap_8 FILLER_72_631 ();
 sg13g2_decap_4 FILLER_72_638 ();
 sg13g2_fill_2 FILLER_72_642 ();
 sg13g2_fill_2 FILLER_72_653 ();
 sg13g2_decap_8 FILLER_72_678 ();
 sg13g2_fill_1 FILLER_72_690 ();
 sg13g2_decap_4 FILLER_72_696 ();
 sg13g2_fill_2 FILLER_72_700 ();
 sg13g2_fill_1 FILLER_72_715 ();
 sg13g2_decap_8 FILLER_72_720 ();
 sg13g2_decap_8 FILLER_72_727 ();
 sg13g2_decap_8 FILLER_72_734 ();
 sg13g2_decap_8 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_748 ();
 sg13g2_decap_8 FILLER_72_755 ();
 sg13g2_decap_8 FILLER_72_762 ();
 sg13g2_decap_8 FILLER_72_769 ();
 sg13g2_decap_8 FILLER_72_776 ();
 sg13g2_decap_8 FILLER_72_783 ();
 sg13g2_decap_8 FILLER_72_790 ();
 sg13g2_decap_8 FILLER_72_797 ();
 sg13g2_decap_8 FILLER_72_804 ();
 sg13g2_decap_8 FILLER_72_811 ();
 sg13g2_decap_8 FILLER_72_818 ();
 sg13g2_decap_8 FILLER_72_825 ();
 sg13g2_decap_8 FILLER_72_832 ();
 sg13g2_decap_8 FILLER_72_839 ();
 sg13g2_decap_8 FILLER_72_846 ();
 sg13g2_decap_8 FILLER_72_853 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_4 FILLER_73_25 ();
 sg13g2_fill_2 FILLER_73_29 ();
 sg13g2_fill_2 FILLER_73_72 ();
 sg13g2_fill_1 FILLER_73_74 ();
 sg13g2_fill_1 FILLER_73_95 ();
 sg13g2_fill_2 FILLER_73_107 ();
 sg13g2_fill_1 FILLER_73_109 ();
 sg13g2_fill_1 FILLER_73_131 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_2 FILLER_73_167 ();
 sg13g2_fill_1 FILLER_73_169 ();
 sg13g2_fill_2 FILLER_73_192 ();
 sg13g2_fill_1 FILLER_73_194 ();
 sg13g2_fill_1 FILLER_73_250 ();
 sg13g2_fill_2 FILLER_73_292 ();
 sg13g2_fill_1 FILLER_73_294 ();
 sg13g2_fill_2 FILLER_73_330 ();
 sg13g2_fill_1 FILLER_73_340 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_decap_8 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_73_414 ();
 sg13g2_decap_8 FILLER_73_421 ();
 sg13g2_decap_8 FILLER_73_428 ();
 sg13g2_decap_8 FILLER_73_435 ();
 sg13g2_fill_2 FILLER_73_442 ();
 sg13g2_decap_8 FILLER_73_449 ();
 sg13g2_decap_8 FILLER_73_456 ();
 sg13g2_fill_2 FILLER_73_542 ();
 sg13g2_decap_8 FILLER_73_557 ();
 sg13g2_fill_2 FILLER_73_564 ();
 sg13g2_fill_2 FILLER_73_580 ();
 sg13g2_decap_8 FILLER_73_611 ();
 sg13g2_decap_8 FILLER_73_618 ();
 sg13g2_fill_1 FILLER_73_625 ();
 sg13g2_decap_8 FILLER_73_652 ();
 sg13g2_decap_8 FILLER_73_659 ();
 sg13g2_decap_8 FILLER_73_670 ();
 sg13g2_decap_4 FILLER_73_677 ();
 sg13g2_fill_1 FILLER_73_681 ();
 sg13g2_decap_8 FILLER_73_685 ();
 sg13g2_fill_2 FILLER_73_692 ();
 sg13g2_fill_1 FILLER_73_694 ();
 sg13g2_decap_4 FILLER_73_699 ();
 sg13g2_fill_2 FILLER_73_703 ();
 sg13g2_decap_8 FILLER_73_731 ();
 sg13g2_decap_8 FILLER_73_738 ();
 sg13g2_decap_8 FILLER_73_745 ();
 sg13g2_decap_8 FILLER_73_752 ();
 sg13g2_decap_8 FILLER_73_759 ();
 sg13g2_decap_8 FILLER_73_766 ();
 sg13g2_decap_8 FILLER_73_773 ();
 sg13g2_decap_8 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_4 FILLER_73_857 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_4 FILLER_74_21 ();
 sg13g2_fill_1 FILLER_74_25 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_109 ();
 sg13g2_fill_1 FILLER_74_143 ();
 sg13g2_decap_4 FILLER_74_156 ();
 sg13g2_fill_1 FILLER_74_160 ();
 sg13g2_fill_2 FILLER_74_174 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_fill_1 FILLER_74_182 ();
 sg13g2_fill_2 FILLER_74_188 ();
 sg13g2_fill_1 FILLER_74_190 ();
 sg13g2_decap_4 FILLER_74_230 ();
 sg13g2_fill_1 FILLER_74_234 ();
 sg13g2_fill_2 FILLER_74_239 ();
 sg13g2_fill_1 FILLER_74_241 ();
 sg13g2_decap_4 FILLER_74_320 ();
 sg13g2_fill_2 FILLER_74_324 ();
 sg13g2_decap_8 FILLER_74_330 ();
 sg13g2_decap_8 FILLER_74_351 ();
 sg13g2_fill_1 FILLER_74_358 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_4 FILLER_74_370 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_fill_2 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_412 ();
 sg13g2_decap_8 FILLER_74_424 ();
 sg13g2_decap_4 FILLER_74_431 ();
 sg13g2_fill_2 FILLER_74_435 ();
 sg13g2_decap_8 FILLER_74_458 ();
 sg13g2_decap_8 FILLER_74_465 ();
 sg13g2_decap_8 FILLER_74_472 ();
 sg13g2_decap_8 FILLER_74_479 ();
 sg13g2_decap_8 FILLER_74_486 ();
 sg13g2_fill_1 FILLER_74_493 ();
 sg13g2_decap_4 FILLER_74_512 ();
 sg13g2_fill_1 FILLER_74_516 ();
 sg13g2_fill_2 FILLER_74_533 ();
 sg13g2_decap_4 FILLER_74_540 ();
 sg13g2_decap_8 FILLER_74_549 ();
 sg13g2_fill_1 FILLER_74_556 ();
 sg13g2_decap_8 FILLER_74_575 ();
 sg13g2_fill_2 FILLER_74_582 ();
 sg13g2_decap_8 FILLER_74_609 ();
 sg13g2_decap_8 FILLER_74_616 ();
 sg13g2_decap_8 FILLER_74_623 ();
 sg13g2_decap_8 FILLER_74_630 ();
 sg13g2_decap_8 FILLER_74_641 ();
 sg13g2_decap_8 FILLER_74_648 ();
 sg13g2_fill_2 FILLER_74_681 ();
 sg13g2_fill_1 FILLER_74_683 ();
 sg13g2_decap_8 FILLER_74_716 ();
 sg13g2_decap_8 FILLER_74_723 ();
 sg13g2_decap_8 FILLER_74_730 ();
 sg13g2_decap_8 FILLER_74_737 ();
 sg13g2_decap_8 FILLER_74_744 ();
 sg13g2_decap_8 FILLER_74_751 ();
 sg13g2_decap_8 FILLER_74_758 ();
 sg13g2_decap_8 FILLER_74_765 ();
 sg13g2_decap_8 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_779 ();
 sg13g2_decap_8 FILLER_74_786 ();
 sg13g2_decap_8 FILLER_74_793 ();
 sg13g2_decap_8 FILLER_74_800 ();
 sg13g2_decap_8 FILLER_74_807 ();
 sg13g2_decap_8 FILLER_74_814 ();
 sg13g2_decap_8 FILLER_74_821 ();
 sg13g2_decap_8 FILLER_74_828 ();
 sg13g2_decap_8 FILLER_74_835 ();
 sg13g2_decap_8 FILLER_74_842 ();
 sg13g2_decap_8 FILLER_74_849 ();
 sg13g2_decap_4 FILLER_74_856 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_4 FILLER_75_49 ();
 sg13g2_fill_2 FILLER_75_53 ();
 sg13g2_decap_8 FILLER_75_58 ();
 sg13g2_decap_8 FILLER_75_65 ();
 sg13g2_decap_4 FILLER_75_72 ();
 sg13g2_fill_1 FILLER_75_76 ();
 sg13g2_fill_2 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_104 ();
 sg13g2_fill_2 FILLER_75_113 ();
 sg13g2_decap_8 FILLER_75_153 ();
 sg13g2_decap_8 FILLER_75_160 ();
 sg13g2_fill_2 FILLER_75_167 ();
 sg13g2_fill_1 FILLER_75_169 ();
 sg13g2_fill_2 FILLER_75_175 ();
 sg13g2_fill_1 FILLER_75_177 ();
 sg13g2_fill_1 FILLER_75_183 ();
 sg13g2_fill_1 FILLER_75_195 ();
 sg13g2_fill_1 FILLER_75_213 ();
 sg13g2_fill_2 FILLER_75_223 ();
 sg13g2_fill_1 FILLER_75_225 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_4 FILLER_75_245 ();
 sg13g2_fill_2 FILLER_75_249 ();
 sg13g2_fill_1 FILLER_75_256 ();
 sg13g2_decap_8 FILLER_75_265 ();
 sg13g2_decap_8 FILLER_75_272 ();
 sg13g2_fill_1 FILLER_75_283 ();
 sg13g2_fill_2 FILLER_75_314 ();
 sg13g2_fill_2 FILLER_75_382 ();
 sg13g2_fill_1 FILLER_75_384 ();
 sg13g2_fill_2 FILLER_75_420 ();
 sg13g2_decap_8 FILLER_75_435 ();
 sg13g2_fill_2 FILLER_75_442 ();
 sg13g2_fill_1 FILLER_75_444 ();
 sg13g2_decap_8 FILLER_75_449 ();
 sg13g2_decap_8 FILLER_75_456 ();
 sg13g2_decap_8 FILLER_75_463 ();
 sg13g2_decap_8 FILLER_75_470 ();
 sg13g2_decap_8 FILLER_75_477 ();
 sg13g2_decap_4 FILLER_75_484 ();
 sg13g2_fill_2 FILLER_75_501 ();
 sg13g2_decap_8 FILLER_75_523 ();
 sg13g2_fill_2 FILLER_75_530 ();
 sg13g2_fill_1 FILLER_75_548 ();
 sg13g2_fill_2 FILLER_75_574 ();
 sg13g2_fill_1 FILLER_75_576 ();
 sg13g2_fill_2 FILLER_75_589 ();
 sg13g2_fill_1 FILLER_75_591 ();
 sg13g2_decap_8 FILLER_75_606 ();
 sg13g2_decap_8 FILLER_75_613 ();
 sg13g2_decap_8 FILLER_75_620 ();
 sg13g2_decap_8 FILLER_75_627 ();
 sg13g2_decap_8 FILLER_75_634 ();
 sg13g2_decap_8 FILLER_75_641 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_decap_8 FILLER_75_655 ();
 sg13g2_decap_8 FILLER_75_662 ();
 sg13g2_decap_8 FILLER_75_669 ();
 sg13g2_decap_8 FILLER_75_676 ();
 sg13g2_decap_8 FILLER_75_683 ();
 sg13g2_decap_8 FILLER_75_690 ();
 sg13g2_decap_4 FILLER_75_697 ();
 sg13g2_fill_1 FILLER_75_701 ();
 sg13g2_decap_8 FILLER_75_707 ();
 sg13g2_decap_8 FILLER_75_714 ();
 sg13g2_decap_8 FILLER_75_721 ();
 sg13g2_decap_8 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_735 ();
 sg13g2_decap_8 FILLER_75_742 ();
 sg13g2_decap_8 FILLER_75_749 ();
 sg13g2_decap_8 FILLER_75_756 ();
 sg13g2_decap_8 FILLER_75_763 ();
 sg13g2_decap_8 FILLER_75_770 ();
 sg13g2_decap_8 FILLER_75_777 ();
 sg13g2_decap_8 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_791 ();
 sg13g2_decap_8 FILLER_75_798 ();
 sg13g2_decap_8 FILLER_75_805 ();
 sg13g2_decap_8 FILLER_75_812 ();
 sg13g2_decap_8 FILLER_75_819 ();
 sg13g2_decap_8 FILLER_75_826 ();
 sg13g2_decap_8 FILLER_75_833 ();
 sg13g2_decap_8 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_75_847 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_fill_2 FILLER_76_70 ();
 sg13g2_fill_1 FILLER_76_72 ();
 sg13g2_fill_2 FILLER_76_99 ();
 sg13g2_fill_1 FILLER_76_101 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_1 FILLER_76_113 ();
 sg13g2_fill_2 FILLER_76_119 ();
 sg13g2_fill_1 FILLER_76_121 ();
 sg13g2_fill_1 FILLER_76_152 ();
 sg13g2_fill_1 FILLER_76_171 ();
 sg13g2_fill_2 FILLER_76_198 ();
 sg13g2_fill_1 FILLER_76_226 ();
 sg13g2_fill_2 FILLER_76_241 ();
 sg13g2_decap_8 FILLER_76_269 ();
 sg13g2_decap_4 FILLER_76_276 ();
 sg13g2_fill_1 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_285 ();
 sg13g2_fill_2 FILLER_76_335 ();
 sg13g2_fill_1 FILLER_76_337 ();
 sg13g2_fill_2 FILLER_76_398 ();
 sg13g2_decap_8 FILLER_76_461 ();
 sg13g2_decap_8 FILLER_76_468 ();
 sg13g2_decap_8 FILLER_76_475 ();
 sg13g2_decap_8 FILLER_76_482 ();
 sg13g2_decap_4 FILLER_76_489 ();
 sg13g2_fill_2 FILLER_76_506 ();
 sg13g2_decap_8 FILLER_76_522 ();
 sg13g2_fill_2 FILLER_76_529 ();
 sg13g2_fill_1 FILLER_76_546 ();
 sg13g2_fill_2 FILLER_76_555 ();
 sg13g2_fill_1 FILLER_76_557 ();
 sg13g2_decap_8 FILLER_76_570 ();
 sg13g2_fill_1 FILLER_76_577 ();
 sg13g2_decap_8 FILLER_76_586 ();
 sg13g2_decap_8 FILLER_76_593 ();
 sg13g2_decap_8 FILLER_76_600 ();
 sg13g2_decap_8 FILLER_76_607 ();
 sg13g2_decap_8 FILLER_76_614 ();
 sg13g2_decap_8 FILLER_76_621 ();
 sg13g2_decap_8 FILLER_76_628 ();
 sg13g2_decap_8 FILLER_76_635 ();
 sg13g2_decap_8 FILLER_76_642 ();
 sg13g2_decap_8 FILLER_76_649 ();
 sg13g2_decap_8 FILLER_76_656 ();
 sg13g2_decap_8 FILLER_76_663 ();
 sg13g2_decap_8 FILLER_76_670 ();
 sg13g2_decap_8 FILLER_76_677 ();
 sg13g2_decap_8 FILLER_76_684 ();
 sg13g2_decap_8 FILLER_76_691 ();
 sg13g2_decap_8 FILLER_76_698 ();
 sg13g2_decap_8 FILLER_76_705 ();
 sg13g2_decap_8 FILLER_76_712 ();
 sg13g2_decap_8 FILLER_76_719 ();
 sg13g2_decap_8 FILLER_76_726 ();
 sg13g2_decap_8 FILLER_76_733 ();
 sg13g2_decap_8 FILLER_76_740 ();
 sg13g2_decap_8 FILLER_76_747 ();
 sg13g2_decap_8 FILLER_76_754 ();
 sg13g2_decap_8 FILLER_76_761 ();
 sg13g2_decap_8 FILLER_76_768 ();
 sg13g2_decap_8 FILLER_76_775 ();
 sg13g2_decap_8 FILLER_76_782 ();
 sg13g2_decap_8 FILLER_76_789 ();
 sg13g2_decap_8 FILLER_76_796 ();
 sg13g2_decap_8 FILLER_76_803 ();
 sg13g2_decap_8 FILLER_76_810 ();
 sg13g2_decap_8 FILLER_76_817 ();
 sg13g2_decap_8 FILLER_76_824 ();
 sg13g2_decap_8 FILLER_76_831 ();
 sg13g2_decap_8 FILLER_76_838 ();
 sg13g2_decap_8 FILLER_76_845 ();
 sg13g2_decap_8 FILLER_76_852 ();
 sg13g2_fill_2 FILLER_76_859 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_4 FILLER_77_77 ();
 sg13g2_fill_2 FILLER_77_81 ();
 sg13g2_fill_2 FILLER_77_87 ();
 sg13g2_decap_4 FILLER_77_120 ();
 sg13g2_decap_4 FILLER_77_129 ();
 sg13g2_fill_1 FILLER_77_133 ();
 sg13g2_decap_4 FILLER_77_161 ();
 sg13g2_fill_1 FILLER_77_216 ();
 sg13g2_fill_2 FILLER_77_226 ();
 sg13g2_decap_4 FILLER_77_262 ();
 sg13g2_fill_1 FILLER_77_297 ();
 sg13g2_decap_4 FILLER_77_342 ();
 sg13g2_fill_1 FILLER_77_346 ();
 sg13g2_decap_4 FILLER_77_368 ();
 sg13g2_decap_8 FILLER_77_377 ();
 sg13g2_decap_8 FILLER_77_384 ();
 sg13g2_decap_4 FILLER_77_391 ();
 sg13g2_decap_4 FILLER_77_425 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_77_439 ();
 sg13g2_decap_8 FILLER_77_450 ();
 sg13g2_decap_8 FILLER_77_457 ();
 sg13g2_decap_8 FILLER_77_464 ();
 sg13g2_decap_8 FILLER_77_471 ();
 sg13g2_decap_8 FILLER_77_478 ();
 sg13g2_decap_8 FILLER_77_485 ();
 sg13g2_decap_8 FILLER_77_492 ();
 sg13g2_decap_8 FILLER_77_499 ();
 sg13g2_decap_8 FILLER_77_506 ();
 sg13g2_decap_8 FILLER_77_513 ();
 sg13g2_decap_8 FILLER_77_520 ();
 sg13g2_decap_8 FILLER_77_527 ();
 sg13g2_decap_8 FILLER_77_534 ();
 sg13g2_decap_8 FILLER_77_541 ();
 sg13g2_decap_8 FILLER_77_548 ();
 sg13g2_decap_8 FILLER_77_555 ();
 sg13g2_decap_8 FILLER_77_562 ();
 sg13g2_decap_8 FILLER_77_569 ();
 sg13g2_decap_8 FILLER_77_576 ();
 sg13g2_decap_8 FILLER_77_583 ();
 sg13g2_decap_8 FILLER_77_590 ();
 sg13g2_decap_8 FILLER_77_597 ();
 sg13g2_decap_8 FILLER_77_604 ();
 sg13g2_decap_8 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_decap_8 FILLER_77_625 ();
 sg13g2_decap_8 FILLER_77_632 ();
 sg13g2_decap_8 FILLER_77_639 ();
 sg13g2_decap_8 FILLER_77_646 ();
 sg13g2_decap_8 FILLER_77_653 ();
 sg13g2_decap_8 FILLER_77_660 ();
 sg13g2_decap_8 FILLER_77_667 ();
 sg13g2_decap_8 FILLER_77_674 ();
 sg13g2_decap_8 FILLER_77_681 ();
 sg13g2_decap_8 FILLER_77_688 ();
 sg13g2_decap_8 FILLER_77_695 ();
 sg13g2_decap_8 FILLER_77_702 ();
 sg13g2_decap_8 FILLER_77_709 ();
 sg13g2_decap_8 FILLER_77_716 ();
 sg13g2_decap_8 FILLER_77_723 ();
 sg13g2_decap_8 FILLER_77_730 ();
 sg13g2_decap_8 FILLER_77_737 ();
 sg13g2_decap_8 FILLER_77_744 ();
 sg13g2_decap_8 FILLER_77_751 ();
 sg13g2_decap_8 FILLER_77_758 ();
 sg13g2_decap_8 FILLER_77_765 ();
 sg13g2_decap_8 FILLER_77_772 ();
 sg13g2_decap_8 FILLER_77_779 ();
 sg13g2_decap_8 FILLER_77_786 ();
 sg13g2_decap_8 FILLER_77_793 ();
 sg13g2_decap_8 FILLER_77_800 ();
 sg13g2_decap_8 FILLER_77_807 ();
 sg13g2_decap_8 FILLER_77_814 ();
 sg13g2_decap_8 FILLER_77_821 ();
 sg13g2_decap_8 FILLER_77_828 ();
 sg13g2_decap_8 FILLER_77_835 ();
 sg13g2_decap_8 FILLER_77_842 ();
 sg13g2_decap_8 FILLER_77_849 ();
 sg13g2_decap_4 FILLER_77_856 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_4 FILLER_78_77 ();
 sg13g2_fill_2 FILLER_78_81 ();
 sg13g2_fill_1 FILLER_78_109 ();
 sg13g2_fill_2 FILLER_78_163 ();
 sg13g2_fill_1 FILLER_78_165 ();
 sg13g2_fill_1 FILLER_78_232 ();
 sg13g2_decap_8 FILLER_78_255 ();
 sg13g2_decap_8 FILLER_78_262 ();
 sg13g2_decap_8 FILLER_78_269 ();
 sg13g2_decap_8 FILLER_78_276 ();
 sg13g2_decap_8 FILLER_78_283 ();
 sg13g2_decap_4 FILLER_78_290 ();
 sg13g2_fill_1 FILLER_78_294 ();
 sg13g2_fill_2 FILLER_78_326 ();
 sg13g2_fill_1 FILLER_78_354 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_78_435 ();
 sg13g2_decap_8 FILLER_78_442 ();
 sg13g2_decap_8 FILLER_78_449 ();
 sg13g2_decap_8 FILLER_78_456 ();
 sg13g2_decap_8 FILLER_78_463 ();
 sg13g2_decap_8 FILLER_78_470 ();
 sg13g2_decap_8 FILLER_78_477 ();
 sg13g2_decap_8 FILLER_78_484 ();
 sg13g2_decap_8 FILLER_78_491 ();
 sg13g2_decap_8 FILLER_78_498 ();
 sg13g2_decap_8 FILLER_78_505 ();
 sg13g2_decap_8 FILLER_78_512 ();
 sg13g2_decap_8 FILLER_78_519 ();
 sg13g2_decap_8 FILLER_78_526 ();
 sg13g2_decap_8 FILLER_78_533 ();
 sg13g2_decap_8 FILLER_78_540 ();
 sg13g2_decap_8 FILLER_78_547 ();
 sg13g2_decap_8 FILLER_78_554 ();
 sg13g2_decap_8 FILLER_78_561 ();
 sg13g2_decap_8 FILLER_78_568 ();
 sg13g2_decap_8 FILLER_78_575 ();
 sg13g2_decap_8 FILLER_78_582 ();
 sg13g2_decap_8 FILLER_78_589 ();
 sg13g2_decap_8 FILLER_78_596 ();
 sg13g2_decap_8 FILLER_78_603 ();
 sg13g2_decap_8 FILLER_78_610 ();
 sg13g2_decap_8 FILLER_78_617 ();
 sg13g2_decap_8 FILLER_78_624 ();
 sg13g2_decap_8 FILLER_78_631 ();
 sg13g2_decap_8 FILLER_78_638 ();
 sg13g2_decap_8 FILLER_78_645 ();
 sg13g2_decap_8 FILLER_78_652 ();
 sg13g2_decap_8 FILLER_78_659 ();
 sg13g2_decap_8 FILLER_78_666 ();
 sg13g2_decap_8 FILLER_78_673 ();
 sg13g2_decap_8 FILLER_78_680 ();
 sg13g2_decap_8 FILLER_78_687 ();
 sg13g2_decap_8 FILLER_78_694 ();
 sg13g2_decap_8 FILLER_78_701 ();
 sg13g2_decap_8 FILLER_78_708 ();
 sg13g2_decap_8 FILLER_78_715 ();
 sg13g2_decap_8 FILLER_78_722 ();
 sg13g2_decap_8 FILLER_78_729 ();
 sg13g2_decap_8 FILLER_78_736 ();
 sg13g2_decap_8 FILLER_78_743 ();
 sg13g2_decap_8 FILLER_78_750 ();
 sg13g2_decap_8 FILLER_78_757 ();
 sg13g2_decap_8 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_771 ();
 sg13g2_decap_8 FILLER_78_778 ();
 sg13g2_decap_8 FILLER_78_785 ();
 sg13g2_decap_8 FILLER_78_792 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_806 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_8 FILLER_78_820 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_4 FILLER_79_91 ();
 sg13g2_fill_1 FILLER_79_95 ();
 sg13g2_fill_1 FILLER_79_108 ();
 sg13g2_decap_4 FILLER_79_113 ();
 sg13g2_fill_2 FILLER_79_117 ();
 sg13g2_decap_8 FILLER_79_128 ();
 sg13g2_fill_2 FILLER_79_135 ();
 sg13g2_decap_8 FILLER_79_150 ();
 sg13g2_decap_8 FILLER_79_166 ();
 sg13g2_decap_4 FILLER_79_173 ();
 sg13g2_fill_2 FILLER_79_181 ();
 sg13g2_decap_4 FILLER_79_191 ();
 sg13g2_fill_2 FILLER_79_195 ();
 sg13g2_decap_8 FILLER_79_201 ();
 sg13g2_fill_2 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_210 ();
 sg13g2_fill_2 FILLER_79_215 ();
 sg13g2_fill_1 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_223 ();
 sg13g2_fill_2 FILLER_79_230 ();
 sg13g2_decap_8 FILLER_79_236 ();
 sg13g2_decap_8 FILLER_79_243 ();
 sg13g2_decap_8 FILLER_79_250 ();
 sg13g2_decap_8 FILLER_79_257 ();
 sg13g2_decap_8 FILLER_79_264 ();
 sg13g2_decap_8 FILLER_79_271 ();
 sg13g2_decap_8 FILLER_79_278 ();
 sg13g2_decap_8 FILLER_79_285 ();
 sg13g2_decap_8 FILLER_79_292 ();
 sg13g2_decap_8 FILLER_79_299 ();
 sg13g2_decap_4 FILLER_79_306 ();
 sg13g2_fill_1 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_4 FILLER_79_329 ();
 sg13g2_fill_2 FILLER_79_333 ();
 sg13g2_decap_4 FILLER_79_348 ();
 sg13g2_fill_1 FILLER_79_352 ();
 sg13g2_decap_4 FILLER_79_362 ();
 sg13g2_decap_8 FILLER_79_379 ();
 sg13g2_decap_4 FILLER_79_386 ();
 sg13g2_fill_1 FILLER_79_390 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_79_409 ();
 sg13g2_decap_4 FILLER_79_416 ();
 sg13g2_decap_8 FILLER_79_424 ();
 sg13g2_decap_8 FILLER_79_431 ();
 sg13g2_decap_8 FILLER_79_438 ();
 sg13g2_decap_8 FILLER_79_445 ();
 sg13g2_decap_8 FILLER_79_452 ();
 sg13g2_decap_8 FILLER_79_459 ();
 sg13g2_decap_8 FILLER_79_466 ();
 sg13g2_decap_8 FILLER_79_473 ();
 sg13g2_decap_8 FILLER_79_480 ();
 sg13g2_decap_8 FILLER_79_487 ();
 sg13g2_decap_8 FILLER_79_494 ();
 sg13g2_decap_8 FILLER_79_501 ();
 sg13g2_decap_8 FILLER_79_508 ();
 sg13g2_decap_8 FILLER_79_515 ();
 sg13g2_decap_8 FILLER_79_522 ();
 sg13g2_decap_8 FILLER_79_529 ();
 sg13g2_decap_8 FILLER_79_536 ();
 sg13g2_decap_8 FILLER_79_543 ();
 sg13g2_decap_8 FILLER_79_550 ();
 sg13g2_decap_8 FILLER_79_557 ();
 sg13g2_decap_8 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_571 ();
 sg13g2_decap_8 FILLER_79_578 ();
 sg13g2_decap_8 FILLER_79_585 ();
 sg13g2_decap_8 FILLER_79_592 ();
 sg13g2_decap_8 FILLER_79_599 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_8 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_620 ();
 sg13g2_decap_8 FILLER_79_627 ();
 sg13g2_decap_8 FILLER_79_634 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_648 ();
 sg13g2_decap_8 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_662 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_8 FILLER_79_676 ();
 sg13g2_decap_8 FILLER_79_683 ();
 sg13g2_decap_8 FILLER_79_690 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_725 ();
 sg13g2_decap_8 FILLER_79_732 ();
 sg13g2_decap_8 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_767 ();
 sg13g2_decap_8 FILLER_79_774 ();
 sg13g2_decap_8 FILLER_79_781 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_4 FILLER_79_858 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_250 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_decap_8 FILLER_80_341 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_decap_8 FILLER_80_355 ();
 sg13g2_decap_8 FILLER_80_362 ();
 sg13g2_decap_8 FILLER_80_369 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_decap_8 FILLER_80_429 ();
 sg13g2_decap_8 FILLER_80_436 ();
 sg13g2_decap_8 FILLER_80_443 ();
 sg13g2_decap_8 FILLER_80_450 ();
 sg13g2_decap_8 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_464 ();
 sg13g2_decap_8 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_478 ();
 sg13g2_decap_8 FILLER_80_485 ();
 sg13g2_decap_8 FILLER_80_492 ();
 sg13g2_decap_8 FILLER_80_499 ();
 sg13g2_decap_8 FILLER_80_506 ();
 sg13g2_decap_8 FILLER_80_513 ();
 sg13g2_decap_8 FILLER_80_520 ();
 sg13g2_decap_8 FILLER_80_527 ();
 sg13g2_decap_8 FILLER_80_534 ();
 sg13g2_decap_8 FILLER_80_541 ();
 sg13g2_decap_8 FILLER_80_548 ();
 sg13g2_decap_8 FILLER_80_555 ();
 sg13g2_decap_8 FILLER_80_562 ();
 sg13g2_decap_8 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_576 ();
 sg13g2_decap_8 FILLER_80_583 ();
 sg13g2_decap_8 FILLER_80_590 ();
 sg13g2_decap_8 FILLER_80_597 ();
 sg13g2_decap_8 FILLER_80_604 ();
 sg13g2_decap_8 FILLER_80_611 ();
 sg13g2_decap_8 FILLER_80_618 ();
 sg13g2_decap_8 FILLER_80_625 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_8 FILLER_80_639 ();
 sg13g2_decap_8 FILLER_80_646 ();
 sg13g2_decap_8 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_660 ();
 sg13g2_decap_8 FILLER_80_667 ();
 sg13g2_decap_8 FILLER_80_674 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_695 ();
 sg13g2_decap_8 FILLER_80_702 ();
 sg13g2_decap_8 FILLER_80_709 ();
 sg13g2_decap_8 FILLER_80_716 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_4 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net277;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
endmodule

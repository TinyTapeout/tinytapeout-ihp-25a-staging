module tt_um_jamesrosssharp_tiny1bitam (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire COMP_OUT;
 wire PWM_OUT;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire clknet_0_clk;
 wire \am_sdr0.count[0] ;
 wire \am_sdr0.count[1] ;
 wire \am_sdr0.count[2] ;
 wire \am_sdr0.count[3] ;
 wire \am_sdr0.count[4] ;
 wire \am_sdr0.count[5] ;
 wire \am_sdr0.count[6] ;
 wire \am_sdr0.count[7] ;
 wire \am_sdr0.det0.alpha_yn_1[0] ;
 wire \am_sdr0.det0.env_det[0] ;
 wire \am_sdr0.det0.env_out[0] ;
 wire \am_sdr0.det0.env_out[1] ;
 wire \am_sdr0.det0.env_out[2] ;
 wire \am_sdr0.det0.env_out[3] ;
 wire \am_sdr0.det0.env_out[4] ;
 wire \am_sdr0.det0.env_out[5] ;
 wire \am_sdr0.det0.env_out[6] ;
 wire \am_sdr0.det0.env_out[7] ;
 wire \am_sdr0.det0.ifreq[1] ;
 wire \am_sdr0.det0.ifreq[2] ;
 wire \am_sdr0.det0.ifreq[3] ;
 wire \am_sdr0.det0.ifreq[4] ;
 wire \am_sdr0.det0.ifreq[5] ;
 wire \am_sdr0.det0.ifreq[6] ;
 wire \am_sdr0.det0.ifreq[7] ;
 wire \am_sdr0.det0.yn_1[10] ;
 wire \am_sdr0.det0.yn_1[11] ;
 wire \am_sdr0.det0.yn_1[12] ;
 wire \am_sdr0.det0.yn_1[13] ;
 wire \am_sdr0.det0.yn_1[14] ;
 wire \am_sdr0.det0.yn_1[15] ;
 wire \am_sdr0.det0.yn_1[16] ;
 wire \am_sdr0.det0.yn_1[17] ;
 wire \am_sdr0.det0.yn_1[18] ;
 wire \am_sdr0.det0.yn_1[19] ;
 wire \am_sdr0.det0.yn_1[1] ;
 wire \am_sdr0.det0.yn_1[2] ;
 wire \am_sdr0.det0.yn_1[3] ;
 wire \am_sdr0.det0.yn_1[4] ;
 wire \am_sdr0.det0.yn_1[5] ;
 wire \am_sdr0.det0.yn_1[6] ;
 wire \am_sdr0.det0.yn_1[7] ;
 wire \am_sdr0.det0.yn_1[8] ;
 wire \am_sdr0.det0.yn_1[9] ;
 wire \am_sdr0.filt0.gain_spi[0] ;
 wire \am_sdr0.filt0.gain_spi[1] ;
 wire \am_sdr0.filt0.gain_spi[2] ;
 wire \am_sdr0.filt0.if_out[0] ;
 wire \am_sdr0.filt0.if_out[1] ;
 wire \am_sdr0.filt0.if_out[2] ;
 wire \am_sdr0.filt0.if_out[3] ;
 wire \am_sdr0.filt0.if_out[4] ;
 wire \am_sdr0.filt0.if_out[5] ;
 wire \am_sdr0.filt0.if_out[6] ;
 wire \am_sdr0.filt0.if_out[7] ;
 wire \am_sdr0.filt0.mul_a1[0] ;
 wire \am_sdr0.filt0.mul_a1[1] ;
 wire \am_sdr0.filt0.mul_a2[1] ;
 wire \am_sdr0.filt0.mul_b2[0] ;
 wire \am_sdr0.filt0.xn_1[0] ;
 wire \am_sdr0.filt0.xn_1[1] ;
 wire \am_sdr0.filt0.xn_1[2] ;
 wire \am_sdr0.filt0.xn_1[3] ;
 wire \am_sdr0.filt0.xn_1[4] ;
 wire \am_sdr0.filt0.xn_1[5] ;
 wire \am_sdr0.filt0.xn_1[6] ;
 wire \am_sdr0.filt0.xn_1[7] ;
 wire \am_sdr0.filt0.xn_2[1] ;
 wire \am_sdr0.filt0.xn_2[2] ;
 wire \am_sdr0.filt0.xn_2[3] ;
 wire \am_sdr0.filt0.xn_2[4] ;
 wire \am_sdr0.filt0.xn_2[5] ;
 wire \am_sdr0.filt0.xn_2[6] ;
 wire \am_sdr0.filt0.xn_2[7] ;
 wire \am_sdr0.filt0.yn_1[10] ;
 wire \am_sdr0.filt0.yn_1[11] ;
 wire \am_sdr0.filt0.yn_1[12] ;
 wire \am_sdr0.filt0.yn_1[13] ;
 wire \am_sdr0.filt0.yn_1[2] ;
 wire \am_sdr0.filt0.yn_1[3] ;
 wire \am_sdr0.filt0.yn_1[4] ;
 wire \am_sdr0.filt0.yn_1[5] ;
 wire \am_sdr0.filt0.yn_1[6] ;
 wire \am_sdr0.filt0.yn_1[7] ;
 wire \am_sdr0.filt0.yn_1[8] ;
 wire \am_sdr0.filt0.yn_1[9] ;
 wire \am_sdr0.filt0.yn_2[10] ;
 wire \am_sdr0.filt0.yn_2[11] ;
 wire \am_sdr0.filt0.yn_2[12] ;
 wire \am_sdr0.filt0.yn_2[13] ;
 wire \am_sdr0.filt0.yn_2[1] ;
 wire \am_sdr0.filt0.yn_2[2] ;
 wire \am_sdr0.filt0.yn_2[3] ;
 wire \am_sdr0.filt0.yn_2[4] ;
 wire \am_sdr0.filt0.yn_2[5] ;
 wire \am_sdr0.filt0.yn_2[6] ;
 wire \am_sdr0.filt0.yn_2[7] ;
 wire \am_sdr0.filt0.yn_2[8] ;
 wire \am_sdr0.filt0.yn_2[9] ;
 wire \am_sdr0.nco0.nco_phase[0] ;
 wire \am_sdr0.nco0.nco_phase[10] ;
 wire \am_sdr0.nco0.nco_phase[11] ;
 wire \am_sdr0.nco0.nco_phase[12] ;
 wire \am_sdr0.nco0.nco_phase[13] ;
 wire \am_sdr0.nco0.nco_phase[14] ;
 wire \am_sdr0.nco0.nco_phase[15] ;
 wire \am_sdr0.nco0.nco_phase[16] ;
 wire \am_sdr0.nco0.nco_phase[17] ;
 wire \am_sdr0.nco0.nco_phase[18] ;
 wire \am_sdr0.nco0.nco_phase[19] ;
 wire \am_sdr0.nco0.nco_phase[1] ;
 wire \am_sdr0.nco0.nco_phase[2] ;
 wire \am_sdr0.nco0.nco_phase[3] ;
 wire \am_sdr0.nco0.nco_phase[4] ;
 wire \am_sdr0.nco0.nco_phase[5] ;
 wire \am_sdr0.nco0.nco_phase[6] ;
 wire \am_sdr0.nco0.nco_phase[7] ;
 wire \am_sdr0.nco0.nco_phase[8] ;
 wire \am_sdr0.nco0.nco_phase[9] ;
 wire \am_sdr0.nco0.phase_inc[0] ;
 wire \am_sdr0.nco0.phase_inc[10] ;
 wire \am_sdr0.nco0.phase_inc[11] ;
 wire \am_sdr0.nco0.phase_inc[12] ;
 wire \am_sdr0.nco0.phase_inc[13] ;
 wire \am_sdr0.nco0.phase_inc[14] ;
 wire \am_sdr0.nco0.phase_inc[15] ;
 wire \am_sdr0.nco0.phase_inc[16] ;
 wire \am_sdr0.nco0.phase_inc[17] ;
 wire \am_sdr0.nco0.phase_inc[18] ;
 wire \am_sdr0.nco0.phase_inc[19] ;
 wire \am_sdr0.nco0.phase_inc[1] ;
 wire \am_sdr0.nco0.phase_inc[2] ;
 wire \am_sdr0.nco0.phase_inc[3] ;
 wire \am_sdr0.nco0.phase_inc[4] ;
 wire \am_sdr0.nco0.phase_inc[5] ;
 wire \am_sdr0.nco0.phase_inc[6] ;
 wire \am_sdr0.nco0.phase_inc[7] ;
 wire \am_sdr0.nco0.phase_inc[8] ;
 wire \am_sdr0.nco0.phase_inc[9] ;
 wire \am_sdr0.nco0.rf_a ;
 wire \am_sdr0.spi0.CS_q ;
 wire \am_sdr0.spi0.CS_qq ;
 wire \am_sdr0.spi0.CS_qqq ;
 wire \am_sdr0.spi0.MOSI_q ;
 wire \am_sdr0.spi0.MOSI_qq ;
 wire \am_sdr0.spi0.SCK_q ;
 wire \am_sdr0.spi0.SCK_qq ;
 wire \am_sdr0.spi0.SCK_qqq ;
 wire \am_sdr0.spi0.state[0] ;
 wire \am_sdr0.spi0.state[1] ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;

 sg13g2_inv_1 _3030_ (.Y(_2127_),
    .A(net246));
 sg13g2_inv_1 _3031_ (.Y(_2128_),
    .A(net251));
 sg13g2_inv_1 _3032_ (.Y(_2129_),
    .A(net261));
 sg13g2_inv_1 _3033_ (.Y(_2130_),
    .A(\am_sdr0.nco0.phase_inc[17] ));
 sg13g2_inv_1 _3034_ (.Y(_2131_),
    .A(\am_sdr0.nco0.phase_inc[16] ));
 sg13g2_inv_1 _3035_ (.Y(_2132_),
    .A(net257));
 sg13g2_inv_1 _3036_ (.Y(_2133_),
    .A(net245));
 sg13g2_inv_1 _3037_ (.Y(_2134_),
    .A(net270));
 sg13g2_inv_1 _3038_ (.Y(_2135_),
    .A(\am_sdr0.nco0.phase_inc[6] ));
 sg13g2_inv_1 _3039_ (.Y(_2136_),
    .A(net232));
 sg13g2_inv_1 _3040_ (.Y(_2137_),
    .A(net271));
 sg13g2_inv_1 _3041_ (.Y(_2138_),
    .A(net273));
 sg13g2_inv_1 _3042_ (.Y(_2139_),
    .A(\am_sdr0.nco0.phase_inc[2] ));
 sg13g2_inv_1 _3043_ (.Y(_2140_),
    .A(\am_sdr0.nco0.phase_inc[1] ));
 sg13g2_inv_1 _3044_ (.Y(_2141_),
    .A(\am_sdr0.nco0.phase_inc[0] ));
 sg13g2_inv_1 _3045_ (.Y(_2142_),
    .A(net231));
 sg13g2_inv_1 _3046_ (.Y(_2143_),
    .A(\am_sdr0.nco0.nco_phase[15] ));
 sg13g2_inv_1 _3047_ (.Y(_2144_),
    .A(net417));
 sg13g2_inv_2 _3048_ (.Y(_2145_),
    .A(net282));
 sg13g2_inv_1 _3049_ (.Y(_2146_),
    .A(net272));
 sg13g2_inv_2 _3050_ (.Y(_2147_),
    .A(net374));
 sg13g2_inv_1 _3051_ (.Y(_2148_),
    .A(net367));
 sg13g2_inv_1 _3052_ (.Y(_2149_),
    .A(net365));
 sg13g2_inv_2 _3053_ (.Y(_2150_),
    .A(net360));
 sg13g2_inv_1 _3054_ (.Y(_2151_),
    .A(net358));
 sg13g2_inv_1 _3055_ (.Y(_2152_),
    .A(net378));
 sg13g2_inv_2 _3056_ (.Y(_2153_),
    .A(net354));
 sg13g2_inv_2 _3057_ (.Y(_2154_),
    .A(net352));
 sg13g2_inv_1 _3058_ (.Y(_2155_),
    .A(net264));
 sg13g2_inv_1 _3059_ (.Y(_2156_),
    .A(\am_sdr0.filt0.xn_2[5] ));
 sg13g2_inv_2 _3060_ (.Y(_2157_),
    .A(\am_sdr0.filt0.mul_b2[0] ));
 sg13g2_inv_1 _3061_ (.Y(_2158_),
    .A(_0016_));
 sg13g2_inv_1 _3062_ (.Y(_2159_),
    .A(_0018_));
 sg13g2_inv_1 _3063_ (.Y(_2160_),
    .A(net346));
 sg13g2_inv_1 _3064_ (.Y(_2161_),
    .A(COMP_OUT));
 sg13g2_inv_1 _3065_ (.Y(_2162_),
    .A(net220));
 sg13g2_inv_1 _3066_ (.Y(_2163_),
    .A(net214));
 sg13g2_inv_1 _3067_ (.Y(_2164_),
    .A(net253));
 sg13g2_inv_1 _3068_ (.Y(_2165_),
    .A(net216));
 sg13g2_inv_1 _3069_ (.Y(_2166_),
    .A(net256));
 sg13g2_inv_1 _3070_ (.Y(_2167_),
    .A(\am_sdr0.count[5] ));
 sg13g2_inv_1 _3071_ (.Y(_2168_),
    .A(net265));
 sg13g2_inv_1 _3072_ (.Y(_2169_),
    .A(net283));
 sg13g2_inv_1 _3073_ (.Y(_2170_),
    .A(net223));
 sg13g2_inv_1 _3074_ (.Y(_2171_),
    .A(\am_sdr0.count[2] ));
 sg13g2_inv_1 _3075_ (.Y(_2172_),
    .A(\am_sdr0.det0.env_out[1] ));
 sg13g2_inv_1 _3076_ (.Y(_2173_),
    .A(net287));
 sg13g2_inv_1 _3077_ (.Y(_2174_),
    .A(\am_sdr0.det0.alpha_yn_1[0] ));
 sg13g2_inv_1 _3078_ (.Y(_2175_),
    .A(\am_sdr0.det0.yn_1[10] ));
 sg13g2_nand2_1 _3079_ (.Y(_2176_),
    .A(\am_sdr0.nco0.phase_inc[16] ),
    .B(\am_sdr0.nco0.nco_phase[16] ));
 sg13g2_xnor2_1 _3080_ (.Y(_2177_),
    .A(\am_sdr0.nco0.phase_inc[16] ),
    .B(\am_sdr0.nco0.nco_phase[16] ));
 sg13g2_nand2_1 _3081_ (.Y(_2178_),
    .A(net281),
    .B(\am_sdr0.nco0.nco_phase[14] ));
 sg13g2_nor2_1 _3082_ (.A(\am_sdr0.nco0.phase_inc[14] ),
    .B(\am_sdr0.nco0.nco_phase[14] ),
    .Y(_2179_));
 sg13g2_xor2_1 _3083_ (.B(net435),
    .A(\am_sdr0.nco0.phase_inc[14] ),
    .X(_2180_));
 sg13g2_nor2_1 _3084_ (.A(\am_sdr0.nco0.phase_inc[13] ),
    .B(\am_sdr0.nco0.nco_phase[13] ),
    .Y(_2181_));
 sg13g2_and2_1 _3085_ (.A(net241),
    .B(\am_sdr0.nco0.nco_phase[12] ),
    .X(_2182_));
 sg13g2_xor2_1 _3086_ (.B(net312),
    .A(net241),
    .X(_2183_));
 sg13g2_nor2_1 _3087_ (.A(net245),
    .B(net316),
    .Y(_2184_));
 sg13g2_nand2_1 _3088_ (.Y(_2185_),
    .A(net245),
    .B(net316));
 sg13g2_xnor2_1 _3089_ (.Y(_2186_),
    .A(net270),
    .B(net314));
 sg13g2_nand2_1 _3090_ (.Y(_2187_),
    .A(net276),
    .B(net300));
 sg13g2_nand2_1 _3091_ (.Y(_2188_),
    .A(net268),
    .B(net304));
 sg13g2_nand2_1 _3092_ (.Y(_2189_),
    .A(net236),
    .B(net322));
 sg13g2_nand2_1 _3093_ (.Y(_2190_),
    .A(net232),
    .B(net429));
 sg13g2_nand2_1 _3094_ (.Y(_2191_),
    .A(net271),
    .B(net318));
 sg13g2_nand2_1 _3095_ (.Y(_2192_),
    .A(net273),
    .B(net323));
 sg13g2_nand2_1 _3096_ (.Y(_2193_),
    .A(net280),
    .B(net432));
 sg13g2_nand2_1 _3097_ (.Y(_2194_),
    .A(net278),
    .B(net325));
 sg13g2_and2_1 _3098_ (.A(net243),
    .B(net228),
    .X(_2195_));
 sg13g2_xor2_1 _3099_ (.B(net325),
    .A(\am_sdr0.nco0.phase_inc[1] ),
    .X(_2196_));
 sg13g2_nand2_1 _3100_ (.Y(_2197_),
    .A(_2195_),
    .B(_2196_));
 sg13g2_xnor2_1 _3101_ (.Y(_2198_),
    .A(\am_sdr0.nco0.phase_inc[2] ),
    .B(net433));
 sg13g2_a21o_1 _3102_ (.A2(_2197_),
    .A1(_2194_),
    .B1(_2198_),
    .X(_2199_));
 sg13g2_xnor2_1 _3103_ (.Y(_2200_),
    .A(\am_sdr0.nco0.phase_inc[3] ),
    .B(net323));
 sg13g2_a21o_1 _3104_ (.A2(_2199_),
    .A1(_2193_),
    .B1(_2200_),
    .X(_2201_));
 sg13g2_xnor2_1 _3105_ (.Y(_2202_),
    .A(\am_sdr0.nco0.phase_inc[4] ),
    .B(net318));
 sg13g2_a21o_1 _3106_ (.A2(_2201_),
    .A1(_2192_),
    .B1(_2202_),
    .X(_2203_));
 sg13g2_xnor2_1 _3107_ (.Y(_2204_),
    .A(\am_sdr0.nco0.phase_inc[5] ),
    .B(\am_sdr0.nco0.nco_phase[5] ));
 sg13g2_a21o_1 _3108_ (.A2(_2203_),
    .A1(_2191_),
    .B1(_2204_),
    .X(_2205_));
 sg13g2_xnor2_1 _3109_ (.Y(_2206_),
    .A(\am_sdr0.nco0.phase_inc[6] ),
    .B(net322));
 sg13g2_a21o_1 _3110_ (.A2(_2205_),
    .A1(_2190_),
    .B1(_2206_),
    .X(_2207_));
 sg13g2_xnor2_1 _3111_ (.Y(_2208_),
    .A(\am_sdr0.nco0.phase_inc[7] ),
    .B(net304));
 sg13g2_a21o_1 _3112_ (.A2(_2207_),
    .A1(_2189_),
    .B1(_2208_),
    .X(_2209_));
 sg13g2_xnor2_1 _3113_ (.Y(_2210_),
    .A(net249),
    .B(\am_sdr0.nco0.nco_phase[8] ));
 sg13g2_a21oi_1 _3114_ (.A1(_2188_),
    .A2(_2209_),
    .Y(_2211_),
    .B1(_2210_));
 sg13g2_a21o_1 _3115_ (.A2(\am_sdr0.nco0.nco_phase[8] ),
    .A1(net249),
    .B1(_2211_),
    .X(_2212_));
 sg13g2_o21ai_1 _3116_ (.B1(_2212_),
    .Y(_2213_),
    .A1(\am_sdr0.nco0.phase_inc[9] ),
    .A2(net300));
 sg13g2_a21oi_1 _3117_ (.A1(_2187_),
    .A2(_2213_),
    .Y(_2214_),
    .B1(_2186_));
 sg13g2_a21oi_1 _3118_ (.A1(net270),
    .A2(net314),
    .Y(_2215_),
    .B1(_2214_));
 sg13g2_o21ai_1 _3119_ (.B1(_2185_),
    .Y(_2216_),
    .A1(_2184_),
    .A2(_2215_));
 sg13g2_a21o_1 _3120_ (.A2(_2216_),
    .A1(_2183_),
    .B1(_2182_),
    .X(_2217_));
 sg13g2_a21oi_1 _3121_ (.A1(\am_sdr0.nco0.phase_inc[13] ),
    .A2(\am_sdr0.nco0.nco_phase[13] ),
    .Y(_2218_),
    .B1(_2217_));
 sg13g2_or2_1 _3122_ (.X(_2219_),
    .B(_2218_),
    .A(_2181_));
 sg13g2_o21ai_1 _3123_ (.B1(_2178_),
    .Y(_2220_),
    .A1(_2179_),
    .A2(_2219_));
 sg13g2_a21oi_1 _3124_ (.A1(\am_sdr0.nco0.phase_inc[15] ),
    .A2(\am_sdr0.nco0.nco_phase[15] ),
    .Y(_2221_),
    .B1(_2220_));
 sg13g2_a21oi_1 _3125_ (.A1(_2132_),
    .A2(_2143_),
    .Y(_2222_),
    .B1(_2221_));
 sg13g2_nand2b_1 _3126_ (.Y(_2223_),
    .B(_2222_),
    .A_N(_2177_));
 sg13g2_xnor2_1 _3127_ (.Y(_2224_),
    .A(\am_sdr0.nco0.phase_inc[17] ),
    .B(\am_sdr0.nco0.nco_phase[17] ));
 sg13g2_a21oi_1 _3128_ (.A1(_2176_),
    .A2(_2223_),
    .Y(_2225_),
    .B1(_2224_));
 sg13g2_a21oi_1 _3129_ (.A1(\am_sdr0.nco0.phase_inc[17] ),
    .A2(\am_sdr0.nco0.nco_phase[17] ),
    .Y(_2226_),
    .B1(_2225_));
 sg13g2_nand2_1 _3130_ (.Y(_2227_),
    .A(\am_sdr0.nco0.phase_inc[18] ),
    .B(\am_sdr0.nco0.nco_phase[18] ));
 sg13g2_xnor2_1 _3131_ (.Y(_2228_),
    .A(\am_sdr0.nco0.phase_inc[18] ),
    .B(\am_sdr0.nco0.nco_phase[18] ));
 sg13g2_or2_1 _3132_ (.X(_2229_),
    .B(_2228_),
    .A(_2226_));
 sg13g2_a21oi_1 _3133_ (.A1(_2226_),
    .A2(_2228_),
    .Y(_2230_),
    .B1(net409));
 sg13g2_nand2_2 _3134_ (.Y(_2231_),
    .A(_2229_),
    .B(_2230_));
 sg13g2_inv_1 _3135_ (.Y(_0178_),
    .A(_2231_));
 sg13g2_nand3_1 _3136_ (.B(_2223_),
    .C(_2224_),
    .A(_2176_),
    .Y(_2232_));
 sg13g2_nor2b_1 _3137_ (.A(_2225_),
    .B_N(_2232_),
    .Y(_2233_));
 sg13g2_nand2_1 _3138_ (.Y(_2234_),
    .A(net425),
    .B(_2233_));
 sg13g2_inv_1 _3139_ (.Y(_0177_),
    .A(_2234_));
 sg13g2_nor2_1 _3140_ (.A(_2231_),
    .B(_2234_),
    .Y(_2235_));
 sg13g2_xnor2_1 _3141_ (.Y(_2236_),
    .A(_2177_),
    .B(_2222_));
 sg13g2_nand2_2 _3142_ (.Y(_2237_),
    .A(net425),
    .B(_2236_));
 sg13g2_inv_1 _3143_ (.Y(_0176_),
    .A(_2237_));
 sg13g2_nand2_1 _3144_ (.Y(_2238_),
    .A(_0177_),
    .B(_0176_));
 sg13g2_a21o_1 _3145_ (.A2(_2238_),
    .A1(_2231_),
    .B1(_2235_),
    .X(_0000_));
 sg13g2_nor2_2 _3146_ (.A(_0177_),
    .B(_0176_),
    .Y(_2239_));
 sg13g2_a21oi_1 _3147_ (.A1(_2231_),
    .A2(_2239_),
    .Y(_2240_),
    .B1(_2235_));
 sg13g2_xnor2_1 _3148_ (.Y(_2241_),
    .A(\am_sdr0.nco0.phase_inc[19] ),
    .B(\am_sdr0.nco0.nco_phase[19] ));
 sg13g2_nand3_1 _3149_ (.B(_2229_),
    .C(_2241_),
    .A(_2227_),
    .Y(_2242_));
 sg13g2_a21o_1 _3150_ (.A2(_2229_),
    .A1(_2227_),
    .B1(_2241_),
    .X(_2243_));
 sg13g2_nand3_1 _3151_ (.B(_2242_),
    .C(_2243_),
    .A(net425),
    .Y(_2244_));
 sg13g2_inv_2 _3152_ (.Y(_0179_),
    .A(_2244_));
 sg13g2_and2_1 _3153_ (.A(_0000_),
    .B(_0179_),
    .X(_2245_));
 sg13g2_nand2_1 _3154_ (.Y(_2246_),
    .A(_2240_),
    .B(_2245_));
 sg13g2_o21ai_1 _3155_ (.B1(_2246_),
    .Y(_0001_),
    .A1(_2240_),
    .A2(_0179_));
 sg13g2_nand2_1 _3156_ (.Y(_2247_),
    .A(_0177_),
    .B(_2237_));
 sg13g2_xnor2_1 _3157_ (.Y(_2248_),
    .A(_0178_),
    .B(_2244_));
 sg13g2_xor2_1 _3158_ (.B(_2248_),
    .A(_2247_),
    .X(_2249_));
 sg13g2_and2_1 _3159_ (.A(_0000_),
    .B(_2249_),
    .X(_0002_));
 sg13g2_nand2_1 _3160_ (.Y(_2250_),
    .A(_2231_),
    .B(_2237_));
 sg13g2_o21ai_1 _3161_ (.B1(_2250_),
    .Y(_2251_),
    .A1(_2231_),
    .A2(_2238_));
 sg13g2_nor2_1 _3162_ (.A(_2245_),
    .B(_2251_),
    .Y(_2252_));
 sg13g2_a21oi_1 _3163_ (.A1(_0179_),
    .A2(_2251_),
    .Y(_0003_),
    .B1(_2252_));
 sg13g2_nor2_1 _3164_ (.A(_0177_),
    .B(_2237_),
    .Y(_2253_));
 sg13g2_nor2_1 _3165_ (.A(_2231_),
    .B(_2253_),
    .Y(_2254_));
 sg13g2_nand2_1 _3166_ (.Y(_2255_),
    .A(_2235_),
    .B(_0179_));
 sg13g2_o21ai_1 _3167_ (.B1(_2255_),
    .Y(_0004_),
    .A1(_2245_),
    .A2(_2254_));
 sg13g2_nand2_1 _3168_ (.Y(_2256_),
    .A(_2239_),
    .B(_0179_));
 sg13g2_and2_1 _3169_ (.A(_2249_),
    .B(_2256_),
    .X(_0005_));
 sg13g2_a21oi_1 _3170_ (.A1(_2231_),
    .A2(_2237_),
    .Y(_2257_),
    .B1(_2253_));
 sg13g2_nand3_1 _3171_ (.B(_0179_),
    .C(_2257_),
    .A(_2233_),
    .Y(_2258_));
 sg13g2_o21ai_1 _3172_ (.B1(_2258_),
    .Y(_0006_),
    .A1(_0179_),
    .A2(_2257_));
 sg13g2_nand2_1 _3173_ (.Y(_2259_),
    .A(_0178_),
    .B(_2239_));
 sg13g2_and2_1 _3174_ (.A(_2248_),
    .B(_2259_),
    .X(_0007_));
 sg13g2_nand2_1 _3175_ (.Y(_2260_),
    .A(net188),
    .B(COMP_OUT));
 sg13g2_xnor2_1 _3176_ (.Y(_0008_),
    .A(net239),
    .B(_2260_));
 sg13g2_nor2_1 _3177_ (.A(net188),
    .B(_0032_),
    .Y(_2261_));
 sg13g2_a21oi_1 _3178_ (.A1(_0020_),
    .A2(_2261_),
    .Y(_2262_),
    .B1(_2161_));
 sg13g2_o21ai_1 _3179_ (.B1(_2262_),
    .Y(_2263_),
    .A1(_0020_),
    .A2(_2261_));
 sg13g2_o21ai_1 _3180_ (.B1(_2263_),
    .Y(_0009_),
    .A1(COMP_OUT),
    .A2(_2162_));
 sg13g2_xor2_1 _3181_ (.B(_2262_),
    .A(net212),
    .X(_0010_));
 sg13g2_nor4_2 _3182_ (.A(net188),
    .B(_0032_),
    .C(_0033_),
    .Y(_2264_),
    .D(net212));
 sg13g2_inv_1 _3183_ (.Y(_2265_),
    .A(_2264_));
 sg13g2_a21oi_1 _3184_ (.A1(_0021_),
    .A2(_2264_),
    .Y(_2266_),
    .B1(_2161_));
 sg13g2_o21ai_1 _3185_ (.B1(_2266_),
    .Y(_2267_),
    .A1(_0021_),
    .A2(_2264_));
 sg13g2_o21ai_1 _3186_ (.B1(_2267_),
    .Y(_0011_),
    .A1(COMP_OUT),
    .A2(_2163_));
 sg13g2_xor2_1 _3187_ (.B(_2266_),
    .A(net206),
    .X(_0012_));
 sg13g2_nand2_1 _3188_ (.Y(_2268_),
    .A(_2161_),
    .B(net201));
 sg13g2_nor3_1 _3189_ (.A(_0035_),
    .B(_0036_),
    .C(_2265_),
    .Y(_2269_));
 sg13g2_a21o_1 _3190_ (.A2(_2269_),
    .A1(_0022_),
    .B1(_2161_),
    .X(_2270_));
 sg13g2_nor2_1 _3191_ (.A(_0022_),
    .B(_2269_),
    .Y(_2271_));
 sg13g2_o21ai_1 _3192_ (.B1(net202),
    .Y(_0013_),
    .A1(_2270_),
    .A2(_2271_));
 sg13g2_xnor2_1 _3193_ (.Y(_0014_),
    .A(net204),
    .B(_2270_));
 sg13g2_nor4_2 _3194_ (.A(\am_sdr0.spi0.state[1] ),
    .B(net293),
    .C(_2142_),
    .Y(_2272_),
    .D(net222));
 sg13g2_nor2b_2 _3195_ (.A(\am_sdr0.spi0.state[1] ),
    .B_N(\am_sdr0.spi0.state[0] ),
    .Y(_2273_));
 sg13g2_nand3b_1 _3196_ (.B(net343),
    .C(\am_sdr0.spi0.SCK_qq ),
    .Y(_2274_),
    .A_N(\am_sdr0.spi0.SCK_qqq ));
 sg13g2_nor2b_1 _3197_ (.A(_2272_),
    .B_N(_2274_),
    .Y(_2275_));
 sg13g2_nand2b_2 _3198_ (.Y(_2276_),
    .B(_2274_),
    .A_N(_2272_));
 sg13g2_nand2_1 _3199_ (.Y(_2277_),
    .A(net420),
    .B(net335));
 sg13g2_and2_1 _3200_ (.A(net421),
    .B(_2273_),
    .X(_2278_));
 sg13g2_nand2_1 _3201_ (.Y(_2279_),
    .A(net209),
    .B(_2278_));
 sg13g2_a22oi_1 _3202_ (.Y(_0040_),
    .B1(net332),
    .B2(net210),
    .A2(net336),
    .A1(_2141_));
 sg13g2_nand2_1 _3203_ (.Y(_2280_),
    .A(net243),
    .B(net339));
 sg13g2_a22oi_1 _3204_ (.Y(_0041_),
    .B1(net331),
    .B2(_2280_),
    .A2(net336),
    .A1(_2140_));
 sg13g2_nand2_1 _3205_ (.Y(_2281_),
    .A(net278),
    .B(net338));
 sg13g2_a22oi_1 _3206_ (.Y(_0042_),
    .B1(net332),
    .B2(_2281_),
    .A2(net336),
    .A1(_2139_));
 sg13g2_nand2_1 _3207_ (.Y(_2282_),
    .A(net280),
    .B(net338));
 sg13g2_a22oi_1 _3208_ (.Y(_0043_),
    .B1(net331),
    .B2(_2282_),
    .A2(net335),
    .A1(_2138_));
 sg13g2_nand2_1 _3209_ (.Y(_2283_),
    .A(net273),
    .B(net338));
 sg13g2_a22oi_1 _3210_ (.Y(_0044_),
    .B1(net331),
    .B2(_2283_),
    .A2(net335),
    .A1(_2137_));
 sg13g2_nand2_1 _3211_ (.Y(_2284_),
    .A(net271),
    .B(net338));
 sg13g2_a22oi_1 _3212_ (.Y(_0045_),
    .B1(net331),
    .B2(_2284_),
    .A2(net335),
    .A1(_2136_));
 sg13g2_nand2_1 _3213_ (.Y(_2285_),
    .A(net232),
    .B(net338));
 sg13g2_a22oi_1 _3214_ (.Y(_0046_),
    .B1(net331),
    .B2(_2285_),
    .A2(net335),
    .A1(_2135_));
 sg13g2_nand3_1 _3215_ (.B(net343),
    .C(_2276_),
    .A(net236),
    .Y(_2286_));
 sg13g2_a21oi_1 _3216_ (.A1(\am_sdr0.nco0.phase_inc[7] ),
    .A2(net335),
    .Y(_2287_),
    .B1(net408));
 sg13g2_nand2_1 _3217_ (.Y(_0047_),
    .A(_2286_),
    .B(_2287_));
 sg13g2_nand3_1 _3218_ (.B(_2273_),
    .C(_2276_),
    .A(net268),
    .Y(_2288_));
 sg13g2_a21oi_1 _3219_ (.A1(net249),
    .A2(net335),
    .Y(_2289_),
    .B1(net408));
 sg13g2_nand2_1 _3220_ (.Y(_0048_),
    .A(net269),
    .B(_2289_));
 sg13g2_nand3_1 _3221_ (.B(net343),
    .C(_2276_),
    .A(net249),
    .Y(_2290_));
 sg13g2_a21oi_1 _3222_ (.A1(\am_sdr0.nco0.phase_inc[9] ),
    .A2(net334),
    .Y(_2291_),
    .B1(net407));
 sg13g2_nand2_1 _3223_ (.Y(_0049_),
    .A(_2290_),
    .B(_2291_));
 sg13g2_nand2_1 _3224_ (.Y(_2292_),
    .A(net276),
    .B(net339));
 sg13g2_a22oi_1 _3225_ (.Y(_0050_),
    .B1(net332),
    .B2(_2292_),
    .A2(net334),
    .A1(_2134_));
 sg13g2_nand2_1 _3226_ (.Y(_2293_),
    .A(net270),
    .B(net339));
 sg13g2_a22oi_1 _3227_ (.Y(_0051_),
    .B1(net332),
    .B2(_2293_),
    .A2(net334),
    .A1(_2133_));
 sg13g2_nand3_1 _3228_ (.B(net343),
    .C(_2276_),
    .A(net245),
    .Y(_2294_));
 sg13g2_a21oi_1 _3229_ (.A1(net241),
    .A2(net334),
    .Y(_2295_),
    .B1(net409));
 sg13g2_nand2_1 _3230_ (.Y(_0052_),
    .A(_2294_),
    .B(_2295_));
 sg13g2_nand3_1 _3231_ (.B(net343),
    .C(_2276_),
    .A(net241),
    .Y(_2296_));
 sg13g2_a21oi_1 _3232_ (.A1(\am_sdr0.nco0.phase_inc[13] ),
    .A2(net337),
    .Y(_2297_),
    .B1(net409));
 sg13g2_nand2_1 _3233_ (.Y(_0053_),
    .A(_2296_),
    .B(_2297_));
 sg13g2_nand3_1 _3234_ (.B(net343),
    .C(_2276_),
    .A(net274),
    .Y(_2298_));
 sg13g2_a21oi_1 _3235_ (.A1(\am_sdr0.nco0.phase_inc[14] ),
    .A2(net337),
    .Y(_2299_),
    .B1(net409));
 sg13g2_nand2_1 _3236_ (.Y(_0054_),
    .A(_2298_),
    .B(_2299_));
 sg13g2_nand2_1 _3237_ (.Y(_2300_),
    .A(net281),
    .B(net339));
 sg13g2_a22oi_1 _3238_ (.Y(_0055_),
    .B1(net331),
    .B2(_2300_),
    .A2(net336),
    .A1(_2132_));
 sg13g2_nand2_1 _3239_ (.Y(_2301_),
    .A(net257),
    .B(net338));
 sg13g2_a22oi_1 _3240_ (.Y(_0056_),
    .B1(net331),
    .B2(_2301_),
    .A2(net336),
    .A1(_2131_));
 sg13g2_nand2_1 _3241_ (.Y(_2302_),
    .A(net259),
    .B(net338));
 sg13g2_a22oi_1 _3242_ (.Y(_0057_),
    .B1(net331),
    .B2(_2302_),
    .A2(net335),
    .A1(_2130_));
 sg13g2_nand2_1 _3243_ (.Y(_2303_),
    .A(net277),
    .B(net339));
 sg13g2_a22oi_1 _3244_ (.Y(_0058_),
    .B1(net332),
    .B2(_2303_),
    .A2(net337),
    .A1(_2129_));
 sg13g2_nand2_1 _3245_ (.Y(_2304_),
    .A(net261),
    .B(net339));
 sg13g2_a22oi_1 _3246_ (.Y(_0059_),
    .B1(net332),
    .B2(_2304_),
    .A2(net334),
    .A1(_2128_));
 sg13g2_nand3_1 _3247_ (.B(net343),
    .C(_2276_),
    .A(net251),
    .Y(_2305_));
 sg13g2_a21oi_1 _3248_ (.A1(\am_sdr0.filt0.gain_spi[0] ),
    .A2(net334),
    .Y(_2306_),
    .B1(net409));
 sg13g2_nand2_1 _3249_ (.Y(_0060_),
    .A(_2305_),
    .B(_2306_));
 sg13g2_nand3_1 _3250_ (.B(net343),
    .C(_2276_),
    .A(net290),
    .Y(_2307_));
 sg13g2_a21oi_1 _3251_ (.A1(\am_sdr0.filt0.gain_spi[1] ),
    .A2(net334),
    .Y(_2308_),
    .B1(net408));
 sg13g2_nand2_1 _3252_ (.Y(_0061_),
    .A(_2307_),
    .B(_2308_));
 sg13g2_nand2_1 _3253_ (.Y(_2309_),
    .A(\am_sdr0.filt0.gain_spi[1] ),
    .B(net339));
 sg13g2_a22oi_1 _3254_ (.Y(_0062_),
    .B1(net332),
    .B2(_2309_),
    .A2(net334),
    .A1(_2127_));
 sg13g2_nand2_1 _3255_ (.Y(_2310_),
    .A(_2142_),
    .B(net222));
 sg13g2_a22oi_1 _3256_ (.Y(_2311_),
    .B1(_2278_),
    .B2(_2310_),
    .A2(net294),
    .A1(net425));
 sg13g2_inv_1 _3257_ (.Y(_0063_),
    .A(net295));
 sg13g2_and3_1 _3258_ (.X(_0064_),
    .A(_2142_),
    .B(net222),
    .C(net338));
 sg13g2_and2_1 _3259_ (.A(net422),
    .B(net191),
    .X(_0065_));
 sg13g2_and2_1 _3260_ (.A(net422),
    .B(net4),
    .X(_0066_));
 sg13g2_and2_1 _3261_ (.A(net425),
    .B(net194),
    .X(_0067_));
 sg13g2_and2_1 _3262_ (.A(net222),
    .B(net425),
    .X(_0068_));
 sg13g2_and2_1 _3263_ (.A(net422),
    .B(net3),
    .X(_0069_));
 sg13g2_nor2_1 _3264_ (.A(_2172_),
    .B(\am_sdr0.count[1] ),
    .Y(_2312_));
 sg13g2_nor2b_1 _3265_ (.A(\am_sdr0.count[0] ),
    .B_N(\am_sdr0.det0.env_out[0] ),
    .Y(_2313_));
 sg13g2_a22oi_1 _3266_ (.Y(_2314_),
    .B1(_2172_),
    .B2(\am_sdr0.count[1] ),
    .A2(\am_sdr0.count[2] ),
    .A1(_2170_));
 sg13g2_o21ai_1 _3267_ (.B1(_2314_),
    .Y(_2315_),
    .A1(_2312_),
    .A2(_2313_));
 sg13g2_a22oi_1 _3268_ (.Y(_2316_),
    .B1(\am_sdr0.det0.env_out[2] ),
    .B2(_2171_),
    .A2(_2169_),
    .A1(\am_sdr0.det0.env_out[3] ));
 sg13g2_nand2b_1 _3269_ (.Y(_2317_),
    .B(\am_sdr0.count[3] ),
    .A_N(\am_sdr0.det0.env_out[3] ));
 sg13g2_o21ai_1 _3270_ (.B1(_2317_),
    .Y(_2318_),
    .A1(_2168_),
    .A2(\am_sdr0.det0.env_out[4] ));
 sg13g2_a21oi_1 _3271_ (.A1(_2315_),
    .A2(_2316_),
    .Y(_2319_),
    .B1(_2318_));
 sg13g2_a221oi_1 _3272_ (.B2(net255),
    .C1(_2319_),
    .B1(_2168_),
    .A1(net256),
    .Y(_2320_),
    .A2(_2167_));
 sg13g2_a21oi_1 _3273_ (.A1(_2166_),
    .A2(net263),
    .Y(_2321_),
    .B1(_2320_));
 sg13g2_o21ai_1 _3274_ (.B1(_2321_),
    .Y(_2322_),
    .A1(net248),
    .A2(_2165_));
 sg13g2_a22oi_1 _3275_ (.Y(_2323_),
    .B1(net248),
    .B2(_2165_),
    .A2(_2164_),
    .A1(net262));
 sg13g2_o21ai_1 _3276_ (.B1(net421),
    .Y(_2324_),
    .A1(net262),
    .A2(_2164_));
 sg13g2_a21oi_1 _3277_ (.A1(_2322_),
    .A2(_2323_),
    .Y(_0070_),
    .B1(_2324_));
 sg13g2_and2_1 _3278_ (.A(net422),
    .B(net192),
    .X(_0071_));
 sg13g2_and2_1 _3279_ (.A(net417),
    .B(net187),
    .X(_0072_));
 sg13g2_o21ai_1 _3280_ (.B1(net417),
    .Y(_2325_),
    .A1(\am_sdr0.count[1] ),
    .A2(net224));
 sg13g2_a21oi_1 _3281_ (.A1(\am_sdr0.count[1] ),
    .A2(net224),
    .Y(_0073_),
    .B1(_2325_));
 sg13g2_a21oi_1 _3282_ (.A1(\am_sdr0.count[1] ),
    .A2(net224),
    .Y(_2326_),
    .B1(net226));
 sg13g2_nand3_1 _3283_ (.B(\am_sdr0.count[1] ),
    .C(net224),
    .A(net226),
    .Y(_2327_));
 sg13g2_nand2_1 _3284_ (.Y(_2328_),
    .A(net418),
    .B(_2327_));
 sg13g2_nor2_1 _3285_ (.A(net227),
    .B(_2328_),
    .Y(_0074_));
 sg13g2_and2_1 _3286_ (.A(_2169_),
    .B(_2327_),
    .X(_2329_));
 sg13g2_nor2_1 _3287_ (.A(_2169_),
    .B(_2327_),
    .Y(_2330_));
 sg13g2_nor3_1 _3288_ (.A(net407),
    .B(_2329_),
    .C(_2330_),
    .Y(_0075_));
 sg13g2_nor3_2 _3289_ (.A(_2168_),
    .B(_2169_),
    .C(_2327_),
    .Y(_2331_));
 sg13g2_o21ai_1 _3290_ (.B1(net419),
    .Y(_2332_),
    .A1(net265),
    .A2(_2330_));
 sg13g2_nor2_1 _3291_ (.A(_2331_),
    .B(net266),
    .Y(_0076_));
 sg13g2_xnor2_1 _3292_ (.Y(_2333_),
    .A(net263),
    .B(_2331_));
 sg13g2_nor2_1 _3293_ (.A(net407),
    .B(_2333_),
    .Y(_0077_));
 sg13g2_a21oi_1 _3294_ (.A1(\am_sdr0.count[5] ),
    .A2(_2331_),
    .Y(_2334_),
    .B1(net216));
 sg13g2_nand3_1 _3295_ (.B(\am_sdr0.count[5] ),
    .C(_2331_),
    .A(net216),
    .Y(_2335_));
 sg13g2_nand2_1 _3296_ (.Y(_2336_),
    .A(net419),
    .B(_2335_));
 sg13g2_nor2_1 _3297_ (.A(net217),
    .B(_2336_),
    .Y(_0078_));
 sg13g2_o21ai_1 _3298_ (.B1(net419),
    .Y(_2337_),
    .A1(_2164_),
    .A2(_2335_));
 sg13g2_a21oi_1 _3299_ (.A1(_2164_),
    .A2(_2335_),
    .Y(_0079_),
    .B1(_2337_));
 sg13g2_nor2_2 _3300_ (.A(\am_sdr0.det0.ifreq[1] ),
    .B(\am_sdr0.det0.env_det[0] ),
    .Y(_2338_));
 sg13g2_nand2b_2 _3301_ (.Y(_2339_),
    .B(_2338_),
    .A_N(\am_sdr0.det0.ifreq[2] ));
 sg13g2_nor2_1 _3302_ (.A(\am_sdr0.det0.ifreq[3] ),
    .B(_2339_),
    .Y(_2340_));
 sg13g2_nor3_1 _3303_ (.A(\am_sdr0.det0.ifreq[4] ),
    .B(\am_sdr0.det0.ifreq[3] ),
    .C(_2339_),
    .Y(_2341_));
 sg13g2_nor2b_1 _3304_ (.A(\am_sdr0.det0.ifreq[5] ),
    .B_N(_2341_),
    .Y(_2342_));
 sg13g2_nand2b_1 _3305_ (.Y(_2343_),
    .B(_2342_),
    .A_N(\am_sdr0.det0.ifreq[6] ));
 sg13g2_a21oi_2 _3306_ (.B1(_0024_),
    .Y(_2344_),
    .A2(_2343_),
    .A1(\am_sdr0.det0.ifreq[7] ));
 sg13g2_and2_1 _3307_ (.A(\am_sdr0.det0.yn_1[3] ),
    .B(\am_sdr0.det0.yn_1[2] ),
    .X(_2345_));
 sg13g2_xor2_1 _3308_ (.B(\am_sdr0.det0.yn_1[2] ),
    .A(\am_sdr0.det0.yn_1[3] ),
    .X(_2346_));
 sg13g2_a21oi_2 _3309_ (.B1(_2345_),
    .Y(_2347_),
    .A2(_2346_),
    .A1(\am_sdr0.det0.yn_1[4] ));
 sg13g2_and2_1 _3310_ (.A(\am_sdr0.det0.yn_1[3] ),
    .B(\am_sdr0.det0.yn_1[4] ),
    .X(_2348_));
 sg13g2_xor2_1 _3311_ (.B(\am_sdr0.det0.yn_1[4] ),
    .A(\am_sdr0.det0.yn_1[3] ),
    .X(_2349_));
 sg13g2_xnor2_1 _3312_ (.Y(_2350_),
    .A(\am_sdr0.det0.yn_1[5] ),
    .B(_2349_));
 sg13g2_nor2_1 _3313_ (.A(_2347_),
    .B(_2350_),
    .Y(_2351_));
 sg13g2_xor2_1 _3314_ (.B(_2350_),
    .A(_2347_),
    .X(_2352_));
 sg13g2_and2_1 _3315_ (.A(net405),
    .B(\am_sdr0.det0.yn_1[7] ),
    .X(_2353_));
 sg13g2_xor2_1 _3316_ (.B(\am_sdr0.det0.yn_1[7] ),
    .A(\am_sdr0.det0.yn_1[6] ),
    .X(_2354_));
 sg13g2_xnor2_1 _3317_ (.Y(_2355_),
    .A(\am_sdr0.det0.yn_1[8] ),
    .B(_2354_));
 sg13g2_inv_1 _3318_ (.Y(_2356_),
    .A(_2355_));
 sg13g2_a21oi_2 _3319_ (.B1(_2351_),
    .Y(_2357_),
    .A2(_2356_),
    .A1(_2352_));
 sg13g2_a21oi_2 _3320_ (.B1(_2348_),
    .Y(_2358_),
    .A2(_2349_),
    .A1(\am_sdr0.det0.yn_1[5] ));
 sg13g2_and2_1 _3321_ (.A(\am_sdr0.det0.yn_1[4] ),
    .B(\am_sdr0.det0.yn_1[5] ),
    .X(_2359_));
 sg13g2_xor2_1 _3322_ (.B(\am_sdr0.det0.yn_1[5] ),
    .A(\am_sdr0.det0.yn_1[4] ),
    .X(_2360_));
 sg13g2_xnor2_1 _3323_ (.Y(_2361_),
    .A(net405),
    .B(_2360_));
 sg13g2_inv_1 _3324_ (.Y(_2362_),
    .A(_2361_));
 sg13g2_nor2_1 _3325_ (.A(_2358_),
    .B(_2361_),
    .Y(_2363_));
 sg13g2_xor2_1 _3326_ (.B(_2361_),
    .A(_2358_),
    .X(_2364_));
 sg13g2_and2_1 _3327_ (.A(net404),
    .B(\am_sdr0.det0.yn_1[8] ),
    .X(_2365_));
 sg13g2_xor2_1 _3328_ (.B(\am_sdr0.det0.yn_1[8] ),
    .A(net404),
    .X(_2366_));
 sg13g2_xnor2_1 _3329_ (.Y(_2367_),
    .A(\am_sdr0.det0.yn_1[9] ),
    .B(_2366_));
 sg13g2_inv_1 _3330_ (.Y(_2368_),
    .A(_2367_));
 sg13g2_xnor2_1 _3331_ (.Y(_2369_),
    .A(_2364_),
    .B(_2368_));
 sg13g2_nor2_1 _3332_ (.A(_2357_),
    .B(_2369_),
    .Y(_2370_));
 sg13g2_xor2_1 _3333_ (.B(_2369_),
    .A(_2357_),
    .X(_2371_));
 sg13g2_and2_1 _3334_ (.A(\am_sdr0.det0.yn_1[9] ),
    .B(\am_sdr0.det0.yn_1[10] ),
    .X(_2372_));
 sg13g2_xor2_1 _3335_ (.B(\am_sdr0.det0.yn_1[10] ),
    .A(\am_sdr0.det0.yn_1[9] ),
    .X(_2373_));
 sg13g2_a21oi_2 _3336_ (.B1(_2372_),
    .Y(_2374_),
    .A2(_2373_),
    .A1(\am_sdr0.det0.yn_1[11] ));
 sg13g2_inv_1 _3337_ (.Y(_2375_),
    .A(_2374_));
 sg13g2_a21oi_2 _3338_ (.B1(_2353_),
    .Y(_2376_),
    .A2(_2354_),
    .A1(\am_sdr0.det0.yn_1[8] ));
 sg13g2_and2_1 _3339_ (.A(\am_sdr0.det0.yn_1[10] ),
    .B(\am_sdr0.det0.yn_1[11] ),
    .X(_2377_));
 sg13g2_xor2_1 _3340_ (.B(\am_sdr0.det0.yn_1[11] ),
    .A(\am_sdr0.det0.yn_1[10] ),
    .X(_2378_));
 sg13g2_xnor2_1 _3341_ (.Y(_2379_),
    .A(\am_sdr0.det0.yn_1[12] ),
    .B(_2378_));
 sg13g2_nor2_1 _3342_ (.A(_2376_),
    .B(_2379_),
    .Y(_2380_));
 sg13g2_xor2_1 _3343_ (.B(_2379_),
    .A(_2376_),
    .X(_2381_));
 sg13g2_xnor2_1 _3344_ (.Y(_2382_),
    .A(_2374_),
    .B(_2381_));
 sg13g2_a21oi_1 _3345_ (.A1(_2371_),
    .A2(_2382_),
    .Y(_2383_),
    .B1(_2370_));
 sg13g2_a21oi_1 _3346_ (.A1(_2364_),
    .A2(_2368_),
    .Y(_2384_),
    .B1(_2363_));
 sg13g2_a21oi_2 _3347_ (.B1(_2359_),
    .Y(_2385_),
    .A2(_2360_),
    .A1(net405));
 sg13g2_nand2_1 _3348_ (.Y(_2386_),
    .A(net405),
    .B(\am_sdr0.det0.yn_1[5] ));
 sg13g2_xor2_1 _3349_ (.B(\am_sdr0.det0.yn_1[5] ),
    .A(net405),
    .X(_2387_));
 sg13g2_nand2_1 _3350_ (.Y(_2388_),
    .A(net404),
    .B(_2387_));
 sg13g2_xnor2_1 _3351_ (.Y(_2389_),
    .A(net404),
    .B(_2387_));
 sg13g2_nor2_1 _3352_ (.A(_2385_),
    .B(_2389_),
    .Y(_2390_));
 sg13g2_xor2_1 _3353_ (.B(_2389_),
    .A(_2385_),
    .X(_2391_));
 sg13g2_and2_1 _3354_ (.A(\am_sdr0.det0.yn_1[9] ),
    .B(\am_sdr0.det0.yn_1[8] ),
    .X(_2392_));
 sg13g2_xor2_1 _3355_ (.B(\am_sdr0.det0.yn_1[8] ),
    .A(\am_sdr0.det0.yn_1[9] ),
    .X(_2393_));
 sg13g2_xnor2_1 _3356_ (.Y(_2394_),
    .A(\am_sdr0.det0.yn_1[10] ),
    .B(_2393_));
 sg13g2_inv_1 _3357_ (.Y(_2395_),
    .A(_2394_));
 sg13g2_xnor2_1 _3358_ (.Y(_2396_),
    .A(_2391_),
    .B(_2395_));
 sg13g2_nor2_1 _3359_ (.A(_2384_),
    .B(_2396_),
    .Y(_2397_));
 sg13g2_xor2_1 _3360_ (.B(_2396_),
    .A(_2384_),
    .X(_2398_));
 sg13g2_a21oi_2 _3361_ (.B1(_2377_),
    .Y(_2399_),
    .A2(_2378_),
    .A1(\am_sdr0.det0.yn_1[12] ));
 sg13g2_inv_1 _3362_ (.Y(_2400_),
    .A(_2399_));
 sg13g2_a21oi_2 _3363_ (.B1(_2365_),
    .Y(_2401_),
    .A2(_2366_),
    .A1(\am_sdr0.det0.yn_1[9] ));
 sg13g2_and2_1 _3364_ (.A(\am_sdr0.det0.yn_1[11] ),
    .B(\am_sdr0.det0.yn_1[12] ),
    .X(_2402_));
 sg13g2_xor2_1 _3365_ (.B(\am_sdr0.det0.yn_1[12] ),
    .A(\am_sdr0.det0.yn_1[11] ),
    .X(_2403_));
 sg13g2_xnor2_1 _3366_ (.Y(_2404_),
    .A(\am_sdr0.det0.yn_1[13] ),
    .B(_2403_));
 sg13g2_nor2_1 _3367_ (.A(_2401_),
    .B(_2404_),
    .Y(_2405_));
 sg13g2_xor2_1 _3368_ (.B(_2404_),
    .A(_2401_),
    .X(_2406_));
 sg13g2_xnor2_1 _3369_ (.Y(_2407_),
    .A(_2399_),
    .B(_2406_));
 sg13g2_xnor2_1 _3370_ (.Y(_2408_),
    .A(_2398_),
    .B(_2407_));
 sg13g2_a21oi_1 _3371_ (.A1(_2375_),
    .A2(_2381_),
    .Y(_2409_),
    .B1(_2380_));
 sg13g2_xor2_1 _3372_ (.B(_2408_),
    .A(_2383_),
    .X(_2410_));
 sg13g2_nand2b_1 _3373_ (.Y(_2411_),
    .B(_2410_),
    .A_N(_2409_));
 sg13g2_o21ai_1 _3374_ (.B1(_2411_),
    .Y(_2412_),
    .A1(_2383_),
    .A2(_2408_));
 sg13g2_a21oi_1 _3375_ (.A1(_2400_),
    .A2(_2406_),
    .Y(_2413_),
    .B1(_2405_));
 sg13g2_a21oi_1 _3376_ (.A1(_2398_),
    .A2(_2407_),
    .Y(_2414_),
    .B1(_2397_));
 sg13g2_a21oi_1 _3377_ (.A1(_2391_),
    .A2(_2395_),
    .Y(_2415_),
    .B1(_2390_));
 sg13g2_and2_2 _3378_ (.A(_2386_),
    .B(_2388_),
    .X(_2416_));
 sg13g2_nand2b_1 _3379_ (.Y(_2417_),
    .B(_2356_),
    .A_N(_2416_));
 sg13g2_xnor2_1 _3380_ (.Y(_2418_),
    .A(_2355_),
    .B(_2416_));
 sg13g2_xnor2_1 _3381_ (.Y(_2419_),
    .A(\am_sdr0.det0.yn_1[11] ),
    .B(_2373_));
 sg13g2_xor2_1 _3382_ (.B(_2419_),
    .A(_2418_),
    .X(_2420_));
 sg13g2_nor2b_1 _3383_ (.A(_2415_),
    .B_N(_2420_),
    .Y(_2421_));
 sg13g2_xnor2_1 _3384_ (.Y(_2422_),
    .A(_2415_),
    .B(_2420_));
 sg13g2_a21oi_2 _3385_ (.B1(_2402_),
    .Y(_2423_),
    .A2(_2403_),
    .A1(\am_sdr0.det0.yn_1[13] ));
 sg13g2_inv_1 _3386_ (.Y(_2424_),
    .A(_2423_));
 sg13g2_a21oi_2 _3387_ (.B1(_2392_),
    .Y(_2425_),
    .A2(_2393_),
    .A1(\am_sdr0.det0.yn_1[10] ));
 sg13g2_inv_1 _3388_ (.Y(_2426_),
    .A(_2425_));
 sg13g2_and2_1 _3389_ (.A(\am_sdr0.det0.yn_1[12] ),
    .B(\am_sdr0.det0.yn_1[13] ),
    .X(_2427_));
 sg13g2_xor2_1 _3390_ (.B(\am_sdr0.det0.yn_1[13] ),
    .A(\am_sdr0.det0.yn_1[12] ),
    .X(_2428_));
 sg13g2_xnor2_1 _3391_ (.Y(_2429_),
    .A(\am_sdr0.det0.yn_1[14] ),
    .B(_2428_));
 sg13g2_nor2_1 _3392_ (.A(_2425_),
    .B(_2429_),
    .Y(_2430_));
 sg13g2_xor2_1 _3393_ (.B(_2429_),
    .A(_2425_),
    .X(_2431_));
 sg13g2_xnor2_1 _3394_ (.Y(_2432_),
    .A(_2423_),
    .B(_2431_));
 sg13g2_xnor2_1 _3395_ (.Y(_2433_),
    .A(_2422_),
    .B(_2432_));
 sg13g2_xor2_1 _3396_ (.B(_2433_),
    .A(_2414_),
    .X(_2434_));
 sg13g2_nand2b_1 _3397_ (.Y(_2435_),
    .B(_2434_),
    .A_N(_2413_));
 sg13g2_xnor2_1 _3398_ (.Y(_2436_),
    .A(_2413_),
    .B(_2434_));
 sg13g2_and2_1 _3399_ (.A(_2412_),
    .B(_2436_),
    .X(_2437_));
 sg13g2_xor2_1 _3400_ (.B(_2436_),
    .A(_2412_),
    .X(_2438_));
 sg13g2_a21oi_1 _3401_ (.A1(\am_sdr0.det0.yn_1[15] ),
    .A2(_2438_),
    .Y(_2439_),
    .B1(_2437_));
 sg13g2_o21ai_1 _3402_ (.B1(_2435_),
    .Y(_2440_),
    .A1(_2414_),
    .A2(_2433_));
 sg13g2_a21oi_1 _3403_ (.A1(_2424_),
    .A2(_2431_),
    .Y(_2441_),
    .B1(_2430_));
 sg13g2_inv_1 _3404_ (.Y(_2442_),
    .A(_2441_));
 sg13g2_a21oi_2 _3405_ (.B1(_2421_),
    .Y(_2443_),
    .A2(_2432_),
    .A1(_2422_));
 sg13g2_o21ai_1 _3406_ (.B1(_2417_),
    .Y(_2444_),
    .A1(_2418_),
    .A2(_2419_));
 sg13g2_or2_1 _3407_ (.X(_2445_),
    .B(_2376_),
    .A(_2367_));
 sg13g2_xnor2_1 _3408_ (.Y(_2446_),
    .A(_2367_),
    .B(_2376_));
 sg13g2_xor2_1 _3409_ (.B(_2446_),
    .A(_2379_),
    .X(_2447_));
 sg13g2_xnor2_1 _3410_ (.Y(_2448_),
    .A(_2444_),
    .B(_2447_));
 sg13g2_a21oi_2 _3411_ (.B1(_2427_),
    .Y(_2449_),
    .A2(_2428_),
    .A1(\am_sdr0.det0.yn_1[14] ));
 sg13g2_and2_1 _3412_ (.A(\am_sdr0.det0.yn_1[13] ),
    .B(\am_sdr0.det0.yn_1[14] ),
    .X(_2450_));
 sg13g2_xor2_1 _3413_ (.B(\am_sdr0.det0.yn_1[14] ),
    .A(\am_sdr0.det0.yn_1[13] ),
    .X(_2451_));
 sg13g2_xnor2_1 _3414_ (.Y(_2452_),
    .A(\am_sdr0.det0.yn_1[15] ),
    .B(_2451_));
 sg13g2_inv_1 _3415_ (.Y(_2453_),
    .A(_2452_));
 sg13g2_xor2_1 _3416_ (.B(_2452_),
    .A(_2374_),
    .X(_2454_));
 sg13g2_nand2b_1 _3417_ (.Y(_2455_),
    .B(_2454_),
    .A_N(_2449_));
 sg13g2_xnor2_1 _3418_ (.Y(_2456_),
    .A(_2449_),
    .B(_2454_));
 sg13g2_nor2b_1 _3419_ (.A(_2448_),
    .B_N(_2456_),
    .Y(_2457_));
 sg13g2_xnor2_1 _3420_ (.Y(_2458_),
    .A(_2448_),
    .B(_2456_));
 sg13g2_nor2b_1 _3421_ (.A(_2443_),
    .B_N(_2458_),
    .Y(_2459_));
 sg13g2_xnor2_1 _3422_ (.Y(_2460_),
    .A(_2443_),
    .B(_2458_));
 sg13g2_xnor2_1 _3423_ (.Y(_2461_),
    .A(_2441_),
    .B(_2460_));
 sg13g2_and2_1 _3424_ (.A(_2440_),
    .B(_2461_),
    .X(_2462_));
 sg13g2_xor2_1 _3425_ (.B(_2461_),
    .A(_2440_),
    .X(_2463_));
 sg13g2_xnor2_1 _3426_ (.Y(_2464_),
    .A(net403),
    .B(_2463_));
 sg13g2_nor2_1 _3427_ (.A(_2439_),
    .B(_2464_),
    .Y(_2465_));
 sg13g2_and2_1 _3428_ (.A(\am_sdr0.det0.yn_1[2] ),
    .B(\am_sdr0.det0.yn_1[1] ),
    .X(_2466_));
 sg13g2_xor2_1 _3429_ (.B(\am_sdr0.det0.yn_1[1] ),
    .A(\am_sdr0.det0.yn_1[2] ),
    .X(_2467_));
 sg13g2_a21oi_2 _3430_ (.B1(_2466_),
    .Y(_2468_),
    .A2(_2467_),
    .A1(\am_sdr0.det0.yn_1[3] ));
 sg13g2_xnor2_1 _3431_ (.Y(_2469_),
    .A(\am_sdr0.det0.yn_1[4] ),
    .B(_2346_));
 sg13g2_nor2_1 _3432_ (.A(_2468_),
    .B(_2469_),
    .Y(_2470_));
 sg13g2_nand2_1 _3433_ (.Y(_2471_),
    .A(_2468_),
    .B(_2469_));
 sg13g2_nand2b_2 _3434_ (.Y(_2472_),
    .B(_2471_),
    .A_N(_2470_));
 sg13g2_nor2_1 _3435_ (.A(_2389_),
    .B(_2472_),
    .Y(_2473_));
 sg13g2_nor2_2 _3436_ (.A(_2470_),
    .B(_2473_),
    .Y(_2474_));
 sg13g2_xnor2_1 _3437_ (.Y(_2475_),
    .A(_2352_),
    .B(_2356_));
 sg13g2_nor2_1 _3438_ (.A(_2474_),
    .B(_2475_),
    .Y(_2476_));
 sg13g2_xor2_1 _3439_ (.B(_2475_),
    .A(_2474_),
    .X(_2477_));
 sg13g2_nor2_1 _3440_ (.A(_2416_),
    .B(_2419_),
    .Y(_2478_));
 sg13g2_xor2_1 _3441_ (.B(_2419_),
    .A(_2416_),
    .X(_2479_));
 sg13g2_xnor2_1 _3442_ (.Y(_2480_),
    .A(_2425_),
    .B(_2479_));
 sg13g2_a21oi_1 _3443_ (.A1(_2477_),
    .A2(_2480_),
    .Y(_2481_),
    .B1(_2476_));
 sg13g2_xnor2_1 _3444_ (.Y(_2482_),
    .A(_2371_),
    .B(_2382_));
 sg13g2_nor2_1 _3445_ (.A(_2481_),
    .B(_2482_),
    .Y(_2483_));
 sg13g2_a21oi_1 _3446_ (.A1(_2426_),
    .A2(_2479_),
    .Y(_2484_),
    .B1(_2478_));
 sg13g2_inv_1 _3447_ (.Y(_2485_),
    .A(_2484_));
 sg13g2_xor2_1 _3448_ (.B(_2482_),
    .A(_2481_),
    .X(_2486_));
 sg13g2_a21oi_1 _3449_ (.A1(_2485_),
    .A2(_2486_),
    .Y(_2487_),
    .B1(_2483_));
 sg13g2_xnor2_1 _3450_ (.Y(_2488_),
    .A(_2409_),
    .B(_2410_));
 sg13g2_nand2b_1 _3451_ (.Y(_2489_),
    .B(_2488_),
    .A_N(_2487_));
 sg13g2_xnor2_1 _3452_ (.Y(_2490_),
    .A(_2487_),
    .B(_2488_));
 sg13g2_nand2_1 _3453_ (.Y(_2491_),
    .A(\am_sdr0.det0.yn_1[14] ),
    .B(_2490_));
 sg13g2_and2_1 _3454_ (.A(_2489_),
    .B(_2491_),
    .X(_2492_));
 sg13g2_xnor2_1 _3455_ (.Y(_2493_),
    .A(\am_sdr0.det0.yn_1[15] ),
    .B(_2438_));
 sg13g2_nor2_1 _3456_ (.A(_2492_),
    .B(_2493_),
    .Y(_2494_));
 sg13g2_inv_1 _3457_ (.Y(_2495_),
    .A(_2494_));
 sg13g2_and2_1 _3458_ (.A(\am_sdr0.det0.yn_1[1] ),
    .B(\am_sdr0.det0.alpha_yn_1[0] ),
    .X(_2496_));
 sg13g2_nand2_1 _3459_ (.Y(_2497_),
    .A(\am_sdr0.det0.yn_1[1] ),
    .B(\am_sdr0.det0.alpha_yn_1[0] ));
 sg13g2_xor2_1 _3460_ (.B(\am_sdr0.det0.alpha_yn_1[0] ),
    .A(\am_sdr0.det0.yn_1[1] ),
    .X(_2498_));
 sg13g2_a21oi_2 _3461_ (.B1(_2496_),
    .Y(_2499_),
    .A2(_2498_),
    .A1(\am_sdr0.det0.yn_1[2] ));
 sg13g2_xnor2_1 _3462_ (.Y(_2500_),
    .A(\am_sdr0.det0.yn_1[3] ),
    .B(_2467_));
 sg13g2_nor2_1 _3463_ (.A(_2499_),
    .B(_2500_),
    .Y(_2501_));
 sg13g2_xor2_1 _3464_ (.B(_2500_),
    .A(_2499_),
    .X(_2502_));
 sg13g2_a21oi_2 _3465_ (.B1(_2501_),
    .Y(_2503_),
    .A2(_2502_),
    .A1(_2362_));
 sg13g2_xor2_1 _3466_ (.B(_2472_),
    .A(_2389_),
    .X(_2504_));
 sg13g2_nor2b_1 _3467_ (.A(_2503_),
    .B_N(_2504_),
    .Y(_2505_));
 sg13g2_xnor2_1 _3468_ (.Y(_2506_),
    .A(_2503_),
    .B(_2504_));
 sg13g2_xor2_1 _3469_ (.B(_2394_),
    .A(_2385_),
    .X(_2507_));
 sg13g2_nand2b_1 _3470_ (.Y(_2508_),
    .B(_2507_),
    .A_N(_2401_));
 sg13g2_xnor2_1 _3471_ (.Y(_2509_),
    .A(_2401_),
    .B(_2507_));
 sg13g2_a21oi_2 _3472_ (.B1(_2505_),
    .Y(_2510_),
    .A2(_2509_),
    .A1(_2506_));
 sg13g2_xnor2_1 _3473_ (.Y(_2511_),
    .A(_2477_),
    .B(_2480_));
 sg13g2_o21ai_1 _3474_ (.B1(_2508_),
    .Y(_2512_),
    .A1(_2385_),
    .A2(_2394_));
 sg13g2_xor2_1 _3475_ (.B(_2511_),
    .A(_2510_),
    .X(_2513_));
 sg13g2_nand2_1 _3476_ (.Y(_2514_),
    .A(_2512_),
    .B(_2513_));
 sg13g2_o21ai_1 _3477_ (.B1(_2514_),
    .Y(_2515_),
    .A1(_2510_),
    .A2(_2511_));
 sg13g2_xnor2_1 _3478_ (.Y(_2516_),
    .A(_2484_),
    .B(_2486_));
 sg13g2_and2_1 _3479_ (.A(_2515_),
    .B(_2516_),
    .X(_2517_));
 sg13g2_xor2_1 _3480_ (.B(_2516_),
    .A(_2515_),
    .X(_2518_));
 sg13g2_a21oi_1 _3481_ (.A1(\am_sdr0.det0.yn_1[13] ),
    .A2(_2518_),
    .Y(_2519_),
    .B1(_2517_));
 sg13g2_xnor2_1 _3482_ (.Y(_2520_),
    .A(\am_sdr0.det0.yn_1[14] ),
    .B(_2490_));
 sg13g2_or2_1 _3483_ (.X(_2521_),
    .B(_2520_),
    .A(_2519_));
 sg13g2_xnor2_1 _3484_ (.Y(_2522_),
    .A(\am_sdr0.det0.yn_1[2] ),
    .B(_2498_));
 sg13g2_a22oi_1 _3485_ (.Y(_2523_),
    .B1(_2497_),
    .B2(_2522_),
    .A2(_2466_),
    .A1(\am_sdr0.det0.alpha_yn_1[0] ));
 sg13g2_a221oi_1 _3486_ (.B2(_2522_),
    .C1(_2350_),
    .B1(_2497_),
    .A1(\am_sdr0.det0.alpha_yn_1[0] ),
    .Y(_2524_),
    .A2(_2466_));
 sg13g2_a21oi_2 _3487_ (.B1(_2524_),
    .Y(_2525_),
    .A2(_2496_),
    .A1(\am_sdr0.det0.yn_1[2] ));
 sg13g2_xnor2_1 _3488_ (.Y(_2526_),
    .A(_2361_),
    .B(_2502_));
 sg13g2_nor2b_1 _3489_ (.A(_2525_),
    .B_N(_2526_),
    .Y(_2527_));
 sg13g2_nor2_1 _3490_ (.A(_2358_),
    .B(_2367_),
    .Y(_2528_));
 sg13g2_xor2_1 _3491_ (.B(_2367_),
    .A(_2358_),
    .X(_2529_));
 sg13g2_nor2b_1 _3492_ (.A(_2376_),
    .B_N(_2529_),
    .Y(_2530_));
 sg13g2_xnor2_1 _3493_ (.Y(_2531_),
    .A(_2376_),
    .B(_2529_));
 sg13g2_xnor2_1 _3494_ (.Y(_2532_),
    .A(_2525_),
    .B(_2526_));
 sg13g2_a21oi_1 _3495_ (.A1(_2531_),
    .A2(_2532_),
    .Y(_2533_),
    .B1(_2527_));
 sg13g2_xnor2_1 _3496_ (.Y(_2534_),
    .A(_2506_),
    .B(_2509_));
 sg13g2_nor2_1 _3497_ (.A(_2528_),
    .B(_2530_),
    .Y(_2535_));
 sg13g2_xor2_1 _3498_ (.B(_2534_),
    .A(_2533_),
    .X(_2536_));
 sg13g2_nand2b_1 _3499_ (.Y(_2537_),
    .B(_2536_),
    .A_N(_2535_));
 sg13g2_o21ai_1 _3500_ (.B1(_2537_),
    .Y(_2538_),
    .A1(_2533_),
    .A2(_2534_));
 sg13g2_xor2_1 _3501_ (.B(_2513_),
    .A(_2512_),
    .X(_2539_));
 sg13g2_and2_1 _3502_ (.A(_2538_),
    .B(_2539_),
    .X(_2540_));
 sg13g2_xor2_1 _3503_ (.B(_2539_),
    .A(_2538_),
    .X(_2541_));
 sg13g2_a21oi_1 _3504_ (.A1(\am_sdr0.det0.yn_1[12] ),
    .A2(_2541_),
    .Y(_2542_),
    .B1(_2540_));
 sg13g2_xnor2_1 _3505_ (.Y(_2543_),
    .A(\am_sdr0.det0.yn_1[13] ),
    .B(_2518_));
 sg13g2_nor2_1 _3506_ (.A(_2542_),
    .B(_2543_),
    .Y(_2544_));
 sg13g2_inv_1 _3507_ (.Y(_2545_),
    .A(_2544_));
 sg13g2_nor2b_1 _3508_ (.A(_2469_),
    .B_N(_2498_),
    .Y(_2546_));
 sg13g2_xnor2_1 _3509_ (.Y(_2547_),
    .A(_2350_),
    .B(_2523_));
 sg13g2_nand2_1 _3510_ (.Y(_2548_),
    .A(_2546_),
    .B(_2547_));
 sg13g2_xor2_1 _3511_ (.B(_2355_),
    .A(_2347_),
    .X(_2549_));
 sg13g2_nand2b_1 _3512_ (.Y(_2550_),
    .B(_2549_),
    .A_N(_2416_));
 sg13g2_xor2_1 _3513_ (.B(_2549_),
    .A(_2416_),
    .X(_2551_));
 sg13g2_xnor2_1 _3514_ (.Y(_2552_),
    .A(_2546_),
    .B(_2547_));
 sg13g2_o21ai_1 _3515_ (.B1(_2548_),
    .Y(_2553_),
    .A1(_2551_),
    .A2(_2552_));
 sg13g2_xnor2_1 _3516_ (.Y(_2554_),
    .A(_2531_),
    .B(_2532_));
 sg13g2_nor2b_1 _3517_ (.A(_2554_),
    .B_N(_2553_),
    .Y(_2555_));
 sg13g2_o21ai_1 _3518_ (.B1(_2550_),
    .Y(_2556_),
    .A1(_2347_),
    .A2(_2355_));
 sg13g2_nand2b_1 _3519_ (.Y(_2557_),
    .B(_2554_),
    .A_N(_2553_));
 sg13g2_xor2_1 _3520_ (.B(_2554_),
    .A(_2553_),
    .X(_2558_));
 sg13g2_a21o_1 _3521_ (.A2(_2557_),
    .A1(_2556_),
    .B1(_2555_),
    .X(_2559_));
 sg13g2_xnor2_1 _3522_ (.Y(_2560_),
    .A(_2535_),
    .B(_2536_));
 sg13g2_and2_1 _3523_ (.A(_2559_),
    .B(_2560_),
    .X(_2561_));
 sg13g2_xor2_1 _3524_ (.B(_2560_),
    .A(_2559_),
    .X(_2562_));
 sg13g2_a21oi_1 _3525_ (.A1(\am_sdr0.det0.yn_1[11] ),
    .A2(_2562_),
    .Y(_2563_),
    .B1(_2561_));
 sg13g2_xnor2_1 _3526_ (.Y(_2564_),
    .A(\am_sdr0.det0.yn_1[12] ),
    .B(_2541_));
 sg13g2_or2_1 _3527_ (.X(_2565_),
    .B(_2564_),
    .A(_2563_));
 sg13g2_or2_2 _3528_ (.X(_2566_),
    .B(_2500_),
    .A(_2174_));
 sg13g2_xnor2_1 _3529_ (.Y(_2567_),
    .A(_2469_),
    .B(_2498_));
 sg13g2_nand2b_1 _3530_ (.Y(_2568_),
    .B(_2567_),
    .A_N(_2566_));
 sg13g2_xnor2_1 _3531_ (.Y(_2569_),
    .A(_2566_),
    .B(_2567_));
 sg13g2_nor2_1 _3532_ (.A(_2389_),
    .B(_2468_),
    .Y(_2570_));
 sg13g2_xnor2_1 _3533_ (.Y(_2571_),
    .A(_2389_),
    .B(_2468_));
 sg13g2_nor2_1 _3534_ (.A(_2385_),
    .B(_2571_),
    .Y(_2572_));
 sg13g2_xor2_1 _3535_ (.B(_2571_),
    .A(_2385_),
    .X(_2573_));
 sg13g2_nand2_1 _3536_ (.Y(_2574_),
    .A(_2569_),
    .B(_2573_));
 sg13g2_and2_1 _3537_ (.A(_2568_),
    .B(_2574_),
    .X(_2575_));
 sg13g2_xnor2_1 _3538_ (.Y(_2576_),
    .A(_2551_),
    .B(_2552_));
 sg13g2_or2_1 _3539_ (.X(_2577_),
    .B(_2576_),
    .A(_2575_));
 sg13g2_nor2_1 _3540_ (.A(_2570_),
    .B(_2572_),
    .Y(_2578_));
 sg13g2_and2_1 _3541_ (.A(_2575_),
    .B(_2576_),
    .X(_2579_));
 sg13g2_xor2_1 _3542_ (.B(_2576_),
    .A(_2575_),
    .X(_2580_));
 sg13g2_o21ai_1 _3543_ (.B1(_2577_),
    .Y(_2581_),
    .A1(_2578_),
    .A2(_2579_));
 sg13g2_xnor2_1 _3544_ (.Y(_2582_),
    .A(_2556_),
    .B(_2558_));
 sg13g2_xnor2_1 _3545_ (.Y(_2583_),
    .A(_2581_),
    .B(_2582_));
 sg13g2_nor2_1 _3546_ (.A(_2175_),
    .B(_2583_),
    .Y(_2584_));
 sg13g2_a21oi_1 _3547_ (.A1(_2581_),
    .A2(_2582_),
    .Y(_2585_),
    .B1(_2584_));
 sg13g2_xnor2_1 _3548_ (.Y(_2586_),
    .A(\am_sdr0.det0.yn_1[11] ),
    .B(_2562_));
 sg13g2_nor2_1 _3549_ (.A(_2585_),
    .B(_2586_),
    .Y(_2587_));
 sg13g2_nor2_1 _3550_ (.A(_2361_),
    .B(_2499_),
    .Y(_2588_));
 sg13g2_xnor2_1 _3551_ (.Y(_2589_),
    .A(_2361_),
    .B(_2499_));
 sg13g2_nor2_1 _3552_ (.A(_2358_),
    .B(_2589_),
    .Y(_2590_));
 sg13g2_xor2_1 _3553_ (.B(_2589_),
    .A(_2358_),
    .X(_2591_));
 sg13g2_nand2_1 _3554_ (.Y(_2592_),
    .A(_2174_),
    .B(_2500_));
 sg13g2_nand2_1 _3555_ (.Y(_2593_),
    .A(_2566_),
    .B(_2592_));
 sg13g2_and3_1 _3556_ (.X(_2594_),
    .A(_2566_),
    .B(_2591_),
    .C(_2592_));
 sg13g2_xor2_1 _3557_ (.B(_2573_),
    .A(_2569_),
    .X(_2595_));
 sg13g2_nand2_1 _3558_ (.Y(_2596_),
    .A(_2594_),
    .B(_2595_));
 sg13g2_nor2_1 _3559_ (.A(_2588_),
    .B(_2590_),
    .Y(_2597_));
 sg13g2_xnor2_1 _3560_ (.Y(_2598_),
    .A(_2594_),
    .B(_2595_));
 sg13g2_o21ai_1 _3561_ (.B1(_2596_),
    .Y(_2599_),
    .A1(_2597_),
    .A2(_2598_));
 sg13g2_xnor2_1 _3562_ (.Y(_2600_),
    .A(_2578_),
    .B(_2580_));
 sg13g2_and2_1 _3563_ (.A(_2599_),
    .B(_2600_),
    .X(_2601_));
 sg13g2_xor2_1 _3564_ (.B(_2600_),
    .A(_2599_),
    .X(_2602_));
 sg13g2_a21oi_1 _3565_ (.A1(\am_sdr0.det0.yn_1[9] ),
    .A2(_2602_),
    .Y(_2603_),
    .B1(_2601_));
 sg13g2_xnor2_1 _3566_ (.Y(_2604_),
    .A(_2175_),
    .B(_2583_));
 sg13g2_or2_1 _3567_ (.X(_2605_),
    .B(_2604_),
    .A(_2603_));
 sg13g2_xor2_1 _3568_ (.B(_2604_),
    .A(_2603_),
    .X(_2606_));
 sg13g2_xnor2_1 _3569_ (.Y(_2607_),
    .A(\am_sdr0.det0.yn_1[9] ),
    .B(_2602_));
 sg13g2_xor2_1 _3570_ (.B(_2593_),
    .A(_2591_),
    .X(_2608_));
 sg13g2_xnor2_1 _3571_ (.Y(_2609_),
    .A(_2350_),
    .B(_2496_));
 sg13g2_nand2b_1 _3572_ (.Y(_2610_),
    .B(_2609_),
    .A_N(_2347_));
 sg13g2_xnor2_1 _3573_ (.Y(_2611_),
    .A(_2347_),
    .B(_2609_));
 sg13g2_nor2b_1 _3574_ (.A(_2522_),
    .B_N(_2611_),
    .Y(_2612_));
 sg13g2_nor2b_1 _3575_ (.A(_2608_),
    .B_N(_2612_),
    .Y(_2613_));
 sg13g2_o21ai_1 _3576_ (.B1(_2610_),
    .Y(_2614_),
    .A1(_2350_),
    .A2(_2497_));
 sg13g2_xnor2_1 _3577_ (.Y(_2615_),
    .A(_2608_),
    .B(_2612_));
 sg13g2_a21oi_1 _3578_ (.A1(_2614_),
    .A2(_2615_),
    .Y(_2616_),
    .B1(_2613_));
 sg13g2_xor2_1 _3579_ (.B(_2598_),
    .A(_2597_),
    .X(_2617_));
 sg13g2_nor2b_1 _3580_ (.A(_2616_),
    .B_N(_2617_),
    .Y(_2618_));
 sg13g2_xnor2_1 _3581_ (.Y(_2619_),
    .A(_2616_),
    .B(_2617_));
 sg13g2_a21oi_1 _3582_ (.A1(\am_sdr0.det0.yn_1[8] ),
    .A2(_2619_),
    .Y(_2620_),
    .B1(_2618_));
 sg13g2_nor2_1 _3583_ (.A(_2607_),
    .B(_2620_),
    .Y(_2621_));
 sg13g2_xor2_1 _3584_ (.B(_2619_),
    .A(\am_sdr0.det0.yn_1[8] ),
    .X(_2622_));
 sg13g2_xnor2_1 _3585_ (.Y(_2623_),
    .A(_2522_),
    .B(_2611_));
 sg13g2_a21oi_1 _3586_ (.A1(_2471_),
    .A2(_2498_),
    .Y(_2624_),
    .B1(_2470_));
 sg13g2_nand2b_1 _3587_ (.Y(_2625_),
    .B(_2623_),
    .A_N(_2624_));
 sg13g2_xor2_1 _3588_ (.B(_2615_),
    .A(_2614_),
    .X(_2626_));
 sg13g2_nor2b_1 _3589_ (.A(_2625_),
    .B_N(_2626_),
    .Y(_2627_));
 sg13g2_xnor2_1 _3590_ (.Y(_2628_),
    .A(_2625_),
    .B(_2626_));
 sg13g2_a21o_1 _3591_ (.A2(_2628_),
    .A1(net404),
    .B1(_2627_),
    .X(_2629_));
 sg13g2_nand2_1 _3592_ (.Y(_2630_),
    .A(_2622_),
    .B(_2629_));
 sg13g2_or2_1 _3593_ (.X(_2631_),
    .B(_2628_),
    .A(net404));
 sg13g2_nand2b_1 _3594_ (.Y(_2632_),
    .B(_2592_),
    .A_N(_2499_));
 sg13g2_xor2_1 _3595_ (.B(_2498_),
    .A(_2472_),
    .X(_2633_));
 sg13g2_a21oi_1 _3596_ (.A1(_2566_),
    .A2(_2632_),
    .Y(_2634_),
    .B1(_2633_));
 sg13g2_xnor2_1 _3597_ (.Y(_2635_),
    .A(_2623_),
    .B(_2624_));
 sg13g2_o21ai_1 _3598_ (.B1(_2634_),
    .Y(_2636_),
    .A1(net405),
    .A2(_2635_));
 sg13g2_nand2_1 _3599_ (.Y(_2637_),
    .A(net405),
    .B(_2635_));
 sg13g2_a22oi_1 _3600_ (.Y(_2638_),
    .B1(_2636_),
    .B2(_2637_),
    .A2(_2628_),
    .A1(net404));
 sg13g2_nand3_1 _3601_ (.B(\am_sdr0.det0.yn_1[5] ),
    .C(net404),
    .A(net405),
    .Y(_2639_));
 sg13g2_o21ai_1 _3602_ (.B1(_2639_),
    .Y(_2640_),
    .A1(_2388_),
    .A2(_2568_));
 sg13g2_a21oi_1 _3603_ (.A1(_2631_),
    .A2(_2638_),
    .Y(_2641_),
    .B1(_2640_));
 sg13g2_nor2_1 _3604_ (.A(_2622_),
    .B(_2629_),
    .Y(_2642_));
 sg13g2_a221oi_1 _3605_ (.B2(_2641_),
    .C1(_2642_),
    .B1(_2630_),
    .A1(_2607_),
    .Y(_2643_),
    .A2(_2620_));
 sg13g2_o21ai_1 _3606_ (.B1(_2606_),
    .Y(_2644_),
    .A1(_2621_),
    .A2(_2643_));
 sg13g2_xnor2_1 _3607_ (.Y(_2645_),
    .A(_2585_),
    .B(_2586_));
 sg13g2_a21oi_1 _3608_ (.A1(_2605_),
    .A2(_2644_),
    .Y(_2646_),
    .B1(_2645_));
 sg13g2_a21o_1 _3609_ (.A2(_2644_),
    .A1(_2605_),
    .B1(_2645_),
    .X(_2647_));
 sg13g2_nor2_1 _3610_ (.A(_2587_),
    .B(_2646_),
    .Y(_2648_));
 sg13g2_xor2_1 _3611_ (.B(_2564_),
    .A(_2563_),
    .X(_2649_));
 sg13g2_o21ai_1 _3612_ (.B1(_2649_),
    .Y(_2650_),
    .A1(_2587_),
    .A2(_2646_));
 sg13g2_xnor2_1 _3613_ (.Y(_2651_),
    .A(_2542_),
    .B(_2543_));
 sg13g2_a21oi_1 _3614_ (.A1(_2565_),
    .A2(_2650_),
    .Y(_2652_),
    .B1(_2651_));
 sg13g2_a21o_1 _3615_ (.A2(_2650_),
    .A1(_2565_),
    .B1(_2651_),
    .X(_2653_));
 sg13g2_xor2_1 _3616_ (.B(_2520_),
    .A(_2519_),
    .X(_2654_));
 sg13g2_inv_1 _3617_ (.Y(_2655_),
    .A(_2654_));
 sg13g2_a21oi_1 _3618_ (.A1(_2545_),
    .A2(_2653_),
    .Y(_2656_),
    .B1(_2655_));
 sg13g2_o21ai_1 _3619_ (.B1(_2654_),
    .Y(_2657_),
    .A1(_2544_),
    .A2(_2652_));
 sg13g2_xnor2_1 _3620_ (.Y(_2658_),
    .A(_2492_),
    .B(_2493_));
 sg13g2_a21o_1 _3621_ (.A2(_2657_),
    .A1(_2521_),
    .B1(_2658_),
    .X(_2659_));
 sg13g2_xor2_1 _3622_ (.B(_2464_),
    .A(_2439_),
    .X(_2660_));
 sg13g2_inv_1 _3623_ (.Y(_2661_),
    .A(_2660_));
 sg13g2_a21oi_2 _3624_ (.B1(_2661_),
    .Y(_2662_),
    .A2(_2659_),
    .A1(_2495_));
 sg13g2_a21oi_1 _3625_ (.A1(net403),
    .A2(_2463_),
    .Y(_2663_),
    .B1(_2462_));
 sg13g2_a21oi_1 _3626_ (.A1(_2442_),
    .A2(_2460_),
    .Y(_2664_),
    .B1(_2459_));
 sg13g2_o21ai_1 _3627_ (.B1(_2455_),
    .Y(_2665_),
    .A1(_2374_),
    .A2(_2452_));
 sg13g2_inv_1 _3628_ (.Y(_2666_),
    .A(_2665_));
 sg13g2_a21o_1 _3629_ (.A2(_2447_),
    .A1(_2444_),
    .B1(_2457_),
    .X(_2667_));
 sg13g2_o21ai_1 _3630_ (.B1(_2445_),
    .Y(_2668_),
    .A1(_2379_),
    .A2(_2446_));
 sg13g2_or2_1 _3631_ (.X(_2669_),
    .B(_2401_),
    .A(_2394_));
 sg13g2_xnor2_1 _3632_ (.Y(_2670_),
    .A(_2394_),
    .B(_2401_));
 sg13g2_xor2_1 _3633_ (.B(_2670_),
    .A(_2404_),
    .X(_2671_));
 sg13g2_nand2_1 _3634_ (.Y(_2672_),
    .A(_2668_),
    .B(_2671_));
 sg13g2_xnor2_1 _3635_ (.Y(_2673_),
    .A(_2668_),
    .B(_2671_));
 sg13g2_a21oi_2 _3636_ (.B1(_2450_),
    .Y(_2674_),
    .A2(_2451_),
    .A1(\am_sdr0.det0.yn_1[15] ));
 sg13g2_and2_1 _3637_ (.A(\am_sdr0.det0.yn_1[14] ),
    .B(\am_sdr0.det0.yn_1[15] ),
    .X(_2675_));
 sg13g2_xor2_1 _3638_ (.B(\am_sdr0.det0.yn_1[15] ),
    .A(\am_sdr0.det0.yn_1[14] ),
    .X(_2676_));
 sg13g2_xnor2_1 _3639_ (.Y(_2677_),
    .A(\am_sdr0.det0.yn_1[16] ),
    .B(_2676_));
 sg13g2_inv_1 _3640_ (.Y(_2678_),
    .A(_2677_));
 sg13g2_xor2_1 _3641_ (.B(_2677_),
    .A(_2399_),
    .X(_2679_));
 sg13g2_nand2b_1 _3642_ (.Y(_2680_),
    .B(_2679_),
    .A_N(_2674_));
 sg13g2_xnor2_1 _3643_ (.Y(_2681_),
    .A(_2674_),
    .B(_2679_));
 sg13g2_inv_1 _3644_ (.Y(_2682_),
    .A(_2681_));
 sg13g2_xnor2_1 _3645_ (.Y(_2683_),
    .A(_2673_),
    .B(_2681_));
 sg13g2_nand2_1 _3646_ (.Y(_2684_),
    .A(_2667_),
    .B(_2683_));
 sg13g2_xnor2_1 _3647_ (.Y(_2685_),
    .A(_2667_),
    .B(_2683_));
 sg13g2_xnor2_1 _3648_ (.Y(_2686_),
    .A(_2665_),
    .B(_2685_));
 sg13g2_nand2b_1 _3649_ (.Y(_2687_),
    .B(_2686_),
    .A_N(_2664_));
 sg13g2_xnor2_1 _3650_ (.Y(_2688_),
    .A(_2664_),
    .B(_2686_));
 sg13g2_nand2_1 _3651_ (.Y(_2689_),
    .A(net402),
    .B(_2688_));
 sg13g2_xnor2_1 _3652_ (.Y(_2690_),
    .A(net402),
    .B(_2688_));
 sg13g2_or2_1 _3653_ (.X(_2691_),
    .B(_2690_),
    .A(_2663_));
 sg13g2_xor2_1 _3654_ (.B(_2690_),
    .A(_2663_),
    .X(_2692_));
 sg13g2_o21ai_1 _3655_ (.B1(_2692_),
    .Y(_2693_),
    .A1(_2465_),
    .A2(_2662_));
 sg13g2_or3_1 _3656_ (.A(_2465_),
    .B(_2662_),
    .C(_2692_),
    .X(_2694_));
 sg13g2_and2_1 _3657_ (.A(_2693_),
    .B(_2694_),
    .X(_2695_));
 sg13g2_nand2_1 _3658_ (.Y(_2696_),
    .A(_2344_),
    .B(_2695_));
 sg13g2_and3_1 _3659_ (.X(_2697_),
    .A(_2495_),
    .B(_2659_),
    .C(_2661_));
 sg13g2_nor2_1 _3660_ (.A(\am_sdr0.det0.ifreq[7] ),
    .B(_2343_),
    .Y(_2698_));
 sg13g2_nor2_2 _3661_ (.A(_0024_),
    .B(_2698_),
    .Y(_2699_));
 sg13g2_nor2_1 _3662_ (.A(net430),
    .B(net330),
    .Y(_2700_));
 sg13g2_xnor2_1 _3663_ (.Y(_2701_),
    .A(\am_sdr0.det0.ifreq[6] ),
    .B(_2342_));
 sg13g2_a21oi_1 _3664_ (.A1(net330),
    .A2(_2701_),
    .Y(_2702_),
    .B1(_2700_));
 sg13g2_nor3_1 _3665_ (.A(_2662_),
    .B(_2697_),
    .C(_2702_),
    .Y(_2703_));
 sg13g2_nand3_1 _3666_ (.B(_2657_),
    .C(_2658_),
    .A(_2521_),
    .Y(_2704_));
 sg13g2_nand2_1 _3667_ (.Y(_2705_),
    .A(_2659_),
    .B(_2704_));
 sg13g2_nor2b_1 _3668_ (.A(_2341_),
    .B_N(\am_sdr0.det0.ifreq[5] ),
    .Y(_2706_));
 sg13g2_or3_1 _3669_ (.A(_0024_),
    .B(_2342_),
    .C(_2706_),
    .X(_2707_));
 sg13g2_o21ai_1 _3670_ (.B1(_2707_),
    .Y(_2708_),
    .A1(_0028_),
    .A2(net330));
 sg13g2_nand3_1 _3671_ (.B(_2704_),
    .C(_2708_),
    .A(_2659_),
    .Y(_2709_));
 sg13g2_nor3_1 _3672_ (.A(_2544_),
    .B(_2652_),
    .C(_2654_),
    .Y(_2710_));
 sg13g2_nor2_1 _3673_ (.A(net441),
    .B(net330),
    .Y(_2711_));
 sg13g2_xnor2_1 _3674_ (.Y(_2712_),
    .A(\am_sdr0.det0.ifreq[4] ),
    .B(_2340_));
 sg13g2_a21oi_1 _3675_ (.A1(net330),
    .A2(_2712_),
    .Y(_2713_),
    .B1(_2711_));
 sg13g2_nor3_1 _3676_ (.A(_2656_),
    .B(_2710_),
    .C(_2713_),
    .Y(_2714_));
 sg13g2_nand3_1 _3677_ (.B(_2650_),
    .C(_2651_),
    .A(_2565_),
    .Y(_2715_));
 sg13g2_nand2_1 _3678_ (.Y(_2716_),
    .A(\am_sdr0.det0.ifreq[3] ),
    .B(_2339_));
 sg13g2_nand3b_1 _3679_ (.B(net330),
    .C(_2716_),
    .Y(_2717_),
    .A_N(_2340_));
 sg13g2_o21ai_1 _3680_ (.B1(_2717_),
    .Y(_2718_),
    .A1(_0026_),
    .A2(net330));
 sg13g2_nand3_1 _3681_ (.B(_2715_),
    .C(_2718_),
    .A(_2653_),
    .Y(_2719_));
 sg13g2_xor2_1 _3682_ (.B(_2649_),
    .A(_2648_),
    .X(_2720_));
 sg13g2_nor2_1 _3683_ (.A(net438),
    .B(_2699_),
    .Y(_2721_));
 sg13g2_xnor2_1 _3684_ (.Y(_2722_),
    .A(\am_sdr0.det0.ifreq[2] ),
    .B(_2338_));
 sg13g2_a21oi_2 _3685_ (.B1(_2721_),
    .Y(_2723_),
    .A2(_2722_),
    .A1(net330));
 sg13g2_nor2_1 _3686_ (.A(_2720_),
    .B(_2723_),
    .Y(_2724_));
 sg13g2_nand3_1 _3687_ (.B(_2644_),
    .C(_2645_),
    .A(_2605_),
    .Y(_2725_));
 sg13g2_nand2_1 _3688_ (.Y(_2726_),
    .A(\am_sdr0.det0.ifreq[1] ),
    .B(\am_sdr0.det0.env_det[0] ));
 sg13g2_nand3b_1 _3689_ (.B(_2699_),
    .C(_2726_),
    .Y(_0184_),
    .A_N(_2338_));
 sg13g2_o21ai_1 _3690_ (.B1(_0184_),
    .Y(_0185_),
    .A1(_0023_),
    .A2(_2699_));
 sg13g2_nand3_1 _3691_ (.B(_2725_),
    .C(_0185_),
    .A(_2647_),
    .Y(_0186_));
 sg13g2_or3_1 _3692_ (.A(_2606_),
    .B(_2621_),
    .C(_2643_),
    .X(_0187_));
 sg13g2_nand2_1 _3693_ (.Y(_0188_),
    .A(_2644_),
    .B(_0187_));
 sg13g2_nand3_1 _3694_ (.B(_2644_),
    .C(_0187_),
    .A(net287),
    .Y(_0189_));
 sg13g2_a21o_1 _3695_ (.A2(_2725_),
    .A1(_2647_),
    .B1(_0185_),
    .X(_0190_));
 sg13g2_nand2_1 _3696_ (.Y(_0191_),
    .A(_0186_),
    .B(_0190_));
 sg13g2_o21ai_1 _3697_ (.B1(_0186_),
    .Y(_0192_),
    .A1(_0189_),
    .A2(_0191_));
 sg13g2_xor2_1 _3698_ (.B(_2723_),
    .A(_2720_),
    .X(_0193_));
 sg13g2_a21oi_1 _3699_ (.A1(_0192_),
    .A2(_0193_),
    .Y(_0194_),
    .B1(_2724_));
 sg13g2_a21o_1 _3700_ (.A2(_2715_),
    .A1(_2653_),
    .B1(_2718_),
    .X(_0195_));
 sg13g2_nand2_1 _3701_ (.Y(_0196_),
    .A(_2719_),
    .B(_0195_));
 sg13g2_o21ai_1 _3702_ (.B1(_2719_),
    .Y(_0197_),
    .A1(_0194_),
    .A2(_0196_));
 sg13g2_o21ai_1 _3703_ (.B1(_2713_),
    .Y(_0198_),
    .A1(_2656_),
    .A2(_2710_));
 sg13g2_nor2b_1 _3704_ (.A(_2714_),
    .B_N(_0198_),
    .Y(_0199_));
 sg13g2_a21oi_2 _3705_ (.B1(_2714_),
    .Y(_0200_),
    .A2(_0199_),
    .A1(_0197_));
 sg13g2_xor2_1 _3706_ (.B(_2708_),
    .A(_2705_),
    .X(_0201_));
 sg13g2_o21ai_1 _3707_ (.B1(_2709_),
    .Y(_0202_),
    .A1(_0200_),
    .A2(_0201_));
 sg13g2_o21ai_1 _3708_ (.B1(_2702_),
    .Y(_0203_),
    .A1(_2662_),
    .A2(_2697_));
 sg13g2_nor2b_1 _3709_ (.A(_2703_),
    .B_N(_0203_),
    .Y(_0204_));
 sg13g2_a21oi_2 _3710_ (.B1(_2703_),
    .Y(_0205_),
    .A2(_0204_),
    .A1(_0202_));
 sg13g2_xnor2_1 _3711_ (.Y(_0206_),
    .A(_2344_),
    .B(_2695_));
 sg13g2_o21ai_1 _3712_ (.B1(_2696_),
    .Y(_0207_),
    .A1(_0205_),
    .A2(_0206_));
 sg13g2_o21ai_1 _3713_ (.B1(_2684_),
    .Y(_0208_),
    .A1(_2666_),
    .A2(_2685_));
 sg13g2_o21ai_1 _3714_ (.B1(_2680_),
    .Y(_0209_),
    .A1(_2399_),
    .A2(_2677_));
 sg13g2_inv_1 _3715_ (.Y(_0210_),
    .A(_0209_));
 sg13g2_o21ai_1 _3716_ (.B1(_2672_),
    .Y(_0211_),
    .A1(_2673_),
    .A2(_2682_));
 sg13g2_o21ai_1 _3717_ (.B1(_2669_),
    .Y(_0212_),
    .A1(_2404_),
    .A2(_2670_));
 sg13g2_or2_1 _3718_ (.X(_0213_),
    .B(_2425_),
    .A(_2419_));
 sg13g2_xnor2_1 _3719_ (.Y(_0214_),
    .A(_2419_),
    .B(_2425_));
 sg13g2_xor2_1 _3720_ (.B(_0214_),
    .A(_2429_),
    .X(_0215_));
 sg13g2_xnor2_1 _3721_ (.Y(_0216_),
    .A(_0212_),
    .B(_0215_));
 sg13g2_a21oi_2 _3722_ (.B1(_2675_),
    .Y(_0217_),
    .A2(_2676_),
    .A1(net403));
 sg13g2_and2_1 _3723_ (.A(\am_sdr0.det0.yn_1[15] ),
    .B(net403),
    .X(_0218_));
 sg13g2_xor2_1 _3724_ (.B(net403),
    .A(\am_sdr0.det0.yn_1[15] ),
    .X(_0219_));
 sg13g2_xnor2_1 _3725_ (.Y(_0220_),
    .A(\am_sdr0.det0.yn_1[17] ),
    .B(_0219_));
 sg13g2_inv_1 _3726_ (.Y(_0221_),
    .A(_0220_));
 sg13g2_xor2_1 _3727_ (.B(_0220_),
    .A(_2423_),
    .X(_0222_));
 sg13g2_nor2b_1 _3728_ (.A(_0217_),
    .B_N(_0222_),
    .Y(_0223_));
 sg13g2_xnor2_1 _3729_ (.Y(_0224_),
    .A(_0217_),
    .B(_0222_));
 sg13g2_nor2b_1 _3730_ (.A(_0216_),
    .B_N(_0224_),
    .Y(_0225_));
 sg13g2_xnor2_1 _3731_ (.Y(_0226_),
    .A(_0216_),
    .B(_0224_));
 sg13g2_nand2_1 _3732_ (.Y(_0227_),
    .A(_0211_),
    .B(_0226_));
 sg13g2_xnor2_1 _3733_ (.Y(_0228_),
    .A(_0211_),
    .B(_0226_));
 sg13g2_xnor2_1 _3734_ (.Y(_0229_),
    .A(_0209_),
    .B(_0228_));
 sg13g2_and2_1 _3735_ (.A(_0208_),
    .B(_0229_),
    .X(_0230_));
 sg13g2_xor2_1 _3736_ (.B(_0229_),
    .A(_0208_),
    .X(_0231_));
 sg13g2_xnor2_1 _3737_ (.Y(_0232_),
    .A(net401),
    .B(_0231_));
 sg13g2_a21oi_1 _3738_ (.A1(_2687_),
    .A2(_2689_),
    .Y(_0233_),
    .B1(_0232_));
 sg13g2_nand3_1 _3739_ (.B(_2689_),
    .C(_0232_),
    .A(_2687_),
    .Y(_0234_));
 sg13g2_nand2b_1 _3740_ (.Y(_0235_),
    .B(_0234_),
    .A_N(_0233_));
 sg13g2_a21o_1 _3741_ (.A2(_2693_),
    .A1(_2691_),
    .B1(_0235_),
    .X(_0236_));
 sg13g2_nand3_1 _3742_ (.B(_2693_),
    .C(_0235_),
    .A(_2691_),
    .Y(_0237_));
 sg13g2_and2_1 _3743_ (.A(_0236_),
    .B(_0237_),
    .X(_0238_));
 sg13g2_and2_1 _3744_ (.A(_0207_),
    .B(_0238_),
    .X(_0239_));
 sg13g2_a21oi_1 _3745_ (.A1(net401),
    .A2(_0231_),
    .Y(_0240_),
    .B1(_0230_));
 sg13g2_o21ai_1 _3746_ (.B1(_0227_),
    .Y(_0241_),
    .A1(_0210_),
    .A2(_0228_));
 sg13g2_a21oi_1 _3747_ (.A1(_2424_),
    .A2(_0221_),
    .Y(_0242_),
    .B1(_0223_));
 sg13g2_a21o_1 _3748_ (.A2(_0215_),
    .A1(_0212_),
    .B1(_0225_),
    .X(_0243_));
 sg13g2_o21ai_1 _3749_ (.B1(_0213_),
    .Y(_0244_),
    .A1(_2429_),
    .A2(_0214_));
 sg13g2_nor2_1 _3750_ (.A(_2374_),
    .B(_2379_),
    .Y(_0245_));
 sg13g2_xor2_1 _3751_ (.B(_2379_),
    .A(_2374_),
    .X(_0246_));
 sg13g2_xnor2_1 _3752_ (.Y(_0247_),
    .A(_2452_),
    .B(_0246_));
 sg13g2_xnor2_1 _3753_ (.Y(_0248_),
    .A(_0244_),
    .B(_0247_));
 sg13g2_a21oi_2 _3754_ (.B1(_0218_),
    .Y(_0249_),
    .A2(_0219_),
    .A1(\am_sdr0.det0.yn_1[17] ));
 sg13g2_inv_1 _3755_ (.Y(_0250_),
    .A(_0249_));
 sg13g2_and2_1 _3756_ (.A(net403),
    .B(net402),
    .X(_0251_));
 sg13g2_xor2_1 _3757_ (.B(net402),
    .A(net403),
    .X(_0252_));
 sg13g2_xnor2_1 _3758_ (.Y(_0253_),
    .A(net400),
    .B(_0252_));
 sg13g2_inv_1 _3759_ (.Y(_0254_),
    .A(_0253_));
 sg13g2_nor2_1 _3760_ (.A(_2449_),
    .B(_0253_),
    .Y(_0255_));
 sg13g2_xor2_1 _3761_ (.B(_0253_),
    .A(_2449_),
    .X(_0256_));
 sg13g2_xnor2_1 _3762_ (.Y(_0257_),
    .A(_0249_),
    .B(_0256_));
 sg13g2_nor2b_1 _3763_ (.A(_0248_),
    .B_N(_0257_),
    .Y(_0258_));
 sg13g2_xnor2_1 _3764_ (.Y(_0259_),
    .A(_0248_),
    .B(_0257_));
 sg13g2_nand2_1 _3765_ (.Y(_0260_),
    .A(_0243_),
    .B(_0259_));
 sg13g2_xnor2_1 _3766_ (.Y(_0261_),
    .A(_0243_),
    .B(_0259_));
 sg13g2_xor2_1 _3767_ (.B(_0261_),
    .A(_0242_),
    .X(_0262_));
 sg13g2_and2_1 _3768_ (.A(_0241_),
    .B(_0262_),
    .X(_0263_));
 sg13g2_xor2_1 _3769_ (.B(_0262_),
    .A(_0241_),
    .X(_0264_));
 sg13g2_xnor2_1 _3770_ (.Y(_0265_),
    .A(net399),
    .B(_0264_));
 sg13g2_and2_1 _3771_ (.A(_0240_),
    .B(_0265_),
    .X(_0266_));
 sg13g2_nor2_1 _3772_ (.A(_0240_),
    .B(_0265_),
    .Y(_0267_));
 sg13g2_nor2_1 _3773_ (.A(_0266_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_nor2b_1 _3774_ (.A(_0233_),
    .B_N(_0236_),
    .Y(_0269_));
 sg13g2_xnor2_1 _3775_ (.Y(_0270_),
    .A(_0268_),
    .B(_0269_));
 sg13g2_nand2_1 _3776_ (.Y(_0271_),
    .A(_0239_),
    .B(_0270_));
 sg13g2_o21ai_1 _3777_ (.B1(_0260_),
    .Y(_0272_),
    .A1(_0242_),
    .A2(_0261_));
 sg13g2_a21oi_2 _3778_ (.B1(_0255_),
    .Y(_0273_),
    .A2(_0256_),
    .A1(_0250_));
 sg13g2_a21o_1 _3779_ (.A2(_0247_),
    .A1(_0244_),
    .B1(_0258_),
    .X(_0274_));
 sg13g2_a21oi_2 _3780_ (.B1(_0245_),
    .Y(_0275_),
    .A2(_0246_),
    .A1(_2453_));
 sg13g2_nor2_1 _3781_ (.A(_2399_),
    .B(_2404_),
    .Y(_0276_));
 sg13g2_xor2_1 _3782_ (.B(_2404_),
    .A(_2399_),
    .X(_0277_));
 sg13g2_xnor2_1 _3783_ (.Y(_0278_),
    .A(_2677_),
    .B(_0277_));
 sg13g2_nor2b_1 _3784_ (.A(_0275_),
    .B_N(_0278_),
    .Y(_0279_));
 sg13g2_xnor2_1 _3785_ (.Y(_0280_),
    .A(_0275_),
    .B(_0278_));
 sg13g2_a21oi_2 _3786_ (.B1(_0251_),
    .Y(_0281_),
    .A2(_0252_),
    .A1(net401));
 sg13g2_inv_1 _3787_ (.Y(_0282_),
    .A(_0281_));
 sg13g2_nand2_1 _3788_ (.Y(_0283_),
    .A(net402),
    .B(net400));
 sg13g2_xor2_1 _3789_ (.B(net400),
    .A(net402),
    .X(_0284_));
 sg13g2_o21ai_1 _3790_ (.B1(net399),
    .Y(_0285_),
    .A1(net402),
    .A2(net400));
 sg13g2_xnor2_1 _3791_ (.Y(_0286_),
    .A(\am_sdr0.det0.yn_1[19] ),
    .B(_0284_));
 sg13g2_inv_1 _3792_ (.Y(_0287_),
    .A(_0286_));
 sg13g2_nor2_1 _3793_ (.A(_2674_),
    .B(_0286_),
    .Y(_0288_));
 sg13g2_xor2_1 _3794_ (.B(_0286_),
    .A(_2674_),
    .X(_0289_));
 sg13g2_xnor2_1 _3795_ (.Y(_0290_),
    .A(_0281_),
    .B(_0289_));
 sg13g2_xnor2_1 _3796_ (.Y(_0291_),
    .A(_0280_),
    .B(_0290_));
 sg13g2_nand2b_1 _3797_ (.Y(_0292_),
    .B(_0274_),
    .A_N(_0291_));
 sg13g2_xor2_1 _3798_ (.B(_0291_),
    .A(_0274_),
    .X(_0293_));
 sg13g2_xor2_1 _3799_ (.B(_0293_),
    .A(_0273_),
    .X(_0294_));
 sg13g2_nand2_1 _3800_ (.Y(_0295_),
    .A(_0272_),
    .B(_0294_));
 sg13g2_xnor2_1 _3801_ (.Y(_0296_),
    .A(_0272_),
    .B(_0294_));
 sg13g2_a21oi_1 _3802_ (.A1(net399),
    .A2(_0264_),
    .Y(_0297_),
    .B1(_0263_));
 sg13g2_nor2_1 _3803_ (.A(_0296_),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_xnor2_1 _3804_ (.Y(_0299_),
    .A(_0296_),
    .B(_0297_));
 sg13g2_inv_1 _3805_ (.Y(_0300_),
    .A(_0299_));
 sg13g2_nor2_1 _3806_ (.A(_0233_),
    .B(_0267_),
    .Y(_0301_));
 sg13g2_a21oi_2 _3807_ (.B1(_0266_),
    .Y(_0302_),
    .A2(_0301_),
    .A1(_0236_));
 sg13g2_xnor2_1 _3808_ (.Y(_0303_),
    .A(_0299_),
    .B(_0302_));
 sg13g2_xnor2_1 _3809_ (.Y(_0304_),
    .A(_0300_),
    .B(_0302_));
 sg13g2_nand4_1 _3810_ (.B(_0238_),
    .C(_0270_),
    .A(_0207_),
    .Y(_0305_),
    .D(_0303_));
 sg13g2_nand2_1 _3811_ (.Y(_0306_),
    .A(net413),
    .B(_0305_));
 sg13g2_a21oi_1 _3812_ (.A1(_0271_),
    .A2(_0304_),
    .Y(_0098_),
    .B1(_0306_));
 sg13g2_a21o_1 _3813_ (.A2(net234),
    .A1(net406),
    .B1(_0098_),
    .X(_0080_));
 sg13g2_o21ai_1 _3814_ (.B1(_0292_),
    .Y(_0307_),
    .A1(_0273_),
    .A2(_0293_));
 sg13g2_a21oi_1 _3815_ (.A1(_0282_),
    .A2(_0289_),
    .Y(_0308_),
    .B1(_0288_));
 sg13g2_a21oi_1 _3816_ (.A1(_0280_),
    .A2(_0290_),
    .Y(_0309_),
    .B1(_0279_));
 sg13g2_a21oi_1 _3817_ (.A1(_2678_),
    .A2(_0277_),
    .Y(_0310_),
    .B1(_0276_));
 sg13g2_nor2_1 _3818_ (.A(_2423_),
    .B(_2429_),
    .Y(_0311_));
 sg13g2_xor2_1 _3819_ (.B(_2429_),
    .A(_2423_),
    .X(_0312_));
 sg13g2_xnor2_1 _3820_ (.Y(_0313_),
    .A(_0220_),
    .B(_0312_));
 sg13g2_nand2b_1 _3821_ (.Y(_0314_),
    .B(_0313_),
    .A_N(_0310_));
 sg13g2_xnor2_1 _3822_ (.Y(_0315_),
    .A(_0310_),
    .B(_0313_));
 sg13g2_inv_1 _3823_ (.Y(_0316_),
    .A(_0315_));
 sg13g2_nand2_2 _3824_ (.Y(_0317_),
    .A(_0283_),
    .B(_0285_));
 sg13g2_and2_1 _3825_ (.A(net400),
    .B(\am_sdr0.det0.yn_1[19] ),
    .X(_0318_));
 sg13g2_nor2_1 _3826_ (.A(net400),
    .B(\am_sdr0.det0.yn_1[19] ),
    .Y(_0319_));
 sg13g2_or2_2 _3827_ (.X(_0320_),
    .B(_0319_),
    .A(_0318_));
 sg13g2_inv_1 _3828_ (.Y(_0321_),
    .A(_0320_));
 sg13g2_nor2_1 _3829_ (.A(_0217_),
    .B(_0320_),
    .Y(_0322_));
 sg13g2_xor2_1 _3830_ (.B(_0320_),
    .A(_0217_),
    .X(_0323_));
 sg13g2_xnor2_1 _3831_ (.Y(_0324_),
    .A(_0317_),
    .B(_0323_));
 sg13g2_xor2_1 _3832_ (.B(_0324_),
    .A(_0315_),
    .X(_0325_));
 sg13g2_xor2_1 _3833_ (.B(_0325_),
    .A(_0309_),
    .X(_0326_));
 sg13g2_nand2b_1 _3834_ (.Y(_0327_),
    .B(_0326_),
    .A_N(_0308_));
 sg13g2_xnor2_1 _3835_ (.Y(_0328_),
    .A(_0308_),
    .B(_0326_));
 sg13g2_nand2_1 _3836_ (.Y(_0329_),
    .A(_0307_),
    .B(_0328_));
 sg13g2_xnor2_1 _3837_ (.Y(_0330_),
    .A(_0307_),
    .B(_0328_));
 sg13g2_nor2_1 _3838_ (.A(_0295_),
    .B(_0330_),
    .Y(_0331_));
 sg13g2_nand2_1 _3839_ (.Y(_0332_),
    .A(_0295_),
    .B(_0330_));
 sg13g2_nor2b_1 _3840_ (.A(_0331_),
    .B_N(_0332_),
    .Y(_0333_));
 sg13g2_a21oi_1 _3841_ (.A1(_0300_),
    .A2(_0302_),
    .Y(_0334_),
    .B1(_0298_));
 sg13g2_xnor2_1 _3842_ (.Y(_0335_),
    .A(_0333_),
    .B(_0334_));
 sg13g2_nand2b_1 _3843_ (.Y(_0336_),
    .B(_0305_),
    .A_N(_0335_));
 sg13g2_nand2b_2 _3844_ (.Y(_0337_),
    .B(_0335_),
    .A_N(_0305_));
 sg13g2_and3_1 _3845_ (.X(_0099_),
    .A(net417),
    .B(_0336_),
    .C(_0337_));
 sg13g2_a21o_1 _3846_ (.A2(net235),
    .A1(net406),
    .B1(_0099_),
    .X(_0081_));
 sg13g2_o21ai_1 _3847_ (.B1(_0327_),
    .Y(_0338_),
    .A1(_0309_),
    .A2(_0325_));
 sg13g2_a21oi_2 _3848_ (.B1(_0322_),
    .Y(_0339_),
    .A2(_0323_),
    .A1(_0317_));
 sg13g2_o21ai_1 _3849_ (.B1(_0314_),
    .Y(_0340_),
    .A1(_0316_),
    .A2(_0324_));
 sg13g2_a21oi_2 _3850_ (.B1(_0311_),
    .Y(_0341_),
    .A2(_0312_),
    .A1(_0221_));
 sg13g2_nor2_1 _3851_ (.A(_2449_),
    .B(_2452_),
    .Y(_0342_));
 sg13g2_xor2_1 _3852_ (.B(_2452_),
    .A(_2449_),
    .X(_0343_));
 sg13g2_xnor2_1 _3853_ (.Y(_0344_),
    .A(_0253_),
    .B(_0343_));
 sg13g2_nor2b_1 _3854_ (.A(_0341_),
    .B_N(_0344_),
    .Y(_0345_));
 sg13g2_xnor2_1 _3855_ (.Y(_0346_),
    .A(_0341_),
    .B(_0344_));
 sg13g2_nor2b_1 _3856_ (.A(net400),
    .B_N(net399),
    .Y(_0347_));
 sg13g2_xnor2_1 _3857_ (.Y(_0348_),
    .A(_0249_),
    .B(_0347_));
 sg13g2_xnor2_1 _3858_ (.Y(_0349_),
    .A(_0346_),
    .B(_0348_));
 sg13g2_nand2b_1 _3859_ (.Y(_0350_),
    .B(_0340_),
    .A_N(_0349_));
 sg13g2_xor2_1 _3860_ (.B(_0349_),
    .A(_0340_),
    .X(_0351_));
 sg13g2_xor2_1 _3861_ (.B(_0351_),
    .A(_0339_),
    .X(_0352_));
 sg13g2_nand2_1 _3862_ (.Y(_0353_),
    .A(_0338_),
    .B(_0352_));
 sg13g2_xnor2_1 _3863_ (.Y(_0354_),
    .A(_0338_),
    .B(_0352_));
 sg13g2_nor2_1 _3864_ (.A(_0329_),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_or2_1 _3865_ (.X(_0356_),
    .B(_0354_),
    .A(_0329_));
 sg13g2_xor2_1 _3866_ (.B(_0354_),
    .A(_0329_),
    .X(_0357_));
 sg13g2_inv_1 _3867_ (.Y(_0358_),
    .A(_0357_));
 sg13g2_nor2b_1 _3868_ (.A(_0299_),
    .B_N(_0333_),
    .Y(_0359_));
 sg13g2_a221oi_1 _3869_ (.B2(_0302_),
    .C1(_0331_),
    .B1(_0359_),
    .A1(_0298_),
    .Y(_0360_),
    .A2(_0332_));
 sg13g2_xnor2_1 _3870_ (.Y(_0361_),
    .A(_0358_),
    .B(_0360_));
 sg13g2_nand2_1 _3871_ (.Y(_0362_),
    .A(_0337_),
    .B(_0361_));
 sg13g2_nor2_1 _3872_ (.A(_0337_),
    .B(_0361_),
    .Y(_0363_));
 sg13g2_nand3b_1 _3873_ (.B(net417),
    .C(_0362_),
    .Y(_0364_),
    .A_N(_0363_));
 sg13g2_inv_1 _3874_ (.Y(_0100_),
    .A(_0364_));
 sg13g2_o21ai_1 _3875_ (.B1(_0364_),
    .Y(_0082_),
    .A1(net417),
    .A2(_2170_));
 sg13g2_o21ai_1 _3876_ (.B1(_0350_),
    .Y(_0365_),
    .A1(_0339_),
    .A2(_0351_));
 sg13g2_a21oi_1 _3877_ (.A1(_0346_),
    .A2(_0348_),
    .Y(_0366_),
    .B1(_0345_));
 sg13g2_a21oi_1 _3878_ (.A1(_0254_),
    .A2(_0343_),
    .Y(_0367_),
    .B1(_0342_));
 sg13g2_nor2_1 _3879_ (.A(_2674_),
    .B(_2677_),
    .Y(_0368_));
 sg13g2_xor2_1 _3880_ (.B(_2677_),
    .A(_2674_),
    .X(_0369_));
 sg13g2_xnor2_1 _3881_ (.Y(_0370_),
    .A(_0286_),
    .B(_0369_));
 sg13g2_nor2b_1 _3882_ (.A(_0367_),
    .B_N(_0370_),
    .Y(_0371_));
 sg13g2_xnor2_1 _3883_ (.Y(_0372_),
    .A(_0367_),
    .B(_0370_));
 sg13g2_xnor2_1 _3884_ (.Y(_0373_),
    .A(_0281_),
    .B(_0372_));
 sg13g2_nor2b_1 _3885_ (.A(_0366_),
    .B_N(_0373_),
    .Y(_0374_));
 sg13g2_xor2_1 _3886_ (.B(_0373_),
    .A(_0366_),
    .X(_0375_));
 sg13g2_o21ai_1 _3887_ (.B1(net399),
    .Y(_0376_),
    .A1(net400),
    .A2(_0250_));
 sg13g2_nor2_1 _3888_ (.A(_0375_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_xnor2_1 _3889_ (.Y(_0378_),
    .A(_0375_),
    .B(_0376_));
 sg13g2_nand2b_1 _3890_ (.Y(_0379_),
    .B(_0365_),
    .A_N(_0378_));
 sg13g2_xor2_1 _3891_ (.B(_0378_),
    .A(_0365_),
    .X(_0380_));
 sg13g2_nor2_1 _3892_ (.A(_0353_),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_xor2_1 _3893_ (.B(_0380_),
    .A(_0353_),
    .X(_0382_));
 sg13g2_o21ai_1 _3894_ (.B1(_0356_),
    .Y(_0383_),
    .A1(_0358_),
    .A2(_0360_));
 sg13g2_xnor2_1 _3895_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_o21ai_1 _3896_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_0337_),
    .A2(_0361_));
 sg13g2_or3_1 _3897_ (.A(_0337_),
    .B(_0361_),
    .C(_0384_),
    .X(_0386_));
 sg13g2_and3_1 _3898_ (.X(_0101_),
    .A(net417),
    .B(_0385_),
    .C(_0386_));
 sg13g2_a21o_1 _3899_ (.A2(net238),
    .A1(net408),
    .B1(_0101_),
    .X(_0083_));
 sg13g2_a21o_1 _3900_ (.A2(_0372_),
    .A1(_0282_),
    .B1(_0371_),
    .X(_0387_));
 sg13g2_a21oi_1 _3901_ (.A1(_0287_),
    .A2(_0369_),
    .Y(_0388_),
    .B1(_0368_));
 sg13g2_nor2_1 _3902_ (.A(_0217_),
    .B(_0220_),
    .Y(_0389_));
 sg13g2_xor2_1 _3903_ (.B(_0220_),
    .A(_0217_),
    .X(_0390_));
 sg13g2_xnor2_1 _3904_ (.Y(_0391_),
    .A(_0320_),
    .B(_0390_));
 sg13g2_nand2b_1 _3905_ (.Y(_0392_),
    .B(_0391_),
    .A_N(_0388_));
 sg13g2_xnor2_1 _3906_ (.Y(_0393_),
    .A(_0388_),
    .B(_0391_));
 sg13g2_nand2_1 _3907_ (.Y(_0394_),
    .A(_0317_),
    .B(_0393_));
 sg13g2_xnor2_1 _3908_ (.Y(_0395_),
    .A(_0317_),
    .B(_0393_));
 sg13g2_nand2b_1 _3909_ (.Y(_0396_),
    .B(_0387_),
    .A_N(_0395_));
 sg13g2_xor2_1 _3910_ (.B(_0395_),
    .A(_0387_),
    .X(_0397_));
 sg13g2_nor2_1 _3911_ (.A(_0374_),
    .B(_0377_),
    .Y(_0398_));
 sg13g2_or2_1 _3912_ (.X(_0399_),
    .B(_0398_),
    .A(_0397_));
 sg13g2_xnor2_1 _3913_ (.Y(_0400_),
    .A(_0397_),
    .B(_0398_));
 sg13g2_nor2_1 _3914_ (.A(_0379_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_xor2_1 _3915_ (.B(_0400_),
    .A(_0379_),
    .X(_0402_));
 sg13g2_nand2_1 _3916_ (.Y(_0403_),
    .A(_0357_),
    .B(_0382_));
 sg13g2_a21oi_1 _3917_ (.A1(_0355_),
    .A2(_0382_),
    .Y(_0404_),
    .B1(_0381_));
 sg13g2_o21ai_1 _3918_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0360_),
    .A2(_0403_));
 sg13g2_xnor2_1 _3919_ (.Y(_0406_),
    .A(_0402_),
    .B(_0405_));
 sg13g2_or4_1 _3920_ (.A(_0337_),
    .B(_0361_),
    .C(_0384_),
    .D(_0406_),
    .X(_0407_));
 sg13g2_nand2_1 _3921_ (.Y(_0408_),
    .A(net417),
    .B(_0407_));
 sg13g2_a21oi_1 _3922_ (.A1(_0386_),
    .A2(_0406_),
    .Y(_0102_),
    .B1(_0408_));
 sg13g2_a21o_1 _3923_ (.A2(net255),
    .A1(net408),
    .B1(_0102_),
    .X(_0084_));
 sg13g2_a21oi_1 _3924_ (.A1(_0402_),
    .A2(_0405_),
    .Y(_0409_),
    .B1(_0401_));
 sg13g2_and2_1 _3925_ (.A(_0392_),
    .B(_0394_),
    .X(_0410_));
 sg13g2_a21oi_1 _3926_ (.A1(_0321_),
    .A2(_0390_),
    .Y(_0411_),
    .B1(_0389_));
 sg13g2_nand2_2 _3927_ (.Y(_0412_),
    .A(_0250_),
    .B(_0254_));
 sg13g2_xor2_1 _3928_ (.B(_0253_),
    .A(_0249_),
    .X(_0413_));
 sg13g2_nand2_1 _3929_ (.Y(_0414_),
    .A(net399),
    .B(_0413_));
 sg13g2_xnor2_1 _3930_ (.Y(_0415_),
    .A(net399),
    .B(_0413_));
 sg13g2_nor2_1 _3931_ (.A(_0411_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_xor2_1 _3932_ (.B(_0415_),
    .A(_0411_),
    .X(_0417_));
 sg13g2_xor2_1 _3933_ (.B(_0417_),
    .A(_0318_),
    .X(_0418_));
 sg13g2_nor2b_1 _3934_ (.A(_0410_),
    .B_N(_0418_),
    .Y(_0419_));
 sg13g2_xnor2_1 _3935_ (.Y(_0420_),
    .A(_0410_),
    .B(_0418_));
 sg13g2_nand2b_1 _3936_ (.Y(_0421_),
    .B(_0420_),
    .A_N(_0396_));
 sg13g2_xnor2_1 _3937_ (.Y(_0422_),
    .A(_0396_),
    .B(_0420_));
 sg13g2_nand2b_1 _3938_ (.Y(_0423_),
    .B(_0422_),
    .A_N(_0399_));
 sg13g2_xor2_1 _3939_ (.B(_0422_),
    .A(_0399_),
    .X(_0424_));
 sg13g2_xnor2_1 _3940_ (.Y(_0425_),
    .A(_0409_),
    .B(_0424_));
 sg13g2_or2_1 _3941_ (.X(_0426_),
    .B(_0425_),
    .A(_0407_));
 sg13g2_nand2_1 _3942_ (.Y(_0427_),
    .A(net419),
    .B(_0426_));
 sg13g2_a21oi_1 _3943_ (.A1(_0407_),
    .A2(_0425_),
    .Y(_0103_),
    .B1(_0427_));
 sg13g2_a21o_1 _3944_ (.A2(net256),
    .A1(net407),
    .B1(_0103_),
    .X(_0085_));
 sg13g2_o21ai_1 _3945_ (.B1(_0423_),
    .Y(_0428_),
    .A1(_0409_),
    .A2(_0424_));
 sg13g2_xnor2_1 _3946_ (.Y(_0429_),
    .A(_0281_),
    .B(_0286_));
 sg13g2_a21oi_2 _3947_ (.B1(_0429_),
    .Y(_0430_),
    .A2(_0414_),
    .A1(_0412_));
 sg13g2_nand3_1 _3948_ (.B(_0414_),
    .C(_0429_),
    .A(_0412_),
    .Y(_0431_));
 sg13g2_nor2b_1 _3949_ (.A(_0430_),
    .B_N(_0431_),
    .Y(_0432_));
 sg13g2_a21oi_1 _3950_ (.A1(_0318_),
    .A2(_0417_),
    .Y(_0433_),
    .B1(_0416_));
 sg13g2_nand2b_1 _3951_ (.Y(_0434_),
    .B(_0432_),
    .A_N(_0433_));
 sg13g2_xnor2_1 _3952_ (.Y(_0435_),
    .A(_0432_),
    .B(_0433_));
 sg13g2_nor2b_1 _3953_ (.A(_0419_),
    .B_N(_0421_),
    .Y(_0436_));
 sg13g2_nor2b_1 _3954_ (.A(_0421_),
    .B_N(_0435_),
    .Y(_0437_));
 sg13g2_nand2_1 _3955_ (.Y(_0438_),
    .A(_0419_),
    .B(_0435_));
 sg13g2_xnor2_1 _3956_ (.Y(_0439_),
    .A(_0435_),
    .B(_0436_));
 sg13g2_xnor2_1 _3957_ (.Y(_0440_),
    .A(_0428_),
    .B(_0439_));
 sg13g2_and2_1 _3958_ (.A(_0426_),
    .B(_0440_),
    .X(_0441_));
 sg13g2_nor2_1 _3959_ (.A(_0426_),
    .B(_0440_),
    .Y(_0442_));
 sg13g2_nor3_1 _3960_ (.A(net407),
    .B(_0441_),
    .C(_0442_),
    .Y(_0104_));
 sg13g2_a21o_1 _3961_ (.A2(net248),
    .A1(net407),
    .B1(_0104_),
    .X(_0086_));
 sg13g2_a21oi_1 _3962_ (.A1(_0428_),
    .A2(_0439_),
    .Y(_0443_),
    .B1(_0437_));
 sg13g2_nand2b_1 _3963_ (.Y(_0444_),
    .B(net403),
    .A_N(net399));
 sg13g2_nor2_1 _3964_ (.A(net402),
    .B(_0319_),
    .Y(_0445_));
 sg13g2_a22oi_1 _3965_ (.Y(_0446_),
    .B1(_0444_),
    .B2(_0445_),
    .A2(_0319_),
    .A1(_0251_));
 sg13g2_nor2b_1 _3966_ (.A(_0446_),
    .B_N(_0430_),
    .Y(_0447_));
 sg13g2_xnor2_1 _3967_ (.Y(_0448_),
    .A(_0430_),
    .B(_0446_));
 sg13g2_nand2_1 _3968_ (.Y(_0449_),
    .A(_0434_),
    .B(_0438_));
 sg13g2_xor2_1 _3969_ (.B(_0449_),
    .A(_0448_),
    .X(_0450_));
 sg13g2_inv_1 _3970_ (.Y(_0451_),
    .A(_0450_));
 sg13g2_xnor2_1 _3971_ (.Y(_0452_),
    .A(_0443_),
    .B(_0450_));
 sg13g2_nand2_1 _3972_ (.Y(_0453_),
    .A(_0442_),
    .B(_0452_));
 sg13g2_o21ai_1 _3973_ (.B1(net419),
    .Y(_0454_),
    .A1(_0442_),
    .A2(_0452_));
 sg13g2_nor2b_1 _3974_ (.A(_0454_),
    .B_N(_0453_),
    .Y(_0105_));
 sg13g2_a21o_1 _3975_ (.A2(net262),
    .A1(net407),
    .B1(_0105_),
    .X(_0087_));
 sg13g2_nand2_1 _3976_ (.Y(_0455_),
    .A(net414),
    .B(_0189_));
 sg13g2_a21oi_1 _3977_ (.A1(_2173_),
    .A2(_0188_),
    .Y(_0088_),
    .B1(_0455_));
 sg13g2_o21ai_1 _3978_ (.B1(net414),
    .Y(_0456_),
    .A1(_0189_),
    .A2(_0191_));
 sg13g2_a21oi_1 _3979_ (.A1(_0189_),
    .A2(_0191_),
    .Y(_0089_),
    .B1(_0456_));
 sg13g2_o21ai_1 _3980_ (.B1(net414),
    .Y(_0457_),
    .A1(_0192_),
    .A2(_0193_));
 sg13g2_a21oi_1 _3981_ (.A1(_0192_),
    .A2(_0193_),
    .Y(_0090_),
    .B1(_0457_));
 sg13g2_o21ai_1 _3982_ (.B1(net414),
    .Y(_0458_),
    .A1(_0194_),
    .A2(_0196_));
 sg13g2_a21oi_1 _3983_ (.A1(_0194_),
    .A2(_0196_),
    .Y(_0091_),
    .B1(_0458_));
 sg13g2_o21ai_1 _3984_ (.B1(net414),
    .Y(_0459_),
    .A1(_0197_),
    .A2(_0199_));
 sg13g2_a21oi_1 _3985_ (.A1(_0197_),
    .A2(_0199_),
    .Y(_0092_),
    .B1(_0459_));
 sg13g2_o21ai_1 _3986_ (.B1(net414),
    .Y(_0460_),
    .A1(_0200_),
    .A2(_0201_));
 sg13g2_a21oi_1 _3987_ (.A1(_0200_),
    .A2(_0201_),
    .Y(_0093_),
    .B1(_0460_));
 sg13g2_o21ai_1 _3988_ (.B1(net414),
    .Y(_0461_),
    .A1(_0202_),
    .A2(_0204_));
 sg13g2_a21oi_1 _3989_ (.A1(_0202_),
    .A2(_0204_),
    .Y(_0094_),
    .B1(_0461_));
 sg13g2_o21ai_1 _3990_ (.B1(net413),
    .Y(_0462_),
    .A1(_0205_),
    .A2(_0206_));
 sg13g2_a21oi_1 _3991_ (.A1(_0205_),
    .A2(_0206_),
    .Y(_0095_),
    .B1(_0462_));
 sg13g2_o21ai_1 _3992_ (.B1(net413),
    .Y(_0463_),
    .A1(_0207_),
    .A2(_0238_));
 sg13g2_nor2_1 _3993_ (.A(_0239_),
    .B(_0463_),
    .Y(_0096_));
 sg13g2_or2_1 _3994_ (.X(_0464_),
    .B(_0270_),
    .A(_0239_));
 sg13g2_and3_1 _3995_ (.X(_0097_),
    .A(net413),
    .B(_0271_),
    .C(_0464_));
 sg13g2_nand3_1 _3996_ (.B(_0435_),
    .C(_0448_),
    .A(_0419_),
    .Y(_0465_));
 sg13g2_o21ai_1 _3997_ (.B1(_0465_),
    .Y(_0466_),
    .A1(_0443_),
    .A2(_0451_));
 sg13g2_nor2_1 _3998_ (.A(_0434_),
    .B(_0446_),
    .Y(_0467_));
 sg13g2_a21oi_1 _3999_ (.A1(_0284_),
    .A2(_0444_),
    .Y(_0468_),
    .B1(_0319_));
 sg13g2_xnor2_1 _4000_ (.Y(_0469_),
    .A(_0447_),
    .B(_0468_));
 sg13g2_xnor2_1 _4001_ (.Y(_0470_),
    .A(_0467_),
    .B(_0469_));
 sg13g2_xnor2_1 _4002_ (.Y(_0471_),
    .A(_0466_),
    .B(_0470_));
 sg13g2_or2_1 _4003_ (.X(_0472_),
    .B(_0471_),
    .A(_0453_));
 sg13g2_o21ai_1 _4004_ (.B1(net419),
    .Y(_0473_),
    .A1(_0453_),
    .A2(_0471_));
 sg13g2_a21oi_1 _4005_ (.A1(_0453_),
    .A2(_0471_),
    .Y(_0106_),
    .B1(_0473_));
 sg13g2_a21oi_1 _4006_ (.A1(_0467_),
    .A2(_0468_),
    .Y(_0474_),
    .B1(_0447_));
 sg13g2_nand2_1 _4007_ (.Y(_0475_),
    .A(_0285_),
    .B(_0474_));
 sg13g2_a21oi_1 _4008_ (.A1(_0466_),
    .A2(_0470_),
    .Y(_0476_),
    .B1(_0475_));
 sg13g2_a21oi_1 _4009_ (.A1(_0472_),
    .A2(_0476_),
    .Y(_0107_),
    .B1(net407));
 sg13g2_nor2_1 _4010_ (.A(\am_sdr0.filt0.gain_spi[1] ),
    .B(\am_sdr0.filt0.gain_spi[0] ),
    .Y(_0477_));
 sg13g2_and2_2 _4011_ (.A(net442),
    .B(_0477_),
    .X(_0478_));
 sg13g2_nand2_2 _4012_ (.Y(_0479_),
    .A(net398),
    .B(\am_sdr0.filt0.mul_a1[1] ));
 sg13g2_xor2_1 _4013_ (.B(\am_sdr0.filt0.mul_a1[1] ),
    .A(net398),
    .X(_0480_));
 sg13g2_xnor2_1 _4014_ (.Y(_0481_),
    .A(net398),
    .B(\am_sdr0.filt0.mul_a1[1] ));
 sg13g2_nand2_1 _4015_ (.Y(_0482_),
    .A(net397),
    .B(_0480_));
 sg13g2_xnor2_1 _4016_ (.Y(_0483_),
    .A(net397),
    .B(_0480_));
 sg13g2_and2_1 _4017_ (.A(\am_sdr0.filt0.yn_1[12] ),
    .B(net381),
    .X(_0484_));
 sg13g2_or2_1 _4018_ (.X(_0485_),
    .B(net381),
    .A(net382));
 sg13g2_nor2b_1 _4019_ (.A(_0484_),
    .B_N(_0485_),
    .Y(_0486_));
 sg13g2_nand2_1 _4020_ (.Y(_0487_),
    .A(net387),
    .B(_0486_));
 sg13g2_nor2_1 _4021_ (.A(_0030_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_nor2b_1 _4022_ (.A(_0030_),
    .B_N(_0484_),
    .Y(_0489_));
 sg13g2_nor2_1 _4023_ (.A(net381),
    .B(net383),
    .Y(_0490_));
 sg13g2_xnor2_1 _4024_ (.Y(_0491_),
    .A(net381),
    .B(net383));
 sg13g2_nand2_1 _4025_ (.Y(_0492_),
    .A(net384),
    .B(_0489_));
 sg13g2_o21ai_1 _4026_ (.B1(_0492_),
    .Y(_0493_),
    .A1(_0489_),
    .A2(_0491_));
 sg13g2_and2_1 _4027_ (.A(_0488_),
    .B(_0493_),
    .X(_0494_));
 sg13g2_xnor2_1 _4028_ (.Y(_0495_),
    .A(_0488_),
    .B(_0493_));
 sg13g2_nor2_1 _4029_ (.A(_0483_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_xor2_1 _4030_ (.B(_0495_),
    .A(_0483_),
    .X(_0497_));
 sg13g2_nand2_1 _4031_ (.Y(_0498_),
    .A(net384),
    .B(net389));
 sg13g2_xnor2_1 _4032_ (.Y(_0499_),
    .A(net387),
    .B(_0486_));
 sg13g2_a21oi_1 _4033_ (.A1(net387),
    .A2(_0485_),
    .Y(_0500_),
    .B1(_0484_));
 sg13g2_xnor2_1 _4034_ (.Y(_0501_),
    .A(_0030_),
    .B(_0500_));
 sg13g2_nor3_1 _4035_ (.A(_0498_),
    .B(_0499_),
    .C(_0501_),
    .Y(_0502_));
 sg13g2_o21ai_1 _4036_ (.B1(_0501_),
    .Y(_0503_),
    .A1(_0498_),
    .A2(_0499_));
 sg13g2_nand2b_1 _4037_ (.Y(_0504_),
    .B(_0503_),
    .A_N(_0502_));
 sg13g2_nor2_1 _4038_ (.A(_0481_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_o21ai_1 _4039_ (.B1(_0497_),
    .Y(_0506_),
    .A1(_0502_),
    .A2(_0505_));
 sg13g2_o21ai_1 _4040_ (.B1(\am_sdr0.filt0.yn_1[13] ),
    .Y(_0507_),
    .A1(net382),
    .A2(net384));
 sg13g2_a221oi_1 _4041_ (.B2(_0507_),
    .C1(_0489_),
    .B1(_0485_),
    .A1(net384),
    .Y(_0508_),
    .A2(_0484_));
 sg13g2_and2_1 _4042_ (.A(net396),
    .B(net397),
    .X(_0509_));
 sg13g2_and2_2 _4043_ (.A(_0480_),
    .B(_0509_),
    .X(_0510_));
 sg13g2_xor2_1 _4044_ (.B(net397),
    .A(net396),
    .X(_0511_));
 sg13g2_xnor2_1 _4045_ (.Y(_0512_),
    .A(_0480_),
    .B(_0511_));
 sg13g2_a21oi_1 _4046_ (.A1(_0482_),
    .A2(_0512_),
    .Y(_0513_),
    .B1(_0510_));
 sg13g2_nor2b_1 _4047_ (.A(_0508_),
    .B_N(_0513_),
    .Y(_0514_));
 sg13g2_xnor2_1 _4048_ (.Y(_0515_),
    .A(_0508_),
    .B(_0513_));
 sg13g2_o21ai_1 _4049_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_0494_),
    .A2(_0496_));
 sg13g2_or3_1 _4050_ (.A(_0494_),
    .B(_0496_),
    .C(_0515_),
    .X(_0517_));
 sg13g2_and2_1 _4051_ (.A(_0516_),
    .B(_0517_),
    .X(_0518_));
 sg13g2_nand2b_1 _4052_ (.Y(_0519_),
    .B(_0518_),
    .A_N(_0506_));
 sg13g2_xnor2_1 _4053_ (.Y(_0520_),
    .A(_0506_),
    .B(_0518_));
 sg13g2_nand2b_1 _4054_ (.Y(_0521_),
    .B(_0520_),
    .A_N(net342));
 sg13g2_nand3_1 _4055_ (.B(net396),
    .C(net397),
    .A(net395),
    .Y(_0522_));
 sg13g2_nor3_2 _4056_ (.A(net395),
    .B(net396),
    .C(net397),
    .Y(_0523_));
 sg13g2_a21o_1 _4057_ (.A2(_0509_),
    .A1(net395),
    .B1(_0523_),
    .X(_0524_));
 sg13g2_nand2_1 _4058_ (.Y(_0525_),
    .A(_0480_),
    .B(_0524_));
 sg13g2_o21ai_1 _4059_ (.B1(net395),
    .Y(_0526_),
    .A1(net396),
    .A2(net397));
 sg13g2_o21ai_1 _4060_ (.B1(_0526_),
    .Y(_0527_),
    .A1(_0481_),
    .A2(_0511_));
 sg13g2_o21ai_1 _4061_ (.B1(_0525_),
    .Y(_0528_),
    .A1(_0523_),
    .A2(_0527_));
 sg13g2_nand2b_1 _4062_ (.Y(_0529_),
    .B(_0528_),
    .A_N(_0507_));
 sg13g2_xnor2_1 _4063_ (.Y(_0530_),
    .A(_0507_),
    .B(_0528_));
 sg13g2_and2_1 _4064_ (.A(_0514_),
    .B(_0530_),
    .X(_0531_));
 sg13g2_xor2_1 _4065_ (.B(_0530_),
    .A(_0514_),
    .X(_0532_));
 sg13g2_xnor2_1 _4066_ (.Y(_0533_),
    .A(_0510_),
    .B(_0532_));
 sg13g2_nor2_1 _4067_ (.A(_0516_),
    .B(_0533_),
    .Y(_0534_));
 sg13g2_inv_1 _4068_ (.Y(_0535_),
    .A(_0534_));
 sg13g2_xor2_1 _4069_ (.B(_0533_),
    .A(_0516_),
    .X(_0536_));
 sg13g2_nand2b_1 _4070_ (.Y(_0537_),
    .B(_0536_),
    .A_N(net342));
 sg13g2_xor2_1 _4071_ (.B(_0536_),
    .A(net342),
    .X(_0538_));
 sg13g2_and3_1 _4072_ (.X(_0539_),
    .A(_0519_),
    .B(_0521_),
    .C(_0538_));
 sg13g2_inv_1 _4073_ (.Y(_0540_),
    .A(_0539_));
 sg13g2_a21oi_1 _4074_ (.A1(_0519_),
    .A2(_0521_),
    .Y(_0541_),
    .B1(_0538_));
 sg13g2_inv_1 _4075_ (.Y(_0542_),
    .A(_0541_));
 sg13g2_nand2_1 _4076_ (.Y(_0543_),
    .A(_0540_),
    .B(_0542_));
 sg13g2_xnor2_1 _4077_ (.Y(_0544_),
    .A(_0481_),
    .B(_0504_));
 sg13g2_nand2_1 _4078_ (.Y(_0545_),
    .A(\am_sdr0.filt0.yn_1[10] ),
    .B(net382));
 sg13g2_xnor2_1 _4079_ (.Y(_0546_),
    .A(net384),
    .B(net389));
 sg13g2_o21ai_1 _4080_ (.B1(_0498_),
    .Y(_0547_),
    .A1(_0545_),
    .A2(_0546_));
 sg13g2_xnor2_1 _4081_ (.Y(_0548_),
    .A(_0499_),
    .B(_0547_));
 sg13g2_nor3_1 _4082_ (.A(_0499_),
    .B(_0545_),
    .C(_0546_),
    .Y(_0549_));
 sg13g2_a21oi_1 _4083_ (.A1(net398),
    .A2(_0548_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_nor2_1 _4084_ (.A(_0544_),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_or3_1 _4085_ (.A(_0497_),
    .B(_0502_),
    .C(_0505_),
    .X(_0552_));
 sg13g2_and2_1 _4086_ (.A(_0506_),
    .B(_0552_),
    .X(_0553_));
 sg13g2_nand2_1 _4087_ (.Y(_0554_),
    .A(_0551_),
    .B(_0553_));
 sg13g2_xnor2_1 _4088_ (.Y(_0555_),
    .A(_0551_),
    .B(_0553_));
 sg13g2_or2_1 _4089_ (.X(_0556_),
    .B(_0555_),
    .A(_0479_));
 sg13g2_xor2_1 _4090_ (.B(_0520_),
    .A(net342),
    .X(_0557_));
 sg13g2_nand3_1 _4091_ (.B(_0556_),
    .C(_0557_),
    .A(_0554_),
    .Y(_0558_));
 sg13g2_and2_1 _4092_ (.A(net387),
    .B(net384),
    .X(_0559_));
 sg13g2_xor2_1 _4093_ (.B(net382),
    .A(\am_sdr0.filt0.yn_1[10] ),
    .X(_0560_));
 sg13g2_xor2_1 _4094_ (.B(_0560_),
    .A(_0559_),
    .X(_0561_));
 sg13g2_and2_1 _4095_ (.A(\am_sdr0.filt0.yn_1[7] ),
    .B(_0561_),
    .X(_0562_));
 sg13g2_xnor2_1 _4096_ (.Y(_0563_),
    .A(\am_sdr0.filt0.yn_1[7] ),
    .B(_0561_));
 sg13g2_nand3_1 _4097_ (.B(net389),
    .C(net392),
    .A(net385),
    .Y(_0564_));
 sg13g2_xnor2_1 _4098_ (.Y(_0565_),
    .A(net387),
    .B(net383));
 sg13g2_a21o_1 _4099_ (.A2(net389),
    .A1(net385),
    .B1(net392),
    .X(_0566_));
 sg13g2_nand2_1 _4100_ (.Y(_0567_),
    .A(_0564_),
    .B(_0566_));
 sg13g2_or2_1 _4101_ (.X(_0568_),
    .B(_0567_),
    .A(_0565_));
 sg13g2_a21o_1 _4102_ (.A2(_0568_),
    .A1(_0564_),
    .B1(_0563_),
    .X(_0569_));
 sg13g2_xor2_1 _4103_ (.B(_0546_),
    .A(_0545_),
    .X(_0570_));
 sg13g2_a21oi_1 _4104_ (.A1(_0559_),
    .A2(_0560_),
    .Y(_0571_),
    .B1(_0562_));
 sg13g2_nand2b_1 _4105_ (.Y(_0572_),
    .B(_0570_),
    .A_N(_0571_));
 sg13g2_xnor2_1 _4106_ (.Y(_0573_),
    .A(_0570_),
    .B(_0571_));
 sg13g2_nand2_1 _4107_ (.Y(_0574_),
    .A(net381),
    .B(_0573_));
 sg13g2_xnor2_1 _4108_ (.Y(_0575_),
    .A(net381),
    .B(_0573_));
 sg13g2_or2_1 _4109_ (.X(_0576_),
    .B(_0575_),
    .A(_0569_));
 sg13g2_xnor2_1 _4110_ (.Y(_0577_),
    .A(net398),
    .B(_0548_));
 sg13g2_a21oi_1 _4111_ (.A1(_0572_),
    .A2(_0574_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_nand3_1 _4112_ (.B(_0574_),
    .C(_0577_),
    .A(_0572_),
    .Y(_0579_));
 sg13g2_nand2b_1 _4113_ (.Y(_0580_),
    .B(_0579_),
    .A_N(_0578_));
 sg13g2_nor2_1 _4114_ (.A(_0576_),
    .B(_0580_),
    .Y(_0581_));
 sg13g2_xor2_1 _4115_ (.B(_0550_),
    .A(_0544_),
    .X(_0582_));
 sg13g2_nand2_1 _4116_ (.Y(_0583_),
    .A(_0578_),
    .B(_0582_));
 sg13g2_and2_1 _4117_ (.A(_0581_),
    .B(_0582_),
    .X(_0584_));
 sg13g2_xnor2_1 _4118_ (.Y(_0585_),
    .A(_0565_),
    .B(_0567_));
 sg13g2_xor2_1 _4119_ (.B(net389),
    .A(net385),
    .X(_0586_));
 sg13g2_nand2_1 _4120_ (.Y(_0587_),
    .A(net394),
    .B(_0586_));
 sg13g2_nor2_1 _4121_ (.A(_0585_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_inv_1 _4122_ (.Y(_0589_),
    .A(_0588_));
 sg13g2_nand3_1 _4123_ (.B(_0564_),
    .C(_0568_),
    .A(_0563_),
    .Y(_0590_));
 sg13g2_nand2_1 _4124_ (.Y(_0591_),
    .A(_0569_),
    .B(_0590_));
 sg13g2_nor2_1 _4125_ (.A(_0589_),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_xor2_1 _4126_ (.B(_0575_),
    .A(_0569_),
    .X(_0593_));
 sg13g2_nand2_1 _4127_ (.Y(_0594_),
    .A(_0592_),
    .B(_0593_));
 sg13g2_xnor2_1 _4128_ (.Y(_0595_),
    .A(_0576_),
    .B(_0580_));
 sg13g2_or2_1 _4129_ (.X(_0596_),
    .B(_0595_),
    .A(_0594_));
 sg13g2_xor2_1 _4130_ (.B(_0593_),
    .A(_0592_),
    .X(_0597_));
 sg13g2_inv_1 _4131_ (.Y(_0598_),
    .A(_0597_));
 sg13g2_xnor2_1 _4132_ (.Y(_0599_),
    .A(_0589_),
    .B(_0591_));
 sg13g2_nand2_1 _4133_ (.Y(_0600_),
    .A(net387),
    .B(\am_sdr0.filt0.yn_1[7] ));
 sg13g2_xnor2_1 _4134_ (.Y(_0601_),
    .A(net394),
    .B(_0586_));
 sg13g2_nor2_1 _4135_ (.A(_0600_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_xor2_1 _4136_ (.B(_0587_),
    .A(_0585_),
    .X(_0603_));
 sg13g2_nand2_1 _4137_ (.Y(_0604_),
    .A(_0602_),
    .B(_0603_));
 sg13g2_xnor2_1 _4138_ (.Y(_0605_),
    .A(_0602_),
    .B(_0603_));
 sg13g2_nand3_1 _4139_ (.B(net392),
    .C(net394),
    .A(net390),
    .Y(_0606_));
 sg13g2_a21o_2 _4140_ (.A2(net394),
    .A1(net390),
    .B1(net392),
    .X(_0607_));
 sg13g2_nand3_1 _4141_ (.B(_0606_),
    .C(_0607_),
    .A(net389),
    .Y(_0608_));
 sg13g2_xor2_1 _4142_ (.B(net390),
    .A(net387),
    .X(_0609_));
 sg13g2_nand2b_1 _4143_ (.Y(_0610_),
    .B(_0609_),
    .A_N(_0608_));
 sg13g2_nor2_2 _4144_ (.A(_2145_),
    .B(_0606_),
    .Y(_0611_));
 sg13g2_xnor2_1 _4145_ (.Y(_0612_),
    .A(_2145_),
    .B(_0606_));
 sg13g2_xor2_1 _4146_ (.B(_0609_),
    .A(_0608_),
    .X(_0613_));
 sg13g2_o21ai_1 _4147_ (.B1(_0610_),
    .Y(_0614_),
    .A1(_0612_),
    .A2(_0613_));
 sg13g2_xor2_1 _4148_ (.B(_0601_),
    .A(_0600_),
    .X(_0615_));
 sg13g2_and2_1 _4149_ (.A(_0614_),
    .B(_0615_),
    .X(_0616_));
 sg13g2_or2_1 _4150_ (.X(_0617_),
    .B(_0615_),
    .A(_0614_));
 sg13g2_xnor2_1 _4151_ (.Y(_0618_),
    .A(_0614_),
    .B(_0615_));
 sg13g2_a21oi_2 _4152_ (.B1(_0616_),
    .Y(_0619_),
    .A2(_0617_),
    .A1(_0611_));
 sg13g2_nor2_1 _4153_ (.A(_0605_),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_a21oi_1 _4154_ (.A1(_0602_),
    .A2(_0603_),
    .Y(_0621_),
    .B1(_0620_));
 sg13g2_nor2_1 _4155_ (.A(_0599_),
    .B(_0604_),
    .Y(_0622_));
 sg13g2_nor3_1 _4156_ (.A(_0599_),
    .B(_0605_),
    .C(_0619_),
    .Y(_0623_));
 sg13g2_xnor2_1 _4157_ (.Y(_0624_),
    .A(_0599_),
    .B(_0621_));
 sg13g2_a21o_1 _4158_ (.A2(_0607_),
    .A1(_0606_),
    .B1(net388),
    .X(_0625_));
 sg13g2_and2_1 _4159_ (.A(_0608_),
    .B(_0625_),
    .X(_0626_));
 sg13g2_xor2_1 _4160_ (.B(_0613_),
    .A(_0612_),
    .X(_0627_));
 sg13g2_and3_1 _4161_ (.X(_0628_),
    .A(net396),
    .B(_0626_),
    .C(_0627_));
 sg13g2_xnor2_1 _4162_ (.Y(_0629_),
    .A(_0611_),
    .B(_0618_));
 sg13g2_and2_1 _4163_ (.A(_0628_),
    .B(_0629_),
    .X(_0630_));
 sg13g2_xor2_1 _4164_ (.B(_0619_),
    .A(_0605_),
    .X(_0631_));
 sg13g2_nor2_1 _4165_ (.A(_0630_),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_or2_1 _4166_ (.X(_0633_),
    .B(_0631_),
    .A(_0630_));
 sg13g2_and2_1 _4167_ (.A(_0630_),
    .B(_0631_),
    .X(_0634_));
 sg13g2_nand2_1 _4168_ (.Y(_0635_),
    .A(\am_sdr0.filt0.mul_a1[1] ),
    .B(\am_sdr0.filt0.yn_1[4] ));
 sg13g2_xnor2_1 _4169_ (.Y(_0636_),
    .A(_2146_),
    .B(_0635_));
 sg13g2_inv_1 _4170_ (.Y(_0637_),
    .A(_0636_));
 sg13g2_or2_1 _4171_ (.X(_0638_),
    .B(net393),
    .A(net390));
 sg13g2_xor2_1 _4172_ (.B(net394),
    .A(net390),
    .X(_0639_));
 sg13g2_nand2b_1 _4173_ (.Y(_0640_),
    .B(_0639_),
    .A_N(_0636_));
 sg13g2_o21ai_1 _4174_ (.B1(_0640_),
    .Y(_0641_),
    .A1(_2146_),
    .A2(_0635_));
 sg13g2_xnor2_1 _4175_ (.Y(_0642_),
    .A(\am_sdr0.filt0.yn_1[3] ),
    .B(_0626_));
 sg13g2_nor2b_1 _4176_ (.A(_0642_),
    .B_N(_0641_),
    .Y(_0643_));
 sg13g2_and2_1 _4177_ (.A(_0627_),
    .B(_0643_),
    .X(_0644_));
 sg13g2_inv_1 _4178_ (.Y(_0645_),
    .A(_0644_));
 sg13g2_xnor2_1 _4179_ (.Y(_0646_),
    .A(_0628_),
    .B(_0629_));
 sg13g2_nor2_1 _4180_ (.A(_0645_),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_xnor2_1 _4181_ (.Y(_0648_),
    .A(_0644_),
    .B(_0646_));
 sg13g2_xnor2_1 _4182_ (.Y(_0649_),
    .A(_0645_),
    .B(_0646_));
 sg13g2_a21o_1 _4183_ (.A2(net397),
    .A1(\am_sdr0.filt0.yn_1[4] ),
    .B1(net396),
    .X(_0650_));
 sg13g2_nand2_1 _4184_ (.Y(_0651_),
    .A(_0522_),
    .B(_0650_));
 sg13g2_a22oi_1 _4185_ (.Y(_0652_),
    .B1(_0650_),
    .B2(net398),
    .A2(_0509_),
    .A1(net395));
 sg13g2_xor2_1 _4186_ (.B(net395),
    .A(\am_sdr0.filt0.mul_a1[1] ),
    .X(_0653_));
 sg13g2_nand2b_1 _4187_ (.Y(_0654_),
    .B(_0653_),
    .A_N(_0652_));
 sg13g2_xnor2_1 _4188_ (.Y(_0655_),
    .A(_0636_),
    .B(_0639_));
 sg13g2_nand2b_2 _4189_ (.Y(_0656_),
    .B(_0655_),
    .A_N(_0654_));
 sg13g2_inv_1 _4190_ (.Y(_0657_),
    .A(_0656_));
 sg13g2_xnor2_1 _4191_ (.Y(_0658_),
    .A(_0652_),
    .B(_0653_));
 sg13g2_and3_1 _4192_ (.X(_0659_),
    .A(net392),
    .B(_0655_),
    .C(_0658_));
 sg13g2_nand3_1 _4193_ (.B(_0655_),
    .C(_0658_),
    .A(net392),
    .Y(_0660_));
 sg13g2_nand2_1 _4194_ (.Y(_0661_),
    .A(_0656_),
    .B(_0660_));
 sg13g2_xor2_1 _4195_ (.B(_0642_),
    .A(_0641_),
    .X(_0662_));
 sg13g2_nor2b_1 _4196_ (.A(_0662_),
    .B_N(_0661_),
    .Y(_0663_));
 sg13g2_a21oi_1 _4197_ (.A1(\am_sdr0.filt0.yn_1[3] ),
    .A2(_0626_),
    .Y(_0664_),
    .B1(_0643_));
 sg13g2_xnor2_1 _4198_ (.Y(_0665_),
    .A(_0627_),
    .B(_0664_));
 sg13g2_a21oi_1 _4199_ (.A1(net392),
    .A2(_0658_),
    .Y(_0666_),
    .B1(_0655_));
 sg13g2_or2_1 _4200_ (.X(_0667_),
    .B(_0666_),
    .A(_0659_));
 sg13g2_o21ai_1 _4201_ (.B1(_0654_),
    .Y(_0668_),
    .A1(_0659_),
    .A2(_0666_));
 sg13g2_xnor2_1 _4202_ (.Y(_0669_),
    .A(net392),
    .B(_0658_));
 sg13g2_xnor2_1 _4203_ (.Y(_0670_),
    .A(net398),
    .B(_0651_));
 sg13g2_and2_1 _4204_ (.A(net393),
    .B(_0670_),
    .X(_0671_));
 sg13g2_nor2b_1 _4205_ (.A(_0669_),
    .B_N(_0671_),
    .Y(_0672_));
 sg13g2_nand2b_1 _4206_ (.Y(_0673_),
    .B(_0671_),
    .A_N(_0669_));
 sg13g2_nand3_1 _4207_ (.B(_0668_),
    .C(_0672_),
    .A(_0656_),
    .Y(_0674_));
 sg13g2_xor2_1 _4208_ (.B(_0662_),
    .A(_0661_),
    .X(_0675_));
 sg13g2_nor2_1 _4209_ (.A(_0674_),
    .B(_0675_),
    .Y(_0676_));
 sg13g2_o21ai_1 _4210_ (.B1(_0665_),
    .Y(_0677_),
    .A1(_0663_),
    .A2(_0676_));
 sg13g2_xor2_1 _4211_ (.B(_0665_),
    .A(_0663_),
    .X(_0678_));
 sg13g2_xnor2_1 _4212_ (.Y(_0679_),
    .A(_0669_),
    .B(_0671_));
 sg13g2_nor2_1 _4213_ (.A(net393),
    .B(_0670_),
    .Y(_0680_));
 sg13g2_xnor2_1 _4214_ (.Y(_0681_),
    .A(net393),
    .B(_0670_));
 sg13g2_nand3_1 _4215_ (.B(\am_sdr0.filt0.yn_1[3] ),
    .C(_0637_),
    .A(\am_sdr0.filt0.mul_a1[1] ),
    .Y(_0682_));
 sg13g2_nor2_1 _4216_ (.A(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_or4_1 _4217_ (.A(_0669_),
    .B(_0671_),
    .C(_0680_),
    .D(_0682_),
    .X(_0684_));
 sg13g2_nand4_1 _4218_ (.B(_0668_),
    .C(_0679_),
    .A(_0656_),
    .Y(_0685_),
    .D(_0683_));
 sg13g2_nand3_1 _4219_ (.B(_2145_),
    .C(\am_sdr0.filt0.yn_1[2] ),
    .A(net398),
    .Y(_0686_));
 sg13g2_or3_1 _4220_ (.A(_0512_),
    .B(_0681_),
    .C(_0686_),
    .X(_0687_));
 sg13g2_xnor2_1 _4221_ (.Y(_0688_),
    .A(_0679_),
    .B(_0683_));
 sg13g2_or2_1 _4222_ (.X(_0689_),
    .B(_0688_),
    .A(_0687_));
 sg13g2_a221oi_1 _4223_ (.B2(_0683_),
    .C1(_0672_),
    .B1(_0679_),
    .A1(_0656_),
    .Y(_0690_),
    .A2(_0668_));
 sg13g2_a221oi_1 _4224_ (.B2(_0684_),
    .C1(_0657_),
    .B1(_0673_),
    .A1(_0654_),
    .Y(_0691_),
    .A2(_0667_));
 sg13g2_or4_1 _4225_ (.A(_0687_),
    .B(_0688_),
    .C(_0690_),
    .D(_0691_),
    .X(_0692_));
 sg13g2_nand2_1 _4226_ (.Y(_0693_),
    .A(_0685_),
    .B(_0692_));
 sg13g2_xnor2_1 _4227_ (.Y(_0694_),
    .A(_0674_),
    .B(_0675_));
 sg13g2_a21oi_1 _4228_ (.A1(_0685_),
    .A2(_0692_),
    .Y(_0695_),
    .B1(_0694_));
 sg13g2_nand2_1 _4229_ (.Y(_0696_),
    .A(_0678_),
    .B(_0695_));
 sg13g2_a21oi_1 _4230_ (.A1(_0677_),
    .A2(_0696_),
    .Y(_0697_),
    .B1(_0649_));
 sg13g2_nor2_1 _4231_ (.A(_0647_),
    .B(_0697_),
    .Y(_0698_));
 sg13g2_a21o_1 _4232_ (.A2(_0647_),
    .A1(_0633_),
    .B1(_0634_),
    .X(_0699_));
 sg13g2_xor2_1 _4233_ (.B(_0631_),
    .A(_0630_),
    .X(_0700_));
 sg13g2_nor4_1 _4234_ (.A(_0632_),
    .B(_0634_),
    .C(_0649_),
    .D(_0677_),
    .Y(_0701_));
 sg13g2_and4_1 _4235_ (.A(_0648_),
    .B(_0678_),
    .C(_0695_),
    .D(_0700_),
    .X(_0702_));
 sg13g2_nor3_2 _4236_ (.A(_0699_),
    .B(_0701_),
    .C(_0702_),
    .Y(_0703_));
 sg13g2_nor2_1 _4237_ (.A(_0624_),
    .B(_0703_),
    .Y(_0704_));
 sg13g2_nor3_1 _4238_ (.A(_0598_),
    .B(_0624_),
    .C(_0703_),
    .Y(_0705_));
 sg13g2_and2_1 _4239_ (.A(_0597_),
    .B(_0622_),
    .X(_0706_));
 sg13g2_nor2_1 _4240_ (.A(_0597_),
    .B(_0622_),
    .Y(_0707_));
 sg13g2_nor2_1 _4241_ (.A(_0623_),
    .B(_0706_),
    .Y(_0708_));
 sg13g2_nor2_1 _4242_ (.A(_0707_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_nor2_1 _4243_ (.A(_0705_),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_xnor2_1 _4244_ (.Y(_0711_),
    .A(_0594_),
    .B(_0595_));
 sg13g2_inv_1 _4245_ (.Y(_0712_),
    .A(_0711_));
 sg13g2_o21ai_1 _4246_ (.B1(_0712_),
    .Y(_0713_),
    .A1(_0705_),
    .A2(_0709_));
 sg13g2_nor2_1 _4247_ (.A(_0578_),
    .B(_0581_),
    .Y(_0714_));
 sg13g2_xor2_1 _4248_ (.B(_0714_),
    .A(_0582_),
    .X(_0715_));
 sg13g2_a21oi_2 _4249_ (.B1(_0715_),
    .Y(_0716_),
    .A2(_0713_),
    .A1(_0596_));
 sg13g2_xor2_1 _4250_ (.B(_0555_),
    .A(net342),
    .X(_0717_));
 sg13g2_nor2b_1 _4251_ (.A(_0583_),
    .B_N(_0717_),
    .Y(_0718_));
 sg13g2_xnor2_1 _4252_ (.Y(_0719_),
    .A(_0583_),
    .B(_0717_));
 sg13g2_o21ai_1 _4253_ (.B1(_0719_),
    .Y(_0720_),
    .A1(_0584_),
    .A2(_0716_));
 sg13g2_a21o_1 _4254_ (.A2(_0556_),
    .A1(_0554_),
    .B1(_0557_),
    .X(_0721_));
 sg13g2_inv_1 _4255_ (.Y(_0722_),
    .A(_0721_));
 sg13g2_nand2_1 _4256_ (.Y(_0723_),
    .A(_0558_),
    .B(_0721_));
 sg13g2_and3_1 _4257_ (.X(_0724_),
    .A(_0558_),
    .B(_0719_),
    .C(_0721_));
 sg13g2_o21ai_1 _4258_ (.B1(_0724_),
    .Y(_0725_),
    .A1(_0584_),
    .A2(_0716_));
 sg13g2_a21oi_2 _4259_ (.B1(_0722_),
    .Y(_0726_),
    .A2(_0718_),
    .A1(_0558_));
 sg13g2_a21o_1 _4260_ (.A2(_0726_),
    .A1(_0725_),
    .B1(_0543_),
    .X(_0727_));
 sg13g2_nand3_1 _4261_ (.B(_0725_),
    .C(_0726_),
    .A(_0543_),
    .Y(_0728_));
 sg13g2_and2_1 _4262_ (.A(_0727_),
    .B(_0728_),
    .X(_0729_));
 sg13g2_and2_1 _4263_ (.A(net367),
    .B(net370),
    .X(_0730_));
 sg13g2_xor2_1 _4264_ (.B(net370),
    .A(net367),
    .X(_0731_));
 sg13g2_a21oi_2 _4265_ (.B1(_0730_),
    .Y(_0732_),
    .A2(_0731_),
    .A1(net365));
 sg13g2_nand2_1 _4266_ (.Y(_0733_),
    .A(net361),
    .B(net355));
 sg13g2_nor2_1 _4267_ (.A(net360),
    .B(net354),
    .Y(_0734_));
 sg13g2_xnor2_1 _4268_ (.Y(_0735_),
    .A(net361),
    .B(net354));
 sg13g2_xnor2_1 _4269_ (.Y(_0736_),
    .A(_2151_),
    .B(_0735_));
 sg13g2_or2_1 _4270_ (.X(_0737_),
    .B(_0736_),
    .A(_0732_));
 sg13g2_and2_1 _4271_ (.A(net360),
    .B(net363),
    .X(_0738_));
 sg13g2_xor2_1 _4272_ (.B(net363),
    .A(net360),
    .X(_0739_));
 sg13g2_a21oi_2 _4273_ (.B1(_0738_),
    .Y(_0740_),
    .A2(_0739_),
    .A1(net358));
 sg13g2_xnor2_1 _4274_ (.Y(_0741_),
    .A(_0732_),
    .B(_0736_));
 sg13g2_o21ai_1 _4275_ (.B1(_0737_),
    .Y(_0742_),
    .A1(_0740_),
    .A2(_0741_));
 sg13g2_nor2b_1 _4276_ (.A(net353),
    .B_N(net351),
    .Y(_0743_));
 sg13g2_nand2_1 _4277_ (.Y(_0744_),
    .A(_0742_),
    .B(_0743_));
 sg13g2_and2_1 _4278_ (.A(net351),
    .B(net352),
    .X(_0745_));
 sg13g2_nand2_1 _4279_ (.Y(_0746_),
    .A(net351),
    .B(net353));
 sg13g2_and2_1 _4280_ (.A(net349),
    .B(net354),
    .X(_0747_));
 sg13g2_a22oi_1 _4281_ (.Y(_0748_),
    .B1(_0745_),
    .B2(net354),
    .A2(_2159_),
    .A1(_2154_));
 sg13g2_xnor2_1 _4282_ (.Y(_0749_),
    .A(_0742_),
    .B(_0743_));
 sg13g2_o21ai_1 _4283_ (.B1(_0744_),
    .Y(_0750_),
    .A1(_0748_),
    .A2(_0749_));
 sg13g2_xnor2_1 _4284_ (.Y(_0751_),
    .A(net366),
    .B(_0731_));
 sg13g2_inv_1 _4285_ (.Y(_0752_),
    .A(_0751_));
 sg13g2_nand2_1 _4286_ (.Y(_0753_),
    .A(net371),
    .B(net376));
 sg13g2_nor2_1 _4287_ (.A(net371),
    .B(net376),
    .Y(_0754_));
 sg13g2_xor2_1 _4288_ (.B(net375),
    .A(net371),
    .X(_0755_));
 sg13g2_xnor2_1 _4289_ (.Y(_0756_),
    .A(net372),
    .B(net375));
 sg13g2_mux2_1 _4290_ (.A0(net372),
    .A1(_0756_),
    .S(net373),
    .X(_0757_));
 sg13g2_nand2_1 _4291_ (.Y(_0758_),
    .A(net373),
    .B(net375));
 sg13g2_nor2_1 _4292_ (.A(net372),
    .B(_0758_),
    .Y(_0759_));
 sg13g2_a21oi_1 _4293_ (.A1(_0752_),
    .A2(_0757_),
    .Y(_0760_),
    .B1(_0759_));
 sg13g2_and2_1 _4294_ (.A(net367),
    .B(net365),
    .X(_0761_));
 sg13g2_xor2_1 _4295_ (.B(net365),
    .A(net367),
    .X(_0762_));
 sg13g2_xor2_1 _4296_ (.B(_0762_),
    .A(net363),
    .X(_0763_));
 sg13g2_nand2_1 _4297_ (.Y(_0764_),
    .A(net372),
    .B(net373));
 sg13g2_nor2_1 _4298_ (.A(net370),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_and2_1 _4299_ (.A(net372),
    .B(net370),
    .X(_0766_));
 sg13g2_xor2_1 _4300_ (.B(net370),
    .A(net372),
    .X(_0767_));
 sg13g2_a21oi_1 _4301_ (.A1(net372),
    .A2(net373),
    .Y(_0768_),
    .B1(_0767_));
 sg13g2_nor2_1 _4302_ (.A(_0765_),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_xor2_1 _4303_ (.B(_0769_),
    .A(_0763_),
    .X(_0770_));
 sg13g2_nor2b_1 _4304_ (.A(_0760_),
    .B_N(_0770_),
    .Y(_0771_));
 sg13g2_xor2_1 _4305_ (.B(_0741_),
    .A(_0740_),
    .X(_0772_));
 sg13g2_xnor2_1 _4306_ (.Y(_0773_),
    .A(_0760_),
    .B(_0770_));
 sg13g2_a21oi_1 _4307_ (.A1(_0772_),
    .A2(_0773_),
    .Y(_0774_),
    .B1(_0771_));
 sg13g2_a21oi_1 _4308_ (.A1(_0763_),
    .A2(_0769_),
    .Y(_0775_),
    .B1(_0765_));
 sg13g2_and2_1 _4309_ (.A(net365),
    .B(net363),
    .X(_0776_));
 sg13g2_xor2_1 _4310_ (.B(net363),
    .A(net365),
    .X(_0777_));
 sg13g2_xnor2_1 _4311_ (.Y(_0778_),
    .A(_2150_),
    .B(_0777_));
 sg13g2_xnor2_1 _4312_ (.Y(_0779_),
    .A(net360),
    .B(_0777_));
 sg13g2_mux2_1 _4313_ (.A0(_0731_),
    .A1(net367),
    .S(_0766_),
    .X(_0780_));
 sg13g2_xnor2_1 _4314_ (.Y(_0781_),
    .A(_0779_),
    .B(_0780_));
 sg13g2_nor2b_1 _4315_ (.A(_0775_),
    .B_N(_0781_),
    .Y(_0782_));
 sg13g2_xnor2_1 _4316_ (.Y(_0783_),
    .A(_0775_),
    .B(_0781_));
 sg13g2_a21oi_1 _4317_ (.A1(net360),
    .A2(net355),
    .Y(_0784_),
    .B1(net358));
 sg13g2_nor2_1 _4318_ (.A(_2150_),
    .B(_2151_),
    .Y(_0785_));
 sg13g2_nor2_2 _4319_ (.A(_0734_),
    .B(_0784_),
    .Y(_0786_));
 sg13g2_a21oi_2 _4320_ (.B1(_0761_),
    .Y(_0787_),
    .A2(_0762_),
    .A1(net363));
 sg13g2_xnor2_1 _4321_ (.Y(_0788_),
    .A(net357),
    .B(net352));
 sg13g2_nand2_1 _4322_ (.Y(_0789_),
    .A(net354),
    .B(_0788_));
 sg13g2_xnor2_1 _4323_ (.Y(_0790_),
    .A(net355),
    .B(_0788_));
 sg13g2_nor2b_1 _4324_ (.A(_0787_),
    .B_N(_0790_),
    .Y(_0791_));
 sg13g2_xor2_1 _4325_ (.B(_0790_),
    .A(_0787_),
    .X(_0792_));
 sg13g2_nor3_1 _4326_ (.A(_0734_),
    .B(_0784_),
    .C(_0792_),
    .Y(_0793_));
 sg13g2_xnor2_1 _4327_ (.Y(_0794_),
    .A(_0786_),
    .B(_0792_));
 sg13g2_xnor2_1 _4328_ (.Y(_0795_),
    .A(_0783_),
    .B(_0794_));
 sg13g2_nor2_1 _4329_ (.A(_0774_),
    .B(_0795_),
    .Y(_0796_));
 sg13g2_xor2_1 _4330_ (.B(_0795_),
    .A(_0774_),
    .X(_0797_));
 sg13g2_xor2_1 _4331_ (.B(_0749_),
    .A(_0748_),
    .X(_0798_));
 sg13g2_a21oi_1 _4332_ (.A1(_0797_),
    .A2(_0798_),
    .Y(_0799_),
    .B1(_0796_));
 sg13g2_nor2_2 _4333_ (.A(_0791_),
    .B(_0793_),
    .Y(_0800_));
 sg13g2_nor2_1 _4334_ (.A(_0746_),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_xnor2_1 _4335_ (.Y(_0802_),
    .A(_0746_),
    .B(_0800_));
 sg13g2_a21oi_1 _4336_ (.A1(_0783_),
    .A2(_0794_),
    .Y(_0803_),
    .B1(_0782_));
 sg13g2_a22oi_1 _4337_ (.Y(_0804_),
    .B1(_0778_),
    .B2(_0780_),
    .A2(_0766_),
    .A1(_2148_));
 sg13g2_xnor2_1 _4338_ (.Y(_0805_),
    .A(net357),
    .B(_0739_));
 sg13g2_mux2_1 _4339_ (.A0(_0762_),
    .A1(net365),
    .S(_0730_),
    .X(_0806_));
 sg13g2_nor2b_1 _4340_ (.A(_0805_),
    .B_N(_0806_),
    .Y(_0807_));
 sg13g2_xnor2_1 _4341_ (.Y(_0808_),
    .A(_0805_),
    .B(_0806_));
 sg13g2_nor2b_1 _4342_ (.A(_0804_),
    .B_N(_0808_),
    .Y(_0809_));
 sg13g2_xnor2_1 _4343_ (.Y(_0810_),
    .A(_0804_),
    .B(_0808_));
 sg13g2_a21oi_2 _4344_ (.B1(_0776_),
    .Y(_0811_),
    .A2(_0777_),
    .A1(net360));
 sg13g2_nor2_1 _4345_ (.A(_2153_),
    .B(_2154_),
    .Y(_0812_));
 sg13g2_xor2_1 _4346_ (.B(net353),
    .A(net355),
    .X(_0813_));
 sg13g2_nor2_1 _4347_ (.A(net349),
    .B(_0812_),
    .Y(_0814_));
 sg13g2_xnor2_1 _4348_ (.Y(_0815_),
    .A(net350),
    .B(_0813_));
 sg13g2_nor2_1 _4349_ (.A(_0811_),
    .B(_0815_),
    .Y(_0816_));
 sg13g2_xnor2_1 _4350_ (.Y(_0817_),
    .A(_0811_),
    .B(_0815_));
 sg13g2_nor2_1 _4351_ (.A(net357),
    .B(_0812_),
    .Y(_0818_));
 sg13g2_a21oi_2 _4352_ (.B1(_0818_),
    .Y(_0819_),
    .A2(_2154_),
    .A1(_2153_));
 sg13g2_nor2b_1 _4353_ (.A(_0817_),
    .B_N(_0819_),
    .Y(_0820_));
 sg13g2_xnor2_1 _4354_ (.Y(_0821_),
    .A(_0817_),
    .B(_0819_));
 sg13g2_xnor2_1 _4355_ (.Y(_0822_),
    .A(_0810_),
    .B(_0821_));
 sg13g2_nor2_1 _4356_ (.A(_0803_),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_xor2_1 _4357_ (.B(_0822_),
    .A(_0803_),
    .X(_0824_));
 sg13g2_nor2b_1 _4358_ (.A(_0802_),
    .B_N(_0824_),
    .Y(_0825_));
 sg13g2_xnor2_1 _4359_ (.Y(_0826_),
    .A(_0802_),
    .B(_0824_));
 sg13g2_nand2b_1 _4360_ (.Y(_0827_),
    .B(_0826_),
    .A_N(_0799_));
 sg13g2_xnor2_1 _4361_ (.Y(_0828_),
    .A(_0799_),
    .B(_0826_));
 sg13g2_nand2_1 _4362_ (.Y(_0829_),
    .A(_0750_),
    .B(_0828_));
 sg13g2_xnor2_1 _4363_ (.Y(_0830_),
    .A(_0750_),
    .B(_0828_));
 sg13g2_xor2_1 _4364_ (.B(_0757_),
    .A(_0751_),
    .X(_0831_));
 sg13g2_xnor2_1 _4365_ (.Y(_0832_),
    .A(_2148_),
    .B(_0767_));
 sg13g2_nand2_1 _4366_ (.Y(_0833_),
    .A(net374),
    .B(net377));
 sg13g2_xnor2_1 _4367_ (.Y(_0834_),
    .A(net374),
    .B(net377));
 sg13g2_nand2b_1 _4368_ (.Y(_0835_),
    .B(net374),
    .A_N(net376));
 sg13g2_mux2_1 _4369_ (.A0(net373),
    .A1(_0834_),
    .S(net375),
    .X(_0836_));
 sg13g2_nand2_2 _4370_ (.Y(_0837_),
    .A(net375),
    .B(net377));
 sg13g2_nor2_1 _4371_ (.A(net373),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_a21oi_1 _4372_ (.A1(_0832_),
    .A2(_0836_),
    .Y(_0839_),
    .B1(_0838_));
 sg13g2_nor2_1 _4373_ (.A(_0831_),
    .B(_0839_),
    .Y(_0840_));
 sg13g2_a21oi_2 _4374_ (.B1(_0766_),
    .Y(_0841_),
    .A2(_0767_),
    .A1(net367));
 sg13g2_inv_1 _4375_ (.Y(_0842_),
    .A(_0841_));
 sg13g2_or2_1 _4376_ (.X(_0843_),
    .B(_0841_),
    .A(_0805_));
 sg13g2_xnor2_1 _4377_ (.Y(_0844_),
    .A(_0805_),
    .B(_0841_));
 sg13g2_xnor2_1 _4378_ (.Y(_0845_),
    .A(_0811_),
    .B(_0844_));
 sg13g2_xnor2_1 _4379_ (.Y(_0846_),
    .A(_0831_),
    .B(_0839_));
 sg13g2_nor2_1 _4380_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_nor2_1 _4381_ (.A(_0840_),
    .B(_0847_),
    .Y(_0848_));
 sg13g2_xnor2_1 _4382_ (.Y(_0849_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_nor2_1 _4383_ (.A(_0848_),
    .B(_0849_),
    .Y(_0850_));
 sg13g2_o21ai_1 _4384_ (.B1(_0843_),
    .Y(_0851_),
    .A1(_0811_),
    .A2(_0844_));
 sg13g2_nand2_1 _4385_ (.Y(_0852_),
    .A(_2153_),
    .B(net352));
 sg13g2_nor2_1 _4386_ (.A(_0747_),
    .B(_0812_),
    .Y(_0853_));
 sg13g2_o21ai_1 _4387_ (.B1(_0852_),
    .Y(_0854_),
    .A1(_0745_),
    .A2(_0853_));
 sg13g2_and2_1 _4388_ (.A(_0851_),
    .B(_0854_),
    .X(_0855_));
 sg13g2_xor2_1 _4389_ (.B(_0854_),
    .A(_0851_),
    .X(_0856_));
 sg13g2_nor2_1 _4390_ (.A(net357),
    .B(_2153_),
    .Y(_0857_));
 sg13g2_nand2_1 _4391_ (.Y(_0858_),
    .A(net357),
    .B(_0812_));
 sg13g2_o21ai_1 _4392_ (.B1(_0858_),
    .Y(_0859_),
    .A1(net354),
    .A2(_0018_));
 sg13g2_xnor2_1 _4393_ (.Y(_0860_),
    .A(_0856_),
    .B(_0859_));
 sg13g2_inv_1 _4394_ (.Y(_0861_),
    .A(_0860_));
 sg13g2_xor2_1 _4395_ (.B(_0849_),
    .A(_0848_),
    .X(_0862_));
 sg13g2_a21oi_1 _4396_ (.A1(_0861_),
    .A2(_0862_),
    .Y(_0863_),
    .B1(_0850_));
 sg13g2_xnor2_1 _4397_ (.Y(_0864_),
    .A(_0797_),
    .B(_0798_));
 sg13g2_or2_1 _4398_ (.X(_0865_),
    .B(_0864_),
    .A(_0863_));
 sg13g2_a21o_1 _4399_ (.A2(_0859_),
    .A1(_0856_),
    .B1(_0855_),
    .X(_0866_));
 sg13g2_xor2_1 _4400_ (.B(_0864_),
    .A(_0863_),
    .X(_0867_));
 sg13g2_nand2_1 _4401_ (.Y(_0868_),
    .A(_0866_),
    .B(_0867_));
 sg13g2_nand3_1 _4402_ (.B(_0865_),
    .C(_0868_),
    .A(_0830_),
    .Y(_0869_));
 sg13g2_a21oi_1 _4403_ (.A1(_0865_),
    .A2(_0868_),
    .Y(_0870_),
    .B1(_0830_));
 sg13g2_inv_1 _4404_ (.Y(_0871_),
    .A(_0870_));
 sg13g2_nand2_1 _4405_ (.Y(_0872_),
    .A(_0869_),
    .B(_0871_));
 sg13g2_xnor2_1 _4406_ (.Y(_0873_),
    .A(_0866_),
    .B(_0867_));
 sg13g2_xor2_1 _4407_ (.B(net373),
    .A(net372),
    .X(_0874_));
 sg13g2_nand2_1 _4408_ (.Y(_0875_),
    .A(net369),
    .B(_0874_));
 sg13g2_xor2_1 _4409_ (.B(_0874_),
    .A(net369),
    .X(_0876_));
 sg13g2_nand2_1 _4410_ (.Y(_0877_),
    .A(net375),
    .B(net378));
 sg13g2_nor2_2 _4411_ (.A(net375),
    .B(net377),
    .Y(_0878_));
 sg13g2_a21o_1 _4412_ (.A2(net377),
    .A1(net375),
    .B1(net378),
    .X(_0879_));
 sg13g2_o21ai_1 _4413_ (.B1(_0877_),
    .Y(_0880_),
    .A1(_0878_),
    .A2(_0879_));
 sg13g2_nand2_2 _4414_ (.Y(_0881_),
    .A(\am_sdr0.filt0.yn_2[1] ),
    .B(net378));
 sg13g2_nor2_2 _4415_ (.A(net376),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_a21oi_2 _4416_ (.B1(_0882_),
    .Y(_0883_),
    .A2(_0880_),
    .A1(_0876_));
 sg13g2_xnor2_1 _4417_ (.Y(_0884_),
    .A(_0832_),
    .B(_0836_));
 sg13g2_nor2_1 _4418_ (.A(_0883_),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_xor2_1 _4419_ (.B(_0884_),
    .A(_0883_),
    .X(_0886_));
 sg13g2_and2_2 _4420_ (.A(_0764_),
    .B(_0875_),
    .X(_0887_));
 sg13g2_nand2b_1 _4421_ (.Y(_0888_),
    .B(_0778_),
    .A_N(_0887_));
 sg13g2_xnor2_1 _4422_ (.Y(_0889_),
    .A(_0779_),
    .B(_0887_));
 sg13g2_xor2_1 _4423_ (.B(_0889_),
    .A(_0787_),
    .X(_0890_));
 sg13g2_a21oi_1 _4424_ (.A1(_0886_),
    .A2(_0890_),
    .Y(_0891_),
    .B1(_0885_));
 sg13g2_xnor2_1 _4425_ (.Y(_0892_),
    .A(_0845_),
    .B(_0846_));
 sg13g2_nor2_1 _4426_ (.A(_0891_),
    .B(_0892_),
    .Y(_0893_));
 sg13g2_nor2_1 _4427_ (.A(_0733_),
    .B(_0788_),
    .Y(_0894_));
 sg13g2_xor2_1 _4428_ (.B(_0788_),
    .A(_0733_),
    .X(_0895_));
 sg13g2_a21oi_1 _4429_ (.A1(net351),
    .A2(_0895_),
    .Y(_0896_),
    .B1(_0894_));
 sg13g2_o21ai_1 _4430_ (.B1(_0888_),
    .Y(_0897_),
    .A1(_0787_),
    .A2(_0889_));
 sg13g2_a21o_1 _4431_ (.A2(_0813_),
    .A1(net357),
    .B1(_0857_),
    .X(_0898_));
 sg13g2_xor2_1 _4432_ (.B(_0898_),
    .A(_0897_),
    .X(_0899_));
 sg13g2_nor2b_1 _4433_ (.A(_0896_),
    .B_N(_0899_),
    .Y(_0900_));
 sg13g2_xnor2_1 _4434_ (.Y(_0901_),
    .A(_0896_),
    .B(_0899_));
 sg13g2_xor2_1 _4435_ (.B(_0892_),
    .A(_0891_),
    .X(_0902_));
 sg13g2_a21oi_1 _4436_ (.A1(_0901_),
    .A2(_0902_),
    .Y(_0903_),
    .B1(_0893_));
 sg13g2_xnor2_1 _4437_ (.Y(_0904_),
    .A(_0860_),
    .B(_0862_));
 sg13g2_nor2b_1 _4438_ (.A(_0903_),
    .B_N(_0904_),
    .Y(_0905_));
 sg13g2_a21o_1 _4439_ (.A2(_0898_),
    .A1(_0897_),
    .B1(_0900_),
    .X(_0906_));
 sg13g2_xnor2_1 _4440_ (.Y(_0907_),
    .A(_0903_),
    .B(_0904_));
 sg13g2_a21oi_1 _4441_ (.A1(_0906_),
    .A2(_0907_),
    .Y(_0908_),
    .B1(_0905_));
 sg13g2_nor2_1 _4442_ (.A(_0873_),
    .B(_0908_),
    .Y(_0909_));
 sg13g2_inv_1 _4443_ (.Y(_0910_),
    .A(_0909_));
 sg13g2_xor2_1 _4444_ (.B(net378),
    .A(net377),
    .X(_0911_));
 sg13g2_xnor2_1 _4445_ (.Y(_0912_),
    .A(net373),
    .B(_0755_));
 sg13g2_nand2b_2 _4446_ (.Y(_0913_),
    .B(_0911_),
    .A_N(_0912_));
 sg13g2_xnor2_1 _4447_ (.Y(_0914_),
    .A(_0876_),
    .B(_0880_));
 sg13g2_nor2_1 _4448_ (.A(_0913_),
    .B(_0914_),
    .Y(_0915_));
 sg13g2_nand2_1 _4449_ (.Y(_0916_),
    .A(_0913_),
    .B(_0914_));
 sg13g2_xnor2_1 _4450_ (.Y(_0917_),
    .A(_0913_),
    .B(_0914_));
 sg13g2_a21oi_2 _4451_ (.B1(_0754_),
    .Y(_0918_),
    .A2(_0753_),
    .A1(_2147_));
 sg13g2_nand2_1 _4452_ (.Y(_0919_),
    .A(_0763_),
    .B(_0918_));
 sg13g2_xnor2_1 _4453_ (.Y(_0920_),
    .A(_0763_),
    .B(_0918_));
 sg13g2_xor2_1 _4454_ (.B(_0920_),
    .A(_0732_),
    .X(_0921_));
 sg13g2_a21oi_1 _4455_ (.A1(_0916_),
    .A2(_0921_),
    .Y(_0922_),
    .B1(_0915_));
 sg13g2_xnor2_1 _4456_ (.Y(_0923_),
    .A(_0886_),
    .B(_0890_));
 sg13g2_nor2_1 _4457_ (.A(_0922_),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_xor2_1 _4458_ (.B(_0923_),
    .A(_0922_),
    .X(_0925_));
 sg13g2_nand2_1 _4459_ (.Y(_0926_),
    .A(net364),
    .B(net359));
 sg13g2_nor2_1 _4460_ (.A(_0735_),
    .B(_0926_),
    .Y(_0927_));
 sg13g2_xor2_1 _4461_ (.B(_0926_),
    .A(_0735_),
    .X(_0928_));
 sg13g2_a21oi_2 _4462_ (.B1(_0927_),
    .Y(_0929_),
    .A2(_0928_),
    .A1(net353));
 sg13g2_o21ai_1 _4463_ (.B1(_0919_),
    .Y(_0930_),
    .A1(_0732_),
    .A2(_0920_));
 sg13g2_xnor2_1 _4464_ (.Y(_0931_),
    .A(net351),
    .B(_0895_));
 sg13g2_nand2b_1 _4465_ (.Y(_0932_),
    .B(_0930_),
    .A_N(_0931_));
 sg13g2_xor2_1 _4466_ (.B(_0931_),
    .A(_0930_),
    .X(_0933_));
 sg13g2_xor2_1 _4467_ (.B(_0933_),
    .A(_0929_),
    .X(_0934_));
 sg13g2_a21oi_1 _4468_ (.A1(_0925_),
    .A2(_0934_),
    .Y(_0935_),
    .B1(_0924_));
 sg13g2_xnor2_1 _4469_ (.Y(_0936_),
    .A(_0901_),
    .B(_0902_));
 sg13g2_nor2_1 _4470_ (.A(_0935_),
    .B(_0936_),
    .Y(_0937_));
 sg13g2_o21ai_1 _4471_ (.B1(_0932_),
    .Y(_0938_),
    .A1(_0929_),
    .A2(_0933_));
 sg13g2_xor2_1 _4472_ (.B(_0936_),
    .A(_0935_),
    .X(_0939_));
 sg13g2_and2_1 _4473_ (.A(_0938_),
    .B(_0939_),
    .X(_0940_));
 sg13g2_xor2_1 _4474_ (.B(_0907_),
    .A(_0906_),
    .X(_0941_));
 sg13g2_nor3_2 _4475_ (.A(_0937_),
    .B(_0940_),
    .C(_0941_),
    .Y(_0942_));
 sg13g2_o21ai_1 _4476_ (.B1(_0941_),
    .Y(_0943_),
    .A1(_0937_),
    .A2(_0940_));
 sg13g2_xor2_1 _4477_ (.B(_0834_),
    .A(net376),
    .X(_0944_));
 sg13g2_nand2b_1 _4478_ (.Y(_0945_),
    .B(net378),
    .A_N(_0944_));
 sg13g2_xnor2_1 _4479_ (.Y(_0946_),
    .A(_0911_),
    .B(_0912_));
 sg13g2_nor2b_1 _4480_ (.A(_0945_),
    .B_N(_0946_),
    .Y(_0947_));
 sg13g2_xnor2_1 _4481_ (.Y(_0948_),
    .A(_0945_),
    .B(_0946_));
 sg13g2_a21oi_2 _4482_ (.B1(_0878_),
    .Y(_0949_),
    .A2(_0837_),
    .A1(_2147_));
 sg13g2_nor2b_1 _4483_ (.A(_0751_),
    .B_N(_0949_),
    .Y(_0950_));
 sg13g2_xnor2_1 _4484_ (.Y(_0951_),
    .A(_0751_),
    .B(_0949_));
 sg13g2_xnor2_1 _4485_ (.Y(_0952_),
    .A(_0841_),
    .B(_0951_));
 sg13g2_a21oi_1 _4486_ (.A1(_0948_),
    .A2(_0952_),
    .Y(_0953_),
    .B1(_0947_));
 sg13g2_xnor2_1 _4487_ (.Y(_0954_),
    .A(_0917_),
    .B(_0921_));
 sg13g2_nor2b_1 _4488_ (.A(_0953_),
    .B_N(_0954_),
    .Y(_0955_));
 sg13g2_xnor2_1 _4489_ (.Y(_0956_),
    .A(_0953_),
    .B(_0954_));
 sg13g2_xor2_1 _4490_ (.B(net359),
    .A(net363),
    .X(_0957_));
 sg13g2_and2_1 _4491_ (.A(net360),
    .B(_0957_),
    .X(_0958_));
 sg13g2_a21oi_1 _4492_ (.A1(net365),
    .A2(net361),
    .Y(_0959_),
    .B1(_0957_));
 sg13g2_a21oi_1 _4493_ (.A1(net366),
    .A2(_0958_),
    .Y(_0960_),
    .B1(_0959_));
 sg13g2_a22oi_1 _4494_ (.Y(_0961_),
    .B1(_0960_),
    .B2(net356),
    .A2(_0958_),
    .A1(net366));
 sg13g2_a21oi_1 _4495_ (.A1(_0842_),
    .A2(_0951_),
    .Y(_0962_),
    .B1(_0950_));
 sg13g2_xnor2_1 _4496_ (.Y(_0963_),
    .A(net353),
    .B(_0928_));
 sg13g2_xor2_1 _4497_ (.B(_0963_),
    .A(_0962_),
    .X(_0964_));
 sg13g2_nand2b_1 _4498_ (.Y(_0965_),
    .B(_0964_),
    .A_N(_0961_));
 sg13g2_xnor2_1 _4499_ (.Y(_0966_),
    .A(_0961_),
    .B(_0964_));
 sg13g2_a21oi_1 _4500_ (.A1(_0956_),
    .A2(_0966_),
    .Y(_0967_),
    .B1(_0955_));
 sg13g2_xnor2_1 _4501_ (.Y(_0968_),
    .A(_0925_),
    .B(_0934_));
 sg13g2_nor2_1 _4502_ (.A(_0967_),
    .B(_0968_),
    .Y(_0969_));
 sg13g2_o21ai_1 _4503_ (.B1(_0965_),
    .Y(_0970_),
    .A1(_0962_),
    .A2(_0963_));
 sg13g2_xor2_1 _4504_ (.B(_0968_),
    .A(_0967_),
    .X(_0971_));
 sg13g2_and2_1 _4505_ (.A(_0970_),
    .B(_0971_),
    .X(_0972_));
 sg13g2_xor2_1 _4506_ (.B(_0939_),
    .A(_0938_),
    .X(_0973_));
 sg13g2_o21ai_1 _4507_ (.B1(_0973_),
    .Y(_0974_),
    .A1(_0969_),
    .A2(_0972_));
 sg13g2_inv_1 _4508_ (.Y(_0975_),
    .A(_0974_));
 sg13g2_o21ai_1 _4509_ (.B1(_0943_),
    .Y(_0976_),
    .A1(_0942_),
    .A2(_0974_));
 sg13g2_xnor2_1 _4510_ (.Y(_0977_),
    .A(_0970_),
    .B(_0971_));
 sg13g2_xnor2_1 _4511_ (.Y(_0978_),
    .A(net378),
    .B(_0944_));
 sg13g2_nor2b_2 _4512_ (.A(_0878_),
    .B_N(_0879_),
    .Y(_0979_));
 sg13g2_nand2_1 _4513_ (.Y(_0980_),
    .A(_0832_),
    .B(_0979_));
 sg13g2_nor2_1 _4514_ (.A(_0832_),
    .B(_0979_),
    .Y(_0981_));
 sg13g2_xor2_1 _4515_ (.B(_0979_),
    .A(_0832_),
    .X(_0982_));
 sg13g2_xnor2_1 _4516_ (.Y(_0983_),
    .A(_0887_),
    .B(_0982_));
 sg13g2_nand2_1 _4517_ (.Y(_0984_),
    .A(_0978_),
    .B(_0983_));
 sg13g2_xnor2_1 _4518_ (.Y(_0985_),
    .A(_0948_),
    .B(_0952_));
 sg13g2_nor2_1 _4519_ (.A(_0984_),
    .B(_0985_),
    .Y(_0986_));
 sg13g2_xor2_1 _4520_ (.B(_0985_),
    .A(_0984_),
    .X(_0987_));
 sg13g2_nand2_1 _4521_ (.Y(_0988_),
    .A(net368),
    .B(net364));
 sg13g2_xor2_1 _4522_ (.B(net362),
    .A(\am_sdr0.filt0.yn_2[7] ),
    .X(_0989_));
 sg13g2_nor2b_1 _4523_ (.A(_0988_),
    .B_N(_0989_),
    .Y(_0990_));
 sg13g2_xnor2_1 _4524_ (.Y(_0991_),
    .A(_0988_),
    .B(_0989_));
 sg13g2_a21oi_1 _4525_ (.A1(\am_sdr0.filt0.yn_2[10] ),
    .A2(_0991_),
    .Y(_0992_),
    .B1(_0990_));
 sg13g2_o21ai_1 _4526_ (.B1(_0980_),
    .Y(_0993_),
    .A1(_0887_),
    .A2(_0981_));
 sg13g2_xnor2_1 _4527_ (.Y(_0994_),
    .A(net356),
    .B(_0960_));
 sg13g2_nor2b_1 _4528_ (.A(_0994_),
    .B_N(_0993_),
    .Y(_0995_));
 sg13g2_xor2_1 _4529_ (.B(_0994_),
    .A(_0993_),
    .X(_0996_));
 sg13g2_nor2_1 _4530_ (.A(_0992_),
    .B(_0996_),
    .Y(_0997_));
 sg13g2_xor2_1 _4531_ (.B(_0996_),
    .A(_0992_),
    .X(_0998_));
 sg13g2_a21oi_1 _4532_ (.A1(_0987_),
    .A2(_0998_),
    .Y(_0999_),
    .B1(_0986_));
 sg13g2_xnor2_1 _4533_ (.Y(_1000_),
    .A(_0956_),
    .B(_0966_));
 sg13g2_nor2_1 _4534_ (.A(_0995_),
    .B(_0997_),
    .Y(_1001_));
 sg13g2_xor2_1 _4535_ (.B(_1000_),
    .A(_0999_),
    .X(_1002_));
 sg13g2_nand2b_1 _4536_ (.Y(_1003_),
    .B(_1002_),
    .A_N(_1001_));
 sg13g2_o21ai_1 _4537_ (.B1(_1003_),
    .Y(_1004_),
    .A1(_0999_),
    .A2(_1000_));
 sg13g2_nand2b_1 _4538_ (.Y(_1005_),
    .B(_0977_),
    .A_N(_1004_));
 sg13g2_nor2b_1 _4539_ (.A(_0977_),
    .B_N(_1004_),
    .Y(_1006_));
 sg13g2_xor2_1 _4540_ (.B(_1002_),
    .A(_1001_),
    .X(_1007_));
 sg13g2_and3_1 _4541_ (.X(_1008_),
    .A(net377),
    .B(net378),
    .C(_0876_));
 sg13g2_xnor2_1 _4542_ (.Y(_1009_),
    .A(_0876_),
    .B(_0881_));
 sg13g2_xnor2_1 _4543_ (.Y(_1010_),
    .A(_0918_),
    .B(_1009_));
 sg13g2_xnor2_1 _4544_ (.Y(_1011_),
    .A(net376),
    .B(_0911_));
 sg13g2_nor2_1 _4545_ (.A(_1010_),
    .B(_1011_),
    .Y(_1012_));
 sg13g2_xnor2_1 _4546_ (.Y(_1013_),
    .A(_0978_),
    .B(_0983_));
 sg13g2_nor3_1 _4547_ (.A(_1010_),
    .B(_1011_),
    .C(_1013_),
    .Y(_1014_));
 sg13g2_xnor2_1 _4548_ (.Y(_1015_),
    .A(_1012_),
    .B(_1013_));
 sg13g2_nand2_1 _4549_ (.Y(_1016_),
    .A(net370),
    .B(net366));
 sg13g2_xor2_1 _4550_ (.B(net364),
    .A(net368),
    .X(_1017_));
 sg13g2_nor2b_1 _4551_ (.A(_1016_),
    .B_N(_1017_),
    .Y(_1018_));
 sg13g2_xnor2_1 _4552_ (.Y(_1019_),
    .A(_1016_),
    .B(_1017_));
 sg13g2_a21oi_1 _4553_ (.A1(net362),
    .A2(_1019_),
    .Y(_1020_),
    .B1(_1018_));
 sg13g2_inv_1 _4554_ (.Y(_1021_),
    .A(_1020_));
 sg13g2_a21oi_1 _4555_ (.A1(_0918_),
    .A2(_1009_),
    .Y(_1022_),
    .B1(_1008_));
 sg13g2_xnor2_1 _4556_ (.Y(_1023_),
    .A(\am_sdr0.filt0.yn_2[10] ),
    .B(_0991_));
 sg13g2_nor2_1 _4557_ (.A(_1022_),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_xor2_1 _4558_ (.B(_1023_),
    .A(_1022_),
    .X(_1025_));
 sg13g2_xnor2_1 _4559_ (.Y(_1026_),
    .A(_1020_),
    .B(_1025_));
 sg13g2_a21oi_1 _4560_ (.A1(_1015_),
    .A2(_1026_),
    .Y(_1027_),
    .B1(_1014_));
 sg13g2_xor2_1 _4561_ (.B(_0998_),
    .A(_0987_),
    .X(_1028_));
 sg13g2_nand2b_1 _4562_ (.Y(_1029_),
    .B(_1028_),
    .A_N(_1027_));
 sg13g2_a21oi_1 _4563_ (.A1(_1021_),
    .A2(_1025_),
    .Y(_1030_),
    .B1(_1024_));
 sg13g2_xnor2_1 _4564_ (.Y(_1031_),
    .A(_1027_),
    .B(_1028_));
 sg13g2_nand2b_1 _4565_ (.Y(_1032_),
    .B(_1031_),
    .A_N(_1030_));
 sg13g2_nand2_1 _4566_ (.Y(_1033_),
    .A(_1029_),
    .B(_1032_));
 sg13g2_a21oi_2 _4567_ (.B1(_1007_),
    .Y(_1034_),
    .A2(_1032_),
    .A1(_1029_));
 sg13g2_nand2b_1 _4568_ (.Y(_1035_),
    .B(_0949_),
    .A_N(_0912_));
 sg13g2_xnor2_1 _4569_ (.Y(_1036_),
    .A(_0912_),
    .B(_0949_));
 sg13g2_nand2_1 _4570_ (.Y(_1037_),
    .A(_0911_),
    .B(_1036_));
 sg13g2_xnor2_1 _4571_ (.Y(_1038_),
    .A(_1010_),
    .B(_1011_));
 sg13g2_nor2_1 _4572_ (.A(_1037_),
    .B(_1038_),
    .Y(_1039_));
 sg13g2_xor2_1 _4573_ (.B(_1038_),
    .A(_1037_),
    .X(_1040_));
 sg13g2_xor2_1 _4574_ (.B(net366),
    .A(net369),
    .X(_1041_));
 sg13g2_nand2_1 _4575_ (.Y(_1042_),
    .A(net371),
    .B(net368));
 sg13g2_and3_1 _4576_ (.X(_1043_),
    .A(\am_sdr0.filt0.yn_2[4] ),
    .B(net368),
    .C(_1041_));
 sg13g2_xnor2_1 _4577_ (.Y(_1044_),
    .A(_1041_),
    .B(_1042_));
 sg13g2_a21oi_1 _4578_ (.A1(net364),
    .A2(_1044_),
    .Y(_1045_),
    .B1(_1043_));
 sg13g2_xnor2_1 _4579_ (.Y(_1046_),
    .A(net362),
    .B(_1019_));
 sg13g2_or2_1 _4580_ (.X(_1047_),
    .B(_1046_),
    .A(_1035_));
 sg13g2_xnor2_1 _4581_ (.Y(_1048_),
    .A(_1035_),
    .B(_1046_));
 sg13g2_xor2_1 _4582_ (.B(_1048_),
    .A(_1045_),
    .X(_1049_));
 sg13g2_a21oi_2 _4583_ (.B1(_1039_),
    .Y(_1050_),
    .A2(_1049_),
    .A1(_1040_));
 sg13g2_xor2_1 _4584_ (.B(_1026_),
    .A(_1015_),
    .X(_1051_));
 sg13g2_nor2b_1 _4585_ (.A(_1050_),
    .B_N(_1051_),
    .Y(_1052_));
 sg13g2_o21ai_1 _4586_ (.B1(_1047_),
    .Y(_1053_),
    .A1(_1045_),
    .A2(_1048_));
 sg13g2_xnor2_1 _4587_ (.Y(_1054_),
    .A(_1050_),
    .B(_1051_));
 sg13g2_a21oi_2 _4588_ (.B1(_1052_),
    .Y(_1055_),
    .A2(_1054_),
    .A1(_1053_));
 sg13g2_xor2_1 _4589_ (.B(_1031_),
    .A(_1030_),
    .X(_1056_));
 sg13g2_nor2_1 _4590_ (.A(_1055_),
    .B(_1056_),
    .Y(_1057_));
 sg13g2_nand2_1 _4591_ (.Y(_1058_),
    .A(_1055_),
    .B(_1056_));
 sg13g2_inv_1 _4592_ (.Y(_1059_),
    .A(_1058_));
 sg13g2_xnor2_1 _4593_ (.Y(_1060_),
    .A(_1053_),
    .B(_1054_));
 sg13g2_xnor2_1 _4594_ (.Y(_1061_),
    .A(_0911_),
    .B(_1036_));
 sg13g2_nand2b_1 _4595_ (.Y(_1062_),
    .B(_0979_),
    .A_N(_0944_));
 sg13g2_xnor2_1 _4596_ (.Y(_1063_),
    .A(_0944_),
    .B(_0979_));
 sg13g2_nand2_1 _4597_ (.Y(_1064_),
    .A(\am_sdr0.filt0.mul_a2[1] ),
    .B(_1063_));
 sg13g2_nor2_1 _4598_ (.A(_1061_),
    .B(_1064_),
    .Y(_1065_));
 sg13g2_xor2_1 _4599_ (.B(_1064_),
    .A(_1061_),
    .X(_1066_));
 sg13g2_xor2_1 _4600_ (.B(net368),
    .A(\am_sdr0.filt0.yn_2[4] ),
    .X(_1067_));
 sg13g2_nand2_1 _4601_ (.Y(_1068_),
    .A(net374),
    .B(net369));
 sg13g2_and3_1 _4602_ (.X(_1069_),
    .A(net374),
    .B(net369),
    .C(_1067_));
 sg13g2_xnor2_1 _4603_ (.Y(_1070_),
    .A(_1067_),
    .B(_1068_));
 sg13g2_a21oi_2 _4604_ (.B1(_1069_),
    .Y(_1071_),
    .A2(_1070_),
    .A1(net366));
 sg13g2_xnor2_1 _4605_ (.Y(_1072_),
    .A(net364),
    .B(_1044_));
 sg13g2_xnor2_1 _4606_ (.Y(_1073_),
    .A(_1062_),
    .B(_1072_));
 sg13g2_or2_1 _4607_ (.X(_1074_),
    .B(_1073_),
    .A(_1071_));
 sg13g2_xor2_1 _4608_ (.B(_1073_),
    .A(_1071_),
    .X(_1075_));
 sg13g2_a21oi_1 _4609_ (.A1(_1066_),
    .A2(_1075_),
    .Y(_1076_),
    .B1(_1065_));
 sg13g2_xnor2_1 _4610_ (.Y(_1077_),
    .A(_1040_),
    .B(_1049_));
 sg13g2_nor2_1 _4611_ (.A(_1076_),
    .B(_1077_),
    .Y(_1078_));
 sg13g2_o21ai_1 _4612_ (.B1(_1074_),
    .Y(_1079_),
    .A1(_1062_),
    .A2(_1072_));
 sg13g2_xor2_1 _4613_ (.B(_1077_),
    .A(_1076_),
    .X(_1080_));
 sg13g2_a21oi_1 _4614_ (.A1(_1079_),
    .A2(_1080_),
    .Y(_1081_),
    .B1(_1078_));
 sg13g2_or2_1 _4615_ (.X(_1082_),
    .B(_1081_),
    .A(_1060_));
 sg13g2_xnor2_1 _4616_ (.Y(_1083_),
    .A(_1060_),
    .B(_1081_));
 sg13g2_xnor2_1 _4617_ (.Y(_1084_),
    .A(\am_sdr0.filt0.mul_a2[1] ),
    .B(_1063_));
 sg13g2_xor2_1 _4618_ (.B(net369),
    .A(net374),
    .X(_1085_));
 sg13g2_nand2b_1 _4619_ (.Y(_1086_),
    .B(_1085_),
    .A_N(_0753_));
 sg13g2_xnor2_1 _4620_ (.Y(_1087_),
    .A(_0753_),
    .B(_1085_));
 sg13g2_nand2_1 _4621_ (.Y(_1088_),
    .A(net368),
    .B(_1087_));
 sg13g2_nand2_1 _4622_ (.Y(_1089_),
    .A(_1086_),
    .B(_1088_));
 sg13g2_nand3_1 _4623_ (.B(net377),
    .C(\am_sdr0.filt0.mul_a2[1] ),
    .A(net376),
    .Y(_1090_));
 sg13g2_xnor2_1 _4624_ (.Y(_1091_),
    .A(net366),
    .B(_1070_));
 sg13g2_nor2_1 _4625_ (.A(_1090_),
    .B(_1091_),
    .Y(_1092_));
 sg13g2_nand2_1 _4626_ (.Y(_1093_),
    .A(_1090_),
    .B(_1091_));
 sg13g2_xnor2_1 _4627_ (.Y(_1094_),
    .A(_1090_),
    .B(_1091_));
 sg13g2_xnor2_1 _4628_ (.Y(_1095_),
    .A(_1089_),
    .B(_1094_));
 sg13g2_nand2b_1 _4629_ (.Y(_1096_),
    .B(_1095_),
    .A_N(_1084_));
 sg13g2_xnor2_1 _4630_ (.Y(_1097_),
    .A(_1066_),
    .B(_1075_));
 sg13g2_nor2_1 _4631_ (.A(_1096_),
    .B(_1097_),
    .Y(_1098_));
 sg13g2_a21oi_1 _4632_ (.A1(_1089_),
    .A2(_1093_),
    .Y(_1099_),
    .B1(_1092_));
 sg13g2_xor2_1 _4633_ (.B(_1097_),
    .A(_1096_),
    .X(_1100_));
 sg13g2_nor2b_1 _4634_ (.A(_1099_),
    .B_N(_1100_),
    .Y(_1101_));
 sg13g2_nor2_1 _4635_ (.A(_1098_),
    .B(_1101_),
    .Y(_1102_));
 sg13g2_xor2_1 _4636_ (.B(_1080_),
    .A(_1079_),
    .X(_1103_));
 sg13g2_nand2b_1 _4637_ (.Y(_1104_),
    .B(_1103_),
    .A_N(_1102_));
 sg13g2_xnor2_1 _4638_ (.Y(_1105_),
    .A(_1084_),
    .B(_1095_));
 sg13g2_nor2_1 _4639_ (.A(_0756_),
    .B(_0833_),
    .Y(_1106_));
 sg13g2_xnor2_1 _4640_ (.Y(_1107_),
    .A(_0755_),
    .B(_0833_));
 sg13g2_a21oi_2 _4641_ (.B1(_1106_),
    .Y(_1108_),
    .A2(_1107_),
    .A1(net369));
 sg13g2_xnor2_1 _4642_ (.Y(_1109_),
    .A(net367),
    .B(_1087_));
 sg13g2_nand2_1 _4643_ (.Y(_1110_),
    .A(_0881_),
    .B(_1011_));
 sg13g2_nand2_1 _4644_ (.Y(_1111_),
    .A(_1090_),
    .B(_1110_));
 sg13g2_xor2_1 _4645_ (.B(_1109_),
    .A(_1108_),
    .X(_1112_));
 sg13g2_nand2b_1 _4646_ (.Y(_1113_),
    .B(_1112_),
    .A_N(_1111_));
 sg13g2_o21ai_1 _4647_ (.B1(_1113_),
    .Y(_1114_),
    .A1(_1108_),
    .A2(_1109_));
 sg13g2_and2_1 _4648_ (.A(_1105_),
    .B(_1114_),
    .X(_1115_));
 sg13g2_xnor2_1 _4649_ (.Y(_1116_),
    .A(_1099_),
    .B(_1100_));
 sg13g2_and2_1 _4650_ (.A(_1115_),
    .B(_1116_),
    .X(_1117_));
 sg13g2_xor2_1 _4651_ (.B(_1114_),
    .A(_1105_),
    .X(_1118_));
 sg13g2_xor2_1 _4652_ (.B(_1112_),
    .A(_1111_),
    .X(_1119_));
 sg13g2_nor2_1 _4653_ (.A(_0834_),
    .B(_0877_),
    .Y(_1120_));
 sg13g2_xor2_1 _4654_ (.B(_0877_),
    .A(_0834_),
    .X(_1121_));
 sg13g2_a21oi_1 _4655_ (.A1(net371),
    .A2(_1121_),
    .Y(_1122_),
    .B1(_1120_));
 sg13g2_xnor2_1 _4656_ (.Y(_1123_),
    .A(net369),
    .B(_1107_));
 sg13g2_nor2_1 _4657_ (.A(_1122_),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_xor2_1 _4658_ (.B(_1123_),
    .A(_1122_),
    .X(_1125_));
 sg13g2_a21oi_2 _4659_ (.B1(_1124_),
    .Y(_1126_),
    .A2(_1125_),
    .A1(_0911_));
 sg13g2_nor2_2 _4660_ (.A(_1119_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_nand2_1 _4661_ (.Y(_1128_),
    .A(_1118_),
    .B(_1127_));
 sg13g2_xor2_1 _4662_ (.B(_1125_),
    .A(_0911_),
    .X(_1129_));
 sg13g2_xnor2_1 _4663_ (.Y(_1130_),
    .A(net371),
    .B(_1121_));
 sg13g2_a22oi_1 _4664_ (.Y(_1131_),
    .B1(_0835_),
    .B2(_1130_),
    .A2(_0758_),
    .A1(_2152_));
 sg13g2_nand2_1 _4665_ (.Y(_1132_),
    .A(_1129_),
    .B(_1131_));
 sg13g2_xnor2_1 _4666_ (.Y(_1133_),
    .A(_1119_),
    .B(_1126_));
 sg13g2_or2_1 _4667_ (.X(_1134_),
    .B(_1133_),
    .A(_1132_));
 sg13g2_nor3_2 _4668_ (.A(_0837_),
    .B(_0874_),
    .C(_0978_),
    .Y(_1135_));
 sg13g2_xor2_1 _4669_ (.B(_1131_),
    .A(_1129_),
    .X(_1136_));
 sg13g2_and2_1 _4670_ (.A(_1135_),
    .B(_1136_),
    .X(_1137_));
 sg13g2_nand3_1 _4671_ (.B(_2147_),
    .C(_0882_),
    .A(net371),
    .Y(_1138_));
 sg13g2_xnor2_1 _4672_ (.Y(_1139_),
    .A(_1135_),
    .B(_1136_));
 sg13g2_and4_1 _4673_ (.A(net371),
    .B(_2147_),
    .C(_0882_),
    .D(_1136_),
    .X(_1140_));
 sg13g2_xor2_1 _4674_ (.B(_1133_),
    .A(_1132_),
    .X(_1141_));
 sg13g2_o21ai_1 _4675_ (.B1(_1141_),
    .Y(_1142_),
    .A1(_1137_),
    .A2(_1140_));
 sg13g2_xnor2_1 _4676_ (.Y(_1143_),
    .A(_1118_),
    .B(_1127_));
 sg13g2_a21o_1 _4677_ (.A2(_1142_),
    .A1(_1134_),
    .B1(_1143_),
    .X(_1144_));
 sg13g2_xnor2_1 _4678_ (.Y(_1145_),
    .A(_1115_),
    .B(_1116_));
 sg13g2_a21oi_2 _4679_ (.B1(_1145_),
    .Y(_1146_),
    .A2(_1144_),
    .A1(_1128_));
 sg13g2_xnor2_1 _4680_ (.Y(_1147_),
    .A(_1102_),
    .B(_1103_));
 sg13g2_o21ai_1 _4681_ (.B1(_1147_),
    .Y(_1148_),
    .A1(_1117_),
    .A2(_1146_));
 sg13g2_a21o_2 _4682_ (.A2(_1148_),
    .A1(_1104_),
    .B1(_1083_),
    .X(_1149_));
 sg13g2_nor2b_1 _4683_ (.A(_1057_),
    .B_N(_1082_),
    .Y(_1150_));
 sg13g2_a21oi_1 _4684_ (.A1(_1149_),
    .A2(_1150_),
    .Y(_1151_),
    .B1(_1059_));
 sg13g2_xor2_1 _4685_ (.B(_1033_),
    .A(_1007_),
    .X(_1152_));
 sg13g2_a221oi_1 _4686_ (.B2(_1150_),
    .C1(_1152_),
    .B1(_1149_),
    .A1(_1055_),
    .Y(_1153_),
    .A2(_1056_));
 sg13g2_xor2_1 _4687_ (.B(_1004_),
    .A(_0977_),
    .X(_1154_));
 sg13g2_or2_1 _4688_ (.X(_1155_),
    .B(_1154_),
    .A(_1152_));
 sg13g2_a221oi_1 _4689_ (.B2(_1150_),
    .C1(_1155_),
    .B1(_1149_),
    .A1(_1055_),
    .Y(_1156_),
    .A2(_1056_));
 sg13g2_a21oi_1 _4690_ (.A1(_1005_),
    .A2(_1034_),
    .Y(_1157_),
    .B1(_1006_));
 sg13g2_inv_1 _4691_ (.Y(_1158_),
    .A(_1157_));
 sg13g2_nand2b_1 _4692_ (.Y(_1159_),
    .B(_1157_),
    .A_N(_0976_));
 sg13g2_nor3_1 _4693_ (.A(_0969_),
    .B(_0972_),
    .C(_0973_),
    .Y(_1160_));
 sg13g2_a21oi_1 _4694_ (.A1(_0943_),
    .A2(_1160_),
    .Y(_1161_),
    .B1(_0942_));
 sg13g2_o21ai_1 _4695_ (.B1(_1161_),
    .Y(_1162_),
    .A1(_1156_),
    .A2(_1159_));
 sg13g2_xnor2_1 _4696_ (.Y(_1163_),
    .A(_0873_),
    .B(_0908_));
 sg13g2_o21ai_1 _4697_ (.B1(_0910_),
    .Y(_1164_),
    .A1(_1162_),
    .A2(_1163_));
 sg13g2_xnor2_1 _4698_ (.Y(_1165_),
    .A(_0872_),
    .B(_1164_));
 sg13g2_nor2_1 _4699_ (.A(_0729_),
    .B(_1165_),
    .Y(_1166_));
 sg13g2_xor2_1 _4700_ (.B(_1165_),
    .A(_0729_),
    .X(_1167_));
 sg13g2_a21oi_1 _4701_ (.A1(net344),
    .A2(_1167_),
    .Y(_1168_),
    .B1(_1166_));
 sg13g2_nor2_1 _4702_ (.A(_0823_),
    .B(_0825_),
    .Y(_1169_));
 sg13g2_o21ai_1 _4703_ (.B1(net350),
    .Y(_1170_),
    .A1(_0816_),
    .A2(_0820_));
 sg13g2_or3_1 _4704_ (.A(net350),
    .B(_0816_),
    .C(_0820_),
    .X(_1171_));
 sg13g2_and2_1 _4705_ (.A(_1170_),
    .B(_1171_),
    .X(_1172_));
 sg13g2_a21oi_1 _4706_ (.A1(_0810_),
    .A2(_0821_),
    .Y(_1173_),
    .B1(_0809_));
 sg13g2_a21oi_1 _4707_ (.A1(_2149_),
    .A2(_0730_),
    .Y(_1174_),
    .B1(_0807_));
 sg13g2_nor2b_1 _4708_ (.A(net363),
    .B_N(_0761_),
    .Y(_1175_));
 sg13g2_nor2_1 _4709_ (.A(_0761_),
    .B(_0777_),
    .Y(_1176_));
 sg13g2_nor2_1 _4710_ (.A(_1175_),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_nor2b_1 _4711_ (.A(_0736_),
    .B_N(_1177_),
    .Y(_1178_));
 sg13g2_xnor2_1 _4712_ (.Y(_1179_),
    .A(_0736_),
    .B(_1177_));
 sg13g2_nor2b_1 _4713_ (.A(_1174_),
    .B_N(_1179_),
    .Y(_1180_));
 sg13g2_xnor2_1 _4714_ (.Y(_1181_),
    .A(_1174_),
    .B(_1179_));
 sg13g2_nor2_1 _4715_ (.A(_2154_),
    .B(_0740_),
    .Y(_1182_));
 sg13g2_xnor2_1 _4716_ (.Y(_1183_),
    .A(net352),
    .B(_0740_));
 sg13g2_a21oi_2 _4717_ (.B1(_0814_),
    .Y(_1184_),
    .A2(_2154_),
    .A1(_2153_));
 sg13g2_xor2_1 _4718_ (.B(_1184_),
    .A(_1183_),
    .X(_1185_));
 sg13g2_xnor2_1 _4719_ (.Y(_1186_),
    .A(_1181_),
    .B(_1185_));
 sg13g2_nor2_1 _4720_ (.A(_1173_),
    .B(_1186_),
    .Y(_1187_));
 sg13g2_xor2_1 _4721_ (.B(_1186_),
    .A(_1173_),
    .X(_1188_));
 sg13g2_xnor2_1 _4722_ (.Y(_1189_),
    .A(_1172_),
    .B(_1188_));
 sg13g2_nor2_1 _4723_ (.A(_1169_),
    .B(_1189_),
    .Y(_1190_));
 sg13g2_xor2_1 _4724_ (.B(_1189_),
    .A(_1169_),
    .X(_1191_));
 sg13g2_and2_1 _4725_ (.A(_0801_),
    .B(_1191_),
    .X(_1192_));
 sg13g2_xnor2_1 _4726_ (.Y(_1193_),
    .A(_0801_),
    .B(_1191_));
 sg13g2_a21oi_1 _4727_ (.A1(_0827_),
    .A2(_0829_),
    .Y(_1194_),
    .B1(_1193_));
 sg13g2_nand3_1 _4728_ (.B(_0829_),
    .C(_1193_),
    .A(_0827_),
    .Y(_1195_));
 sg13g2_inv_1 _4729_ (.Y(_1196_),
    .A(_1195_));
 sg13g2_nor2_1 _4730_ (.A(_1194_),
    .B(_1196_),
    .Y(_1197_));
 sg13g2_nand3b_1 _4731_ (.B(_0871_),
    .C(_0869_),
    .Y(_1198_),
    .A_N(_1163_));
 sg13g2_a21oi_1 _4732_ (.A1(_0869_),
    .A2(_0909_),
    .Y(_1199_),
    .B1(_0870_));
 sg13g2_o21ai_1 _4733_ (.B1(_1199_),
    .Y(_1200_),
    .A1(_1162_),
    .A2(_1198_));
 sg13g2_xnor2_1 _4734_ (.Y(_1201_),
    .A(_1197_),
    .B(_1200_));
 sg13g2_a21o_1 _4735_ (.A2(_0532_),
    .A1(_0510_),
    .B1(_0531_),
    .X(_1202_));
 sg13g2_nand3_1 _4736_ (.B(_0480_),
    .C(_0511_),
    .A(net395),
    .Y(_1203_));
 sg13g2_nand2_1 _4737_ (.Y(_1204_),
    .A(_0481_),
    .B(_0523_));
 sg13g2_o21ai_1 _4738_ (.B1(_1204_),
    .Y(_1205_),
    .A1(_0481_),
    .A2(_0526_));
 sg13g2_xor2_1 _4739_ (.B(net393),
    .A(net380),
    .X(_1206_));
 sg13g2_nand2b_1 _4740_ (.Y(_1207_),
    .B(_1206_),
    .A_N(_1205_));
 sg13g2_xnor2_1 _4741_ (.Y(_1208_),
    .A(_1205_),
    .B(_1206_));
 sg13g2_nand2b_1 _4742_ (.Y(_1209_),
    .B(_1208_),
    .A_N(_0529_));
 sg13g2_xnor2_1 _4743_ (.Y(_1210_),
    .A(_0529_),
    .B(_1208_));
 sg13g2_inv_1 _4744_ (.Y(_1211_),
    .A(_1210_));
 sg13g2_xnor2_1 _4745_ (.Y(_1212_),
    .A(_1203_),
    .B(_1210_));
 sg13g2_xnor2_1 _4746_ (.Y(_1213_),
    .A(_1202_),
    .B(_1212_));
 sg13g2_nor2_1 _4747_ (.A(net342),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_xnor2_1 _4748_ (.Y(_1215_),
    .A(net342),
    .B(_1213_));
 sg13g2_nand3_1 _4749_ (.B(_0537_),
    .C(_1215_),
    .A(_0535_),
    .Y(_1216_));
 sg13g2_inv_1 _4750_ (.Y(_1217_),
    .A(_1216_));
 sg13g2_a21oi_1 _4751_ (.A1(_0535_),
    .A2(_0537_),
    .Y(_1218_),
    .B1(_1215_));
 sg13g2_nor2_1 _4752_ (.A(_1217_),
    .B(_1218_),
    .Y(_1219_));
 sg13g2_nand3_1 _4753_ (.B(_0727_),
    .C(_1219_),
    .A(_0542_),
    .Y(_1220_));
 sg13g2_a21o_1 _4754_ (.A2(_0727_),
    .A1(_0542_),
    .B1(_1219_),
    .X(_1221_));
 sg13g2_nand3_1 _4755_ (.B(_1220_),
    .C(_1221_),
    .A(_1201_),
    .Y(_1222_));
 sg13g2_a21o_1 _4756_ (.A2(_1221_),
    .A1(_1220_),
    .B1(_1201_),
    .X(_1223_));
 sg13g2_and3_1 _4757_ (.X(_1224_),
    .A(net345),
    .B(_1222_),
    .C(_1223_));
 sg13g2_nand3_1 _4758_ (.B(_1222_),
    .C(_1223_),
    .A(net344),
    .Y(_1225_));
 sg13g2_a21oi_1 _4759_ (.A1(_1222_),
    .A2(_1223_),
    .Y(_1226_),
    .B1(net344));
 sg13g2_or3_1 _4760_ (.A(_1168_),
    .B(_1224_),
    .C(_1226_),
    .X(_1227_));
 sg13g2_nand2b_1 _4761_ (.Y(_1228_),
    .B(\am_sdr0.filt0.xn_2[5] ),
    .A_N(\am_sdr0.filt0.xn_2[3] ));
 sg13g2_nor2b_1 _4762_ (.A(\am_sdr0.filt0.xn_2[4] ),
    .B_N(\am_sdr0.filt0.xn_2[6] ),
    .Y(_1229_));
 sg13g2_xnor2_1 _4763_ (.Y(_1230_),
    .A(\am_sdr0.filt0.xn_2[6] ),
    .B(\am_sdr0.filt0.xn_2[4] ));
 sg13g2_nand2b_1 _4764_ (.Y(_1231_),
    .B(_1230_),
    .A_N(_1228_));
 sg13g2_xnor2_1 _4765_ (.Y(_1232_),
    .A(_1228_),
    .B(_1230_));
 sg13g2_nand2_1 _4766_ (.Y(_1233_),
    .A(\am_sdr0.filt0.xn_2[7] ),
    .B(_1232_));
 sg13g2_nand2_1 _4767_ (.Y(_1234_),
    .A(_2156_),
    .B(_1229_));
 sg13g2_xnor2_1 _4768_ (.Y(_1235_),
    .A(\am_sdr0.filt0.xn_2[5] ),
    .B(_1229_));
 sg13g2_inv_1 _4769_ (.Y(_1236_),
    .A(_1235_));
 sg13g2_a21oi_2 _4770_ (.B1(_1236_),
    .Y(_1237_),
    .A2(_1233_),
    .A1(_1231_));
 sg13g2_a21oi_1 _4771_ (.A1(\am_sdr0.filt0.xn_2[7] ),
    .A2(_2156_),
    .Y(_1238_),
    .B1(\am_sdr0.filt0.xn_2[6] ));
 sg13g2_nand3_1 _4772_ (.B(\am_sdr0.filt0.xn_2[6] ),
    .C(_2156_),
    .A(\am_sdr0.filt0.xn_2[7] ),
    .Y(_1239_));
 sg13g2_nand2b_1 _4773_ (.Y(_1240_),
    .B(_1239_),
    .A_N(_1238_));
 sg13g2_o21ai_1 _4774_ (.B1(_1234_),
    .Y(_1241_),
    .A1(_2156_),
    .A2(_0015_));
 sg13g2_and2_1 _4775_ (.A(_1240_),
    .B(_1241_),
    .X(_1242_));
 sg13g2_xor2_1 _4776_ (.B(_1241_),
    .A(_1240_),
    .X(_1243_));
 sg13g2_and2_1 _4777_ (.A(_1237_),
    .B(_1243_),
    .X(_1244_));
 sg13g2_xnor2_1 _4778_ (.Y(_1245_),
    .A(\am_sdr0.filt0.xn_2[7] ),
    .B(_1232_));
 sg13g2_xnor2_1 _4779_ (.Y(_1246_),
    .A(\am_sdr0.filt0.xn_2[5] ),
    .B(\am_sdr0.filt0.xn_2[3] ));
 sg13g2_nor2b_1 _4780_ (.A(\am_sdr0.filt0.xn_2[2] ),
    .B_N(\am_sdr0.filt0.xn_2[4] ),
    .Y(_1247_));
 sg13g2_nand2_1 _4781_ (.Y(_1248_),
    .A(_1246_),
    .B(_1247_));
 sg13g2_xor2_1 _4782_ (.B(_1247_),
    .A(_1246_),
    .X(_1249_));
 sg13g2_nand2_1 _4783_ (.Y(_1250_),
    .A(\am_sdr0.filt0.xn_2[6] ),
    .B(_1249_));
 sg13g2_a21oi_2 _4784_ (.B1(_1245_),
    .Y(_1251_),
    .A2(_1250_),
    .A1(_1248_));
 sg13g2_nand3_1 _4785_ (.B(_1233_),
    .C(_1236_),
    .A(_1231_),
    .Y(_1252_));
 sg13g2_nor2b_1 _4786_ (.A(_1237_),
    .B_N(_1252_),
    .Y(_1253_));
 sg13g2_nand2_1 _4787_ (.Y(_1254_),
    .A(_1251_),
    .B(_1253_));
 sg13g2_nand3_1 _4788_ (.B(_1248_),
    .C(_1250_),
    .A(_1245_),
    .Y(_1255_));
 sg13g2_nand2b_1 _4789_ (.Y(_1256_),
    .B(_1255_),
    .A_N(_1251_));
 sg13g2_xnor2_1 _4790_ (.Y(_1257_),
    .A(\am_sdr0.filt0.xn_2[6] ),
    .B(_1249_));
 sg13g2_xnor2_1 _4791_ (.Y(_1258_),
    .A(\am_sdr0.filt0.xn_2[4] ),
    .B(\am_sdr0.filt0.xn_2[2] ));
 sg13g2_nor2b_1 _4792_ (.A(\am_sdr0.filt0.xn_2[1] ),
    .B_N(\am_sdr0.filt0.xn_2[3] ),
    .Y(_1259_));
 sg13g2_nand2_1 _4793_ (.Y(_1260_),
    .A(_1258_),
    .B(_1259_));
 sg13g2_xor2_1 _4794_ (.B(_1259_),
    .A(_1258_),
    .X(_1261_));
 sg13g2_nand2_1 _4795_ (.Y(_1262_),
    .A(\am_sdr0.filt0.xn_2[5] ),
    .B(_1261_));
 sg13g2_a21oi_2 _4796_ (.B1(_1257_),
    .Y(_1263_),
    .A2(_1262_),
    .A1(_1260_));
 sg13g2_nor2b_1 _4797_ (.A(_1256_),
    .B_N(_1263_),
    .Y(_1264_));
 sg13g2_nand3_1 _4798_ (.B(_1260_),
    .C(_1262_),
    .A(_1257_),
    .Y(_1265_));
 sg13g2_nand2b_1 _4799_ (.Y(_1266_),
    .B(_1265_),
    .A_N(_1263_));
 sg13g2_xnor2_1 _4800_ (.Y(_1267_),
    .A(\am_sdr0.filt0.xn_2[5] ),
    .B(_1261_));
 sg13g2_xnor2_1 _4801_ (.Y(_1268_),
    .A(\am_sdr0.filt0.xn_2[3] ),
    .B(\am_sdr0.filt0.xn_2[1] ));
 sg13g2_nand2_1 _4802_ (.Y(_1269_),
    .A(_2157_),
    .B(_1268_));
 sg13g2_xnor2_1 _4803_ (.Y(_1270_),
    .A(\am_sdr0.filt0.mul_b2[0] ),
    .B(_1268_));
 sg13g2_nand2_1 _4804_ (.Y(_1271_),
    .A(\am_sdr0.filt0.xn_2[4] ),
    .B(_1270_));
 sg13g2_a21oi_1 _4805_ (.A1(_1269_),
    .A2(_1271_),
    .Y(_1272_),
    .B1(_1267_));
 sg13g2_inv_1 _4806_ (.Y(_1273_),
    .A(_1272_));
 sg13g2_nand3_1 _4807_ (.B(_1269_),
    .C(_1271_),
    .A(_1267_),
    .Y(_1274_));
 sg13g2_nand2_1 _4808_ (.Y(_1275_),
    .A(_1273_),
    .B(_1274_));
 sg13g2_inv_1 _4809_ (.Y(_1276_),
    .A(_1275_));
 sg13g2_xnor2_1 _4810_ (.Y(_1277_),
    .A(\am_sdr0.filt0.xn_2[4] ),
    .B(_1270_));
 sg13g2_nand2_1 _4811_ (.Y(_1278_),
    .A(\am_sdr0.filt0.xn_2[2] ),
    .B(\am_sdr0.filt0.mul_b2[0] ));
 sg13g2_nor2_1 _4812_ (.A(_1277_),
    .B(_1278_),
    .Y(_1279_));
 sg13g2_xor2_1 _4813_ (.B(_1278_),
    .A(_1277_),
    .X(_1280_));
 sg13g2_xnor2_1 _4814_ (.Y(_1281_),
    .A(\am_sdr0.filt0.xn_2[1] ),
    .B(\am_sdr0.filt0.mul_b2[0] ));
 sg13g2_nor2_1 _4815_ (.A(\am_sdr0.filt0.xn_2[2] ),
    .B(_2157_),
    .Y(_1282_));
 sg13g2_a21o_1 _4816_ (.A2(_1281_),
    .A1(\am_sdr0.filt0.xn_2[2] ),
    .B1(_1282_),
    .X(_1283_));
 sg13g2_and2_1 _4817_ (.A(\am_sdr0.filt0.xn_2[2] ),
    .B(\am_sdr0.filt0.xn_2[1] ),
    .X(_1284_));
 sg13g2_a22oi_1 _4818_ (.Y(_1285_),
    .B1(_1284_),
    .B2(_2157_),
    .A2(_1283_),
    .A1(\am_sdr0.filt0.xn_2[3] ));
 sg13g2_nor2b_1 _4819_ (.A(_1285_),
    .B_N(_1280_),
    .Y(_1286_));
 sg13g2_nand3b_1 _4820_ (.B(\am_sdr0.filt0.xn_2[1] ),
    .C(_1282_),
    .Y(_1287_),
    .A_N(\am_sdr0.filt0.xn_2[3] ));
 sg13g2_inv_1 _4821_ (.Y(_1288_),
    .A(_1287_));
 sg13g2_xnor2_1 _4822_ (.Y(_1289_),
    .A(_1280_),
    .B(_1285_));
 sg13g2_a21oi_1 _4823_ (.A1(_1288_),
    .A2(_1289_),
    .Y(_1290_),
    .B1(_1286_));
 sg13g2_xnor2_1 _4824_ (.Y(_1291_),
    .A(_1275_),
    .B(_1279_));
 sg13g2_nor2b_1 _4825_ (.A(_1290_),
    .B_N(_1291_),
    .Y(_1292_));
 sg13g2_a21oi_1 _4826_ (.A1(_1276_),
    .A2(_1279_),
    .Y(_1293_),
    .B1(_1292_));
 sg13g2_xnor2_1 _4827_ (.Y(_1294_),
    .A(_1266_),
    .B(_1272_));
 sg13g2_nand2b_1 _4828_ (.Y(_1295_),
    .B(_1294_),
    .A_N(_1293_));
 sg13g2_o21ai_1 _4829_ (.B1(_1295_),
    .Y(_1296_),
    .A1(_1266_),
    .A2(_1273_));
 sg13g2_xnor2_1 _4830_ (.Y(_1297_),
    .A(_1256_),
    .B(_1263_));
 sg13g2_a21oi_1 _4831_ (.A1(_1296_),
    .A2(_1297_),
    .Y(_1298_),
    .B1(_1264_));
 sg13g2_xnor2_1 _4832_ (.Y(_1299_),
    .A(_1251_),
    .B(_1253_));
 sg13g2_o21ai_1 _4833_ (.B1(_1254_),
    .Y(_1300_),
    .A1(_1298_),
    .A2(_1299_));
 sg13g2_xor2_1 _4834_ (.B(_1243_),
    .A(_1237_),
    .X(_1301_));
 sg13g2_a21oi_1 _4835_ (.A1(_1300_),
    .A2(_1301_),
    .Y(_1302_),
    .B1(_1244_));
 sg13g2_o21ai_1 _4836_ (.B1(\am_sdr0.filt0.xn_2[6] ),
    .Y(_1303_),
    .A1(\am_sdr0.filt0.xn_2[7] ),
    .A2(_0015_));
 sg13g2_nand2_1 _4837_ (.Y(_1304_),
    .A(\am_sdr0.filt0.xn_2[7] ),
    .B(_0015_));
 sg13g2_nor2b_1 _4838_ (.A(_1303_),
    .B_N(_1304_),
    .Y(_1305_));
 sg13g2_nor2_1 _4839_ (.A(_1238_),
    .B(_1305_),
    .Y(_1306_));
 sg13g2_nand2b_1 _4840_ (.Y(_1307_),
    .B(_1242_),
    .A_N(_1306_));
 sg13g2_xnor2_1 _4841_ (.Y(_1308_),
    .A(_1242_),
    .B(_1306_));
 sg13g2_nand2b_1 _4842_ (.Y(_1309_),
    .B(_1308_),
    .A_N(_1302_));
 sg13g2_o21ai_1 _4843_ (.B1(_1303_),
    .Y(_1310_),
    .A1(\am_sdr0.filt0.xn_2[5] ),
    .A2(_1304_));
 sg13g2_a21o_1 _4844_ (.A2(_1304_),
    .A1(_1238_),
    .B1(_1310_),
    .X(_1311_));
 sg13g2_nand3_1 _4845_ (.B(_1309_),
    .C(_1311_),
    .A(_1307_),
    .Y(_1312_));
 sg13g2_inv_1 _4846_ (.Y(_1313_),
    .A(net328));
 sg13g2_o21ai_1 _4847_ (.B1(_1168_),
    .Y(_1314_),
    .A1(_1224_),
    .A2(_1226_));
 sg13g2_nand3_1 _4848_ (.B(net327),
    .C(_1314_),
    .A(_1227_),
    .Y(_1315_));
 sg13g2_nand2_1 _4849_ (.Y(_1316_),
    .A(_1222_),
    .B(_1225_));
 sg13g2_o21ai_1 _4850_ (.B1(_1209_),
    .Y(_1317_),
    .A1(_1203_),
    .A2(_1211_));
 sg13g2_nor2_1 _4851_ (.A(_0481_),
    .B(_0522_),
    .Y(_1318_));
 sg13g2_nand2_2 _4852_ (.Y(_1319_),
    .A(net395),
    .B(_0510_));
 sg13g2_nand2_2 _4853_ (.Y(_1320_),
    .A(_1204_),
    .B(_1319_));
 sg13g2_xor2_1 _4854_ (.B(net393),
    .A(net391),
    .X(_1321_));
 sg13g2_nand2_1 _4855_ (.Y(_1322_),
    .A(net379),
    .B(net391));
 sg13g2_o21ai_1 _4856_ (.B1(_1322_),
    .Y(_1323_),
    .A1(net380),
    .A2(_1321_));
 sg13g2_xnor2_1 _4857_ (.Y(_1324_),
    .A(_1320_),
    .B(_1323_));
 sg13g2_nor2_1 _4858_ (.A(_1207_),
    .B(_1324_),
    .Y(_1325_));
 sg13g2_xor2_1 _4859_ (.B(_1324_),
    .A(_1207_),
    .X(_1326_));
 sg13g2_xnor2_1 _4860_ (.Y(_1327_),
    .A(_1318_),
    .B(_1326_));
 sg13g2_nand2b_1 _4861_ (.Y(_1328_),
    .B(_1317_),
    .A_N(_1327_));
 sg13g2_xor2_1 _4862_ (.B(_1327_),
    .A(_1317_),
    .X(_1329_));
 sg13g2_xor2_1 _4863_ (.B(_1329_),
    .A(net342),
    .X(_1330_));
 sg13g2_a21oi_1 _4864_ (.A1(_1202_),
    .A2(_1212_),
    .Y(_1331_),
    .B1(_1214_));
 sg13g2_nor2b_1 _4865_ (.A(_1331_),
    .B_N(_1330_),
    .Y(_1332_));
 sg13g2_xnor2_1 _4866_ (.Y(_1333_),
    .A(_1330_),
    .B(_1331_));
 sg13g2_a21oi_1 _4867_ (.A1(_0541_),
    .A2(_1216_),
    .Y(_1334_),
    .B1(_1218_));
 sg13g2_and2_1 _4868_ (.A(_0726_),
    .B(_1334_),
    .X(_1335_));
 sg13g2_o21ai_1 _4869_ (.B1(_1216_),
    .Y(_1336_),
    .A1(_0540_),
    .A2(_1218_));
 sg13g2_a21oi_2 _4870_ (.B1(_1336_),
    .Y(_1337_),
    .A2(_1335_),
    .A1(_0725_));
 sg13g2_xnor2_1 _4871_ (.Y(_1338_),
    .A(_1333_),
    .B(_1337_));
 sg13g2_inv_1 _4872_ (.Y(_1339_),
    .A(_1338_));
 sg13g2_a21oi_1 _4873_ (.A1(_1172_),
    .A2(_1188_),
    .Y(_1340_),
    .B1(_1187_));
 sg13g2_a21oi_1 _4874_ (.A1(_1183_),
    .A2(_1184_),
    .Y(_1341_),
    .B1(_1182_));
 sg13g2_nand2b_1 _4875_ (.Y(_1342_),
    .B(net349),
    .A_N(_1341_));
 sg13g2_inv_1 _4876_ (.Y(_1343_),
    .A(_1342_));
 sg13g2_xnor2_1 _4877_ (.Y(_1344_),
    .A(net350),
    .B(_1341_));
 sg13g2_a21o_1 _4878_ (.A2(_1185_),
    .A1(_1181_),
    .B1(_1180_),
    .X(_1345_));
 sg13g2_nor2_1 _4879_ (.A(_1175_),
    .B(_1178_),
    .Y(_1346_));
 sg13g2_nor2_1 _4880_ (.A(_0739_),
    .B(_0776_),
    .Y(_1347_));
 sg13g2_a21oi_1 _4881_ (.A1(_2150_),
    .A2(_0776_),
    .Y(_1348_),
    .B1(_1347_));
 sg13g2_xnor2_1 _4882_ (.Y(_1349_),
    .A(_0790_),
    .B(_1348_));
 sg13g2_nor2_1 _4883_ (.A(_1346_),
    .B(_1349_),
    .Y(_1350_));
 sg13g2_xnor2_1 _4884_ (.Y(_1351_),
    .A(_1346_),
    .B(_1349_));
 sg13g2_nor2b_2 _4885_ (.A(_0018_),
    .B_N(net348),
    .Y(_1352_));
 sg13g2_nand2_2 _4886_ (.Y(_1353_),
    .A(net350),
    .B(_2159_));
 sg13g2_xnor2_1 _4887_ (.Y(_1354_),
    .A(net348),
    .B(_0018_));
 sg13g2_xor2_1 _4888_ (.B(_0018_),
    .A(net348),
    .X(_1355_));
 sg13g2_xnor2_1 _4889_ (.Y(_1356_),
    .A(_0786_),
    .B(_1354_));
 sg13g2_nor2_1 _4890_ (.A(_1351_),
    .B(_1356_),
    .Y(_1357_));
 sg13g2_xnor2_1 _4891_ (.Y(_1358_),
    .A(_1351_),
    .B(_1356_));
 sg13g2_nor2b_1 _4892_ (.A(_1358_),
    .B_N(_1345_),
    .Y(_1359_));
 sg13g2_xnor2_1 _4893_ (.Y(_1360_),
    .A(_1345_),
    .B(_1358_));
 sg13g2_xnor2_1 _4894_ (.Y(_1361_),
    .A(_1344_),
    .B(_1360_));
 sg13g2_nor2_1 _4895_ (.A(_1340_),
    .B(_1361_),
    .Y(_1362_));
 sg13g2_xor2_1 _4896_ (.B(_1361_),
    .A(_1340_),
    .X(_1363_));
 sg13g2_nor2b_1 _4897_ (.A(_1170_),
    .B_N(_1363_),
    .Y(_1364_));
 sg13g2_xnor2_1 _4898_ (.Y(_1365_),
    .A(_1170_),
    .B(_1363_));
 sg13g2_nor3_2 _4899_ (.A(_1190_),
    .B(_1192_),
    .C(_1365_),
    .Y(_1366_));
 sg13g2_o21ai_1 _4900_ (.B1(_1365_),
    .Y(_1367_),
    .A1(_1190_),
    .A2(_1192_));
 sg13g2_nor2b_1 _4901_ (.A(_1366_),
    .B_N(_1367_),
    .Y(_1368_));
 sg13g2_a21oi_1 _4902_ (.A1(_1197_),
    .A2(_1200_),
    .Y(_1369_),
    .B1(_1194_));
 sg13g2_xnor2_1 _4903_ (.Y(_1370_),
    .A(_1368_),
    .B(_1369_));
 sg13g2_nor2_1 _4904_ (.A(_1339_),
    .B(_1370_),
    .Y(_1371_));
 sg13g2_xnor2_1 _4905_ (.Y(_1372_),
    .A(_1338_),
    .B(_1370_));
 sg13g2_xnor2_1 _4906_ (.Y(_1373_),
    .A(net347),
    .B(_1372_));
 sg13g2_and2_1 _4907_ (.A(_1316_),
    .B(_1373_),
    .X(_1374_));
 sg13g2_xor2_1 _4908_ (.B(_1373_),
    .A(_1316_),
    .X(_1375_));
 sg13g2_xnor2_1 _4909_ (.Y(_1376_),
    .A(net327),
    .B(_1375_));
 sg13g2_a21oi_1 _4910_ (.A1(_1227_),
    .A2(_1315_),
    .Y(_1377_),
    .B1(_1376_));
 sg13g2_and3_1 _4911_ (.X(_1378_),
    .A(_1227_),
    .B(_1315_),
    .C(_1376_));
 sg13g2_or2_1 _4912_ (.X(_1379_),
    .B(_1378_),
    .A(_1377_));
 sg13g2_nor2_1 _4913_ (.A(_0975_),
    .B(_1160_),
    .Y(_1380_));
 sg13g2_o21ai_1 _4914_ (.B1(_1380_),
    .Y(_1381_),
    .A1(_1156_),
    .A2(_1158_));
 sg13g2_or3_1 _4915_ (.A(_1156_),
    .B(_1158_),
    .C(_1380_),
    .X(_1382_));
 sg13g2_nand3_1 _4916_ (.B(_0713_),
    .C(_0715_),
    .A(_0596_),
    .Y(_1383_));
 sg13g2_nor2b_1 _4917_ (.A(_0716_),
    .B_N(_1383_),
    .Y(_1384_));
 sg13g2_a21oi_2 _4918_ (.B1(_1384_),
    .Y(_1385_),
    .A2(_1382_),
    .A1(_1381_));
 sg13g2_and3_2 _4919_ (.X(_1386_),
    .A(_1381_),
    .B(_1382_),
    .C(_1384_));
 sg13g2_nor2_1 _4920_ (.A(_2155_),
    .B(\am_sdr0.filt0.if_out[5] ),
    .Y(_1387_));
 sg13g2_nand3b_1 _4921_ (.B(_1387_),
    .C(\am_sdr0.filt0.if_out[6] ),
    .Y(_1388_),
    .A_N(\am_sdr0.filt0.if_out[4] ));
 sg13g2_nand2_1 _4922_ (.Y(_1389_),
    .A(\am_sdr0.filt0.if_out[6] ),
    .B(\am_sdr0.filt0.if_out[4] ));
 sg13g2_nand4_1 _4923_ (.B(\am_sdr0.filt0.if_out[6] ),
    .C(\am_sdr0.filt0.if_out[5] ),
    .A(_2155_),
    .Y(_1390_),
    .D(\am_sdr0.filt0.if_out[4] ));
 sg13g2_o21ai_1 _4924_ (.B1(_1390_),
    .Y(_1391_),
    .A1(\am_sdr0.filt0.if_out[6] ),
    .A2(_1387_));
 sg13g2_nand2b_1 _4925_ (.Y(_1392_),
    .B(_1388_),
    .A_N(_1391_));
 sg13g2_nand2_1 _4926_ (.Y(_1393_),
    .A(\am_sdr0.filt0.if_out[4] ),
    .B(\am_sdr0.filt0.if_out[2] ));
 sg13g2_xor2_1 _4927_ (.B(\am_sdr0.filt0.if_out[2] ),
    .A(\am_sdr0.filt0.if_out[4] ),
    .X(_1394_));
 sg13g2_nand2_1 _4928_ (.Y(_1395_),
    .A(\am_sdr0.filt0.if_out[3] ),
    .B(\am_sdr0.filt0.if_out[1] ));
 sg13g2_nand3_1 _4929_ (.B(\am_sdr0.filt0.if_out[1] ),
    .C(_1394_),
    .A(\am_sdr0.filt0.if_out[3] ),
    .Y(_1396_));
 sg13g2_nor2_1 _4930_ (.A(\am_sdr0.filt0.if_out[5] ),
    .B(_1396_),
    .Y(_1397_));
 sg13g2_xor2_1 _4931_ (.B(\am_sdr0.filt0.if_out[1] ),
    .A(\am_sdr0.filt0.if_out[3] ),
    .X(_1398_));
 sg13g2_nand2_1 _4932_ (.Y(_1399_),
    .A(\am_sdr0.filt0.if_out[2] ),
    .B(\am_sdr0.filt0.if_out[0] ));
 sg13g2_nand3_1 _4933_ (.B(\am_sdr0.filt0.if_out[0] ),
    .C(_1398_),
    .A(\am_sdr0.filt0.if_out[2] ),
    .Y(_1400_));
 sg13g2_nor2_1 _4934_ (.A(\am_sdr0.filt0.if_out[4] ),
    .B(_1400_),
    .Y(_1401_));
 sg13g2_nand2_1 _4935_ (.Y(_1402_),
    .A(\am_sdr0.filt0.if_out[5] ),
    .B(\am_sdr0.filt0.if_out[3] ));
 sg13g2_xor2_1 _4936_ (.B(\am_sdr0.filt0.if_out[3] ),
    .A(\am_sdr0.filt0.if_out[5] ),
    .X(_1403_));
 sg13g2_nand2_1 _4937_ (.Y(_1404_),
    .A(_1393_),
    .B(_1396_));
 sg13g2_xnor2_1 _4938_ (.Y(_1405_),
    .A(_1403_),
    .B(_1404_));
 sg13g2_inv_1 _4939_ (.Y(_1406_),
    .A(_1405_));
 sg13g2_a21oi_1 _4940_ (.A1(_1401_),
    .A2(_1406_),
    .Y(_1407_),
    .B1(_1397_));
 sg13g2_xor2_1 _4941_ (.B(\am_sdr0.filt0.if_out[4] ),
    .A(\am_sdr0.filt0.if_out[6] ),
    .X(_1408_));
 sg13g2_nand2b_1 _4942_ (.Y(_1409_),
    .B(_1403_),
    .A_N(_1393_));
 sg13g2_nand2_1 _4943_ (.Y(_1410_),
    .A(_1402_),
    .B(_1409_));
 sg13g2_xnor2_1 _4944_ (.Y(_1411_),
    .A(_1408_),
    .B(_1410_));
 sg13g2_nor2_1 _4945_ (.A(_1407_),
    .B(_1411_),
    .Y(_1412_));
 sg13g2_nor2_1 _4946_ (.A(\am_sdr0.filt0.if_out[6] ),
    .B(_1409_),
    .Y(_1413_));
 sg13g2_nor2_1 _4947_ (.A(_1412_),
    .B(_1413_),
    .Y(_1414_));
 sg13g2_xor2_1 _4948_ (.B(\am_sdr0.filt0.if_out[5] ),
    .A(\am_sdr0.filt0.if_out[7] ),
    .X(_1415_));
 sg13g2_nand2b_1 _4949_ (.Y(_1416_),
    .B(_1408_),
    .A_N(_1402_));
 sg13g2_nand2_1 _4950_ (.Y(_1417_),
    .A(_1389_),
    .B(_1416_));
 sg13g2_xnor2_1 _4951_ (.Y(_1418_),
    .A(_1415_),
    .B(_1417_));
 sg13g2_nor2_1 _4952_ (.A(_1414_),
    .B(_1418_),
    .Y(_1419_));
 sg13g2_nor2_1 _4953_ (.A(\am_sdr0.filt0.if_out[7] ),
    .B(_1416_),
    .Y(_1420_));
 sg13g2_nor2_1 _4954_ (.A(_1419_),
    .B(_1420_),
    .Y(_1421_));
 sg13g2_o21ai_1 _4955_ (.B1(\am_sdr0.filt0.if_out[7] ),
    .Y(_1422_),
    .A1(\am_sdr0.filt0.if_out[6] ),
    .A2(\am_sdr0.filt0.if_out[5] ));
 sg13g2_o21ai_1 _4956_ (.B1(_1422_),
    .Y(_1423_),
    .A1(_1392_),
    .A2(_1421_));
 sg13g2_nor2b_1 _4957_ (.A(_1423_),
    .B_N(_1390_),
    .Y(_1424_));
 sg13g2_or3_1 _4958_ (.A(_1385_),
    .B(_1386_),
    .C(_1424_),
    .X(_1425_));
 sg13g2_nor2b_1 _4959_ (.A(_1385_),
    .B_N(_1425_),
    .Y(_1426_));
 sg13g2_or3_1 _4960_ (.A(_0584_),
    .B(_0716_),
    .C(_0719_),
    .X(_1427_));
 sg13g2_and2_1 _4961_ (.A(_0720_),
    .B(_1427_),
    .X(_1428_));
 sg13g2_nand2b_1 _4962_ (.Y(_1429_),
    .B(_0943_),
    .A_N(_0942_));
 sg13g2_nand2_1 _4963_ (.Y(_1430_),
    .A(_0974_),
    .B(_1381_));
 sg13g2_xnor2_1 _4964_ (.Y(_1431_),
    .A(_1429_),
    .B(_1430_));
 sg13g2_nor2_1 _4965_ (.A(_1428_),
    .B(_1431_),
    .Y(_1432_));
 sg13g2_xor2_1 _4966_ (.B(_1431_),
    .A(_1428_),
    .X(_1433_));
 sg13g2_xnor2_1 _4967_ (.Y(_1434_),
    .A(net347),
    .B(_1433_));
 sg13g2_nor2b_1 _4968_ (.A(_1426_),
    .B_N(_1434_),
    .Y(_1435_));
 sg13g2_xnor2_1 _4969_ (.Y(_1436_),
    .A(_1302_),
    .B(_1308_));
 sg13g2_xnor2_1 _4970_ (.Y(_1437_),
    .A(_1426_),
    .B(_1434_));
 sg13g2_a21o_2 _4971_ (.A2(_1437_),
    .A1(_1436_),
    .B1(_1435_),
    .X(_1438_));
 sg13g2_inv_1 _4972_ (.Y(_1439_),
    .A(_1438_));
 sg13g2_a21o_1 _4973_ (.A2(_1433_),
    .A1(net345),
    .B1(_1432_),
    .X(_1440_));
 sg13g2_xnor2_1 _4974_ (.Y(_1441_),
    .A(_1162_),
    .B(_1163_));
 sg13g2_nor2b_1 _4975_ (.A(_0718_),
    .B_N(_0720_),
    .Y(_1442_));
 sg13g2_xnor2_1 _4976_ (.Y(_1443_),
    .A(_0723_),
    .B(_1442_));
 sg13g2_and2_1 _4977_ (.A(_1441_),
    .B(_1443_),
    .X(_1444_));
 sg13g2_xor2_1 _4978_ (.B(_1443_),
    .A(_1441_),
    .X(_1445_));
 sg13g2_xnor2_1 _4979_ (.Y(_1446_),
    .A(net347),
    .B(_1445_));
 sg13g2_nand2_1 _4980_ (.Y(_1447_),
    .A(_1440_),
    .B(_1446_));
 sg13g2_xnor2_1 _4981_ (.Y(_1448_),
    .A(_1440_),
    .B(_1446_));
 sg13g2_xnor2_1 _4982_ (.Y(_1449_),
    .A(net329),
    .B(_1448_));
 sg13g2_xnor2_1 _4983_ (.Y(_1450_),
    .A(_1151_),
    .B(_1152_));
 sg13g2_nor2_1 _4984_ (.A(_0706_),
    .B(_0707_),
    .Y(_1451_));
 sg13g2_nor2_1 _4985_ (.A(_0623_),
    .B(_0704_),
    .Y(_1452_));
 sg13g2_xnor2_1 _4986_ (.Y(_1453_),
    .A(_1451_),
    .B(_1452_));
 sg13g2_nor2_1 _4987_ (.A(_1450_),
    .B(_1453_),
    .Y(_1454_));
 sg13g2_xnor2_1 _4988_ (.Y(_1455_),
    .A(_1414_),
    .B(_1418_));
 sg13g2_inv_1 _4989_ (.Y(_1456_),
    .A(_1455_));
 sg13g2_xor2_1 _4990_ (.B(_1453_),
    .A(_1450_),
    .X(_1457_));
 sg13g2_a21oi_1 _4991_ (.A1(_1456_),
    .A2(_1457_),
    .Y(_1458_),
    .B1(_1454_));
 sg13g2_xnor2_1 _4992_ (.Y(_1459_),
    .A(_1392_),
    .B(_1421_));
 sg13g2_inv_1 _4993_ (.Y(_1460_),
    .A(_1459_));
 sg13g2_xnor2_1 _4994_ (.Y(_1461_),
    .A(_0710_),
    .B(_0711_));
 sg13g2_or3_1 _4995_ (.A(_1034_),
    .B(_1153_),
    .C(_1154_),
    .X(_1462_));
 sg13g2_o21ai_1 _4996_ (.B1(_1154_),
    .Y(_1463_),
    .A1(_1034_),
    .A2(_1153_));
 sg13g2_nand3_1 _4997_ (.B(_1462_),
    .C(_1463_),
    .A(_1461_),
    .Y(_1464_));
 sg13g2_a21oi_1 _4998_ (.A1(_1462_),
    .A2(_1463_),
    .Y(_1465_),
    .B1(_1461_));
 sg13g2_a21o_1 _4999_ (.A2(_1463_),
    .A1(_1462_),
    .B1(_1461_),
    .X(_1466_));
 sg13g2_and3_1 _5000_ (.X(_1467_),
    .A(_1460_),
    .B(_1464_),
    .C(_1466_));
 sg13g2_a21oi_1 _5001_ (.A1(_1464_),
    .A2(_1466_),
    .Y(_1468_),
    .B1(_1460_));
 sg13g2_nor3_1 _5002_ (.A(_1458_),
    .B(_1467_),
    .C(_1468_),
    .Y(_1469_));
 sg13g2_xor2_1 _5003_ (.B(_1299_),
    .A(_1298_),
    .X(_1470_));
 sg13g2_o21ai_1 _5004_ (.B1(_1458_),
    .Y(_1471_),
    .A1(_1467_),
    .A2(_1468_));
 sg13g2_nor2b_1 _5005_ (.A(_1469_),
    .B_N(_1471_),
    .Y(_1472_));
 sg13g2_a21oi_1 _5006_ (.A1(_1470_),
    .A2(_1471_),
    .Y(_1473_),
    .B1(_1469_));
 sg13g2_xnor2_1 _5007_ (.Y(_1474_),
    .A(_1300_),
    .B(_1301_));
 sg13g2_inv_1 _5008_ (.Y(_1475_),
    .A(_1474_));
 sg13g2_o21ai_1 _5009_ (.B1(_1464_),
    .Y(_1476_),
    .A1(_1459_),
    .A2(_1465_));
 sg13g2_o21ai_1 _5010_ (.B1(_1424_),
    .Y(_1477_),
    .A1(_1385_),
    .A2(_1386_));
 sg13g2_nand3_1 _5011_ (.B(_1476_),
    .C(_1477_),
    .A(_1425_),
    .Y(_1478_));
 sg13g2_a21o_1 _5012_ (.A2(_1477_),
    .A1(_1425_),
    .B1(_1476_),
    .X(_1479_));
 sg13g2_and3_1 _5013_ (.X(_1480_),
    .A(_1475_),
    .B(_1478_),
    .C(_1479_));
 sg13g2_nand3_1 _5014_ (.B(_1478_),
    .C(_1479_),
    .A(_1475_),
    .Y(_1481_));
 sg13g2_a21oi_1 _5015_ (.A1(_1478_),
    .A2(_1479_),
    .Y(_1482_),
    .B1(_1475_));
 sg13g2_nor3_1 _5016_ (.A(_1473_),
    .B(_1480_),
    .C(_1482_),
    .Y(_1483_));
 sg13g2_o21ai_1 _5017_ (.B1(_1473_),
    .Y(_1484_),
    .A1(_1480_),
    .A2(_1482_));
 sg13g2_xor2_1 _5018_ (.B(_1472_),
    .A(_1470_),
    .X(_1485_));
 sg13g2_xnor2_1 _5019_ (.Y(_1486_),
    .A(_0624_),
    .B(_0703_));
 sg13g2_nor2_1 _5020_ (.A(_1057_),
    .B(_1059_),
    .Y(_1487_));
 sg13g2_a21o_1 _5021_ (.A2(_1149_),
    .A1(_1082_),
    .B1(_1487_),
    .X(_1488_));
 sg13g2_nand3_1 _5022_ (.B(_1149_),
    .C(_1487_),
    .A(_1082_),
    .Y(_1489_));
 sg13g2_nand3_1 _5023_ (.B(_1488_),
    .C(_1489_),
    .A(_1486_),
    .Y(_1490_));
 sg13g2_xnor2_1 _5024_ (.Y(_1491_),
    .A(_1407_),
    .B(_1411_));
 sg13g2_inv_1 _5025_ (.Y(_1492_),
    .A(_1491_));
 sg13g2_a21o_1 _5026_ (.A2(_1489_),
    .A1(_1488_),
    .B1(_1486_),
    .X(_1493_));
 sg13g2_nand3_1 _5027_ (.B(_1492_),
    .C(_1493_),
    .A(_1490_),
    .Y(_1494_));
 sg13g2_nand2_1 _5028_ (.Y(_1495_),
    .A(_1490_),
    .B(_1494_));
 sg13g2_xnor2_1 _5029_ (.Y(_1496_),
    .A(_1455_),
    .B(_1457_));
 sg13g2_nand2_1 _5030_ (.Y(_1497_),
    .A(_1495_),
    .B(_1496_));
 sg13g2_xnor2_1 _5031_ (.Y(_1498_),
    .A(_1296_),
    .B(_1297_));
 sg13g2_xnor2_1 _5032_ (.Y(_1499_),
    .A(_1495_),
    .B(_1496_));
 sg13g2_o21ai_1 _5033_ (.B1(_1497_),
    .Y(_1500_),
    .A1(_1498_),
    .A2(_1499_));
 sg13g2_nand2_1 _5034_ (.Y(_1501_),
    .A(_1485_),
    .B(_1500_));
 sg13g2_xor2_1 _5035_ (.B(_1499_),
    .A(_1498_),
    .X(_1502_));
 sg13g2_nand3_1 _5036_ (.B(_1104_),
    .C(_1148_),
    .A(_1083_),
    .Y(_1503_));
 sg13g2_xnor2_1 _5037_ (.Y(_1504_),
    .A(_0698_),
    .B(_0700_));
 sg13g2_a21oi_1 _5038_ (.A1(_1149_),
    .A2(_1503_),
    .Y(_1505_),
    .B1(_1504_));
 sg13g2_xor2_1 _5039_ (.B(_1405_),
    .A(_1401_),
    .X(_1506_));
 sg13g2_and3_1 _5040_ (.X(_1507_),
    .A(_1149_),
    .B(_1503_),
    .C(_1504_));
 sg13g2_or3_1 _5041_ (.A(_1505_),
    .B(_1506_),
    .C(_1507_),
    .X(_1508_));
 sg13g2_nand2b_1 _5042_ (.Y(_1509_),
    .B(_1508_),
    .A_N(_1505_));
 sg13g2_a21o_1 _5043_ (.A2(_1493_),
    .A1(_1490_),
    .B1(_1492_),
    .X(_1510_));
 sg13g2_nand3_1 _5044_ (.B(_1509_),
    .C(_1510_),
    .A(_1494_),
    .Y(_1511_));
 sg13g2_xnor2_1 _5045_ (.Y(_1512_),
    .A(_1293_),
    .B(_1294_));
 sg13g2_a21o_1 _5046_ (.A2(_1510_),
    .A1(_1494_),
    .B1(_1509_),
    .X(_1513_));
 sg13g2_nand3_1 _5047_ (.B(_1512_),
    .C(_1513_),
    .A(_1511_),
    .Y(_1514_));
 sg13g2_nand2_1 _5048_ (.Y(_1515_),
    .A(_1511_),
    .B(_1514_));
 sg13g2_and2_1 _5049_ (.A(_1502_),
    .B(_1515_),
    .X(_1516_));
 sg13g2_xor2_1 _5050_ (.B(_1515_),
    .A(_1502_),
    .X(_1517_));
 sg13g2_a21o_1 _5051_ (.A2(_1513_),
    .A1(_1511_),
    .B1(_1512_),
    .X(_1518_));
 sg13g2_nand3_1 _5052_ (.B(_0677_),
    .C(_0696_),
    .A(_0649_),
    .Y(_1519_));
 sg13g2_nor2b_1 _5053_ (.A(_0697_),
    .B_N(_1519_),
    .Y(_1520_));
 sg13g2_or3_1 _5054_ (.A(_1117_),
    .B(_1146_),
    .C(_1147_),
    .X(_1521_));
 sg13g2_a21oi_1 _5055_ (.A1(_1148_),
    .A2(_1521_),
    .Y(_1522_),
    .B1(_1520_));
 sg13g2_a21o_1 _5056_ (.A2(_1521_),
    .A1(_1148_),
    .B1(_1520_),
    .X(_1523_));
 sg13g2_nand3_1 _5057_ (.B(_1520_),
    .C(_1521_),
    .A(_1148_),
    .Y(_1524_));
 sg13g2_nand2_1 _5058_ (.Y(_1525_),
    .A(_1395_),
    .B(_1400_));
 sg13g2_xor2_1 _5059_ (.B(_1525_),
    .A(_1394_),
    .X(_1526_));
 sg13g2_and3_1 _5060_ (.X(_1527_),
    .A(_1523_),
    .B(_1524_),
    .C(_1526_));
 sg13g2_or2_1 _5061_ (.X(_1528_),
    .B(_1527_),
    .A(_1522_));
 sg13g2_o21ai_1 _5062_ (.B1(_1506_),
    .Y(_1529_),
    .A1(_1505_),
    .A2(_1507_));
 sg13g2_nand3_1 _5063_ (.B(_1528_),
    .C(_1529_),
    .A(_1508_),
    .Y(_1530_));
 sg13g2_a21oi_1 _5064_ (.A1(_1508_),
    .A2(_1529_),
    .Y(_1531_),
    .B1(_1528_));
 sg13g2_a21o_1 _5065_ (.A2(_1529_),
    .A1(_1508_),
    .B1(_1528_),
    .X(_1532_));
 sg13g2_xnor2_1 _5066_ (.Y(_1533_),
    .A(_1290_),
    .B(_1291_));
 sg13g2_inv_1 _5067_ (.Y(_1534_),
    .A(_1533_));
 sg13g2_and3_1 _5068_ (.X(_1535_),
    .A(_1530_),
    .B(_1532_),
    .C(_1533_));
 sg13g2_o21ai_1 _5069_ (.B1(_1530_),
    .Y(_1536_),
    .A1(_1531_),
    .A2(_1534_));
 sg13g2_nand3_1 _5070_ (.B(_1518_),
    .C(_1536_),
    .A(_1514_),
    .Y(_1537_));
 sg13g2_a21oi_1 _5071_ (.A1(_1514_),
    .A2(_1518_),
    .Y(_1538_),
    .B1(_1536_));
 sg13g2_a21oi_1 _5072_ (.A1(_1530_),
    .A2(_1532_),
    .Y(_1539_),
    .B1(_1533_));
 sg13g2_and3_1 _5073_ (.X(_1540_),
    .A(_1128_),
    .B(_1144_),
    .C(_1145_));
 sg13g2_nor2_1 _5074_ (.A(_0676_),
    .B(_0695_),
    .Y(_1541_));
 sg13g2_xor2_1 _5075_ (.B(_1541_),
    .A(_0678_),
    .X(_1542_));
 sg13g2_o21ai_1 _5076_ (.B1(_1542_),
    .Y(_1543_),
    .A1(_1146_),
    .A2(_1540_));
 sg13g2_xnor2_1 _5077_ (.Y(_1544_),
    .A(_1398_),
    .B(_1399_));
 sg13g2_or3_1 _5078_ (.A(_1146_),
    .B(_1540_),
    .C(_1542_),
    .X(_1545_));
 sg13g2_nand3_1 _5079_ (.B(_1544_),
    .C(_1545_),
    .A(_1543_),
    .Y(_1546_));
 sg13g2_and2_1 _5080_ (.A(_1543_),
    .B(_1546_),
    .X(_1547_));
 sg13g2_a21oi_1 _5081_ (.A1(_1523_),
    .A2(_1524_),
    .Y(_1548_),
    .B1(_1526_));
 sg13g2_nor3_1 _5082_ (.A(_1527_),
    .B(_1547_),
    .C(_1548_),
    .Y(_1549_));
 sg13g2_or3_1 _5083_ (.A(_1527_),
    .B(_1547_),
    .C(_1548_),
    .X(_1550_));
 sg13g2_xnor2_1 _5084_ (.Y(_1551_),
    .A(_1287_),
    .B(_1289_));
 sg13g2_o21ai_1 _5085_ (.B1(_1547_),
    .Y(_1552_),
    .A1(_1527_),
    .A2(_1548_));
 sg13g2_and3_1 _5086_ (.X(_1553_),
    .A(_1550_),
    .B(_1551_),
    .C(_1552_));
 sg13g2_nor2_1 _5087_ (.A(_1549_),
    .B(_1553_),
    .Y(_1554_));
 sg13g2_nor3_1 _5088_ (.A(_1535_),
    .B(_1539_),
    .C(_1554_),
    .Y(_1555_));
 sg13g2_nand3_1 _5089_ (.B(_1142_),
    .C(_1143_),
    .A(_1134_),
    .Y(_1556_));
 sg13g2_xnor2_1 _5090_ (.Y(_1557_),
    .A(_0693_),
    .B(_0694_));
 sg13g2_a21o_1 _5091_ (.A2(_1556_),
    .A1(_1144_),
    .B1(_1557_),
    .X(_1558_));
 sg13g2_nand3_1 _5092_ (.B(_1556_),
    .C(_1557_),
    .A(_1144_),
    .Y(_1559_));
 sg13g2_xor2_1 _5093_ (.B(\am_sdr0.filt0.if_out[0] ),
    .A(\am_sdr0.filt0.if_out[2] ),
    .X(_1560_));
 sg13g2_nand3_1 _5094_ (.B(_1559_),
    .C(_1560_),
    .A(_1558_),
    .Y(_1561_));
 sg13g2_nand2_1 _5095_ (.Y(_1562_),
    .A(_1558_),
    .B(_1561_));
 sg13g2_a21o_1 _5096_ (.A2(_1545_),
    .A1(_1543_),
    .B1(_1544_),
    .X(_1563_));
 sg13g2_nand3_1 _5097_ (.B(_1562_),
    .C(_1563_),
    .A(_1546_),
    .Y(_1564_));
 sg13g2_nand2_1 _5098_ (.Y(_1565_),
    .A(\am_sdr0.filt0.xn_2[1] ),
    .B(_1278_));
 sg13g2_nand2_1 _5099_ (.Y(_1566_),
    .A(_1283_),
    .B(_1565_));
 sg13g2_xor2_1 _5100_ (.B(_1566_),
    .A(\am_sdr0.filt0.xn_2[3] ),
    .X(_1567_));
 sg13g2_inv_1 _5101_ (.Y(_1568_),
    .A(_1567_));
 sg13g2_a21o_1 _5102_ (.A2(_1563_),
    .A1(_1546_),
    .B1(_1562_),
    .X(_1569_));
 sg13g2_nand3_1 _5103_ (.B(_1568_),
    .C(_1569_),
    .A(_1564_),
    .Y(_1570_));
 sg13g2_and2_1 _5104_ (.A(_1564_),
    .B(_1570_),
    .X(_1571_));
 sg13g2_a21oi_1 _5105_ (.A1(_1550_),
    .A2(_1552_),
    .Y(_1572_),
    .B1(_1551_));
 sg13g2_o21ai_1 _5106_ (.B1(_1571_),
    .Y(_1573_),
    .A1(_1553_),
    .A2(_1572_));
 sg13g2_nor3_1 _5107_ (.A(_1553_),
    .B(_1571_),
    .C(_1572_),
    .Y(_1574_));
 sg13g2_a21o_1 _5108_ (.A2(_1569_),
    .A1(_1564_),
    .B1(_1568_),
    .X(_1575_));
 sg13g2_xor2_1 _5109_ (.B(_0688_),
    .A(_0687_),
    .X(_1576_));
 sg13g2_xnor2_1 _5110_ (.Y(_1577_),
    .A(_1138_),
    .B(_1139_));
 sg13g2_nor2b_1 _5111_ (.A(_1576_),
    .B_N(_1577_),
    .Y(_1578_));
 sg13g2_xnor2_1 _5112_ (.Y(_1579_),
    .A(_1576_),
    .B(_1577_));
 sg13g2_a21oi_1 _5113_ (.A1(\am_sdr0.filt0.if_out[0] ),
    .A2(_1579_),
    .Y(_1580_),
    .B1(_1578_));
 sg13g2_o21ai_1 _5114_ (.B1(_0689_),
    .Y(_1581_),
    .A1(_0690_),
    .A2(_0691_));
 sg13g2_nand2_2 _5115_ (.Y(_1582_),
    .A(_0692_),
    .B(_1581_));
 sg13g2_or3_1 _5116_ (.A(_1137_),
    .B(_1140_),
    .C(_1141_),
    .X(_1583_));
 sg13g2_and2_1 _5117_ (.A(_1142_),
    .B(_1583_),
    .X(_1584_));
 sg13g2_nand2b_1 _5118_ (.Y(_1585_),
    .B(_1584_),
    .A_N(_1582_));
 sg13g2_xor2_1 _5119_ (.B(_1584_),
    .A(_1582_),
    .X(_1586_));
 sg13g2_nand2b_1 _5120_ (.Y(_1587_),
    .B(_1586_),
    .A_N(_1580_));
 sg13g2_xor2_1 _5121_ (.B(_1586_),
    .A(_1580_),
    .X(_1588_));
 sg13g2_or2_1 _5122_ (.X(_1589_),
    .B(_1588_),
    .A(_1281_));
 sg13g2_xor2_1 _5123_ (.B(_1579_),
    .A(\am_sdr0.filt0.if_out[0] ),
    .X(_1590_));
 sg13g2_a21oi_1 _5124_ (.A1(\am_sdr0.filt0.if_out[1] ),
    .A2(_1590_),
    .Y(_1591_),
    .B1(_2157_));
 sg13g2_a21oi_1 _5125_ (.A1(\am_sdr0.filt0.mul_b2[0] ),
    .A2(_2158_),
    .Y(_1592_),
    .B1(\am_sdr0.filt0.if_out[1] ));
 sg13g2_nand2b_1 _5126_ (.Y(_1593_),
    .B(_1592_),
    .A_N(_1590_));
 sg13g2_o21ai_1 _5127_ (.B1(_1593_),
    .Y(_1594_),
    .A1(_2158_),
    .A2(_1591_));
 sg13g2_xnor2_1 _5128_ (.Y(_1595_),
    .A(_1281_),
    .B(_1588_));
 sg13g2_xnor2_1 _5129_ (.Y(_1596_),
    .A(\am_sdr0.filt0.if_out[1] ),
    .B(\am_sdr0.filt0.mul_b2[0] ));
 sg13g2_nand2_1 _5130_ (.Y(_1597_),
    .A(_1590_),
    .B(_1596_));
 sg13g2_a21o_1 _5131_ (.A2(_1597_),
    .A1(_1595_),
    .B1(_1594_),
    .X(_1598_));
 sg13g2_nand3_1 _5132_ (.B(_1589_),
    .C(_1598_),
    .A(_1587_),
    .Y(_1599_));
 sg13g2_a21o_1 _5133_ (.A2(_1559_),
    .A1(_1558_),
    .B1(_1560_),
    .X(_1600_));
 sg13g2_nand3_1 _5134_ (.B(_1585_),
    .C(_1600_),
    .A(_1561_),
    .Y(_1601_));
 sg13g2_a21o_1 _5135_ (.A2(_1600_),
    .A1(_1561_),
    .B1(_1585_),
    .X(_1602_));
 sg13g2_xnor2_1 _5136_ (.Y(_1603_),
    .A(\am_sdr0.filt0.xn_2[2] ),
    .B(\am_sdr0.filt0.xn_2[1] ));
 sg13g2_a21oi_2 _5137_ (.B1(_1282_),
    .Y(_1604_),
    .A2(_1603_),
    .A1(_2157_));
 sg13g2_nand3_1 _5138_ (.B(_1602_),
    .C(_1604_),
    .A(_1601_),
    .Y(_1605_));
 sg13g2_a21o_1 _5139_ (.A2(_1602_),
    .A1(_1601_),
    .B1(_1604_),
    .X(_1606_));
 sg13g2_a221oi_1 _5140_ (.B2(_1597_),
    .C1(_1594_),
    .B1(_1595_),
    .A1(_1587_),
    .Y(_1607_),
    .A2(_1589_));
 sg13g2_a21o_1 _5141_ (.A2(_1606_),
    .A1(_1605_),
    .B1(_1607_),
    .X(_1608_));
 sg13g2_and2_1 _5142_ (.A(_1601_),
    .B(_1605_),
    .X(_1609_));
 sg13g2_a22oi_1 _5143_ (.Y(_1610_),
    .B1(_1599_),
    .B2(_1608_),
    .A2(_1575_),
    .A1(_1570_));
 sg13g2_nand4_1 _5144_ (.B(_1575_),
    .C(_1599_),
    .A(_1570_),
    .Y(_1611_),
    .D(_1608_));
 sg13g2_a21oi_1 _5145_ (.A1(_1609_),
    .A2(_1611_),
    .Y(_1612_),
    .B1(_1610_));
 sg13g2_a21o_1 _5146_ (.A2(_1612_),
    .A1(_1573_),
    .B1(_1574_),
    .X(_1613_));
 sg13g2_o21ai_1 _5147_ (.B1(_1554_),
    .Y(_1614_),
    .A1(_1535_),
    .A2(_1539_));
 sg13g2_a21oi_1 _5148_ (.A1(_1613_),
    .A2(_1614_),
    .Y(_1615_),
    .B1(_1555_));
 sg13g2_o21ai_1 _5149_ (.B1(_1537_),
    .Y(_1616_),
    .A1(_1538_),
    .A2(_1615_));
 sg13g2_a21oi_1 _5150_ (.A1(_1517_),
    .A2(_1616_),
    .Y(_1617_),
    .B1(_1516_));
 sg13g2_xnor2_1 _5151_ (.Y(_1618_),
    .A(_1485_),
    .B(_1500_));
 sg13g2_or2_1 _5152_ (.X(_1619_),
    .B(_1618_),
    .A(_1617_));
 sg13g2_nand2_1 _5153_ (.Y(_1620_),
    .A(_1501_),
    .B(_1619_));
 sg13g2_a21oi_1 _5154_ (.A1(_1485_),
    .A2(_1500_),
    .Y(_1621_),
    .B1(_1483_));
 sg13g2_o21ai_1 _5155_ (.B1(_1621_),
    .Y(_1622_),
    .A1(_1617_),
    .A2(_1618_));
 sg13g2_nand2_1 _5156_ (.Y(_1623_),
    .A(_1484_),
    .B(_1622_));
 sg13g2_xnor2_1 _5157_ (.Y(_1624_),
    .A(_1436_),
    .B(_1437_));
 sg13g2_nand2_1 _5158_ (.Y(_1625_),
    .A(_1478_),
    .B(_1481_));
 sg13g2_nor2b_2 _5159_ (.A(_1624_),
    .B_N(_1625_),
    .Y(_1626_));
 sg13g2_xnor2_1 _5160_ (.Y(_1627_),
    .A(_1624_),
    .B(_1625_));
 sg13g2_nand3_1 _5161_ (.B(_1622_),
    .C(_1627_),
    .A(_1484_),
    .Y(_1628_));
 sg13g2_nor2b_1 _5162_ (.A(_1449_),
    .B_N(_1438_),
    .Y(_1629_));
 sg13g2_nor2_1 _5163_ (.A(_1626_),
    .B(_1629_),
    .Y(_1630_));
 sg13g2_xor2_1 _5164_ (.B(_1449_),
    .A(_1438_),
    .X(_1631_));
 sg13g2_a22oi_1 _5165_ (.Y(_1632_),
    .B1(_1628_),
    .B2(_1630_),
    .A2(_1449_),
    .A1(_1439_));
 sg13g2_a21o_1 _5166_ (.A2(_1445_),
    .A1(net345),
    .B1(_1444_),
    .X(_1633_));
 sg13g2_xnor2_1 _5167_ (.Y(_1634_),
    .A(net347),
    .B(_1167_));
 sg13g2_nand2_1 _5168_ (.Y(_1635_),
    .A(_1633_),
    .B(_1634_));
 sg13g2_xnor2_1 _5169_ (.Y(_1636_),
    .A(_1633_),
    .B(_1634_));
 sg13g2_o21ai_1 _5170_ (.B1(_1635_),
    .Y(_1637_),
    .A1(net329),
    .A2(_1636_));
 sg13g2_a21o_1 _5171_ (.A2(_1314_),
    .A1(_1227_),
    .B1(net327),
    .X(_1638_));
 sg13g2_and3_1 _5172_ (.X(_1639_),
    .A(_1315_),
    .B(_1637_),
    .C(_1638_));
 sg13g2_nand3_1 _5173_ (.B(_1637_),
    .C(_1638_),
    .A(_1315_),
    .Y(_1640_));
 sg13g2_a21o_1 _5174_ (.A2(_1638_),
    .A1(_1315_),
    .B1(_1637_),
    .X(_1641_));
 sg13g2_and2_1 _5175_ (.A(_1640_),
    .B(_1641_),
    .X(_1642_));
 sg13g2_xnor2_1 _5176_ (.Y(_1643_),
    .A(net326),
    .B(_1636_));
 sg13g2_o21ai_1 _5177_ (.B1(_1447_),
    .Y(_1644_),
    .A1(net328),
    .A2(_1448_));
 sg13g2_and2_1 _5178_ (.A(_1643_),
    .B(_1644_),
    .X(_1645_));
 sg13g2_xor2_1 _5179_ (.B(_1644_),
    .A(_1643_),
    .X(_1646_));
 sg13g2_nand3_1 _5180_ (.B(_1641_),
    .C(_1646_),
    .A(_1640_),
    .Y(_1647_));
 sg13g2_a221oi_1 _5181_ (.B2(_1630_),
    .C1(_1647_),
    .B1(_1628_),
    .A1(_1439_),
    .Y(_1648_),
    .A2(_1449_));
 sg13g2_and2_1 _5182_ (.A(_1641_),
    .B(_1645_),
    .X(_1649_));
 sg13g2_nor3_1 _5183_ (.A(_1639_),
    .B(_1648_),
    .C(_1649_),
    .Y(_1650_));
 sg13g2_nor2_1 _5184_ (.A(_1379_),
    .B(_1650_),
    .Y(_1651_));
 sg13g2_xor2_1 _5185_ (.B(_1650_),
    .A(_1379_),
    .X(_1652_));
 sg13g2_nand2_1 _5186_ (.Y(_1653_),
    .A(_0478_),
    .B(_1652_));
 sg13g2_nand2_1 _5187_ (.Y(_1654_),
    .A(\am_sdr0.filt0.gain_spi[0] ),
    .B(net440));
 sg13g2_nor2_2 _5188_ (.A(net437),
    .B(_1654_),
    .Y(_1655_));
 sg13g2_a21oi_1 _5189_ (.A1(_1632_),
    .A2(_1646_),
    .Y(_1656_),
    .B1(_1645_));
 sg13g2_xnor2_1 _5190_ (.Y(_1657_),
    .A(_1642_),
    .B(_1656_));
 sg13g2_nand2_1 _5191_ (.Y(_1658_),
    .A(\am_sdr0.filt0.gain_spi[1] ),
    .B(_0017_));
 sg13g2_and3_2 _5192_ (.X(_1659_),
    .A(\am_sdr0.filt0.gain_spi[1] ),
    .B(\am_sdr0.filt0.gain_spi[0] ),
    .C(_0017_));
 sg13g2_nor2b_1 _5193_ (.A(_1626_),
    .B_N(_1628_),
    .Y(_1660_));
 sg13g2_xnor2_1 _5194_ (.Y(_1661_),
    .A(_1631_),
    .B(_1660_));
 sg13g2_inv_1 _5195_ (.Y(_1662_),
    .A(_1661_));
 sg13g2_and2_2 _5196_ (.A(net246),
    .B(_0477_),
    .X(_1663_));
 sg13g2_nand2_1 _5197_ (.Y(_1664_),
    .A(net246),
    .B(_0477_));
 sg13g2_nor2_2 _5198_ (.A(net439),
    .B(_1663_),
    .Y(_1665_));
 sg13g2_nand2b_1 _5199_ (.Y(_1666_),
    .B(_1664_),
    .A_N(_0017_));
 sg13g2_xnor2_1 _5200_ (.Y(_1667_),
    .A(_1623_),
    .B(_1627_));
 sg13g2_a22oi_1 _5201_ (.Y(_1668_),
    .B1(_1663_),
    .B2(_1667_),
    .A2(_1662_),
    .A1(_1659_));
 sg13g2_nor2_2 _5202_ (.A(\am_sdr0.filt0.gain_spi[0] ),
    .B(_1658_),
    .Y(_1669_));
 sg13g2_xor2_1 _5203_ (.B(_1646_),
    .A(_1632_),
    .X(_1670_));
 sg13g2_a22oi_1 _5204_ (.Y(_1671_),
    .B1(_1669_),
    .B2(_1670_),
    .A2(_1657_),
    .A1(_1655_));
 sg13g2_and3_1 _5205_ (.X(_1672_),
    .A(_1666_),
    .B(_1668_),
    .C(_1671_));
 sg13g2_nor2b_1 _5206_ (.A(_1483_),
    .B_N(_1484_),
    .Y(_1673_));
 sg13g2_xnor2_1 _5207_ (.Y(_1674_),
    .A(_1620_),
    .B(_1673_));
 sg13g2_a221oi_1 _5208_ (.B2(_1665_),
    .C1(net406),
    .B1(_1674_),
    .A1(_1653_),
    .Y(_0108_),
    .A2(_1672_));
 sg13g2_nor2_1 _5209_ (.A(_1377_),
    .B(_1651_),
    .Y(_1675_));
 sg13g2_a21oi_1 _5210_ (.A1(net326),
    .A2(_1375_),
    .Y(_1676_),
    .B1(_1374_));
 sg13g2_a21o_1 _5211_ (.A2(_1375_),
    .A1(net326),
    .B1(_1374_),
    .X(_1677_));
 sg13g2_a21o_1 _5212_ (.A2(_1372_),
    .A1(net345),
    .B1(_1371_),
    .X(_1678_));
 sg13g2_a21oi_1 _5213_ (.A1(_1344_),
    .A2(_1360_),
    .Y(_1679_),
    .B1(_1359_));
 sg13g2_o21ai_1 _5214_ (.B1(_1354_),
    .Y(_1680_),
    .A1(net348),
    .A2(_0786_));
 sg13g2_a21oi_1 _5215_ (.A1(net348),
    .A2(_0786_),
    .Y(_1681_),
    .B1(_1680_));
 sg13g2_nor2_1 _5216_ (.A(_1350_),
    .B(_1357_),
    .Y(_1682_));
 sg13g2_a22oi_1 _5217_ (.Y(_1683_),
    .B1(_0790_),
    .B2(_1348_),
    .A2(_0776_),
    .A1(_2150_));
 sg13g2_a21oi_1 _5218_ (.A1(_2150_),
    .A2(_2151_),
    .Y(_1684_),
    .B1(_0958_));
 sg13g2_nor2b_1 _5219_ (.A(_0815_),
    .B_N(_1684_),
    .Y(_1685_));
 sg13g2_xnor2_1 _5220_ (.Y(_1686_),
    .A(_0815_),
    .B(_1684_));
 sg13g2_nor2b_1 _5221_ (.A(_1683_),
    .B_N(_1686_),
    .Y(_1687_));
 sg13g2_xnor2_1 _5222_ (.Y(_1688_),
    .A(_1683_),
    .B(_1686_));
 sg13g2_xnor2_1 _5223_ (.Y(_1689_),
    .A(_0819_),
    .B(_1688_));
 sg13g2_nor2_1 _5224_ (.A(_1682_),
    .B(_1689_),
    .Y(_1690_));
 sg13g2_xor2_1 _5225_ (.B(_1689_),
    .A(_1682_),
    .X(_1691_));
 sg13g2_xnor2_1 _5226_ (.Y(_1692_),
    .A(_1681_),
    .B(_1691_));
 sg13g2_nor2_1 _5227_ (.A(_1679_),
    .B(_1692_),
    .Y(_1693_));
 sg13g2_xor2_1 _5228_ (.B(_1692_),
    .A(_1679_),
    .X(_1694_));
 sg13g2_xnor2_1 _5229_ (.Y(_1695_),
    .A(_1342_),
    .B(_1694_));
 sg13g2_nor2_1 _5230_ (.A(_1362_),
    .B(_1364_),
    .Y(_1696_));
 sg13g2_nor2b_1 _5231_ (.A(_1696_),
    .B_N(_1695_),
    .Y(_1697_));
 sg13g2_xnor2_1 _5232_ (.Y(_1698_),
    .A(_1695_),
    .B(_1696_));
 sg13g2_nand2b_1 _5233_ (.Y(_1699_),
    .B(_1194_),
    .A_N(_1366_));
 sg13g2_and3_1 _5234_ (.X(_1700_),
    .A(_1199_),
    .B(_1367_),
    .C(_1699_));
 sg13g2_o21ai_1 _5235_ (.B1(_1700_),
    .Y(_1701_),
    .A1(_1162_),
    .A2(_1198_));
 sg13g2_o21ai_1 _5236_ (.B1(_1367_),
    .Y(_1702_),
    .A1(_1196_),
    .A2(_1366_));
 sg13g2_nand2_1 _5237_ (.Y(_1703_),
    .A(_1701_),
    .B(_1702_));
 sg13g2_nand3_1 _5238_ (.B(_1701_),
    .C(_1702_),
    .A(_1698_),
    .Y(_1704_));
 sg13g2_xor2_1 _5239_ (.B(_1703_),
    .A(_1698_),
    .X(_1705_));
 sg13g2_o21ai_1 _5240_ (.B1(_1328_),
    .Y(_1706_),
    .A1(net341),
    .A2(_1329_));
 sg13g2_a21oi_1 _5241_ (.A1(_1318_),
    .A2(_1326_),
    .Y(_1707_),
    .B1(_1325_));
 sg13g2_nand3_1 _5242_ (.B(net391),
    .C(net393),
    .A(net380),
    .Y(_1708_));
 sg13g2_o21ai_1 _5243_ (.B1(_1708_),
    .Y(_1709_),
    .A1(_1320_),
    .A2(_1323_));
 sg13g2_nor2_1 _5244_ (.A(net391),
    .B(_0639_),
    .Y(_1710_));
 sg13g2_a21oi_1 _5245_ (.A1(net390),
    .A2(net391),
    .Y(_1711_),
    .B1(_1710_));
 sg13g2_nand2_2 _5246_ (.Y(_1712_),
    .A(net380),
    .B(_1711_));
 sg13g2_nand3_1 _5247_ (.B(net390),
    .C(_1321_),
    .A(net380),
    .Y(_1713_));
 sg13g2_o21ai_1 _5248_ (.B1(_1713_),
    .Y(_1714_),
    .A1(net379),
    .A2(_1711_));
 sg13g2_inv_1 _5249_ (.Y(_1715_),
    .A(_1714_));
 sg13g2_o21ai_1 _5250_ (.B1(_1715_),
    .Y(_1716_),
    .A1(_1321_),
    .A2(_1712_));
 sg13g2_xnor2_1 _5251_ (.Y(_1717_),
    .A(_1320_),
    .B(_1716_));
 sg13g2_nand2b_1 _5252_ (.Y(_1718_),
    .B(_1709_),
    .A_N(_1717_));
 sg13g2_xor2_1 _5253_ (.B(_1717_),
    .A(_1709_),
    .X(_1719_));
 sg13g2_xnor2_1 _5254_ (.Y(_1720_),
    .A(_1319_),
    .B(_1719_));
 sg13g2_xor2_1 _5255_ (.B(_1720_),
    .A(_1707_),
    .X(_1721_));
 sg13g2_nand2b_1 _5256_ (.Y(_1722_),
    .B(_1721_),
    .A_N(net341));
 sg13g2_xnor2_1 _5257_ (.Y(_1723_),
    .A(net341),
    .B(_1721_));
 sg13g2_and2_1 _5258_ (.A(_1706_),
    .B(_1723_),
    .X(_1724_));
 sg13g2_or2_1 _5259_ (.X(_1725_),
    .B(_1723_),
    .A(_1706_));
 sg13g2_nor2b_1 _5260_ (.A(_1724_),
    .B_N(_1725_),
    .Y(_1726_));
 sg13g2_a21oi_1 _5261_ (.A1(_1333_),
    .A2(_1337_),
    .Y(_1727_),
    .B1(_1332_));
 sg13g2_xor2_1 _5262_ (.B(_1727_),
    .A(_1726_),
    .X(_1728_));
 sg13g2_nand2_1 _5263_ (.Y(_1729_),
    .A(_1705_),
    .B(_1728_));
 sg13g2_xnor2_1 _5264_ (.Y(_1730_),
    .A(_1705_),
    .B(_1728_));
 sg13g2_xnor2_1 _5265_ (.Y(_1731_),
    .A(net344),
    .B(_1730_));
 sg13g2_nand2_1 _5266_ (.Y(_1732_),
    .A(_1678_),
    .B(_1731_));
 sg13g2_xnor2_1 _5267_ (.Y(_1733_),
    .A(_1678_),
    .B(_1731_));
 sg13g2_xnor2_1 _5268_ (.Y(_1734_),
    .A(net326),
    .B(_1733_));
 sg13g2_xnor2_1 _5269_ (.Y(_1735_),
    .A(net328),
    .B(_1733_));
 sg13g2_nor2_1 _5270_ (.A(_1676_),
    .B(_1735_),
    .Y(_1736_));
 sg13g2_nand2_1 _5271_ (.Y(_1737_),
    .A(_1677_),
    .B(_1734_));
 sg13g2_nor2_1 _5272_ (.A(_1677_),
    .B(_1734_),
    .Y(_1738_));
 sg13g2_nor2_1 _5273_ (.A(_1736_),
    .B(_1738_),
    .Y(_1739_));
 sg13g2_xor2_1 _5274_ (.B(_1739_),
    .A(_1675_),
    .X(_1740_));
 sg13g2_nand2b_1 _5275_ (.Y(_1741_),
    .B(_0478_),
    .A_N(_1740_));
 sg13g2_a22oi_1 _5276_ (.Y(_1742_),
    .B1(_1670_),
    .B2(_1659_),
    .A2(_1663_),
    .A1(_1662_));
 sg13g2_a22oi_1 _5277_ (.Y(_1743_),
    .B1(_1657_),
    .B2(_1669_),
    .A2(_1655_),
    .A1(_1652_));
 sg13g2_nand4_1 _5278_ (.B(_1741_),
    .C(_1742_),
    .A(net333),
    .Y(_1744_),
    .D(_1743_));
 sg13g2_o21ai_1 _5279_ (.B1(net411),
    .Y(_1745_),
    .A1(_1666_),
    .A2(_1667_));
 sg13g2_nor2b_1 _5280_ (.A(_1745_),
    .B_N(_1744_),
    .Y(_0109_));
 sg13g2_o21ai_1 _5281_ (.B1(_1729_),
    .Y(_1746_),
    .A1(net347),
    .A2(_1730_));
 sg13g2_o21ai_1 _5282_ (.B1(_1722_),
    .Y(_1747_),
    .A1(_1707_),
    .A2(_1720_));
 sg13g2_o21ai_1 _5283_ (.B1(_1718_),
    .Y(_1748_),
    .A1(_1319_),
    .A2(_1719_));
 sg13g2_o21ai_1 _5284_ (.B1(_1713_),
    .Y(_1749_),
    .A1(_1320_),
    .A2(_1716_));
 sg13g2_o21ai_1 _5285_ (.B1(_0606_),
    .Y(_1750_),
    .A1(net391),
    .A2(_0638_));
 sg13g2_xor2_1 _5286_ (.B(net388),
    .A(net379),
    .X(_1751_));
 sg13g2_nor2_1 _5287_ (.A(_1750_),
    .B(_1751_),
    .Y(_1752_));
 sg13g2_xor2_1 _5288_ (.B(_1751_),
    .A(_1750_),
    .X(_1753_));
 sg13g2_xnor2_1 _5289_ (.Y(_1754_),
    .A(_1712_),
    .B(_1753_));
 sg13g2_xnor2_1 _5290_ (.Y(_1755_),
    .A(_0481_),
    .B(_0524_));
 sg13g2_nor2_1 _5291_ (.A(_0606_),
    .B(_1755_),
    .Y(_1756_));
 sg13g2_nand2_1 _5292_ (.Y(_1757_),
    .A(_0606_),
    .B(_1755_));
 sg13g2_nand2b_1 _5293_ (.Y(_1758_),
    .B(_1757_),
    .A_N(_1756_));
 sg13g2_a21oi_2 _5294_ (.B1(_0523_),
    .Y(_1759_),
    .A2(_0522_),
    .A1(_0481_));
 sg13g2_xor2_1 _5295_ (.B(_1759_),
    .A(_1758_),
    .X(_1760_));
 sg13g2_or2_1 _5296_ (.X(_1761_),
    .B(_1760_),
    .A(_1754_));
 sg13g2_xor2_1 _5297_ (.B(_1760_),
    .A(_1754_),
    .X(_1762_));
 sg13g2_nand2_1 _5298_ (.Y(_1763_),
    .A(_1749_),
    .B(_1762_));
 sg13g2_xnor2_1 _5299_ (.Y(_1764_),
    .A(_1749_),
    .B(_1762_));
 sg13g2_xnor2_1 _5300_ (.Y(_1765_),
    .A(_1319_),
    .B(_1764_));
 sg13g2_nand2b_1 _5301_ (.Y(_1766_),
    .B(_1748_),
    .A_N(_1765_));
 sg13g2_xor2_1 _5302_ (.B(_1765_),
    .A(_1748_),
    .X(_1767_));
 sg13g2_xor2_1 _5303_ (.B(_1767_),
    .A(net341),
    .X(_1768_));
 sg13g2_nand2_1 _5304_ (.Y(_1769_),
    .A(_1747_),
    .B(_1768_));
 sg13g2_xnor2_1 _5305_ (.Y(_1770_),
    .A(_1747_),
    .B(_1768_));
 sg13g2_and2_1 _5306_ (.A(_1333_),
    .B(_1726_),
    .X(_1771_));
 sg13g2_a221oi_1 _5307_ (.B2(_1337_),
    .C1(_1724_),
    .B1(_1771_),
    .A1(_1332_),
    .Y(_1772_),
    .A2(_1725_));
 sg13g2_xor2_1 _5308_ (.B(_1772_),
    .A(_1770_),
    .X(_1773_));
 sg13g2_nor2b_1 _5309_ (.A(_1697_),
    .B_N(_1704_),
    .Y(_1774_));
 sg13g2_a21oi_1 _5310_ (.A1(_1343_),
    .A2(_1694_),
    .Y(_1775_),
    .B1(_1693_));
 sg13g2_a21o_1 _5311_ (.A2(_0786_),
    .A1(net348),
    .B1(_1352_),
    .X(_1776_));
 sg13g2_a21oi_1 _5312_ (.A1(_1681_),
    .A2(_1691_),
    .Y(_1777_),
    .B1(_1690_));
 sg13g2_a21oi_1 _5313_ (.A1(_0819_),
    .A2(_1688_),
    .Y(_1778_),
    .B1(_1687_));
 sg13g2_a21oi_1 _5314_ (.A1(net358),
    .A2(_0735_),
    .Y(_1779_),
    .B1(_0857_));
 sg13g2_nor2_1 _5315_ (.A(_2154_),
    .B(_1779_),
    .Y(_1780_));
 sg13g2_xnor2_1 _5316_ (.Y(_1781_),
    .A(net352),
    .B(_1779_));
 sg13g2_a21oi_1 _5317_ (.A1(_2151_),
    .A2(_0738_),
    .Y(_1782_),
    .B1(_1685_));
 sg13g2_nor2b_1 _5318_ (.A(_1782_),
    .B_N(_1781_),
    .Y(_1783_));
 sg13g2_xnor2_1 _5319_ (.Y(_1784_),
    .A(_1781_),
    .B(_1782_));
 sg13g2_xnor2_1 _5320_ (.Y(_1785_),
    .A(_1184_),
    .B(_1784_));
 sg13g2_nor2_1 _5321_ (.A(_1778_),
    .B(_1785_),
    .Y(_1786_));
 sg13g2_xor2_1 _5322_ (.B(_1785_),
    .A(_1778_),
    .X(_1787_));
 sg13g2_xnor2_1 _5323_ (.Y(_1788_),
    .A(_1354_),
    .B(_1787_));
 sg13g2_nor2_1 _5324_ (.A(_1777_),
    .B(_1788_),
    .Y(_1789_));
 sg13g2_xor2_1 _5325_ (.B(_1788_),
    .A(_1777_),
    .X(_1790_));
 sg13g2_xnor2_1 _5326_ (.Y(_1791_),
    .A(_1776_),
    .B(_1790_));
 sg13g2_nor2_1 _5327_ (.A(_1775_),
    .B(_1791_),
    .Y(_1792_));
 sg13g2_xor2_1 _5328_ (.B(_1791_),
    .A(_1775_),
    .X(_1793_));
 sg13g2_xor2_1 _5329_ (.B(_1793_),
    .A(_1774_),
    .X(_1794_));
 sg13g2_nand2b_1 _5330_ (.Y(_1795_),
    .B(_1794_),
    .A_N(_1773_));
 sg13g2_xor2_1 _5331_ (.B(_1794_),
    .A(_1773_),
    .X(_1796_));
 sg13g2_xnor2_1 _5332_ (.Y(_1797_),
    .A(net344),
    .B(_1796_));
 sg13g2_nand2_1 _5333_ (.Y(_1798_),
    .A(_1746_),
    .B(_1797_));
 sg13g2_xnor2_1 _5334_ (.Y(_1799_),
    .A(_1746_),
    .B(_1797_));
 sg13g2_xnor2_1 _5335_ (.Y(_1800_),
    .A(net327),
    .B(_1799_));
 sg13g2_o21ai_1 _5336_ (.B1(_1732_),
    .Y(_1801_),
    .A1(net329),
    .A2(_1733_));
 sg13g2_and2_1 _5337_ (.A(_1800_),
    .B(_1801_),
    .X(_1802_));
 sg13g2_nand2_1 _5338_ (.Y(_1803_),
    .A(_1800_),
    .B(_1801_));
 sg13g2_xnor2_1 _5339_ (.Y(_1804_),
    .A(_1800_),
    .B(_1801_));
 sg13g2_a221oi_1 _5340_ (.B2(_1735_),
    .C1(_1376_),
    .B1(_1676_),
    .A1(_1227_),
    .Y(_1805_),
    .A2(_1315_));
 sg13g2_or4_1 _5341_ (.A(_1639_),
    .B(_1649_),
    .C(_1736_),
    .D(_1805_),
    .X(_1806_));
 sg13g2_a21oi_1 _5342_ (.A1(_1378_),
    .A2(_1737_),
    .Y(_1807_),
    .B1(_1738_));
 sg13g2_o21ai_1 _5343_ (.B1(_1807_),
    .Y(_1808_),
    .A1(_1648_),
    .A2(_1806_));
 sg13g2_xor2_1 _5344_ (.B(_1808_),
    .A(_1804_),
    .X(_1809_));
 sg13g2_nand2b_1 _5345_ (.Y(_1810_),
    .B(_1655_),
    .A_N(_1740_));
 sg13g2_a22oi_1 _5346_ (.Y(_1811_),
    .B1(_1663_),
    .B2(_1670_),
    .A2(_1659_),
    .A1(_1657_));
 sg13g2_a22oi_1 _5347_ (.Y(_1812_),
    .B1(_1809_),
    .B2(_0478_),
    .A2(_1669_),
    .A1(_1652_));
 sg13g2_and3_1 _5348_ (.X(_1813_),
    .A(net333),
    .B(_1811_),
    .C(_1812_));
 sg13g2_a221oi_1 _5349_ (.B2(_1813_),
    .C1(net406),
    .B1(_1810_),
    .A1(_1661_),
    .Y(_0110_),
    .A2(_1665_));
 sg13g2_and2_1 _5350_ (.A(net411),
    .B(_1657_),
    .X(_0122_));
 sg13g2_nand2_1 _5351_ (.Y(_1814_),
    .A(_1663_),
    .B(_0122_));
 sg13g2_o21ai_1 _5352_ (.B1(_1798_),
    .Y(_1815_),
    .A1(net329),
    .A2(_1799_));
 sg13g2_o21ai_1 _5353_ (.B1(_1795_),
    .Y(_1816_),
    .A1(net346),
    .A2(_1796_));
 sg13g2_nand2_1 _5354_ (.Y(_1817_),
    .A(_1698_),
    .B(_1793_));
 sg13g2_a21oi_1 _5355_ (.A1(_1697_),
    .A2(_1793_),
    .Y(_1818_),
    .B1(_1792_));
 sg13g2_o21ai_1 _5356_ (.B1(_1818_),
    .Y(_1819_),
    .A1(_1703_),
    .A2(_1817_));
 sg13g2_a21oi_1 _5357_ (.A1(_1776_),
    .A2(_1790_),
    .Y(_1820_),
    .B1(_1789_));
 sg13g2_a21oi_1 _5358_ (.A1(_1354_),
    .A2(_1787_),
    .Y(_1821_),
    .B1(_1786_));
 sg13g2_a21oi_1 _5359_ (.A1(_1184_),
    .A2(_1784_),
    .Y(_1822_),
    .B1(_1783_));
 sg13g2_a21oi_1 _5360_ (.A1(_2153_),
    .A2(_0785_),
    .Y(_1823_),
    .B1(_1780_));
 sg13g2_xor2_1 _5361_ (.B(_0852_),
    .A(net349),
    .X(_1824_));
 sg13g2_mux2_1 _5362_ (.A0(net349),
    .A1(_1824_),
    .S(_0789_),
    .X(_1825_));
 sg13g2_nor2_1 _5363_ (.A(_1823_),
    .B(_1825_),
    .Y(_1826_));
 sg13g2_xor2_1 _5364_ (.B(_1825_),
    .A(_1823_),
    .X(_1827_));
 sg13g2_xnor2_1 _5365_ (.Y(_1828_),
    .A(net348),
    .B(_1827_));
 sg13g2_nor2_1 _5366_ (.A(_1822_),
    .B(_1828_),
    .Y(_1829_));
 sg13g2_xor2_1 _5367_ (.B(_1828_),
    .A(_1822_),
    .X(_1830_));
 sg13g2_xnor2_1 _5368_ (.Y(_1831_),
    .A(_1355_),
    .B(_1830_));
 sg13g2_nor2b_1 _5369_ (.A(_1821_),
    .B_N(_1831_),
    .Y(_1832_));
 sg13g2_xnor2_1 _5370_ (.Y(_1833_),
    .A(_1821_),
    .B(_1831_));
 sg13g2_xnor2_1 _5371_ (.Y(_1834_),
    .A(_1352_),
    .B(_1833_));
 sg13g2_nor2_1 _5372_ (.A(_1820_),
    .B(_1834_),
    .Y(_1835_));
 sg13g2_xor2_1 _5373_ (.B(_1834_),
    .A(_1820_),
    .X(_1836_));
 sg13g2_xnor2_1 _5374_ (.Y(_1837_),
    .A(_1819_),
    .B(_1836_));
 sg13g2_o21ai_1 _5375_ (.B1(_1769_),
    .Y(_1838_),
    .A1(_1770_),
    .A2(_1772_));
 sg13g2_o21ai_1 _5376_ (.B1(_1766_),
    .Y(_1839_),
    .A1(net341),
    .A2(_1767_));
 sg13g2_o21ai_1 _5377_ (.B1(_1763_),
    .Y(_1840_),
    .A1(_1319_),
    .A2(_1764_));
 sg13g2_a21oi_2 _5378_ (.B1(_1756_),
    .Y(_1841_),
    .A2(_1759_),
    .A1(_1757_));
 sg13g2_o21ai_1 _5379_ (.B1(_1761_),
    .Y(_1842_),
    .A1(_1712_),
    .A2(_1753_));
 sg13g2_nand2_1 _5380_ (.Y(_1843_),
    .A(net386),
    .B(net388));
 sg13g2_xor2_1 _5381_ (.B(net388),
    .A(net386),
    .X(_1844_));
 sg13g2_nor2_1 _5382_ (.A(net379),
    .B(_1844_),
    .Y(_1845_));
 sg13g2_a21o_1 _5383_ (.A2(net386),
    .A1(net379),
    .B1(_1845_),
    .X(_1846_));
 sg13g2_xor2_1 _5384_ (.B(_1846_),
    .A(_1752_),
    .X(_1847_));
 sg13g2_xor2_1 _5385_ (.B(_1847_),
    .A(_1760_),
    .X(_1848_));
 sg13g2_xnor2_1 _5386_ (.Y(_1849_),
    .A(_1842_),
    .B(_1848_));
 sg13g2_nor2_1 _5387_ (.A(_1841_),
    .B(_1849_),
    .Y(_1850_));
 sg13g2_xor2_1 _5388_ (.B(_1849_),
    .A(_1841_),
    .X(_1851_));
 sg13g2_nand2_1 _5389_ (.Y(_1852_),
    .A(_1840_),
    .B(_1851_));
 sg13g2_xnor2_1 _5390_ (.Y(_1853_),
    .A(_1840_),
    .B(_1851_));
 sg13g2_xor2_1 _5391_ (.B(_1853_),
    .A(net340),
    .X(_1854_));
 sg13g2_and2_1 _5392_ (.A(_1839_),
    .B(_1854_),
    .X(_1855_));
 sg13g2_xor2_1 _5393_ (.B(_1854_),
    .A(_1839_),
    .X(_1856_));
 sg13g2_xnor2_1 _5394_ (.Y(_1857_),
    .A(_1838_),
    .B(_1856_));
 sg13g2_and2_1 _5395_ (.A(_1837_),
    .B(_1857_),
    .X(_1858_));
 sg13g2_xor2_1 _5396_ (.B(_1857_),
    .A(_1837_),
    .X(_1859_));
 sg13g2_xnor2_1 _5397_ (.Y(_1860_),
    .A(net346),
    .B(_1859_));
 sg13g2_nand2_1 _5398_ (.Y(_1861_),
    .A(_1816_),
    .B(_1860_));
 sg13g2_xnor2_1 _5399_ (.Y(_1862_),
    .A(_1816_),
    .B(_1860_));
 sg13g2_xnor2_1 _5400_ (.Y(_1863_),
    .A(net326),
    .B(_1862_));
 sg13g2_and2_1 _5401_ (.A(_1815_),
    .B(_1863_),
    .X(_1864_));
 sg13g2_or2_1 _5402_ (.X(_1865_),
    .B(_1863_),
    .A(_1815_));
 sg13g2_xnor2_1 _5403_ (.Y(_1866_),
    .A(_1815_),
    .B(_1863_));
 sg13g2_o21ai_1 _5404_ (.B1(_1803_),
    .Y(_1867_),
    .A1(_1804_),
    .A2(_1808_));
 sg13g2_xnor2_1 _5405_ (.Y(_1868_),
    .A(_1866_),
    .B(_1867_));
 sg13g2_nand2_1 _5406_ (.Y(_1869_),
    .A(_1655_),
    .B(_1809_));
 sg13g2_nand2b_1 _5407_ (.Y(_1870_),
    .B(_1669_),
    .A_N(_1740_));
 sg13g2_a22oi_1 _5408_ (.Y(_1871_),
    .B1(_1868_),
    .B2(_0478_),
    .A2(_1659_),
    .A1(_1652_));
 sg13g2_and4_1 _5409_ (.A(net333),
    .B(_1869_),
    .C(_1870_),
    .D(_1871_),
    .X(_1872_));
 sg13g2_o21ai_1 _5410_ (.B1(net411),
    .Y(_1873_),
    .A1(net333),
    .A2(_1670_));
 sg13g2_o21ai_1 _5411_ (.B1(_1814_),
    .Y(_0111_),
    .A1(_1872_),
    .A2(_1873_));
 sg13g2_a21o_2 _5412_ (.A2(_1859_),
    .A1(net344),
    .B1(_1858_),
    .X(_1874_));
 sg13g2_a21o_1 _5413_ (.A2(_1856_),
    .A1(_1838_),
    .B1(_1855_),
    .X(_1875_));
 sg13g2_o21ai_1 _5414_ (.B1(_1852_),
    .Y(_1876_),
    .A1(net340),
    .A2(_1853_));
 sg13g2_a21oi_1 _5415_ (.A1(_1842_),
    .A2(_1848_),
    .Y(_1877_),
    .B1(_1850_));
 sg13g2_nand2_1 _5416_ (.Y(_1878_),
    .A(net386),
    .B(_1751_));
 sg13g2_or2_1 _5417_ (.X(_1879_),
    .B(_1878_),
    .A(_1750_));
 sg13g2_o21ai_1 _5418_ (.B1(_1879_),
    .Y(_1880_),
    .A1(_1760_),
    .A2(_1847_));
 sg13g2_nand3_1 _5419_ (.B(net386),
    .C(net388),
    .A(net379),
    .Y(_1881_));
 sg13g2_o21ai_1 _5420_ (.B1(_1881_),
    .Y(_1882_),
    .A1(_1750_),
    .A2(_1846_));
 sg13g2_nand2_2 _5421_ (.Y(_1883_),
    .A(_0607_),
    .B(_0638_));
 sg13g2_inv_1 _5422_ (.Y(_1884_),
    .A(_1883_));
 sg13g2_xnor2_1 _5423_ (.Y(_1885_),
    .A(net391),
    .B(_0639_));
 sg13g2_nor2_1 _5424_ (.A(_1843_),
    .B(_1885_),
    .Y(_1886_));
 sg13g2_xor2_1 _5425_ (.B(_1885_),
    .A(_1843_),
    .X(_1887_));
 sg13g2_xnor2_1 _5426_ (.Y(_1888_),
    .A(_1884_),
    .B(_1887_));
 sg13g2_inv_1 _5427_ (.Y(_1889_),
    .A(_1888_));
 sg13g2_xnor2_1 _5428_ (.Y(_1890_),
    .A(net385),
    .B(_1845_));
 sg13g2_xor2_1 _5429_ (.B(_1890_),
    .A(_1888_),
    .X(_1891_));
 sg13g2_nand2b_1 _5430_ (.Y(_1892_),
    .B(_1882_),
    .A_N(_1891_));
 sg13g2_xnor2_1 _5431_ (.Y(_1893_),
    .A(_1882_),
    .B(_1891_));
 sg13g2_inv_1 _5432_ (.Y(_1894_),
    .A(_1893_));
 sg13g2_xnor2_1 _5433_ (.Y(_1895_),
    .A(_1760_),
    .B(_1893_));
 sg13g2_nand2_1 _5434_ (.Y(_1896_),
    .A(_1880_),
    .B(_1895_));
 sg13g2_xnor2_1 _5435_ (.Y(_1897_),
    .A(_1880_),
    .B(_1895_));
 sg13g2_xor2_1 _5436_ (.B(_1897_),
    .A(_1841_),
    .X(_1898_));
 sg13g2_nand2b_1 _5437_ (.Y(_1899_),
    .B(_1898_),
    .A_N(_1877_));
 sg13g2_xnor2_1 _5438_ (.Y(_1900_),
    .A(_1877_),
    .B(_1898_));
 sg13g2_nand2b_1 _5439_ (.Y(_1901_),
    .B(_1900_),
    .A_N(net340));
 sg13g2_xnor2_1 _5440_ (.Y(_1902_),
    .A(net340),
    .B(_1900_));
 sg13g2_and2_1 _5441_ (.A(_1876_),
    .B(_1902_),
    .X(_1903_));
 sg13g2_xnor2_1 _5442_ (.Y(_1904_),
    .A(_1876_),
    .B(_1902_));
 sg13g2_inv_1 _5443_ (.Y(_1905_),
    .A(_1904_));
 sg13g2_xnor2_1 _5444_ (.Y(_1906_),
    .A(_1875_),
    .B(_1905_));
 sg13g2_inv_1 _5445_ (.Y(_1907_),
    .A(_1906_));
 sg13g2_a21oi_1 _5446_ (.A1(_1819_),
    .A2(_1836_),
    .Y(_1908_),
    .B1(_1835_));
 sg13g2_a21oi_1 _5447_ (.A1(_1352_),
    .A2(_1833_),
    .Y(_1909_),
    .B1(_1832_));
 sg13g2_a21oi_1 _5448_ (.A1(_1354_),
    .A2(_1830_),
    .Y(_1910_),
    .B1(_1829_));
 sg13g2_a21oi_1 _5449_ (.A1(net348),
    .A2(_1827_),
    .Y(_1911_),
    .B1(_1826_));
 sg13g2_o21ai_1 _5450_ (.B1(_0747_),
    .Y(_1912_),
    .A1(net357),
    .A2(_2154_));
 sg13g2_nand3_1 _5451_ (.B(net354),
    .C(_2154_),
    .A(net357),
    .Y(_1913_));
 sg13g2_nand3b_1 _5452_ (.B(_0852_),
    .C(_1913_),
    .Y(_1914_),
    .A_N(net349));
 sg13g2_nand2_1 _5453_ (.Y(_1915_),
    .A(_1912_),
    .B(_1914_));
 sg13g2_nor2_1 _5454_ (.A(_1911_),
    .B(_1915_),
    .Y(_1916_));
 sg13g2_xor2_1 _5455_ (.B(_1915_),
    .A(_1911_),
    .X(_1917_));
 sg13g2_xnor2_1 _5456_ (.Y(_1918_),
    .A(_1354_),
    .B(_1917_));
 sg13g2_nor2_1 _5457_ (.A(_1910_),
    .B(_1918_),
    .Y(_1919_));
 sg13g2_xor2_1 _5458_ (.B(_1918_),
    .A(_1910_),
    .X(_1920_));
 sg13g2_xnor2_1 _5459_ (.Y(_1921_),
    .A(_1353_),
    .B(_1920_));
 sg13g2_nand2b_1 _5460_ (.Y(_1922_),
    .B(_1921_),
    .A_N(_1909_));
 sg13g2_xnor2_1 _5461_ (.Y(_1923_),
    .A(_1909_),
    .B(_1921_));
 sg13g2_inv_1 _5462_ (.Y(_1924_),
    .A(_1923_));
 sg13g2_xnor2_1 _5463_ (.Y(_1925_),
    .A(_1908_),
    .B(_1923_));
 sg13g2_xnor2_1 _5464_ (.Y(_1926_),
    .A(_1906_),
    .B(_1925_));
 sg13g2_nand2_1 _5465_ (.Y(_1927_),
    .A(net344),
    .B(_1926_));
 sg13g2_xnor2_1 _5466_ (.Y(_1928_),
    .A(net346),
    .B(_1926_));
 sg13g2_nand2_1 _5467_ (.Y(_1929_),
    .A(_1874_),
    .B(_1928_));
 sg13g2_xnor2_1 _5468_ (.Y(_1930_),
    .A(_1874_),
    .B(_1928_));
 sg13g2_xnor2_1 _5469_ (.Y(_1931_),
    .A(net326),
    .B(_1930_));
 sg13g2_o21ai_1 _5470_ (.B1(_1861_),
    .Y(_1932_),
    .A1(net328),
    .A2(_1862_));
 sg13g2_nand2_1 _5471_ (.Y(_1933_),
    .A(_1931_),
    .B(_1932_));
 sg13g2_inv_1 _5472_ (.Y(_1934_),
    .A(_1933_));
 sg13g2_xor2_1 _5473_ (.B(_1932_),
    .A(_1931_),
    .X(_1935_));
 sg13g2_or2_1 _5474_ (.X(_1936_),
    .B(_1866_),
    .A(_1804_));
 sg13g2_a21oi_1 _5475_ (.A1(_1802_),
    .A2(_1865_),
    .Y(_1937_),
    .B1(_1864_));
 sg13g2_o21ai_1 _5476_ (.B1(_1937_),
    .Y(_1938_),
    .A1(_1808_),
    .A2(_1936_));
 sg13g2_xor2_1 _5477_ (.B(_1938_),
    .A(_1935_),
    .X(_1939_));
 sg13g2_nand2b_1 _5478_ (.Y(_1940_),
    .B(_1659_),
    .A_N(_1740_));
 sg13g2_nand2_1 _5479_ (.Y(_1941_),
    .A(_1669_),
    .B(_1809_));
 sg13g2_a21oi_1 _5480_ (.A1(_0478_),
    .A2(_1939_),
    .Y(_1942_),
    .B1(_1665_));
 sg13g2_a22oi_1 _5481_ (.Y(_1943_),
    .B1(_1868_),
    .B2(_1655_),
    .A2(_1663_),
    .A1(_1652_));
 sg13g2_nand4_1 _5482_ (.B(_1941_),
    .C(_1942_),
    .A(_1940_),
    .Y(_1944_),
    .D(_1943_));
 sg13g2_o21ai_1 _5483_ (.B1(net411),
    .Y(_1945_),
    .A1(_1657_),
    .A2(net333));
 sg13g2_nor2b_1 _5484_ (.A(_1945_),
    .B_N(_1944_),
    .Y(_0112_));
 sg13g2_a21oi_1 _5485_ (.A1(_1935_),
    .A2(_1938_),
    .Y(_1946_),
    .B1(_1934_));
 sg13g2_o21ai_1 _5486_ (.B1(_1929_),
    .Y(_1947_),
    .A1(net328),
    .A2(_1930_));
 sg13g2_o21ai_1 _5487_ (.B1(_1927_),
    .Y(_1948_),
    .A1(_1907_),
    .A2(_1925_));
 sg13g2_o21ai_1 _5488_ (.B1(_1922_),
    .Y(_1949_),
    .A1(_1908_),
    .A2(_1924_));
 sg13g2_a21oi_1 _5489_ (.A1(_1352_),
    .A2(_1920_),
    .Y(_1950_),
    .B1(_1919_));
 sg13g2_a21o_1 _5490_ (.A2(_0747_),
    .A1(net352),
    .B1(_0814_),
    .X(_1951_));
 sg13g2_inv_1 _5491_ (.Y(_1952_),
    .A(_1951_));
 sg13g2_nand2_1 _5492_ (.Y(_1953_),
    .A(_2159_),
    .B(_1824_));
 sg13g2_nand2_1 _5493_ (.Y(_1954_),
    .A(_1912_),
    .B(_1953_));
 sg13g2_xnor2_1 _5494_ (.Y(_1955_),
    .A(_1952_),
    .B(_1954_));
 sg13g2_a21oi_1 _5495_ (.A1(_1354_),
    .A2(_1917_),
    .Y(_1956_),
    .B1(_1916_));
 sg13g2_nor2_1 _5496_ (.A(_1955_),
    .B(_1956_),
    .Y(_1957_));
 sg13g2_xnor2_1 _5497_ (.Y(_1958_),
    .A(_1955_),
    .B(_1956_));
 sg13g2_nor2_1 _5498_ (.A(_1353_),
    .B(_1958_),
    .Y(_1959_));
 sg13g2_xnor2_1 _5499_ (.Y(_1960_),
    .A(_1353_),
    .B(_1958_));
 sg13g2_xor2_1 _5500_ (.B(_1960_),
    .A(_1950_),
    .X(_1961_));
 sg13g2_xor2_1 _5501_ (.B(_1961_),
    .A(_1949_),
    .X(_1962_));
 sg13g2_o21ai_1 _5502_ (.B1(_1896_),
    .Y(_1963_),
    .A1(_1841_),
    .A2(_1897_));
 sg13g2_o21ai_1 _5503_ (.B1(_1892_),
    .Y(_1964_),
    .A1(_1760_),
    .A2(_1894_));
 sg13g2_and2_1 _5504_ (.A(net379),
    .B(_1844_),
    .X(_1965_));
 sg13g2_a22oi_1 _5505_ (.Y(_1966_),
    .B1(_1965_),
    .B2(net385),
    .A2(_1890_),
    .A1(_1889_));
 sg13g2_and2_1 _5506_ (.A(net385),
    .B(net386),
    .X(_1967_));
 sg13g2_xor2_1 _5507_ (.B(net386),
    .A(net385),
    .X(_1968_));
 sg13g2_a21oi_1 _5508_ (.A1(net388),
    .A2(_1968_),
    .Y(_1969_),
    .B1(_1967_));
 sg13g2_or2_1 _5509_ (.X(_1970_),
    .B(_1969_),
    .A(_1885_));
 sg13g2_xnor2_1 _5510_ (.Y(_1971_),
    .A(_1885_),
    .B(_1969_));
 sg13g2_or2_1 _5511_ (.X(_1972_),
    .B(_1971_),
    .A(_1883_));
 sg13g2_xnor2_1 _5512_ (.Y(_1973_),
    .A(_1883_),
    .B(_1971_));
 sg13g2_xor2_1 _5513_ (.B(_1968_),
    .A(net388),
    .X(_1974_));
 sg13g2_mux2_1 _5514_ (.A0(_0491_),
    .A1(net383),
    .S(_1974_),
    .X(_1975_));
 sg13g2_xor2_1 _5515_ (.B(_1975_),
    .A(_1973_),
    .X(_1976_));
 sg13g2_nor2b_1 _5516_ (.A(_1966_),
    .B_N(_1976_),
    .Y(_1977_));
 sg13g2_xnor2_1 _5517_ (.Y(_1978_),
    .A(_1966_),
    .B(_1976_));
 sg13g2_a21oi_1 _5518_ (.A1(_1884_),
    .A2(_1887_),
    .Y(_1979_),
    .B1(_1886_));
 sg13g2_nor2_1 _5519_ (.A(_1755_),
    .B(_1979_),
    .Y(_1980_));
 sg13g2_xor2_1 _5520_ (.B(_1979_),
    .A(_1755_),
    .X(_1981_));
 sg13g2_xnor2_1 _5521_ (.Y(_1982_),
    .A(_1759_),
    .B(_1981_));
 sg13g2_inv_1 _5522_ (.Y(_1983_),
    .A(_1982_));
 sg13g2_xnor2_1 _5523_ (.Y(_1984_),
    .A(_1978_),
    .B(_1983_));
 sg13g2_nand2b_1 _5524_ (.Y(_1985_),
    .B(_1964_),
    .A_N(_1984_));
 sg13g2_xnor2_1 _5525_ (.Y(_1986_),
    .A(_1964_),
    .B(_1984_));
 sg13g2_inv_1 _5526_ (.Y(_1987_),
    .A(_1986_));
 sg13g2_xnor2_1 _5527_ (.Y(_1988_),
    .A(_1841_),
    .B(_1986_));
 sg13g2_nand2_1 _5528_ (.Y(_1989_),
    .A(_1963_),
    .B(_1988_));
 sg13g2_xnor2_1 _5529_ (.Y(_1990_),
    .A(_1963_),
    .B(_1988_));
 sg13g2_xor2_1 _5530_ (.B(_1990_),
    .A(net340),
    .X(_1991_));
 sg13g2_nand2_1 _5531_ (.Y(_1992_),
    .A(_1899_),
    .B(_1901_));
 sg13g2_nor2_1 _5532_ (.A(_1991_),
    .B(_1992_),
    .Y(_1993_));
 sg13g2_xor2_1 _5533_ (.B(_1992_),
    .A(_1991_),
    .X(_1994_));
 sg13g2_a21oi_1 _5534_ (.A1(_1875_),
    .A2(_1905_),
    .Y(_1995_),
    .B1(_1903_));
 sg13g2_xnor2_1 _5535_ (.Y(_1996_),
    .A(_1994_),
    .B(_1995_));
 sg13g2_or2_1 _5536_ (.X(_1997_),
    .B(_1996_),
    .A(_1962_));
 sg13g2_xnor2_1 _5537_ (.Y(_1998_),
    .A(_1962_),
    .B(_1996_));
 sg13g2_xnor2_1 _5538_ (.Y(_1999_),
    .A(net344),
    .B(_1998_));
 sg13g2_nand2_2 _5539_ (.Y(_2000_),
    .A(_1948_),
    .B(_1999_));
 sg13g2_xnor2_1 _5540_ (.Y(_2001_),
    .A(_1948_),
    .B(_1999_));
 sg13g2_xnor2_1 _5541_ (.Y(_2002_),
    .A(net326),
    .B(_2001_));
 sg13g2_nor2_1 _5542_ (.A(_1947_),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_xnor2_1 _5543_ (.Y(_2004_),
    .A(_1947_),
    .B(_2002_));
 sg13g2_xor2_1 _5544_ (.B(_2004_),
    .A(_1946_),
    .X(_2005_));
 sg13g2_a21oi_1 _5545_ (.A1(_1659_),
    .A2(_1809_),
    .Y(_2006_),
    .B1(_1665_));
 sg13g2_o21ai_1 _5546_ (.B1(_2006_),
    .Y(_2007_),
    .A1(_1664_),
    .A2(_1740_));
 sg13g2_a22oi_1 _5547_ (.Y(_2008_),
    .B1(_1939_),
    .B2(_1655_),
    .A2(_1868_),
    .A1(_1669_));
 sg13g2_a21oi_1 _5548_ (.A1(_0478_),
    .A2(_2005_),
    .Y(_2009_),
    .B1(_2007_));
 sg13g2_o21ai_1 _5549_ (.B1(net411),
    .Y(_2010_),
    .A1(_1652_),
    .A2(net333));
 sg13g2_a21oi_1 _5550_ (.A1(_2008_),
    .A2(_2009_),
    .Y(_0113_),
    .B1(_2010_));
 sg13g2_o21ai_1 _5551_ (.B1(_2000_),
    .Y(_2011_),
    .A1(net328),
    .A2(_2001_));
 sg13g2_a21oi_1 _5552_ (.A1(net352),
    .A2(_1352_),
    .Y(_2012_),
    .B1(_0747_));
 sg13g2_a21oi_1 _5553_ (.A1(_1952_),
    .A2(_1954_),
    .Y(_2013_),
    .B1(net349));
 sg13g2_nor2b_1 _5554_ (.A(_2013_),
    .B_N(_2012_),
    .Y(_2014_));
 sg13g2_o21ai_1 _5555_ (.B1(_2014_),
    .Y(_2015_),
    .A1(_1957_),
    .A2(_1959_));
 sg13g2_or3_1 _5556_ (.A(_1957_),
    .B(_1959_),
    .C(_2014_),
    .X(_2016_));
 sg13g2_nand2_1 _5557_ (.Y(_2017_),
    .A(_2015_),
    .B(_2016_));
 sg13g2_o21ai_1 _5558_ (.B1(_2017_),
    .Y(_2018_),
    .A1(_1950_),
    .A2(_1960_));
 sg13g2_a21o_1 _5559_ (.A2(_1961_),
    .A1(_1949_),
    .B1(_2018_),
    .X(_2019_));
 sg13g2_o21ai_1 _5560_ (.B1(_1989_),
    .Y(_2020_),
    .A1(net340),
    .A2(_1990_));
 sg13g2_o21ai_1 _5561_ (.B1(_1985_),
    .Y(_2021_),
    .A1(_1841_),
    .A2(_1987_));
 sg13g2_a21oi_1 _5562_ (.A1(_1759_),
    .A2(_1981_),
    .Y(_2022_),
    .B1(_1980_));
 sg13g2_a21oi_1 _5563_ (.A1(_1978_),
    .A2(_1983_),
    .Y(_2023_),
    .B1(_1977_));
 sg13g2_nand3_1 _5564_ (.B(net383),
    .C(_1974_),
    .A(net380),
    .Y(_2024_));
 sg13g2_o21ai_1 _5565_ (.B1(_2024_),
    .Y(_2025_),
    .A1(_1973_),
    .A2(_1975_));
 sg13g2_nand2_1 _5566_ (.Y(_2026_),
    .A(net382),
    .B(_1974_));
 sg13g2_or2_1 _5567_ (.X(_2027_),
    .B(_2026_),
    .A(_0491_));
 sg13g2_xnor2_1 _5568_ (.Y(_2028_),
    .A(net382),
    .B(_1974_));
 sg13g2_o21ai_1 _5569_ (.B1(_0485_),
    .Y(_2029_),
    .A1(net384),
    .A2(_0484_));
 sg13g2_nor2_1 _5570_ (.A(_2028_),
    .B(_2029_),
    .Y(_2030_));
 sg13g2_a21oi_1 _5571_ (.A1(_0490_),
    .A2(_2028_),
    .Y(_2031_),
    .B1(_2030_));
 sg13g2_nand2_1 _5572_ (.Y(_2032_),
    .A(_2027_),
    .B(_2031_));
 sg13g2_xor2_1 _5573_ (.B(_2032_),
    .A(_1973_),
    .X(_2033_));
 sg13g2_nand2_1 _5574_ (.Y(_2034_),
    .A(_2025_),
    .B(_2033_));
 sg13g2_xnor2_1 _5575_ (.Y(_2035_),
    .A(_2025_),
    .B(_2033_));
 sg13g2_nand3_1 _5576_ (.B(_1970_),
    .C(_1972_),
    .A(_1755_),
    .Y(_2036_));
 sg13g2_a21o_1 _5577_ (.A2(_1972_),
    .A1(_1970_),
    .B1(_1755_),
    .X(_2037_));
 sg13g2_and2_1 _5578_ (.A(_2036_),
    .B(_2037_),
    .X(_2038_));
 sg13g2_xnor2_1 _5579_ (.Y(_2039_),
    .A(_1759_),
    .B(_2038_));
 sg13g2_xnor2_1 _5580_ (.Y(_2040_),
    .A(_2035_),
    .B(_2039_));
 sg13g2_xor2_1 _5581_ (.B(_2040_),
    .A(_2023_),
    .X(_2041_));
 sg13g2_nand2b_1 _5582_ (.Y(_2042_),
    .B(_2041_),
    .A_N(_2022_));
 sg13g2_xnor2_1 _5583_ (.Y(_2043_),
    .A(_2022_),
    .B(_2041_));
 sg13g2_nand2_1 _5584_ (.Y(_2044_),
    .A(_2021_),
    .B(_2043_));
 sg13g2_xnor2_1 _5585_ (.Y(_2045_),
    .A(_2021_),
    .B(_2043_));
 sg13g2_xor2_1 _5586_ (.B(_2045_),
    .A(net340),
    .X(_2046_));
 sg13g2_nand2_1 _5587_ (.Y(_2047_),
    .A(_2020_),
    .B(_2046_));
 sg13g2_xnor2_1 _5588_ (.Y(_2048_),
    .A(_2020_),
    .B(_2046_));
 sg13g2_a221oi_1 _5589_ (.B2(_1992_),
    .C1(_1903_),
    .B1(_1991_),
    .A1(_1875_),
    .Y(_2049_),
    .A2(_1905_));
 sg13g2_or3_1 _5590_ (.A(_1993_),
    .B(_2048_),
    .C(_2049_),
    .X(_2050_));
 sg13g2_o21ai_1 _5591_ (.B1(_2048_),
    .Y(_2051_),
    .A1(_1993_),
    .A2(_2049_));
 sg13g2_a21oi_1 _5592_ (.A1(_2050_),
    .A2(_2051_),
    .Y(_2052_),
    .B1(_2019_));
 sg13g2_nand3_1 _5593_ (.B(_2050_),
    .C(_2051_),
    .A(_2019_),
    .Y(_2053_));
 sg13g2_nor2b_1 _5594_ (.A(_2052_),
    .B_N(_2053_),
    .Y(_2054_));
 sg13g2_nand2_1 _5595_ (.Y(_2055_),
    .A(net346),
    .B(_2052_));
 sg13g2_xnor2_1 _5596_ (.Y(_2056_),
    .A(net346),
    .B(_2054_));
 sg13g2_o21ai_1 _5597_ (.B1(_1997_),
    .Y(_2057_),
    .A1(net346),
    .A2(_1998_));
 sg13g2_and2_1 _5598_ (.A(_2056_),
    .B(_2057_),
    .X(_2058_));
 sg13g2_xor2_1 _5599_ (.B(_2057_),
    .A(_2056_),
    .X(_2059_));
 sg13g2_xnor2_1 _5600_ (.Y(_2060_),
    .A(net328),
    .B(_2059_));
 sg13g2_and2_1 _5601_ (.A(_2011_),
    .B(_2060_),
    .X(_2061_));
 sg13g2_xnor2_1 _5602_ (.Y(_2062_),
    .A(_2011_),
    .B(_2060_));
 sg13g2_a221oi_1 _5603_ (.B2(_2002_),
    .C1(_1934_),
    .B1(_1947_),
    .A1(_1935_),
    .Y(_2063_),
    .A2(_1938_));
 sg13g2_nor2_1 _5604_ (.A(_2003_),
    .B(_2063_),
    .Y(_2064_));
 sg13g2_nor3_1 _5605_ (.A(_2003_),
    .B(_2062_),
    .C(_2063_),
    .Y(_2065_));
 sg13g2_xnor2_1 _5606_ (.Y(_2066_),
    .A(_2062_),
    .B(_2064_));
 sg13g2_nand2_1 _5607_ (.Y(_2067_),
    .A(_1669_),
    .B(_1939_));
 sg13g2_a221oi_1 _5608_ (.B2(_1659_),
    .C1(_1665_),
    .B1(_1868_),
    .A1(_1663_),
    .Y(_2068_),
    .A2(_1809_));
 sg13g2_nand2_1 _5609_ (.Y(_2069_),
    .A(_2067_),
    .B(_2068_));
 sg13g2_a221oi_1 _5610_ (.B2(_0478_),
    .C1(_2069_),
    .B1(_2066_),
    .A1(_1655_),
    .Y(_2070_),
    .A2(_2005_));
 sg13g2_a21oi_1 _5611_ (.A1(_1665_),
    .A2(_1740_),
    .Y(_2071_),
    .B1(net406));
 sg13g2_nor2b_1 _5612_ (.A(_2070_),
    .B_N(_2071_),
    .Y(_0114_));
 sg13g2_a21oi_1 _5613_ (.A1(net326),
    .A2(_2059_),
    .Y(_2072_),
    .B1(_2058_));
 sg13g2_o21ai_1 _5614_ (.B1(_2055_),
    .Y(_2073_),
    .A1(net346),
    .A2(_2053_));
 sg13g2_nand2_1 _5615_ (.Y(_2074_),
    .A(_2047_),
    .B(_2050_));
 sg13g2_o21ai_1 _5616_ (.B1(_2034_),
    .Y(_2075_),
    .A1(_2035_),
    .A2(_2039_));
 sg13g2_nand2b_1 _5617_ (.Y(_2076_),
    .B(_1759_),
    .A_N(_2037_));
 sg13g2_o21ai_1 _5618_ (.B1(_2076_),
    .Y(_2077_),
    .A1(_1759_),
    .A2(_2036_));
 sg13g2_mux2_1 _5619_ (.A0(_2031_),
    .A1(_2027_),
    .S(_1973_),
    .X(_2078_));
 sg13g2_nor3_1 _5620_ (.A(net382),
    .B(net383),
    .C(_1974_),
    .Y(_2079_));
 sg13g2_nand2b_1 _5621_ (.Y(_2080_),
    .B(net383),
    .A_N(net380));
 sg13g2_a21oi_1 _5622_ (.A1(net381),
    .A2(_2026_),
    .Y(_2081_),
    .B1(_2079_));
 sg13g2_o21ai_1 _5623_ (.B1(_2081_),
    .Y(_2082_),
    .A1(_2026_),
    .A2(_2080_));
 sg13g2_xnor2_1 _5624_ (.Y(_2083_),
    .A(net341),
    .B(_2012_));
 sg13g2_xnor2_1 _5625_ (.Y(_2084_),
    .A(_2082_),
    .B(_2083_));
 sg13g2_xnor2_1 _5626_ (.Y(_2085_),
    .A(_2078_),
    .B(_2084_));
 sg13g2_xnor2_1 _5627_ (.Y(_2086_),
    .A(_2077_),
    .B(_2085_));
 sg13g2_xnor2_1 _5628_ (.Y(_2087_),
    .A(_2075_),
    .B(_2086_));
 sg13g2_o21ai_1 _5629_ (.B1(_2042_),
    .Y(_2088_),
    .A1(_2023_),
    .A2(_2040_));
 sg13g2_xnor2_1 _5630_ (.Y(_2089_),
    .A(_2087_),
    .B(_2088_));
 sg13g2_xnor2_1 _5631_ (.Y(_2090_),
    .A(_2015_),
    .B(_2089_));
 sg13g2_o21ai_1 _5632_ (.B1(_2044_),
    .Y(_2091_),
    .A1(net340),
    .A2(_2045_));
 sg13g2_xnor2_1 _5633_ (.Y(_2092_),
    .A(_2090_),
    .B(_2091_));
 sg13g2_xnor2_1 _5634_ (.Y(_2093_),
    .A(net328),
    .B(_2092_));
 sg13g2_xnor2_1 _5635_ (.Y(_2094_),
    .A(_2074_),
    .B(_2093_));
 sg13g2_xnor2_1 _5636_ (.Y(_2095_),
    .A(_2073_),
    .B(_2094_));
 sg13g2_xnor2_1 _5637_ (.Y(_2096_),
    .A(_2072_),
    .B(_2095_));
 sg13g2_or3_1 _5638_ (.A(_2061_),
    .B(_2065_),
    .C(_2096_),
    .X(_2097_));
 sg13g2_o21ai_1 _5639_ (.B1(_2096_),
    .Y(_2098_),
    .A1(_2061_),
    .A2(_2065_));
 sg13g2_nand3_1 _5640_ (.B(_2097_),
    .C(_2098_),
    .A(_0478_),
    .Y(_2099_));
 sg13g2_a22oi_1 _5641_ (.Y(_2100_),
    .B1(_1939_),
    .B2(_1659_),
    .A2(_1868_),
    .A1(_1663_));
 sg13g2_nand2_1 _5642_ (.Y(_2101_),
    .A(net333),
    .B(_2100_));
 sg13g2_a221oi_1 _5643_ (.B2(_1655_),
    .C1(_2101_),
    .B1(_2066_),
    .A1(_1669_),
    .Y(_2102_),
    .A2(_2005_));
 sg13g2_o21ai_1 _5644_ (.B1(net412),
    .Y(_2103_),
    .A1(net333),
    .A2(_1809_));
 sg13g2_a21oi_1 _5645_ (.A1(_2099_),
    .A2(_2102_),
    .Y(_0115_),
    .B1(_2103_));
 sg13g2_o21ai_1 _5646_ (.B1(net426),
    .Y(_2104_),
    .A1(_1517_),
    .A2(_1616_));
 sg13g2_a21oi_1 _5647_ (.A1(_1517_),
    .A2(_1616_),
    .Y(_0116_),
    .B1(_2104_));
 sg13g2_nand2_1 _5648_ (.Y(_2105_),
    .A(_1617_),
    .B(_1618_));
 sg13g2_and3_1 _5649_ (.X(_0117_),
    .A(net426),
    .B(_1619_),
    .C(_2105_));
 sg13g2_nor2_1 _5650_ (.A(net410),
    .B(_1674_),
    .Y(_0118_));
 sg13g2_and2_1 _5651_ (.A(net418),
    .B(_1667_),
    .X(_0119_));
 sg13g2_nor2_1 _5652_ (.A(net410),
    .B(_1661_),
    .Y(_0120_));
 sg13g2_and2_1 _5653_ (.A(net411),
    .B(_1670_),
    .X(_0121_));
 sg13g2_and2_1 _5654_ (.A(net411),
    .B(_1652_),
    .X(_0123_));
 sg13g2_nor2_1 _5655_ (.A(net406),
    .B(_1740_),
    .Y(_0124_));
 sg13g2_and2_1 _5656_ (.A(net412),
    .B(_1809_),
    .X(_0125_));
 sg13g2_and2_1 _5657_ (.A(net412),
    .B(_1868_),
    .X(_0126_));
 sg13g2_and2_1 _5658_ (.A(net411),
    .B(_1939_),
    .X(_0127_));
 sg13g2_and2_1 _5659_ (.A(net412),
    .B(_2005_),
    .X(_0128_));
 sg13g2_and2_1 _5660_ (.A(net412),
    .B(_2066_),
    .X(_0129_));
 sg13g2_and2_1 _5661_ (.A(net416),
    .B(net219),
    .X(_0130_));
 sg13g2_and2_1 _5662_ (.A(net416),
    .B(net321),
    .X(_0131_));
 sg13g2_nor2_1 _5663_ (.A(net406),
    .B(_2146_),
    .Y(_0132_));
 sg13g2_and2_1 _5664_ (.A(net415),
    .B(net396),
    .X(_0133_));
 sg13g2_nor2_1 _5665_ (.A(net406),
    .B(_2145_),
    .Y(_0134_));
 sg13g2_and2_1 _5666_ (.A(net415),
    .B(net393),
    .X(_0135_));
 sg13g2_and2_1 _5667_ (.A(net415),
    .B(net391),
    .X(_0136_));
 sg13g2_and2_1 _5668_ (.A(net415),
    .B(net390),
    .X(_0137_));
 sg13g2_and2_1 _5669_ (.A(net416),
    .B(net388),
    .X(_0138_));
 sg13g2_and2_1 _5670_ (.A(net416),
    .B(net386),
    .X(_0139_));
 sg13g2_and2_1 _5671_ (.A(net415),
    .B(net385),
    .X(_0140_));
 sg13g2_and2_1 _5672_ (.A(net415),
    .B(net383),
    .X(_0141_));
 sg13g2_and2_1 _5673_ (.A(net415),
    .B(net382),
    .X(_0142_));
 sg13g2_and2_1 _5674_ (.A(net415),
    .B(net379),
    .X(_0143_));
 sg13g2_and2_1 _5675_ (.A(net423),
    .B(net288),
    .X(_0144_));
 sg13g2_and2_1 _5676_ (.A(net424),
    .B(net311),
    .X(_0145_));
 sg13g2_and2_1 _5677_ (.A(net422),
    .B(net292),
    .X(_0146_));
 sg13g2_and2_1 _5678_ (.A(net423),
    .B(net289),
    .X(_0147_));
 sg13g2_and2_1 _5679_ (.A(net424),
    .B(net307),
    .X(_0148_));
 sg13g2_and2_1 _5680_ (.A(net424),
    .B(net297),
    .X(_0149_));
 sg13g2_and2_1 _5681_ (.A(net424),
    .B(net286),
    .X(_0150_));
 sg13g2_nor2_1 _5682_ (.A(net409),
    .B(_2155_),
    .Y(_0151_));
 sg13g2_and2_1 _5683_ (.A(net423),
    .B(net200),
    .X(_0152_));
 sg13g2_and2_1 _5684_ (.A(net424),
    .B(net197),
    .X(_0153_));
 sg13g2_and2_1 _5685_ (.A(net423),
    .B(net196),
    .X(_0154_));
 sg13g2_and2_1 _5686_ (.A(net423),
    .B(net193),
    .X(_0155_));
 sg13g2_and2_1 _5687_ (.A(net424),
    .B(net195),
    .X(_0156_));
 sg13g2_and2_1 _5688_ (.A(net424),
    .B(net189),
    .X(_0157_));
 sg13g2_and2_1 _5689_ (.A(net424),
    .B(net190),
    .X(_0158_));
 sg13g2_and2_1 _5690_ (.A(net425),
    .B(net199),
    .X(_0159_));
 sg13g2_o21ai_1 _5691_ (.B1(net420),
    .Y(_2106_),
    .A1(\am_sdr0.nco0.phase_inc[0] ),
    .A2(net228));
 sg13g2_nor2_1 _5692_ (.A(_2195_),
    .B(net229),
    .Y(_0160_));
 sg13g2_o21ai_1 _5693_ (.B1(net420),
    .Y(_2107_),
    .A1(_2195_),
    .A2(net428));
 sg13g2_nor2b_1 _5694_ (.A(_2107_),
    .B_N(_2197_),
    .Y(_0161_));
 sg13g2_nand3_1 _5695_ (.B(_2197_),
    .C(_2198_),
    .A(_2194_),
    .Y(_2108_));
 sg13g2_and3_1 _5696_ (.X(_0162_),
    .A(net420),
    .B(_2199_),
    .C(_2108_));
 sg13g2_nand3_1 _5697_ (.B(_2199_),
    .C(_2200_),
    .A(_2193_),
    .Y(_2109_));
 sg13g2_and3_1 _5698_ (.X(_0163_),
    .A(net421),
    .B(_2201_),
    .C(_2109_));
 sg13g2_nand3_1 _5699_ (.B(_2201_),
    .C(_2202_),
    .A(_2192_),
    .Y(_2110_));
 sg13g2_and3_1 _5700_ (.X(_0164_),
    .A(net420),
    .B(_2203_),
    .C(net324));
 sg13g2_nand3_1 _5701_ (.B(_2203_),
    .C(_2204_),
    .A(_2191_),
    .Y(_2111_));
 sg13g2_and3_1 _5702_ (.X(_0165_),
    .A(net420),
    .B(_2205_),
    .C(net319));
 sg13g2_nand3_1 _5703_ (.B(_2205_),
    .C(_2206_),
    .A(_2190_),
    .Y(_2112_));
 sg13g2_and3_1 _5704_ (.X(_0166_),
    .A(net419),
    .B(_2207_),
    .C(_2112_));
 sg13g2_nand3_1 _5705_ (.B(_2207_),
    .C(_2208_),
    .A(_2189_),
    .Y(_2113_));
 sg13g2_and3_1 _5706_ (.X(_0167_),
    .A(net419),
    .B(_2209_),
    .C(_2113_));
 sg13g2_and3_1 _5707_ (.X(_2114_),
    .A(_2188_),
    .B(_2209_),
    .C(_2210_));
 sg13g2_nor3_1 _5708_ (.A(net408),
    .B(_2211_),
    .C(net305),
    .Y(_0168_));
 sg13g2_xor2_1 _5709_ (.B(net300),
    .A(net276),
    .X(_2115_));
 sg13g2_o21ai_1 _5710_ (.B1(net420),
    .Y(_2116_),
    .A1(_2212_),
    .A2(_2115_));
 sg13g2_a21oi_1 _5711_ (.A1(_2212_),
    .A2(_2115_),
    .Y(_0169_),
    .B1(_2116_));
 sg13g2_nand3_1 _5712_ (.B(_2187_),
    .C(_2213_),
    .A(_2186_),
    .Y(_2117_));
 sg13g2_nand2_1 _5713_ (.Y(_2118_),
    .A(net418),
    .B(_2117_));
 sg13g2_nor2_1 _5714_ (.A(net315),
    .B(_2118_),
    .Y(_0170_));
 sg13g2_nand2b_1 _5715_ (.Y(_2119_),
    .B(_2185_),
    .A_N(_2184_));
 sg13g2_o21ai_1 _5716_ (.B1(net418),
    .Y(_2120_),
    .A1(_2215_),
    .A2(_2119_));
 sg13g2_a21oi_1 _5717_ (.A1(_2215_),
    .A2(_2119_),
    .Y(_0171_),
    .B1(_2120_));
 sg13g2_o21ai_1 _5718_ (.B1(net418),
    .Y(_2121_),
    .A1(_2183_),
    .A2(_2216_));
 sg13g2_a21oi_1 _5719_ (.A1(_2183_),
    .A2(_2216_),
    .Y(_0172_),
    .B1(_2121_));
 sg13g2_xor2_1 _5720_ (.B(net308),
    .A(net274),
    .X(_2122_));
 sg13g2_o21ai_1 _5721_ (.B1(net418),
    .Y(_2123_),
    .A1(_2217_),
    .A2(_2122_));
 sg13g2_a21oi_1 _5722_ (.A1(_2217_),
    .A2(_2122_),
    .Y(_0173_),
    .B1(_2123_));
 sg13g2_xnor2_1 _5723_ (.Y(_2124_),
    .A(net436),
    .B(_2219_));
 sg13g2_and2_1 _5724_ (.A(net418),
    .B(_2124_),
    .X(_0174_));
 sg13g2_xor2_1 _5725_ (.B(net298),
    .A(net257),
    .X(_2125_));
 sg13g2_o21ai_1 _5726_ (.B1(net420),
    .Y(_2126_),
    .A1(_2220_),
    .A2(_2125_));
 sg13g2_a21oi_1 _5727_ (.A1(_2220_),
    .A2(_2125_),
    .Y(_0175_),
    .B1(_2126_));
 sg13g2_and2_1 _5728_ (.A(net422),
    .B(net1),
    .X(_0180_));
 sg13g2_and2_1 _5729_ (.A(net422),
    .B(net2),
    .X(_0181_));
 sg13g2_and2_1 _5730_ (.A(net208),
    .B(net425),
    .X(_0182_));
 sg13g2_and2_1 _5731_ (.A(net422),
    .B(net198),
    .X(_0183_));
 sg13g2_dfrbp_1 _5732_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net58),
    .D(net211),
    .Q_N(_2857_),
    .Q(\am_sdr0.nco0.phase_inc[0] ));
 sg13g2_dfrbp_1 _5733_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net44),
    .D(net244),
    .Q_N(_2856_),
    .Q(\am_sdr0.nco0.phase_inc[1] ));
 sg13g2_dfrbp_1 _5734_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net42),
    .D(net279),
    .Q_N(_2855_),
    .Q(\am_sdr0.nco0.phase_inc[2] ));
 sg13g2_dfrbp_1 _5735_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net40),
    .D(_0043_),
    .Q_N(_2854_),
    .Q(\am_sdr0.nco0.phase_inc[3] ));
 sg13g2_dfrbp_1 _5736_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net38),
    .D(_0044_),
    .Q_N(_2853_),
    .Q(\am_sdr0.nco0.phase_inc[4] ));
 sg13g2_dfrbp_1 _5737_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net36),
    .D(_0045_),
    .Q_N(_2852_),
    .Q(\am_sdr0.nco0.phase_inc[5] ));
 sg13g2_dfrbp_1 _5738_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net34),
    .D(net233),
    .Q_N(_2851_),
    .Q(\am_sdr0.nco0.phase_inc[6] ));
 sg13g2_dfrbp_1 _5739_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net32),
    .D(net237),
    .Q_N(_2850_),
    .Q(\am_sdr0.nco0.phase_inc[7] ));
 sg13g2_dfrbp_1 _5740_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net30),
    .D(_0048_),
    .Q_N(_2849_),
    .Q(\am_sdr0.nco0.phase_inc[8] ));
 sg13g2_dfrbp_1 _5741_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net28),
    .D(net250),
    .Q_N(_2848_),
    .Q(\am_sdr0.nco0.phase_inc[9] ));
 sg13g2_dfrbp_1 _5742_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net186),
    .D(_0050_),
    .Q_N(_2847_),
    .Q(\am_sdr0.nco0.phase_inc[10] ));
 sg13g2_dfrbp_1 _5743_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net184),
    .D(_0051_),
    .Q_N(_2846_),
    .Q(\am_sdr0.nco0.phase_inc[11] ));
 sg13g2_dfrbp_1 _5744_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net182),
    .D(_0052_),
    .Q_N(_2845_),
    .Q(\am_sdr0.nco0.phase_inc[12] ));
 sg13g2_dfrbp_1 _5745_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net180),
    .D(net242),
    .Q_N(_2844_),
    .Q(\am_sdr0.nco0.phase_inc[13] ));
 sg13g2_dfrbp_1 _5746_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net178),
    .D(net275),
    .Q_N(_2843_),
    .Q(\am_sdr0.nco0.phase_inc[14] ));
 sg13g2_dfrbp_1 _5747_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net176),
    .D(_0055_),
    .Q_N(_2842_),
    .Q(\am_sdr0.nco0.phase_inc[15] ));
 sg13g2_dfrbp_1 _5748_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net174),
    .D(net258),
    .Q_N(_2841_),
    .Q(\am_sdr0.nco0.phase_inc[16] ));
 sg13g2_dfrbp_1 _5749_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net172),
    .D(net260),
    .Q_N(_2840_),
    .Q(\am_sdr0.nco0.phase_inc[17] ));
 sg13g2_dfrbp_1 _5750_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net170),
    .D(_0058_),
    .Q_N(_2839_),
    .Q(\am_sdr0.nco0.phase_inc[18] ));
 sg13g2_dfrbp_1 _5751_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net168),
    .D(_0059_),
    .Q_N(_2838_),
    .Q(\am_sdr0.nco0.phase_inc[19] ));
 sg13g2_dfrbp_1 _5752_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net166),
    .D(net252),
    .Q_N(_2837_),
    .Q(\am_sdr0.filt0.gain_spi[0] ));
 sg13g2_dfrbp_1 _5753_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net164),
    .D(net291),
    .Q_N(_2836_),
    .Q(\am_sdr0.filt0.gain_spi[1] ));
 sg13g2_dfrbp_1 _5754_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net162),
    .D(net247),
    .Q_N(_0017_),
    .Q(\am_sdr0.filt0.gain_spi[2] ));
 sg13g2_dfrbp_1 _5755_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net160),
    .D(_0063_),
    .Q_N(_2835_),
    .Q(\am_sdr0.spi0.state[0] ));
 sg13g2_dfrbp_1 _5756_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net158),
    .D(_0064_),
    .Q_N(_2834_),
    .Q(\am_sdr0.spi0.state[1] ));
 sg13g2_dfrbp_1 _5757_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net156),
    .D(_0065_),
    .Q_N(_2833_),
    .Q(COMP_OUT));
 sg13g2_dfrbp_1 _5758_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net155),
    .D(_0066_),
    .Q_N(_2832_),
    .Q(\am_sdr0.spi0.CS_q ));
 sg13g2_dfrbp_1 _5759_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net146),
    .D(_0067_),
    .Q_N(_2831_),
    .Q(\am_sdr0.spi0.CS_qq ));
 sg13g2_dfrbp_1 _5760_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net145),
    .D(_0068_),
    .Q_N(_2830_),
    .Q(\am_sdr0.spi0.CS_qqq ));
 sg13g2_dfrbp_1 _5761_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net144),
    .D(_0069_),
    .Q_N(_2829_),
    .Q(\am_sdr0.spi0.SCK_q ));
 sg13g2_dfrbp_1 _5762_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net59),
    .D(_0070_),
    .Q_N(_2858_),
    .Q(PWM_OUT));
 sg13g2_dfrbp_1 _5763_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net60),
    .D(_0000_),
    .Q_N(_2859_),
    .Q(_0031_));
 sg13g2_dfrbp_1 _5764_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net61),
    .D(_0001_),
    .Q_N(_2860_),
    .Q(_0032_));
 sg13g2_dfrbp_1 _5765_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net62),
    .D(_0002_),
    .Q_N(_0020_),
    .Q(_0033_));
 sg13g2_dfrbp_1 _5766_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net63),
    .D(_0003_),
    .Q_N(_2861_),
    .Q(_0034_));
 sg13g2_dfrbp_1 _5767_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net64),
    .D(_0004_),
    .Q_N(_0021_),
    .Q(_0035_));
 sg13g2_dfrbp_1 _5768_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net65),
    .D(_0005_),
    .Q_N(_2862_),
    .Q(_0036_));
 sg13g2_dfrbp_1 _5769_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net147),
    .D(_0006_),
    .Q_N(_0022_),
    .Q(_0037_));
 sg13g2_dfrbp_1 _5770_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net143),
    .D(_0007_),
    .Q_N(_2828_),
    .Q(_0038_));
 sg13g2_dfrbp_1 _5771_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net142),
    .D(_0071_),
    .Q_N(_2827_),
    .Q(\am_sdr0.spi0.MOSI_qq ));
 sg13g2_dfrbp_1 _5772_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net141),
    .D(_0072_),
    .Q_N(_0039_),
    .Q(\am_sdr0.count[0] ));
 sg13g2_dfrbp_1 _5773_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net140),
    .D(net225),
    .Q_N(_2826_),
    .Q(\am_sdr0.count[1] ));
 sg13g2_dfrbp_1 _5774_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net139),
    .D(_0074_),
    .Q_N(_2825_),
    .Q(\am_sdr0.count[2] ));
 sg13g2_dfrbp_1 _5775_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net138),
    .D(_0075_),
    .Q_N(_2824_),
    .Q(\am_sdr0.count[3] ));
 sg13g2_dfrbp_1 _5776_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net137),
    .D(net267),
    .Q_N(_2823_),
    .Q(\am_sdr0.count[4] ));
 sg13g2_dfrbp_1 _5777_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net136),
    .D(_0077_),
    .Q_N(_2822_),
    .Q(\am_sdr0.count[5] ));
 sg13g2_dfrbp_1 _5778_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net135),
    .D(net218),
    .Q_N(_2821_),
    .Q(\am_sdr0.count[6] ));
 sg13g2_dfrbp_1 _5779_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net134),
    .D(net254),
    .Q_N(_2820_),
    .Q(\am_sdr0.count[7] ));
 sg13g2_dfrbp_1 _5780_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net133),
    .D(_0080_),
    .Q_N(_2819_),
    .Q(\am_sdr0.det0.env_out[0] ));
 sg13g2_dfrbp_1 _5781_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net132),
    .D(_0081_),
    .Q_N(_2818_),
    .Q(\am_sdr0.det0.env_out[1] ));
 sg13g2_dfrbp_1 _5782_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net131),
    .D(_0082_),
    .Q_N(_2817_),
    .Q(\am_sdr0.det0.env_out[2] ));
 sg13g2_dfrbp_1 _5783_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net130),
    .D(_0083_),
    .Q_N(_2816_),
    .Q(\am_sdr0.det0.env_out[3] ));
 sg13g2_dfrbp_1 _5784_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net129),
    .D(_0084_),
    .Q_N(_2815_),
    .Q(\am_sdr0.det0.env_out[4] ));
 sg13g2_dfrbp_1 _5785_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net128),
    .D(_0085_),
    .Q_N(_2814_),
    .Q(\am_sdr0.det0.env_out[5] ));
 sg13g2_dfrbp_1 _5786_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net127),
    .D(_0086_),
    .Q_N(_2813_),
    .Q(\am_sdr0.det0.env_out[6] ));
 sg13g2_dfrbp_1 _5787_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net126),
    .D(_0087_),
    .Q_N(_2812_),
    .Q(\am_sdr0.det0.env_out[7] ));
 sg13g2_dfrbp_1 _5788_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net125),
    .D(_0088_),
    .Q_N(_2811_),
    .Q(\am_sdr0.det0.alpha_yn_1[0] ));
 sg13g2_dfrbp_1 _5789_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net124),
    .D(_0089_),
    .Q_N(_2810_),
    .Q(\am_sdr0.det0.yn_1[1] ));
 sg13g2_dfrbp_1 _5790_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net123),
    .D(_0090_),
    .Q_N(_2809_),
    .Q(\am_sdr0.det0.yn_1[2] ));
 sg13g2_dfrbp_1 _5791_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net122),
    .D(_0091_),
    .Q_N(_2808_),
    .Q(\am_sdr0.det0.yn_1[3] ));
 sg13g2_dfrbp_1 _5792_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net121),
    .D(_0092_),
    .Q_N(_2807_),
    .Q(\am_sdr0.det0.yn_1[4] ));
 sg13g2_dfrbp_1 _5793_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net120),
    .D(_0093_),
    .Q_N(_2806_),
    .Q(\am_sdr0.det0.yn_1[5] ));
 sg13g2_dfrbp_1 _5794_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net119),
    .D(_0094_),
    .Q_N(_2805_),
    .Q(\am_sdr0.det0.yn_1[6] ));
 sg13g2_dfrbp_1 _5795_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net118),
    .D(net431),
    .Q_N(_2804_),
    .Q(\am_sdr0.det0.yn_1[7] ));
 sg13g2_dfrbp_1 _5796_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net117),
    .D(_0096_),
    .Q_N(_2803_),
    .Q(\am_sdr0.det0.yn_1[8] ));
 sg13g2_dfrbp_1 _5797_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net116),
    .D(_0097_),
    .Q_N(_2802_),
    .Q(\am_sdr0.det0.yn_1[9] ));
 sg13g2_dfrbp_1 _5798_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net115),
    .D(_0098_),
    .Q_N(_2801_),
    .Q(\am_sdr0.det0.yn_1[10] ));
 sg13g2_dfrbp_1 _5799_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net114),
    .D(_0099_),
    .Q_N(_2800_),
    .Q(\am_sdr0.det0.yn_1[11] ));
 sg13g2_dfrbp_1 _5800_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net113),
    .D(_0100_),
    .Q_N(_2799_),
    .Q(\am_sdr0.det0.yn_1[12] ));
 sg13g2_dfrbp_1 _5801_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net112),
    .D(_0101_),
    .Q_N(_2798_),
    .Q(\am_sdr0.det0.yn_1[13] ));
 sg13g2_dfrbp_1 _5802_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net111),
    .D(_0102_),
    .Q_N(_2797_),
    .Q(\am_sdr0.det0.yn_1[14] ));
 sg13g2_dfrbp_1 _5803_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net110),
    .D(_0103_),
    .Q_N(_2796_),
    .Q(\am_sdr0.det0.yn_1[15] ));
 sg13g2_dfrbp_1 _5804_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net109),
    .D(_0104_),
    .Q_N(_2795_),
    .Q(\am_sdr0.det0.yn_1[16] ));
 sg13g2_dfrbp_1 _5805_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net108),
    .D(_0105_),
    .Q_N(_2794_),
    .Q(\am_sdr0.det0.yn_1[17] ));
 sg13g2_dfrbp_1 _5806_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net107),
    .D(_0106_),
    .Q_N(_2793_),
    .Q(\am_sdr0.det0.yn_1[18] ));
 sg13g2_dfrbp_1 _5807_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net106),
    .D(_0107_),
    .Q_N(_2792_),
    .Q(\am_sdr0.det0.yn_1[19] ));
 sg13g2_dfrbp_1 _5808_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net105),
    .D(_0108_),
    .Q_N(_2791_),
    .Q(\am_sdr0.det0.env_det[0] ));
 sg13g2_dfrbp_1 _5809_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net104),
    .D(_0109_),
    .Q_N(_0023_),
    .Q(\am_sdr0.det0.ifreq[1] ));
 sg13g2_dfrbp_1 _5810_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net103),
    .D(_0110_),
    .Q_N(_0025_),
    .Q(\am_sdr0.det0.ifreq[2] ));
 sg13g2_dfrbp_1 _5811_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net102),
    .D(_0111_),
    .Q_N(_0026_),
    .Q(\am_sdr0.det0.ifreq[3] ));
 sg13g2_dfrbp_1 _5812_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net101),
    .D(_0112_),
    .Q_N(_0027_),
    .Q(\am_sdr0.det0.ifreq[4] ));
 sg13g2_dfrbp_1 _5813_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net100),
    .D(_0113_),
    .Q_N(_0028_),
    .Q(\am_sdr0.det0.ifreq[5] ));
 sg13g2_dfrbp_1 _5814_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net99),
    .D(_0114_),
    .Q_N(_0029_),
    .Q(\am_sdr0.det0.ifreq[6] ));
 sg13g2_dfrbp_1 _5815_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net98),
    .D(_0115_),
    .Q_N(_0024_),
    .Q(\am_sdr0.det0.ifreq[7] ));
 sg13g2_dfrbp_1 _5816_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net97),
    .D(_0116_),
    .Q_N(_2790_),
    .Q(\am_sdr0.filt0.mul_a1[0] ));
 sg13g2_dfrbp_1 _5817_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net96),
    .D(_0117_),
    .Q_N(_2789_),
    .Q(\am_sdr0.filt0.mul_a1[1] ));
 sg13g2_dfrbp_1 _5818_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net95),
    .D(_0118_),
    .Q_N(_2788_),
    .Q(\am_sdr0.filt0.yn_1[2] ));
 sg13g2_dfrbp_1 _5819_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net94),
    .D(_0119_),
    .Q_N(_2787_),
    .Q(\am_sdr0.filt0.yn_1[3] ));
 sg13g2_dfrbp_1 _5820_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net93),
    .D(_0120_),
    .Q_N(_2786_),
    .Q(\am_sdr0.filt0.yn_1[4] ));
 sg13g2_dfrbp_1 _5821_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net92),
    .D(_0121_),
    .Q_N(_2785_),
    .Q(\am_sdr0.filt0.yn_1[5] ));
 sg13g2_dfrbp_1 _5822_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net91),
    .D(_0122_),
    .Q_N(_2784_),
    .Q(\am_sdr0.filt0.yn_1[6] ));
 sg13g2_dfrbp_1 _5823_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net90),
    .D(_0123_),
    .Q_N(_2783_),
    .Q(\am_sdr0.filt0.yn_1[7] ));
 sg13g2_dfrbp_1 _5824_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net89),
    .D(_0124_),
    .Q_N(_2782_),
    .Q(\am_sdr0.filt0.yn_1[8] ));
 sg13g2_dfrbp_1 _5825_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net88),
    .D(_0125_),
    .Q_N(_2781_),
    .Q(\am_sdr0.filt0.yn_1[9] ));
 sg13g2_dfrbp_1 _5826_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net87),
    .D(_0126_),
    .Q_N(_0030_),
    .Q(\am_sdr0.filt0.yn_1[10] ));
 sg13g2_dfrbp_1 _5827_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net86),
    .D(_0127_),
    .Q_N(_2780_),
    .Q(\am_sdr0.filt0.yn_1[11] ));
 sg13g2_dfrbp_1 _5828_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net85),
    .D(_0128_),
    .Q_N(_2779_),
    .Q(\am_sdr0.filt0.yn_1[12] ));
 sg13g2_dfrbp_1 _5829_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net84),
    .D(_0129_),
    .Q_N(_2778_),
    .Q(\am_sdr0.filt0.yn_1[13] ));
 sg13g2_dfrbp_1 _5830_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net83),
    .D(_0130_),
    .Q_N(_2777_),
    .Q(\am_sdr0.filt0.mul_a2[1] ));
 sg13g2_dfrbp_1 _5831_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net82),
    .D(_0131_),
    .Q_N(_2776_),
    .Q(\am_sdr0.filt0.yn_2[1] ));
 sg13g2_dfrbp_1 _5832_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net81),
    .D(_0132_),
    .Q_N(_2775_),
    .Q(\am_sdr0.filt0.yn_2[2] ));
 sg13g2_dfrbp_1 _5833_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net80),
    .D(_0133_),
    .Q_N(_2774_),
    .Q(\am_sdr0.filt0.yn_2[3] ));
 sg13g2_dfrbp_1 _5834_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net79),
    .D(_0134_),
    .Q_N(_2773_),
    .Q(\am_sdr0.filt0.yn_2[4] ));
 sg13g2_dfrbp_1 _5835_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net78),
    .D(_0135_),
    .Q_N(_2772_),
    .Q(\am_sdr0.filt0.yn_2[5] ));
 sg13g2_dfrbp_1 _5836_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net77),
    .D(_0136_),
    .Q_N(_2771_),
    .Q(\am_sdr0.filt0.yn_2[6] ));
 sg13g2_dfrbp_1 _5837_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net76),
    .D(_0137_),
    .Q_N(_2770_),
    .Q(\am_sdr0.filt0.yn_2[7] ));
 sg13g2_dfrbp_1 _5838_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net75),
    .D(_0138_),
    .Q_N(_2769_),
    .Q(\am_sdr0.filt0.yn_2[8] ));
 sg13g2_dfrbp_1 _5839_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net74),
    .D(_0139_),
    .Q_N(_2768_),
    .Q(\am_sdr0.filt0.yn_2[9] ));
 sg13g2_dfrbp_1 _5840_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net73),
    .D(_0140_),
    .Q_N(_2767_),
    .Q(\am_sdr0.filt0.yn_2[10] ));
 sg13g2_dfrbp_1 _5841_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net72),
    .D(_0141_),
    .Q_N(_2766_),
    .Q(\am_sdr0.filt0.yn_2[11] ));
 sg13g2_dfrbp_1 _5842_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net71),
    .D(_0142_),
    .Q_N(_2765_),
    .Q(\am_sdr0.filt0.yn_2[12] ));
 sg13g2_dfrbp_1 _5843_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net70),
    .D(_0143_),
    .Q_N(_0018_),
    .Q(\am_sdr0.filt0.yn_2[13] ));
 sg13g2_dfrbp_1 _5844_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net69),
    .D(_0144_),
    .Q_N(_2764_),
    .Q(\am_sdr0.filt0.xn_1[0] ));
 sg13g2_dfrbp_1 _5845_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net68),
    .D(_0145_),
    .Q_N(_2763_),
    .Q(\am_sdr0.filt0.xn_1[1] ));
 sg13g2_dfrbp_1 _5846_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net67),
    .D(_0146_),
    .Q_N(_2762_),
    .Q(\am_sdr0.filt0.xn_1[2] ));
 sg13g2_dfrbp_1 _5847_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net66),
    .D(_0147_),
    .Q_N(_2761_),
    .Q(\am_sdr0.filt0.xn_1[3] ));
 sg13g2_dfrbp_1 _5848_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net57),
    .D(_0148_),
    .Q_N(_2760_),
    .Q(\am_sdr0.filt0.xn_1[4] ));
 sg13g2_dfrbp_1 _5849_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net56),
    .D(_0149_),
    .Q_N(_2759_),
    .Q(\am_sdr0.filt0.xn_1[5] ));
 sg13g2_dfrbp_1 _5850_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net55),
    .D(_0150_),
    .Q_N(_2758_),
    .Q(\am_sdr0.filt0.xn_1[6] ));
 sg13g2_dfrbp_1 _5851_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net148),
    .D(_0151_),
    .Q_N(_2863_),
    .Q(\am_sdr0.filt0.xn_1[7] ));
 sg13g2_dfrbp_1 _5852_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net149),
    .D(net188),
    .Q_N(_2864_),
    .Q(\am_sdr0.filt0.if_out[0] ));
 sg13g2_dfrbp_1 _5853_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net150),
    .D(net240),
    .Q_N(_0016_),
    .Q(\am_sdr0.filt0.if_out[1] ));
 sg13g2_dfrbp_1 _5854_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net151),
    .D(net221),
    .Q_N(_2865_),
    .Q(\am_sdr0.filt0.if_out[2] ));
 sg13g2_dfrbp_1 _5855_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net152),
    .D(net213),
    .Q_N(_2866_),
    .Q(\am_sdr0.filt0.if_out[3] ));
 sg13g2_dfrbp_1 _5856_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net153),
    .D(net215),
    .Q_N(_2867_),
    .Q(\am_sdr0.filt0.if_out[4] ));
 sg13g2_dfrbp_1 _5857_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net154),
    .D(net207),
    .Q_N(_2868_),
    .Q(\am_sdr0.filt0.if_out[5] ));
 sg13g2_dfrbp_1 _5858_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net157),
    .D(net203),
    .Q_N(_2869_),
    .Q(\am_sdr0.filt0.if_out[6] ));
 sg13g2_dfrbp_1 _5859_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net54),
    .D(net205),
    .Q_N(_0019_),
    .Q(\am_sdr0.filt0.if_out[7] ));
 sg13g2_dfrbp_1 _5860_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net53),
    .D(_0152_),
    .Q_N(_2757_),
    .Q(\am_sdr0.filt0.mul_b2[0] ));
 sg13g2_dfrbp_1 _5861_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net52),
    .D(_0153_),
    .Q_N(_2756_),
    .Q(\am_sdr0.filt0.xn_2[1] ));
 sg13g2_dfrbp_1 _5862_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net51),
    .D(_0154_),
    .Q_N(_2755_),
    .Q(\am_sdr0.filt0.xn_2[2] ));
 sg13g2_dfrbp_1 _5863_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net50),
    .D(_0155_),
    .Q_N(_2754_),
    .Q(\am_sdr0.filt0.xn_2[3] ));
 sg13g2_dfrbp_1 _5864_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net49),
    .D(_0156_),
    .Q_N(_2753_),
    .Q(\am_sdr0.filt0.xn_2[4] ));
 sg13g2_dfrbp_1 _5865_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net48),
    .D(_0157_),
    .Q_N(_2752_),
    .Q(\am_sdr0.filt0.xn_2[5] ));
 sg13g2_dfrbp_1 _5866_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net47),
    .D(_0158_),
    .Q_N(_2751_),
    .Q(\am_sdr0.filt0.xn_2[6] ));
 sg13g2_dfrbp_1 _5867_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net46),
    .D(_0159_),
    .Q_N(_0015_),
    .Q(\am_sdr0.filt0.xn_2[7] ));
 sg13g2_dfrbp_1 _5868_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net45),
    .D(net230),
    .Q_N(_2750_),
    .Q(\am_sdr0.nco0.nco_phase[0] ));
 sg13g2_dfrbp_1 _5869_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net43),
    .D(_0161_),
    .Q_N(_2749_),
    .Q(\am_sdr0.nco0.nco_phase[1] ));
 sg13g2_dfrbp_1 _5870_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net41),
    .D(_0162_),
    .Q_N(_2748_),
    .Q(\am_sdr0.nco0.nco_phase[2] ));
 sg13g2_dfrbp_1 _5871_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net39),
    .D(_0163_),
    .Q_N(_2747_),
    .Q(\am_sdr0.nco0.nco_phase[3] ));
 sg13g2_dfrbp_1 _5872_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net37),
    .D(_0164_),
    .Q_N(_2746_),
    .Q(\am_sdr0.nco0.nco_phase[4] ));
 sg13g2_dfrbp_1 _5873_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net35),
    .D(_0165_),
    .Q_N(_2745_),
    .Q(\am_sdr0.nco0.nco_phase[5] ));
 sg13g2_dfrbp_1 _5874_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net33),
    .D(_0166_),
    .Q_N(_2744_),
    .Q(\am_sdr0.nco0.nco_phase[6] ));
 sg13g2_dfrbp_1 _5875_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net31),
    .D(_0167_),
    .Q_N(_2743_),
    .Q(\am_sdr0.nco0.nco_phase[7] ));
 sg13g2_dfrbp_1 _5876_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net29),
    .D(net306),
    .Q_N(_2742_),
    .Q(\am_sdr0.nco0.nco_phase[8] ));
 sg13g2_dfrbp_1 _5877_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net27),
    .D(net301),
    .Q_N(_2741_),
    .Q(\am_sdr0.nco0.nco_phase[9] ));
 sg13g2_dfrbp_1 _5878_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net185),
    .D(_0170_),
    .Q_N(_2740_),
    .Q(\am_sdr0.nco0.nco_phase[10] ));
 sg13g2_dfrbp_1 _5879_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net183),
    .D(_0171_),
    .Q_N(_2739_),
    .Q(\am_sdr0.nco0.nco_phase[11] ));
 sg13g2_dfrbp_1 _5880_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net181),
    .D(net313),
    .Q_N(_2738_),
    .Q(\am_sdr0.nco0.nco_phase[12] ));
 sg13g2_dfrbp_1 _5881_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net179),
    .D(net309),
    .Q_N(_2737_),
    .Q(\am_sdr0.nco0.nco_phase[13] ));
 sg13g2_dfrbp_1 _5882_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net177),
    .D(_0174_),
    .Q_N(_2736_),
    .Q(\am_sdr0.nco0.nco_phase[14] ));
 sg13g2_dfrbp_1 _5883_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net175),
    .D(net299),
    .Q_N(_2735_),
    .Q(\am_sdr0.nco0.nco_phase[15] ));
 sg13g2_dfrbp_1 _5884_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net173),
    .D(_0176_),
    .Q_N(_2734_),
    .Q(\am_sdr0.nco0.nco_phase[16] ));
 sg13g2_dfrbp_1 _5885_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net171),
    .D(_0177_),
    .Q_N(_2733_),
    .Q(\am_sdr0.nco0.nco_phase[17] ));
 sg13g2_dfrbp_1 _5886_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net169),
    .D(_0178_),
    .Q_N(_2732_),
    .Q(\am_sdr0.nco0.nco_phase[18] ));
 sg13g2_dfrbp_1 _5887_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net167),
    .D(_0179_),
    .Q_N(_2731_),
    .Q(\am_sdr0.nco0.nco_phase[19] ));
 sg13g2_dfrbp_1 _5888_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net165),
    .D(_0180_),
    .Q_N(_2730_),
    .Q(\am_sdr0.nco0.rf_a ));
 sg13g2_dfrbp_1 _5889_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net163),
    .D(_0181_),
    .Q_N(_2729_),
    .Q(\am_sdr0.spi0.MOSI_q ));
 sg13g2_dfrbp_1 _5890_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net161),
    .D(_0182_),
    .Q_N(_2728_),
    .Q(\am_sdr0.spi0.SCK_qqq ));
 sg13g2_dfrbp_1 _5891_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net159),
    .D(_0183_),
    .Q_N(_2727_),
    .Q(\am_sdr0.spi0.SCK_qq ));
 sg13g2_tiehi _5741__28 (.L_HI(net28));
 sg13g2_tiehi _5876__29 (.L_HI(net29));
 sg13g2_tiehi _5740__30 (.L_HI(net30));
 sg13g2_tiehi _5875__31 (.L_HI(net31));
 sg13g2_tiehi _5739__32 (.L_HI(net32));
 sg13g2_tiehi _5874__33 (.L_HI(net33));
 sg13g2_tiehi _5738__34 (.L_HI(net34));
 sg13g2_tiehi _5873__35 (.L_HI(net35));
 sg13g2_tiehi _5737__36 (.L_HI(net36));
 sg13g2_tiehi _5872__37 (.L_HI(net37));
 sg13g2_tiehi _5736__38 (.L_HI(net38));
 sg13g2_tiehi _5871__39 (.L_HI(net39));
 sg13g2_tiehi _5735__40 (.L_HI(net40));
 sg13g2_tiehi _5870__41 (.L_HI(net41));
 sg13g2_tiehi _5734__42 (.L_HI(net42));
 sg13g2_tiehi _5869__43 (.L_HI(net43));
 sg13g2_tiehi _5733__44 (.L_HI(net44));
 sg13g2_tiehi _5868__45 (.L_HI(net45));
 sg13g2_tiehi _5867__46 (.L_HI(net46));
 sg13g2_tiehi _5866__47 (.L_HI(net47));
 sg13g2_tiehi _5865__48 (.L_HI(net48));
 sg13g2_tiehi _5864__49 (.L_HI(net49));
 sg13g2_tiehi _5863__50 (.L_HI(net50));
 sg13g2_tiehi _5862__51 (.L_HI(net51));
 sg13g2_tiehi _5861__52 (.L_HI(net52));
 sg13g2_tiehi _5860__53 (.L_HI(net53));
 sg13g2_tiehi _5859__54 (.L_HI(net54));
 sg13g2_tiehi _5850__55 (.L_HI(net55));
 sg13g2_tiehi _5849__56 (.L_HI(net56));
 sg13g2_tiehi _5848__57 (.L_HI(net57));
 sg13g2_tiehi _5732__58 (.L_HI(net58));
 sg13g2_tiehi _5762__59 (.L_HI(net59));
 sg13g2_tiehi _5763__60 (.L_HI(net60));
 sg13g2_tiehi _5764__61 (.L_HI(net61));
 sg13g2_tiehi _5765__62 (.L_HI(net62));
 sg13g2_tiehi _5766__63 (.L_HI(net63));
 sg13g2_tiehi _5767__64 (.L_HI(net64));
 sg13g2_tiehi _5768__65 (.L_HI(net65));
 sg13g2_tiehi _5847__66 (.L_HI(net66));
 sg13g2_tiehi _5846__67 (.L_HI(net67));
 sg13g2_tiehi _5845__68 (.L_HI(net68));
 sg13g2_tiehi _5844__69 (.L_HI(net69));
 sg13g2_tiehi _5843__70 (.L_HI(net70));
 sg13g2_tiehi _5842__71 (.L_HI(net71));
 sg13g2_tiehi _5841__72 (.L_HI(net72));
 sg13g2_tiehi _5840__73 (.L_HI(net73));
 sg13g2_tiehi _5839__74 (.L_HI(net74));
 sg13g2_tiehi _5838__75 (.L_HI(net75));
 sg13g2_tiehi _5837__76 (.L_HI(net76));
 sg13g2_tiehi _5836__77 (.L_HI(net77));
 sg13g2_tiehi _5835__78 (.L_HI(net78));
 sg13g2_tiehi _5834__79 (.L_HI(net79));
 sg13g2_tiehi _5833__80 (.L_HI(net80));
 sg13g2_tiehi _5832__81 (.L_HI(net81));
 sg13g2_tiehi _5831__82 (.L_HI(net82));
 sg13g2_tiehi _5830__83 (.L_HI(net83));
 sg13g2_tiehi _5829__84 (.L_HI(net84));
 sg13g2_tiehi _5828__85 (.L_HI(net85));
 sg13g2_tiehi _5827__86 (.L_HI(net86));
 sg13g2_tiehi _5826__87 (.L_HI(net87));
 sg13g2_tiehi _5825__88 (.L_HI(net88));
 sg13g2_tiehi _5824__89 (.L_HI(net89));
 sg13g2_tiehi _5823__90 (.L_HI(net90));
 sg13g2_tiehi _5822__91 (.L_HI(net91));
 sg13g2_tiehi _5821__92 (.L_HI(net92));
 sg13g2_tiehi _5820__93 (.L_HI(net93));
 sg13g2_tiehi _5819__94 (.L_HI(net94));
 sg13g2_tiehi _5818__95 (.L_HI(net95));
 sg13g2_tiehi _5817__96 (.L_HI(net96));
 sg13g2_tiehi _5816__97 (.L_HI(net97));
 sg13g2_tiehi _5815__98 (.L_HI(net98));
 sg13g2_tiehi _5814__99 (.L_HI(net99));
 sg13g2_tiehi _5813__100 (.L_HI(net100));
 sg13g2_tiehi _5812__101 (.L_HI(net101));
 sg13g2_tiehi _5811__102 (.L_HI(net102));
 sg13g2_tiehi _5810__103 (.L_HI(net103));
 sg13g2_tiehi _5809__104 (.L_HI(net104));
 sg13g2_tiehi _5808__105 (.L_HI(net105));
 sg13g2_tiehi _5807__106 (.L_HI(net106));
 sg13g2_tiehi _5806__107 (.L_HI(net107));
 sg13g2_tiehi _5805__108 (.L_HI(net108));
 sg13g2_tiehi _5804__109 (.L_HI(net109));
 sg13g2_tiehi _5803__110 (.L_HI(net110));
 sg13g2_tiehi _5802__111 (.L_HI(net111));
 sg13g2_tiehi _5801__112 (.L_HI(net112));
 sg13g2_tiehi _5800__113 (.L_HI(net113));
 sg13g2_tiehi _5799__114 (.L_HI(net114));
 sg13g2_tiehi _5798__115 (.L_HI(net115));
 sg13g2_tiehi _5797__116 (.L_HI(net116));
 sg13g2_tiehi _5796__117 (.L_HI(net117));
 sg13g2_tiehi _5795__118 (.L_HI(net118));
 sg13g2_tiehi _5794__119 (.L_HI(net119));
 sg13g2_tiehi _5793__120 (.L_HI(net120));
 sg13g2_tiehi _5792__121 (.L_HI(net121));
 sg13g2_tiehi _5791__122 (.L_HI(net122));
 sg13g2_tiehi _5790__123 (.L_HI(net123));
 sg13g2_tiehi _5789__124 (.L_HI(net124));
 sg13g2_tiehi _5788__125 (.L_HI(net125));
 sg13g2_tiehi _5787__126 (.L_HI(net126));
 sg13g2_tiehi _5786__127 (.L_HI(net127));
 sg13g2_tiehi _5785__128 (.L_HI(net128));
 sg13g2_tiehi _5784__129 (.L_HI(net129));
 sg13g2_tiehi _5783__130 (.L_HI(net130));
 sg13g2_tiehi _5782__131 (.L_HI(net131));
 sg13g2_tiehi _5781__132 (.L_HI(net132));
 sg13g2_tiehi _5780__133 (.L_HI(net133));
 sg13g2_tiehi _5779__134 (.L_HI(net134));
 sg13g2_tiehi _5778__135 (.L_HI(net135));
 sg13g2_tiehi _5777__136 (.L_HI(net136));
 sg13g2_tiehi _5776__137 (.L_HI(net137));
 sg13g2_tiehi _5775__138 (.L_HI(net138));
 sg13g2_tiehi _5774__139 (.L_HI(net139));
 sg13g2_tiehi _5773__140 (.L_HI(net140));
 sg13g2_tiehi _5772__141 (.L_HI(net141));
 sg13g2_tiehi _5771__142 (.L_HI(net142));
 sg13g2_tiehi _5770__143 (.L_HI(net143));
 sg13g2_tiehi _5761__144 (.L_HI(net144));
 sg13g2_tiehi _5760__145 (.L_HI(net145));
 sg13g2_tiehi _5759__146 (.L_HI(net146));
 sg13g2_tiehi _5769__147 (.L_HI(net147));
 sg13g2_tiehi _5851__148 (.L_HI(net148));
 sg13g2_tiehi _5852__149 (.L_HI(net149));
 sg13g2_tiehi _5853__150 (.L_HI(net150));
 sg13g2_tiehi _5854__151 (.L_HI(net151));
 sg13g2_tiehi _5855__152 (.L_HI(net152));
 sg13g2_tiehi _5856__153 (.L_HI(net153));
 sg13g2_tiehi _5857__154 (.L_HI(net154));
 sg13g2_tiehi _5758__155 (.L_HI(net155));
 sg13g2_tiehi _5757__156 (.L_HI(net156));
 sg13g2_tiehi _5858__157 (.L_HI(net157));
 sg13g2_tiehi _5756__158 (.L_HI(net158));
 sg13g2_tiehi _5891__159 (.L_HI(net159));
 sg13g2_tiehi _5755__160 (.L_HI(net160));
 sg13g2_tiehi _5890__161 (.L_HI(net161));
 sg13g2_tiehi _5754__162 (.L_HI(net162));
 sg13g2_tiehi _5889__163 (.L_HI(net163));
 sg13g2_tiehi _5753__164 (.L_HI(net164));
 sg13g2_tiehi _5888__165 (.L_HI(net165));
 sg13g2_tiehi _5752__166 (.L_HI(net166));
 sg13g2_tiehi _5887__167 (.L_HI(net167));
 sg13g2_tiehi _5751__168 (.L_HI(net168));
 sg13g2_tiehi _5886__169 (.L_HI(net169));
 sg13g2_tiehi _5750__170 (.L_HI(net170));
 sg13g2_tiehi _5885__171 (.L_HI(net171));
 sg13g2_tiehi _5749__172 (.L_HI(net172));
 sg13g2_tiehi _5884__173 (.L_HI(net173));
 sg13g2_tiehi _5748__174 (.L_HI(net174));
 sg13g2_tiehi _5883__175 (.L_HI(net175));
 sg13g2_tiehi _5747__176 (.L_HI(net176));
 sg13g2_tiehi _5882__177 (.L_HI(net177));
 sg13g2_tiehi _5746__178 (.L_HI(net178));
 sg13g2_tiehi _5881__179 (.L_HI(net179));
 sg13g2_tiehi _5745__180 (.L_HI(net180));
 sg13g2_tiehi _5880__181 (.L_HI(net181));
 sg13g2_tiehi _5744__182 (.L_HI(net182));
 sg13g2_tiehi _5879__183 (.L_HI(net183));
 sg13g2_tiehi _5743__184 (.L_HI(net184));
 sg13g2_tiehi _5878__185 (.L_HI(net185));
 sg13g2_tiehi _5742__186 (.L_HI(net186));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_6 (.L_LO(net6));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_7 (.L_LO(net7));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_8 (.L_LO(net8));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_9 (.L_LO(net9));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_10 (.L_LO(net10));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_11 (.L_LO(net11));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_12 (.L_LO(net12));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_13 (.L_LO(net13));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_14 (.L_LO(net14));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_15 (.L_LO(net15));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_16 (.L_LO(net16));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_17 (.L_LO(net17));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_18 (.L_LO(net18));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_19 (.L_LO(net19));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_20 (.L_LO(net20));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_21 (.L_LO(net21));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_22 (.L_LO(net22));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_23 (.L_LO(net23));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_24 (.L_LO(net24));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_25 (.L_LO(net25));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_26 (.L_LO(net26));
 sg13g2_tiehi _5877__27 (.L_HI(net27));
 sg13g2_buf_1 _6074_ (.A(COMP_OUT),
    .X(uo_out[0]));
 sg13g2_buf_2 _6075_ (.A(PWM_OUT),
    .X(uo_out[1]));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_1313_));
 sg13g2_buf_1 fanout327 (.A(_1313_),
    .X(net327));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_1312_));
 sg13g2_buf_2 fanout329 (.A(_1312_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_2699_),
    .X(net330));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(net332));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_2277_));
 sg13g2_buf_2 fanout333 (.A(_1666_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(net337),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(net337),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net337),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_2275_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(net339),
    .X(net338));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_2278_));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(net341));
 sg13g2_buf_2 fanout341 (.A(_0479_),
    .X(net341));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(_0479_));
 sg13g2_buf_2 fanout343 (.A(_2273_),
    .X(net343));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_2160_));
 sg13g2_buf_1 fanout345 (.A(_2160_),
    .X(net345));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(net347));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_0019_));
 sg13g2_buf_2 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(net350),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(\am_sdr0.filt0.yn_2[13] ),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(\am_sdr0.filt0.yn_2[12] ),
    .X(net353));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(net356));
 sg13g2_buf_2 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_1 fanout356 (.A(\am_sdr0.filt0.yn_2[11] ),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(net359),
    .X(net357));
 sg13g2_buf_1 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(\am_sdr0.filt0.yn_2[10] ),
    .X(net359));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(net361));
 sg13g2_buf_2 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(\am_sdr0.filt0.yn_2[9] ),
    .X(net362));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(net364));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(\am_sdr0.filt0.yn_2[8] ));
 sg13g2_buf_2 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(\am_sdr0.filt0.yn_2[7] ));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(\am_sdr0.filt0.yn_2[6] ));
 sg13g2_buf_2 fanout368 (.A(\am_sdr0.filt0.yn_2[6] ),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(net370));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(\am_sdr0.filt0.yn_2[5] ));
 sg13g2_buf_2 fanout371 (.A(\am_sdr0.filt0.yn_2[4] ),
    .X(net371));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(\am_sdr0.filt0.yn_2[4] ));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(\am_sdr0.filt0.yn_2[3] ));
 sg13g2_buf_2 fanout374 (.A(\am_sdr0.filt0.yn_2[3] ),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(\am_sdr0.filt0.yn_2[2] ));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(\am_sdr0.filt0.yn_2[1] ));
 sg13g2_buf_4 fanout378 (.X(net378),
    .A(\am_sdr0.filt0.mul_a2[1] ));
 sg13g2_buf_2 fanout379 (.A(net380),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(net381),
    .X(net380));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(\am_sdr0.filt0.yn_1[13] ));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(net285));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(net284));
 sg13g2_buf_2 fanout384 (.A(\am_sdr0.filt0.yn_1[11] ),
    .X(net384));
 sg13g2_buf_4 fanout385 (.X(net385),
    .A(net317));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(net296));
 sg13g2_buf_2 fanout387 (.A(\am_sdr0.filt0.yn_1[9] ),
    .X(net387));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(net302));
 sg13g2_buf_2 fanout389 (.A(\am_sdr0.filt0.yn_1[8] ),
    .X(net389));
 sg13g2_buf_4 fanout390 (.X(net390),
    .A(net434));
 sg13g2_buf_4 fanout391 (.X(net391),
    .A(net303));
 sg13g2_buf_2 fanout392 (.A(\am_sdr0.filt0.yn_1[6] ),
    .X(net392));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(net310));
 sg13g2_buf_2 fanout394 (.A(\am_sdr0.filt0.yn_1[5] ),
    .X(net394));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(\am_sdr0.filt0.yn_1[4] ));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(net320));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(\am_sdr0.filt0.yn_1[2] ));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(\am_sdr0.filt0.mul_a1[0] ));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(\am_sdr0.det0.yn_1[19] ));
 sg13g2_buf_2 fanout400 (.A(net401),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(\am_sdr0.det0.yn_1[18] ),
    .X(net401));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(\am_sdr0.det0.yn_1[17] ));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(\am_sdr0.det0.yn_1[16] ));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(\am_sdr0.det0.yn_1[7] ));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(\am_sdr0.det0.yn_1[6] ));
 sg13g2_buf_2 fanout406 (.A(net410),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(net410),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_2144_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(net412),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(net413),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(net427));
 sg13g2_buf_2 fanout415 (.A(net416),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(net427),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(net418),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(net427),
    .X(net418));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(net421));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(net421));
 sg13g2_buf_2 fanout421 (.A(net427),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(net426),
    .X(net422));
 sg13g2_buf_1 fanout423 (.A(net426),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(net426),
    .X(net424));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(net426));
 sg13g2_buf_2 fanout426 (.A(net427),
    .X(net426));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_jamesrosssharp_tiny1bitam_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0039_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0031_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold3 (.A(\am_sdr0.filt0.xn_1[5] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold4 (.A(\am_sdr0.filt0.xn_1[6] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold5 (.A(\am_sdr0.nco0.rf_a ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold6 (.A(\am_sdr0.spi0.MOSI_q ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold7 (.A(\am_sdr0.filt0.xn_1[3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold8 (.A(\am_sdr0.spi0.CS_q ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold9 (.A(\am_sdr0.filt0.xn_1[4] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold10 (.A(\am_sdr0.filt0.xn_1[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold11 (.A(\am_sdr0.filt0.xn_1[1] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold12 (.A(\am_sdr0.spi0.SCK_q ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold13 (.A(\am_sdr0.filt0.xn_1[7] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold14 (.A(\am_sdr0.filt0.xn_1[0] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0037_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold16 (.A(_2268_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0013_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0038_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0014_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0036_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0012_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold22 (.A(\am_sdr0.spi0.SCK_qq ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold23 (.A(\am_sdr0.spi0.MOSI_qq ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold24 (.A(_2279_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0040_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0034_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0010_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0035_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0011_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold30 (.A(\am_sdr0.count[6] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold31 (.A(_2334_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0078_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold33 (.A(\am_sdr0.filt0.mul_a1[0] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0033_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0009_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold36 (.A(\am_sdr0.spi0.CS_qq ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold37 (.A(\am_sdr0.det0.env_out[2] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold38 (.A(\am_sdr0.count[0] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0073_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold40 (.A(\am_sdr0.count[2] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold41 (.A(_2326_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold42 (.A(\am_sdr0.nco0.nco_phase[0] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold43 (.A(_2106_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0160_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold45 (.A(\am_sdr0.spi0.CS_qqq ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold46 (.A(\am_sdr0.nco0.phase_inc[5] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0046_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold48 (.A(\am_sdr0.det0.env_out[0] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold49 (.A(\am_sdr0.det0.env_out[1] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold50 (.A(\am_sdr0.nco0.phase_inc[6] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0047_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold52 (.A(\am_sdr0.det0.env_out[3] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0032_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0008_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold55 (.A(\am_sdr0.nco0.phase_inc[12] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0053_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold57 (.A(\am_sdr0.nco0.phase_inc[0] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0041_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold59 (.A(\am_sdr0.nco0.phase_inc[11] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold60 (.A(\am_sdr0.filt0.gain_spi[2] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0062_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold62 (.A(\am_sdr0.det0.env_out[6] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold63 (.A(\am_sdr0.nco0.phase_inc[8] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0049_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold65 (.A(\am_sdr0.nco0.phase_inc[19] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0060_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold67 (.A(\am_sdr0.count[7] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0079_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold69 (.A(\am_sdr0.det0.env_out[4] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold70 (.A(\am_sdr0.det0.env_out[5] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold71 (.A(\am_sdr0.nco0.phase_inc[15] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0056_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold73 (.A(\am_sdr0.nco0.phase_inc[16] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0057_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold75 (.A(\am_sdr0.nco0.phase_inc[18] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold76 (.A(\am_sdr0.det0.env_out[7] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold77 (.A(\am_sdr0.count[5] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold78 (.A(\am_sdr0.filt0.if_out[7] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold79 (.A(\am_sdr0.count[4] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold80 (.A(_2332_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0076_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold82 (.A(\am_sdr0.nco0.phase_inc[7] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold83 (.A(_2288_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold84 (.A(\am_sdr0.nco0.phase_inc[10] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold85 (.A(\am_sdr0.nco0.phase_inc[4] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold86 (.A(\am_sdr0.filt0.yn_1[2] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold87 (.A(\am_sdr0.nco0.phase_inc[3] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold88 (.A(\am_sdr0.nco0.phase_inc[13] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0054_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold90 (.A(\am_sdr0.nco0.phase_inc[9] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold91 (.A(\am_sdr0.nco0.phase_inc[17] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold92 (.A(\am_sdr0.nco0.phase_inc[1] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0042_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold94 (.A(\am_sdr0.nco0.phase_inc[2] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold95 (.A(\am_sdr0.nco0.phase_inc[14] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold96 (.A(\am_sdr0.filt0.yn_1[4] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold97 (.A(\am_sdr0.count[3] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold98 (.A(\am_sdr0.filt0.yn_1[11] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold99 (.A(\am_sdr0.filt0.yn_1[12] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold100 (.A(\am_sdr0.filt0.if_out[6] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold101 (.A(\am_sdr0.det0.env_det[0] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold102 (.A(\am_sdr0.filt0.if_out[0] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold103 (.A(\am_sdr0.filt0.if_out[3] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold104 (.A(\am_sdr0.filt0.gain_spi[0] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0061_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold106 (.A(\am_sdr0.filt0.if_out[2] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold107 (.A(\am_sdr0.spi0.state[0] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold108 (.A(_2272_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold109 (.A(_2311_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold110 (.A(\am_sdr0.filt0.yn_1[9] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold111 (.A(\am_sdr0.filt0.if_out[5] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold112 (.A(\am_sdr0.nco0.nco_phase[15] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0175_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold114 (.A(\am_sdr0.nco0.nco_phase[9] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0169_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold116 (.A(\am_sdr0.filt0.yn_1[8] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold117 (.A(\am_sdr0.filt0.yn_1[6] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold118 (.A(\am_sdr0.nco0.nco_phase[7] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold119 (.A(_2114_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0168_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold121 (.A(\am_sdr0.filt0.if_out[4] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold122 (.A(\am_sdr0.nco0.nco_phase[13] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0173_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold124 (.A(\am_sdr0.filt0.yn_1[5] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold125 (.A(\am_sdr0.filt0.if_out[1] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold126 (.A(\am_sdr0.nco0.nco_phase[12] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0172_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold128 (.A(\am_sdr0.nco0.nco_phase[10] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold129 (.A(_2214_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold130 (.A(\am_sdr0.nco0.nco_phase[11] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold131 (.A(\am_sdr0.filt0.yn_1[10] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold132 (.A(\am_sdr0.nco0.nco_phase[4] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold133 (.A(_2111_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold134 (.A(\am_sdr0.filt0.yn_1[3] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold135 (.A(\am_sdr0.filt0.mul_a1[1] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold136 (.A(\am_sdr0.nco0.nco_phase[6] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold137 (.A(\am_sdr0.nco0.nco_phase[3] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold138 (.A(_2110_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold139 (.A(\am_sdr0.nco0.nco_phase[1] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold140 (.A(_2196_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold141 (.A(\am_sdr0.nco0.nco_phase[5] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0029_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0095_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold144 (.A(\am_sdr0.nco0.nco_phase[2] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold145 (.A(\am_sdr0.nco0.nco_phase[2] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold146 (.A(\am_sdr0.filt0.yn_1[7] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold147 (.A(\am_sdr0.nco0.nco_phase[14] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold148 (.A(_2180_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold149 (.A(\am_sdr0.filt0.gain_spi[1] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0025_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0017_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0017_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0027_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0017_),
    .X(net442));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_4 FILLER_0_189 ();
 sg13g2_fill_1 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_fill_2 FILLER_0_219 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_4 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_4 FILLER_0_262 ();
 sg13g2_fill_2 FILLER_0_266 ();
 sg13g2_decap_4 FILLER_0_273 ();
 sg13g2_fill_1 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_fill_2 FILLER_0_296 ();
 sg13g2_fill_1 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_4 FILLER_0_310 ();
 sg13g2_fill_2 FILLER_0_314 ();
 sg13g2_fill_2 FILLER_0_320 ();
 sg13g2_fill_2 FILLER_0_326 ();
 sg13g2_fill_1 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_333 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_decap_8 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_4 FILLER_1_182 ();
 sg13g2_fill_1 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_232 ();
 sg13g2_decap_4 FILLER_1_239 ();
 sg13g2_fill_1 FILLER_1_259 ();
 sg13g2_fill_2 FILLER_1_273 ();
 sg13g2_fill_2 FILLER_1_288 ();
 sg13g2_fill_2 FILLER_1_298 ();
 sg13g2_fill_1 FILLER_1_300 ();
 sg13g2_fill_1 FILLER_1_314 ();
 sg13g2_fill_1 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_4 FILLER_2_168 ();
 sg13g2_fill_2 FILLER_2_172 ();
 sg13g2_fill_2 FILLER_2_195 ();
 sg13g2_fill_1 FILLER_2_197 ();
 sg13g2_fill_2 FILLER_2_205 ();
 sg13g2_fill_1 FILLER_2_207 ();
 sg13g2_fill_2 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_fill_2 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_170 ();
 sg13g2_fill_2 FILLER_3_193 ();
 sg13g2_decap_4 FILLER_3_235 ();
 sg13g2_fill_1 FILLER_3_239 ();
 sg13g2_fill_1 FILLER_3_279 ();
 sg13g2_fill_2 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_324 ();
 sg13g2_fill_2 FILLER_3_338 ();
 sg13g2_fill_1 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_fill_2 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_198 ();
 sg13g2_fill_1 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_fill_1 FILLER_4_216 ();
 sg13g2_decap_8 FILLER_4_230 ();
 sg13g2_decap_8 FILLER_4_237 ();
 sg13g2_decap_8 FILLER_4_244 ();
 sg13g2_fill_1 FILLER_4_260 ();
 sg13g2_decap_4 FILLER_4_270 ();
 sg13g2_fill_1 FILLER_4_274 ();
 sg13g2_fill_2 FILLER_4_279 ();
 sg13g2_fill_1 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_fill_2 FILLER_4_319 ();
 sg13g2_decap_4 FILLER_4_326 ();
 sg13g2_fill_1 FILLER_4_330 ();
 sg13g2_decap_4 FILLER_4_335 ();
 sg13g2_fill_1 FILLER_4_339 ();
 sg13g2_fill_2 FILLER_4_350 ();
 sg13g2_decap_4 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_4 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_172 ();
 sg13g2_fill_2 FILLER_5_204 ();
 sg13g2_fill_1 FILLER_5_206 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_fill_2 FILLER_5_266 ();
 sg13g2_fill_2 FILLER_5_281 ();
 sg13g2_fill_1 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_fill_2 FILLER_5_311 ();
 sg13g2_fill_1 FILLER_5_313 ();
 sg13g2_decap_4 FILLER_5_335 ();
 sg13g2_fill_1 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_4 FILLER_6_185 ();
 sg13g2_fill_2 FILLER_6_189 ();
 sg13g2_decap_4 FILLER_6_203 ();
 sg13g2_fill_2 FILLER_6_220 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_fill_2 FILLER_6_236 ();
 sg13g2_fill_1 FILLER_6_238 ();
 sg13g2_fill_2 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_276 ();
 sg13g2_fill_2 FILLER_6_283 ();
 sg13g2_fill_1 FILLER_6_289 ();
 sg13g2_fill_2 FILLER_6_333 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_fill_2 FILLER_6_341 ();
 sg13g2_fill_1 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_fill_1 FILLER_7_161 ();
 sg13g2_fill_1 FILLER_7_183 ();
 sg13g2_decap_8 FILLER_7_192 ();
 sg13g2_fill_2 FILLER_7_207 ();
 sg13g2_decap_4 FILLER_7_213 ();
 sg13g2_fill_1 FILLER_7_217 ();
 sg13g2_fill_2 FILLER_7_230 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_fill_2 FILLER_7_249 ();
 sg13g2_fill_1 FILLER_7_251 ();
 sg13g2_decap_4 FILLER_7_275 ();
 sg13g2_fill_2 FILLER_7_358 ();
 sg13g2_fill_1 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_4 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_decap_4 FILLER_8_177 ();
 sg13g2_fill_2 FILLER_8_202 ();
 sg13g2_fill_2 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_235 ();
 sg13g2_fill_2 FILLER_8_241 ();
 sg13g2_fill_1 FILLER_8_243 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_4 FILLER_8_256 ();
 sg13g2_fill_2 FILLER_8_293 ();
 sg13g2_fill_1 FILLER_8_322 ();
 sg13g2_decap_4 FILLER_8_331 ();
 sg13g2_fill_1 FILLER_8_335 ();
 sg13g2_fill_2 FILLER_8_358 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_60 ();
 sg13g2_fill_1 FILLER_9_78 ();
 sg13g2_fill_2 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_90 ();
 sg13g2_decap_8 FILLER_9_97 ();
 sg13g2_decap_8 FILLER_9_104 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_decap_8 FILLER_9_118 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_132 ();
 sg13g2_decap_8 FILLER_9_139 ();
 sg13g2_decap_8 FILLER_9_146 ();
 sg13g2_fill_2 FILLER_9_174 ();
 sg13g2_fill_1 FILLER_9_176 ();
 sg13g2_decap_4 FILLER_9_190 ();
 sg13g2_fill_2 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_fill_2 FILLER_9_228 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_236 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_4 FILLER_9_273 ();
 sg13g2_fill_2 FILLER_9_304 ();
 sg13g2_fill_1 FILLER_9_306 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_4 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_332 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_4 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_56 ();
 sg13g2_fill_2 FILLER_10_83 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_4 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_164 ();
 sg13g2_decap_4 FILLER_10_179 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_fill_2 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_4 FILLER_10_249 ();
 sg13g2_fill_2 FILLER_10_253 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_fill_1 FILLER_10_287 ();
 sg13g2_decap_4 FILLER_10_296 ();
 sg13g2_fill_1 FILLER_10_300 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_fill_2 FILLER_10_314 ();
 sg13g2_fill_1 FILLER_10_316 ();
 sg13g2_fill_2 FILLER_10_346 ();
 sg13g2_fill_1 FILLER_10_348 ();
 sg13g2_fill_1 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_55 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_decap_8 FILLER_11_117 ();
 sg13g2_decap_8 FILLER_11_124 ();
 sg13g2_decap_8 FILLER_11_131 ();
 sg13g2_decap_8 FILLER_11_138 ();
 sg13g2_decap_8 FILLER_11_145 ();
 sg13g2_decap_4 FILLER_11_152 ();
 sg13g2_fill_2 FILLER_11_156 ();
 sg13g2_fill_2 FILLER_11_192 ();
 sg13g2_fill_2 FILLER_11_204 ();
 sg13g2_decap_4 FILLER_11_224 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_decap_4 FILLER_11_233 ();
 sg13g2_fill_1 FILLER_11_237 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_decap_4 FILLER_11_276 ();
 sg13g2_fill_2 FILLER_11_284 ();
 sg13g2_fill_1 FILLER_11_303 ();
 sg13g2_fill_1 FILLER_11_308 ();
 sg13g2_fill_1 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_28 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_1 FILLER_12_54 ();
 sg13g2_fill_2 FILLER_12_87 ();
 sg13g2_fill_1 FILLER_12_94 ();
 sg13g2_decap_8 FILLER_12_108 ();
 sg13g2_decap_8 FILLER_12_115 ();
 sg13g2_decap_8 FILLER_12_122 ();
 sg13g2_decap_8 FILLER_12_129 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_150 ();
 sg13g2_fill_2 FILLER_12_171 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_234 ();
 sg13g2_fill_1 FILLER_12_236 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_fill_1 FILLER_12_273 ();
 sg13g2_fill_1 FILLER_12_278 ();
 sg13g2_fill_2 FILLER_12_300 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_decap_4 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_61 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_143 ();
 sg13g2_decap_8 FILLER_13_150 ();
 sg13g2_fill_2 FILLER_13_157 ();
 sg13g2_fill_1 FILLER_13_159 ();
 sg13g2_fill_1 FILLER_13_194 ();
 sg13g2_fill_2 FILLER_13_203 ();
 sg13g2_fill_1 FILLER_13_218 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_decap_4 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_254 ();
 sg13g2_decap_4 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_4 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_48 ();
 sg13g2_fill_2 FILLER_14_57 ();
 sg13g2_fill_1 FILLER_14_59 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_decap_4 FILLER_14_88 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_decap_8 FILLER_14_106 ();
 sg13g2_decap_4 FILLER_14_113 ();
 sg13g2_decap_8 FILLER_14_143 ();
 sg13g2_decap_8 FILLER_14_150 ();
 sg13g2_fill_2 FILLER_14_157 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_2 FILLER_14_187 ();
 sg13g2_fill_1 FILLER_14_189 ();
 sg13g2_fill_1 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_4 FILLER_14_253 ();
 sg13g2_fill_2 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_4 FILLER_14_328 ();
 sg13g2_fill_1 FILLER_14_332 ();
 sg13g2_fill_2 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_136 ();
 sg13g2_decap_8 FILLER_15_143 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_decap_4 FILLER_15_176 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_decap_8 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_194 ();
 sg13g2_decap_8 FILLER_15_201 ();
 sg13g2_decap_4 FILLER_15_208 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_fill_2 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_decap_4 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_358 ();
 sg13g2_fill_1 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_41 ();
 sg13g2_fill_1 FILLER_16_50 ();
 sg13g2_fill_2 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_66 ();
 sg13g2_fill_2 FILLER_16_83 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_decap_8 FILLER_16_113 ();
 sg13g2_decap_8 FILLER_16_120 ();
 sg13g2_decap_8 FILLER_16_127 ();
 sg13g2_decap_8 FILLER_16_134 ();
 sg13g2_decap_4 FILLER_16_141 ();
 sg13g2_fill_2 FILLER_16_145 ();
 sg13g2_decap_4 FILLER_16_170 ();
 sg13g2_decap_4 FILLER_16_192 ();
 sg13g2_fill_2 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_209 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_247 ();
 sg13g2_fill_1 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_262 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_fill_2 FILLER_16_304 ();
 sg13g2_fill_1 FILLER_16_306 ();
 sg13g2_fill_1 FILLER_16_324 ();
 sg13g2_decap_4 FILLER_16_347 ();
 sg13g2_fill_2 FILLER_16_351 ();
 sg13g2_fill_2 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_fill_2 FILLER_17_75 ();
 sg13g2_fill_1 FILLER_17_96 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_225 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_fill_2 FILLER_17_294 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_decap_4 FILLER_18_73 ();
 sg13g2_fill_2 FILLER_18_92 ();
 sg13g2_fill_2 FILLER_18_115 ();
 sg13g2_decap_4 FILLER_18_139 ();
 sg13g2_fill_2 FILLER_18_143 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_fill_2 FILLER_18_168 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_189 ();
 sg13g2_fill_2 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_decap_4 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_2 FILLER_18_269 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_fill_2 FILLER_18_339 ();
 sg13g2_decap_4 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_47 ();
 sg13g2_fill_2 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_100 ();
 sg13g2_fill_2 FILLER_19_114 ();
 sg13g2_fill_1 FILLER_19_116 ();
 sg13g2_fill_1 FILLER_19_122 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_decap_4 FILLER_19_186 ();
 sg13g2_fill_2 FILLER_19_190 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_4 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_246 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_fill_2 FILLER_19_342 ();
 sg13g2_decap_4 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_fill_1 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_4 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_54 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_fill_2 FILLER_20_74 ();
 sg13g2_fill_2 FILLER_20_89 ();
 sg13g2_decap_8 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_108 ();
 sg13g2_decap_4 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_143 ();
 sg13g2_decap_8 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_157 ();
 sg13g2_decap_8 FILLER_20_164 ();
 sg13g2_decap_8 FILLER_20_176 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_decap_8 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_277 ();
 sg13g2_decap_4 FILLER_20_283 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_333 ();
 sg13g2_fill_1 FILLER_20_335 ();
 sg13g2_decap_4 FILLER_20_356 ();
 sg13g2_fill_2 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_374 ();
 sg13g2_decap_4 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_58 ();
 sg13g2_decap_4 FILLER_21_65 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_4 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_127 ();
 sg13g2_fill_2 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_136 ();
 sg13g2_decap_8 FILLER_21_141 ();
 sg13g2_decap_8 FILLER_21_148 ();
 sg13g2_decap_4 FILLER_21_155 ();
 sg13g2_fill_1 FILLER_21_159 ();
 sg13g2_fill_2 FILLER_21_173 ();
 sg13g2_decap_8 FILLER_21_192 ();
 sg13g2_decap_4 FILLER_21_199 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_decap_4 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_245 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_272 ();
 sg13g2_decap_8 FILLER_21_279 ();
 sg13g2_decap_4 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_fill_2 FILLER_21_323 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_decap_4 FILLER_21_352 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_2 FILLER_21_366 ();
 sg13g2_fill_2 FILLER_21_385 ();
 sg13g2_fill_1 FILLER_21_395 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_decap_8 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_57 ();
 sg13g2_fill_2 FILLER_22_72 ();
 sg13g2_fill_2 FILLER_22_79 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_125 ();
 sg13g2_fill_2 FILLER_22_152 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_189 ();
 sg13g2_fill_1 FILLER_22_199 ();
 sg13g2_decap_4 FILLER_22_204 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_281 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_309 ();
 sg13g2_fill_1 FILLER_22_311 ();
 sg13g2_decap_4 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_fill_1 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_decap_4 FILLER_23_37 ();
 sg13g2_fill_2 FILLER_23_41 ();
 sg13g2_decap_4 FILLER_23_56 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_fill_2 FILLER_23_94 ();
 sg13g2_fill_1 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_decap_4 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_fill_2 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_fill_2 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_4 FILLER_23_371 ();
 sg13g2_fill_2 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_decap_4 FILLER_24_44 ();
 sg13g2_fill_2 FILLER_24_48 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_107 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_4 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_142 ();
 sg13g2_decap_4 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_decap_4 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_decap_4 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_decap_4 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_decap_4 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_334 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_decap_4 FILLER_24_373 ();
 sg13g2_decap_4 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_391 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_18 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_1 FILLER_25_46 ();
 sg13g2_fill_2 FILLER_25_55 ();
 sg13g2_decap_4 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_93 ();
 sg13g2_fill_2 FILLER_25_103 ();
 sg13g2_fill_1 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_176 ();
 sg13g2_fill_2 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_234 ();
 sg13g2_decap_8 FILLER_25_241 ();
 sg13g2_decap_4 FILLER_25_248 ();
 sg13g2_fill_2 FILLER_25_288 ();
 sg13g2_decap_4 FILLER_25_316 ();
 sg13g2_fill_2 FILLER_25_333 ();
 sg13g2_fill_1 FILLER_25_376 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_45 ();
 sg13g2_decap_4 FILLER_26_53 ();
 sg13g2_fill_2 FILLER_26_57 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_76 ();
 sg13g2_fill_2 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_decap_4 FILLER_26_94 ();
 sg13g2_decap_8 FILLER_26_111 ();
 sg13g2_decap_4 FILLER_26_118 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_4 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_decap_4 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_decap_4 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_334 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_29 ();
 sg13g2_fill_2 FILLER_27_33 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_decap_8 FILLER_27_71 ();
 sg13g2_fill_1 FILLER_27_78 ();
 sg13g2_decap_8 FILLER_27_87 ();
 sg13g2_fill_2 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_decap_4 FILLER_27_134 ();
 sg13g2_decap_8 FILLER_27_146 ();
 sg13g2_decap_8 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_160 ();
 sg13g2_decap_8 FILLER_27_167 ();
 sg13g2_decap_4 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_261 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_4 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_4 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_391 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_33 ();
 sg13g2_decap_4 FILLER_28_40 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_111 ();
 sg13g2_fill_1 FILLER_28_120 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_4 FILLER_28_229 ();
 sg13g2_decap_8 FILLER_28_283 ();
 sg13g2_decap_4 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_4 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_decap_4 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_fill_2 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_43 ();
 sg13g2_fill_1 FILLER_29_66 ();
 sg13g2_decap_4 FILLER_29_71 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_fill_2 FILLER_29_122 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_decap_4 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_208 ();
 sg13g2_decap_4 FILLER_29_226 ();
 sg13g2_fill_2 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_decap_4 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_decap_4 FILLER_29_290 ();
 sg13g2_decap_4 FILLER_29_320 ();
 sg13g2_decap_4 FILLER_29_363 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_16 ();
 sg13g2_fill_2 FILLER_30_30 ();
 sg13g2_fill_1 FILLER_30_32 ();
 sg13g2_fill_1 FILLER_30_53 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_4 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_156 ();
 sg13g2_decap_4 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_185 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_215 ();
 sg13g2_decap_4 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_decap_8 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_fill_2 FILLER_30_363 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_9 ();
 sg13g2_fill_1 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_40 ();
 sg13g2_fill_1 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_64 ();
 sg13g2_fill_2 FILLER_31_68 ();
 sg13g2_fill_2 FILLER_31_83 ();
 sg13g2_decap_8 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_181 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_fill_2 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_234 ();
 sg13g2_fill_1 FILLER_31_241 ();
 sg13g2_fill_2 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_decap_8 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_4 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_decap_4 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_decap_4 FILLER_31_373 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_43 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_2 FILLER_32_55 ();
 sg13g2_decap_8 FILLER_32_76 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_160 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_255 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_393 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_18 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_decap_4 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_decap_8 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_fill_2 FILLER_33_100 ();
 sg13g2_fill_1 FILLER_33_102 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_fill_1 FILLER_33_120 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_decap_4 FILLER_33_161 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_decap_4 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_217 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_decap_4 FILLER_33_229 ();
 sg13g2_fill_2 FILLER_33_233 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_23 ();
 sg13g2_decap_4 FILLER_34_43 ();
 sg13g2_decap_4 FILLER_34_60 ();
 sg13g2_fill_2 FILLER_34_64 ();
 sg13g2_decap_4 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_decap_4 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_fill_2 FILLER_34_211 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_246 ();
 sg13g2_decap_4 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_262 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_fill_2 FILLER_34_299 ();
 sg13g2_decap_8 FILLER_34_316 ();
 sg13g2_decap_4 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_decap_4 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_23 ();
 sg13g2_fill_1 FILLER_35_25 ();
 sg13g2_decap_4 FILLER_35_36 ();
 sg13g2_fill_1 FILLER_35_40 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_51 ();
 sg13g2_decap_8 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_92 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_decap_8 FILLER_35_104 ();
 sg13g2_decap_8 FILLER_35_111 ();
 sg13g2_decap_4 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_122 ();
 sg13g2_fill_1 FILLER_35_128 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_decap_4 FILLER_35_191 ();
 sg13g2_decap_4 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_257 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_341 ();
 sg13g2_decap_8 FILLER_35_348 ();
 sg13g2_decap_8 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_decap_8 FILLER_35_369 ();
 sg13g2_decap_4 FILLER_35_376 ();
 sg13g2_fill_1 FILLER_35_380 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_decap_4 FILLER_36_13 ();
 sg13g2_fill_1 FILLER_36_17 ();
 sg13g2_fill_2 FILLER_36_48 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_decap_4 FILLER_36_82 ();
 sg13g2_fill_2 FILLER_36_97 ();
 sg13g2_fill_1 FILLER_36_99 ();
 sg13g2_decap_8 FILLER_36_115 ();
 sg13g2_fill_1 FILLER_36_122 ();
 sg13g2_fill_2 FILLER_36_143 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_fill_1 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_279 ();
 sg13g2_decap_8 FILLER_36_286 ();
 sg13g2_decap_8 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_decap_4 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_decap_4 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_356 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_fill_1 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_4 FILLER_36_391 ();
 sg13g2_fill_1 FILLER_36_395 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_fill_1 FILLER_37_17 ();
 sg13g2_decap_8 FILLER_37_26 ();
 sg13g2_decap_8 FILLER_37_33 ();
 sg13g2_fill_1 FILLER_37_40 ();
 sg13g2_decap_8 FILLER_37_44 ();
 sg13g2_decap_8 FILLER_37_51 ();
 sg13g2_fill_2 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_66 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_decap_8 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_296 ();
 sg13g2_decap_8 FILLER_37_306 ();
 sg13g2_decap_8 FILLER_37_313 ();
 sg13g2_decap_4 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_324 ();
 sg13g2_decap_4 FILLER_37_329 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_53 ();
 sg13g2_fill_2 FILLER_38_72 ();
 sg13g2_decap_8 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_2 FILLER_38_144 ();
 sg13g2_fill_1 FILLER_38_146 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_170 ();
 sg13g2_decap_4 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_decap_8 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_fill_2 FILLER_38_233 ();
 sg13g2_fill_1 FILLER_38_235 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_decap_4 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_323 ();
 sg13g2_fill_2 FILLER_38_353 ();
 sg13g2_fill_2 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_1 FILLER_39_16 ();
 sg13g2_fill_2 FILLER_39_49 ();
 sg13g2_fill_1 FILLER_39_51 ();
 sg13g2_fill_2 FILLER_39_77 ();
 sg13g2_fill_1 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_4 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_116 ();
 sg13g2_fill_2 FILLER_39_130 ();
 sg13g2_fill_2 FILLER_39_148 ();
 sg13g2_fill_1 FILLER_39_150 ();
 sg13g2_fill_1 FILLER_39_156 ();
 sg13g2_decap_8 FILLER_39_174 ();
 sg13g2_decap_8 FILLER_39_181 ();
 sg13g2_fill_1 FILLER_39_188 ();
 sg13g2_fill_2 FILLER_39_213 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_313 ();
 sg13g2_fill_1 FILLER_39_315 ();
 sg13g2_fill_2 FILLER_39_356 ();
 sg13g2_fill_1 FILLER_39_371 ();
 sg13g2_fill_2 FILLER_39_376 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_65 ();
 sg13g2_decap_8 FILLER_40_72 ();
 sg13g2_decap_8 FILLER_40_79 ();
 sg13g2_fill_1 FILLER_40_86 ();
 sg13g2_fill_1 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_decap_4 FILLER_40_200 ();
 sg13g2_fill_1 FILLER_40_231 ();
 sg13g2_fill_1 FILLER_40_249 ();
 sg13g2_decap_8 FILLER_40_269 ();
 sg13g2_decap_4 FILLER_40_276 ();
 sg13g2_fill_2 FILLER_40_280 ();
 sg13g2_fill_2 FILLER_40_287 ();
 sg13g2_fill_1 FILLER_40_289 ();
 sg13g2_fill_1 FILLER_40_321 ();
 sg13g2_decap_8 FILLER_40_340 ();
 sg13g2_decap_4 FILLER_40_347 ();
 sg13g2_fill_2 FILLER_40_351 ();
 sg13g2_fill_2 FILLER_40_357 ();
 sg13g2_fill_1 FILLER_40_359 ();
 sg13g2_decap_8 FILLER_40_368 ();
 sg13g2_decap_4 FILLER_40_375 ();
 sg13g2_fill_1 FILLER_40_379 ();
 sg13g2_fill_1 FILLER_40_388 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_2 ();
 sg13g2_fill_2 FILLER_41_16 ();
 sg13g2_decap_8 FILLER_41_31 ();
 sg13g2_decap_8 FILLER_41_46 ();
 sg13g2_decap_4 FILLER_41_53 ();
 sg13g2_fill_1 FILLER_41_57 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_fill_2 FILLER_41_77 ();
 sg13g2_fill_1 FILLER_41_79 ();
 sg13g2_decap_8 FILLER_41_110 ();
 sg13g2_fill_2 FILLER_41_117 ();
 sg13g2_fill_1 FILLER_41_127 ();
 sg13g2_decap_8 FILLER_41_145 ();
 sg13g2_decap_4 FILLER_41_152 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_decap_4 FILLER_41_162 ();
 sg13g2_fill_1 FILLER_41_166 ();
 sg13g2_decap_8 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_fill_2 FILLER_41_195 ();
 sg13g2_fill_1 FILLER_41_206 ();
 sg13g2_decap_4 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_219 ();
 sg13g2_fill_2 FILLER_41_234 ();
 sg13g2_fill_2 FILLER_41_244 ();
 sg13g2_fill_1 FILLER_41_258 ();
 sg13g2_decap_8 FILLER_41_271 ();
 sg13g2_decap_8 FILLER_41_278 ();
 sg13g2_decap_8 FILLER_41_285 ();
 sg13g2_decap_8 FILLER_41_292 ();
 sg13g2_fill_2 FILLER_41_299 ();
 sg13g2_decap_8 FILLER_41_305 ();
 sg13g2_decap_8 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_319 ();
 sg13g2_fill_1 FILLER_41_321 ();
 sg13g2_decap_8 FILLER_41_346 ();
 sg13g2_fill_2 FILLER_41_353 ();
 sg13g2_fill_1 FILLER_41_355 ();
 sg13g2_fill_2 FILLER_41_387 ();
 sg13g2_fill_1 FILLER_41_389 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_4 ();
 sg13g2_decap_8 FILLER_42_25 ();
 sg13g2_decap_8 FILLER_42_32 ();
 sg13g2_fill_2 FILLER_42_39 ();
 sg13g2_fill_2 FILLER_42_46 ();
 sg13g2_fill_1 FILLER_42_60 ();
 sg13g2_decap_4 FILLER_42_73 ();
 sg13g2_fill_1 FILLER_42_77 ();
 sg13g2_fill_2 FILLER_42_82 ();
 sg13g2_fill_2 FILLER_42_110 ();
 sg13g2_decap_8 FILLER_42_138 ();
 sg13g2_fill_1 FILLER_42_145 ();
 sg13g2_fill_2 FILLER_42_171 ();
 sg13g2_decap_4 FILLER_42_199 ();
 sg13g2_decap_8 FILLER_42_212 ();
 sg13g2_fill_2 FILLER_42_219 ();
 sg13g2_decap_4 FILLER_42_234 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_decap_4 FILLER_42_272 ();
 sg13g2_fill_2 FILLER_42_285 ();
 sg13g2_decap_8 FILLER_42_292 ();
 sg13g2_decap_8 FILLER_42_299 ();
 sg13g2_fill_2 FILLER_42_306 ();
 sg13g2_decap_8 FILLER_42_312 ();
 sg13g2_decap_8 FILLER_42_319 ();
 sg13g2_decap_8 FILLER_42_326 ();
 sg13g2_decap_8 FILLER_42_333 ();
 sg13g2_decap_4 FILLER_42_340 ();
 sg13g2_fill_2 FILLER_42_357 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_9 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_37 ();
 sg13g2_fill_2 FILLER_43_44 ();
 sg13g2_fill_1 FILLER_43_56 ();
 sg13g2_fill_2 FILLER_43_62 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_decap_4 FILLER_43_107 ();
 sg13g2_fill_2 FILLER_43_111 ();
 sg13g2_decap_8 FILLER_43_127 ();
 sg13g2_fill_1 FILLER_43_134 ();
 sg13g2_fill_2 FILLER_43_144 ();
 sg13g2_fill_1 FILLER_43_181 ();
 sg13g2_fill_2 FILLER_43_207 ();
 sg13g2_decap_8 FILLER_43_214 ();
 sg13g2_fill_2 FILLER_43_221 ();
 sg13g2_fill_1 FILLER_43_223 ();
 sg13g2_decap_8 FILLER_43_228 ();
 sg13g2_decap_8 FILLER_43_235 ();
 sg13g2_fill_1 FILLER_43_250 ();
 sg13g2_decap_4 FILLER_43_257 ();
 sg13g2_fill_2 FILLER_43_261 ();
 sg13g2_fill_2 FILLER_43_276 ();
 sg13g2_fill_2 FILLER_43_295 ();
 sg13g2_fill_2 FILLER_43_331 ();
 sg13g2_fill_1 FILLER_43_333 ();
 sg13g2_decap_4 FILLER_43_338 ();
 sg13g2_fill_1 FILLER_43_342 ();
 sg13g2_fill_2 FILLER_43_372 ();
 sg13g2_fill_1 FILLER_43_374 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_fill_2 FILLER_44_21 ();
 sg13g2_fill_1 FILLER_44_23 ();
 sg13g2_fill_1 FILLER_44_37 ();
 sg13g2_fill_2 FILLER_44_51 ();
 sg13g2_fill_2 FILLER_44_70 ();
 sg13g2_fill_1 FILLER_44_78 ();
 sg13g2_decap_8 FILLER_44_88 ();
 sg13g2_fill_2 FILLER_44_147 ();
 sg13g2_fill_1 FILLER_44_149 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_fill_1 FILLER_44_226 ();
 sg13g2_fill_2 FILLER_44_248 ();
 sg13g2_fill_2 FILLER_44_276 ();
 sg13g2_fill_2 FILLER_44_286 ();
 sg13g2_fill_2 FILLER_44_296 ();
 sg13g2_fill_1 FILLER_44_298 ();
 sg13g2_decap_4 FILLER_44_376 ();
 sg13g2_fill_2 FILLER_44_380 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_fill_2 FILLER_45_21 ();
 sg13g2_fill_2 FILLER_45_48 ();
 sg13g2_fill_2 FILLER_45_59 ();
 sg13g2_decap_4 FILLER_45_73 ();
 sg13g2_decap_8 FILLER_45_81 ();
 sg13g2_decap_4 FILLER_45_88 ();
 sg13g2_fill_2 FILLER_45_92 ();
 sg13g2_decap_8 FILLER_45_124 ();
 sg13g2_decap_4 FILLER_45_131 ();
 sg13g2_fill_2 FILLER_45_135 ();
 sg13g2_decap_8 FILLER_45_145 ();
 sg13g2_fill_2 FILLER_45_152 ();
 sg13g2_fill_1 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_203 ();
 sg13g2_fill_1 FILLER_45_205 ();
 sg13g2_fill_1 FILLER_45_238 ();
 sg13g2_decap_4 FILLER_45_318 ();
 sg13g2_fill_1 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_331 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_356 ();
 sg13g2_decap_8 FILLER_45_384 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_20 ();
 sg13g2_fill_2 FILLER_46_27 ();
 sg13g2_fill_1 FILLER_46_29 ();
 sg13g2_decap_8 FILLER_46_48 ();
 sg13g2_decap_4 FILLER_46_55 ();
 sg13g2_fill_1 FILLER_46_59 ();
 sg13g2_decap_4 FILLER_46_76 ();
 sg13g2_fill_2 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_142 ();
 sg13g2_decap_8 FILLER_46_173 ();
 sg13g2_decap_8 FILLER_46_180 ();
 sg13g2_fill_1 FILLER_46_187 ();
 sg13g2_decap_4 FILLER_46_196 ();
 sg13g2_fill_1 FILLER_46_200 ();
 sg13g2_fill_1 FILLER_46_267 ();
 sg13g2_fill_1 FILLER_46_273 ();
 sg13g2_fill_2 FILLER_46_284 ();
 sg13g2_fill_2 FILLER_46_302 ();
 sg13g2_decap_4 FILLER_46_309 ();
 sg13g2_fill_1 FILLER_46_313 ();
 sg13g2_decap_8 FILLER_46_353 ();
 sg13g2_decap_8 FILLER_46_360 ();
 sg13g2_fill_2 FILLER_46_380 ();
 sg13g2_fill_1 FILLER_46_382 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_35 ();
 sg13g2_fill_2 FILLER_47_43 ();
 sg13g2_fill_1 FILLER_47_45 ();
 sg13g2_decap_8 FILLER_47_51 ();
 sg13g2_decap_8 FILLER_47_58 ();
 sg13g2_decap_4 FILLER_47_73 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_fill_2 FILLER_47_95 ();
 sg13g2_fill_1 FILLER_47_97 ();
 sg13g2_fill_2 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_234 ();
 sg13g2_decap_8 FILLER_47_267 ();
 sg13g2_fill_2 FILLER_47_274 ();
 sg13g2_fill_1 FILLER_47_276 ();
 sg13g2_fill_2 FILLER_47_281 ();
 sg13g2_fill_1 FILLER_47_283 ();
 sg13g2_fill_2 FILLER_47_288 ();
 sg13g2_fill_1 FILLER_47_290 ();
 sg13g2_decap_4 FILLER_47_318 ();
 sg13g2_decap_4 FILLER_47_327 ();
 sg13g2_fill_1 FILLER_47_387 ();
 sg13g2_fill_2 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_24 ();
 sg13g2_fill_2 FILLER_48_32 ();
 sg13g2_fill_2 FILLER_48_42 ();
 sg13g2_fill_1 FILLER_48_44 ();
 sg13g2_fill_2 FILLER_48_58 ();
 sg13g2_fill_1 FILLER_48_110 ();
 sg13g2_fill_1 FILLER_48_139 ();
 sg13g2_decap_8 FILLER_48_174 ();
 sg13g2_fill_2 FILLER_48_181 ();
 sg13g2_fill_1 FILLER_48_183 ();
 sg13g2_fill_2 FILLER_48_192 ();
 sg13g2_fill_1 FILLER_48_194 ();
 sg13g2_decap_4 FILLER_48_256 ();
 sg13g2_decap_4 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_282 ();
 sg13g2_decap_4 FILLER_48_289 ();
 sg13g2_fill_1 FILLER_48_293 ();
 sg13g2_fill_2 FILLER_48_322 ();
 sg13g2_fill_2 FILLER_48_359 ();
 sg13g2_fill_1 FILLER_48_361 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_9 ();
 sg13g2_fill_1 FILLER_49_23 ();
 sg13g2_decap_4 FILLER_49_82 ();
 sg13g2_fill_1 FILLER_49_86 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_4 FILLER_49_98 ();
 sg13g2_fill_1 FILLER_49_124 ();
 sg13g2_fill_1 FILLER_49_166 ();
 sg13g2_decap_8 FILLER_49_184 ();
 sg13g2_decap_8 FILLER_49_191 ();
 sg13g2_decap_8 FILLER_49_198 ();
 sg13g2_fill_1 FILLER_49_209 ();
 sg13g2_decap_8 FILLER_49_219 ();
 sg13g2_decap_4 FILLER_49_226 ();
 sg13g2_decap_4 FILLER_49_233 ();
 sg13g2_fill_2 FILLER_49_241 ();
 sg13g2_fill_1 FILLER_49_243 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_fill_2 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_fill_2 FILLER_49_304 ();
 sg13g2_fill_1 FILLER_49_306 ();
 sg13g2_fill_2 FILLER_49_319 ();
 sg13g2_fill_2 FILLER_49_344 ();
 sg13g2_decap_8 FILLER_49_362 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_fill_2 FILLER_49_389 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_23 ();
 sg13g2_fill_2 FILLER_50_48 ();
 sg13g2_fill_2 FILLER_50_58 ();
 sg13g2_fill_1 FILLER_50_60 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_84 ();
 sg13g2_fill_1 FILLER_50_86 ();
 sg13g2_fill_1 FILLER_50_136 ();
 sg13g2_fill_2 FILLER_50_156 ();
 sg13g2_fill_1 FILLER_50_192 ();
 sg13g2_decap_8 FILLER_50_197 ();
 sg13g2_decap_8 FILLER_50_204 ();
 sg13g2_decap_4 FILLER_50_211 ();
 sg13g2_fill_2 FILLER_50_215 ();
 sg13g2_fill_2 FILLER_50_241 ();
 sg13g2_fill_1 FILLER_50_243 ();
 sg13g2_decap_4 FILLER_50_252 ();
 sg13g2_fill_1 FILLER_50_256 ();
 sg13g2_decap_8 FILLER_50_277 ();
 sg13g2_fill_2 FILLER_50_284 ();
 sg13g2_decap_8 FILLER_50_299 ();
 sg13g2_decap_8 FILLER_50_306 ();
 sg13g2_decap_4 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_decap_4 FILLER_50_349 ();
 sg13g2_fill_1 FILLER_50_353 ();
 sg13g2_fill_2 FILLER_50_358 ();
 sg13g2_fill_1 FILLER_50_360 ();
 sg13g2_fill_2 FILLER_50_386 ();
 sg13g2_fill_1 FILLER_50_388 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_31 ();
 sg13g2_decap_4 FILLER_51_38 ();
 sg13g2_decap_4 FILLER_51_47 ();
 sg13g2_fill_1 FILLER_51_51 ();
 sg13g2_fill_1 FILLER_51_56 ();
 sg13g2_fill_2 FILLER_51_65 ();
 sg13g2_fill_2 FILLER_51_101 ();
 sg13g2_decap_8 FILLER_51_107 ();
 sg13g2_fill_1 FILLER_51_114 ();
 sg13g2_decap_8 FILLER_51_212 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_fill_1 FILLER_51_240 ();
 sg13g2_decap_4 FILLER_51_249 ();
 sg13g2_decap_4 FILLER_51_260 ();
 sg13g2_fill_2 FILLER_51_264 ();
 sg13g2_fill_2 FILLER_51_271 ();
 sg13g2_fill_1 FILLER_51_285 ();
 sg13g2_decap_8 FILLER_51_304 ();
 sg13g2_decap_8 FILLER_51_311 ();
 sg13g2_fill_2 FILLER_51_318 ();
 sg13g2_fill_2 FILLER_51_332 ();
 sg13g2_fill_1 FILLER_51_334 ();
 sg13g2_decap_8 FILLER_51_339 ();
 sg13g2_fill_2 FILLER_51_372 ();
 sg13g2_fill_2 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_4 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_4 ();
 sg13g2_fill_2 FILLER_52_13 ();
 sg13g2_decap_8 FILLER_52_38 ();
 sg13g2_decap_8 FILLER_52_45 ();
 sg13g2_decap_8 FILLER_52_52 ();
 sg13g2_decap_8 FILLER_52_59 ();
 sg13g2_decap_8 FILLER_52_66 ();
 sg13g2_decap_4 FILLER_52_80 ();
 sg13g2_fill_2 FILLER_52_84 ();
 sg13g2_decap_4 FILLER_52_90 ();
 sg13g2_fill_1 FILLER_52_101 ();
 sg13g2_fill_2 FILLER_52_106 ();
 sg13g2_fill_2 FILLER_52_132 ();
 sg13g2_fill_2 FILLER_52_201 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_fill_1 FILLER_52_230 ();
 sg13g2_fill_1 FILLER_52_261 ();
 sg13g2_fill_1 FILLER_52_298 ();
 sg13g2_fill_2 FILLER_52_307 ();
 sg13g2_fill_1 FILLER_52_309 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_decap_4 FILLER_52_349 ();
 sg13g2_fill_2 FILLER_52_353 ();
 sg13g2_fill_1 FILLER_52_368 ();
 sg13g2_fill_2 FILLER_52_384 ();
 sg13g2_fill_1 FILLER_52_386 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_4 ();
 sg13g2_decap_8 FILLER_53_13 ();
 sg13g2_decap_4 FILLER_53_20 ();
 sg13g2_fill_1 FILLER_53_24 ();
 sg13g2_decap_4 FILLER_53_38 ();
 sg13g2_fill_2 FILLER_53_47 ();
 sg13g2_decap_8 FILLER_53_53 ();
 sg13g2_decap_8 FILLER_53_60 ();
 sg13g2_decap_4 FILLER_53_87 ();
 sg13g2_fill_1 FILLER_53_130 ();
 sg13g2_fill_1 FILLER_53_140 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_2 FILLER_53_243 ();
 sg13g2_fill_2 FILLER_53_288 ();
 sg13g2_fill_1 FILLER_53_290 ();
 sg13g2_decap_8 FILLER_53_325 ();
 sg13g2_fill_2 FILLER_53_332 ();
 sg13g2_fill_1 FILLER_53_334 ();
 sg13g2_decap_8 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_366 ();
 sg13g2_fill_1 FILLER_53_373 ();
 sg13g2_decap_4 FILLER_53_379 ();
 sg13g2_decap_8 FILLER_53_400 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_4 ();
 sg13g2_fill_2 FILLER_54_17 ();
 sg13g2_decap_4 FILLER_54_27 ();
 sg13g2_fill_2 FILLER_54_60 ();
 sg13g2_fill_1 FILLER_54_62 ();
 sg13g2_fill_1 FILLER_54_71 ();
 sg13g2_decap_4 FILLER_54_98 ();
 sg13g2_fill_1 FILLER_54_143 ();
 sg13g2_fill_2 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_221 ();
 sg13g2_fill_2 FILLER_54_233 ();
 sg13g2_fill_1 FILLER_54_235 ();
 sg13g2_fill_1 FILLER_54_258 ();
 sg13g2_fill_2 FILLER_54_293 ();
 sg13g2_decap_8 FILLER_54_300 ();
 sg13g2_fill_2 FILLER_54_307 ();
 sg13g2_fill_1 FILLER_54_313 ();
 sg13g2_decap_8 FILLER_54_329 ();
 sg13g2_decap_8 FILLER_54_336 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_decap_4 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_fill_2 FILLER_54_392 ();
 sg13g2_fill_1 FILLER_54_394 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_fill_2 FILLER_55_48 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_fill_2 FILLER_55_80 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_fill_2 FILLER_55_190 ();
 sg13g2_fill_2 FILLER_55_201 ();
 sg13g2_fill_1 FILLER_55_203 ();
 sg13g2_decap_4 FILLER_55_208 ();
 sg13g2_fill_1 FILLER_55_212 ();
 sg13g2_decap_4 FILLER_55_221 ();
 sg13g2_fill_2 FILLER_55_225 ();
 sg13g2_decap_8 FILLER_55_236 ();
 sg13g2_fill_2 FILLER_55_243 ();
 sg13g2_fill_1 FILLER_55_245 ();
 sg13g2_fill_2 FILLER_55_254 ();
 sg13g2_decap_8 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_288 ();
 sg13g2_decap_8 FILLER_55_293 ();
 sg13g2_decap_8 FILLER_55_300 ();
 sg13g2_decap_8 FILLER_55_307 ();
 sg13g2_fill_1 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_320 ();
 sg13g2_fill_2 FILLER_55_337 ();
 sg13g2_decap_8 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_368 ();
 sg13g2_decap_8 FILLER_55_374 ();
 sg13g2_decap_8 FILLER_55_381 ();
 sg13g2_fill_2 FILLER_55_388 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_31 ();
 sg13g2_decap_4 FILLER_56_38 ();
 sg13g2_fill_1 FILLER_56_42 ();
 sg13g2_fill_2 FILLER_56_51 ();
 sg13g2_fill_1 FILLER_56_53 ();
 sg13g2_decap_4 FILLER_56_73 ();
 sg13g2_fill_2 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_114 ();
 sg13g2_fill_2 FILLER_56_169 ();
 sg13g2_fill_1 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_208 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_241 ();
 sg13g2_decap_4 FILLER_56_248 ();
 sg13g2_fill_2 FILLER_56_252 ();
 sg13g2_decap_4 FILLER_56_258 ();
 sg13g2_fill_2 FILLER_56_266 ();
 sg13g2_decap_8 FILLER_56_272 ();
 sg13g2_decap_8 FILLER_56_279 ();
 sg13g2_fill_1 FILLER_56_295 ();
 sg13g2_fill_2 FILLER_56_323 ();
 sg13g2_fill_1 FILLER_56_352 ();
 sg13g2_fill_2 FILLER_56_365 ();
 sg13g2_fill_1 FILLER_56_367 ();
 sg13g2_decap_4 FILLER_56_380 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_2 FILLER_57_35 ();
 sg13g2_fill_2 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_68 ();
 sg13g2_decap_8 FILLER_57_75 ();
 sg13g2_decap_8 FILLER_57_82 ();
 sg13g2_fill_2 FILLER_57_89 ();
 sg13g2_fill_1 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_140 ();
 sg13g2_fill_2 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_198 ();
 sg13g2_fill_1 FILLER_57_200 ();
 sg13g2_fill_1 FILLER_57_215 ();
 sg13g2_fill_2 FILLER_57_230 ();
 sg13g2_decap_4 FILLER_57_258 ();
 sg13g2_fill_2 FILLER_57_280 ();
 sg13g2_fill_1 FILLER_57_282 ();
 sg13g2_fill_2 FILLER_57_288 ();
 sg13g2_fill_1 FILLER_57_290 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_fill_2 FILLER_57_347 ();
 sg13g2_fill_2 FILLER_57_388 ();
 sg13g2_fill_1 FILLER_57_390 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_24 ();
 sg13g2_fill_2 FILLER_58_64 ();
 sg13g2_decap_4 FILLER_58_74 ();
 sg13g2_fill_1 FILLER_58_78 ();
 sg13g2_fill_1 FILLER_58_113 ();
 sg13g2_fill_1 FILLER_58_141 ();
 sg13g2_fill_2 FILLER_58_156 ();
 sg13g2_fill_1 FILLER_58_158 ();
 sg13g2_fill_2 FILLER_58_174 ();
 sg13g2_fill_1 FILLER_58_176 ();
 sg13g2_decap_4 FILLER_58_238 ();
 sg13g2_fill_1 FILLER_58_242 ();
 sg13g2_decap_8 FILLER_58_247 ();
 sg13g2_fill_1 FILLER_58_306 ();
 sg13g2_fill_1 FILLER_58_345 ();
 sg13g2_fill_2 FILLER_58_361 ();
 sg13g2_decap_4 FILLER_58_405 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_11 ();
 sg13g2_decap_4 FILLER_59_16 ();
 sg13g2_fill_2 FILLER_59_20 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_4 FILLER_59_49 ();
 sg13g2_fill_1 FILLER_59_53 ();
 sg13g2_fill_1 FILLER_59_59 ();
 sg13g2_fill_2 FILLER_59_68 ();
 sg13g2_fill_1 FILLER_59_70 ();
 sg13g2_fill_1 FILLER_59_132 ();
 sg13g2_fill_2 FILLER_59_171 ();
 sg13g2_fill_1 FILLER_59_178 ();
 sg13g2_fill_1 FILLER_59_192 ();
 sg13g2_fill_2 FILLER_59_202 ();
 sg13g2_fill_1 FILLER_59_204 ();
 sg13g2_fill_1 FILLER_59_219 ();
 sg13g2_decap_8 FILLER_59_246 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_fill_1 FILLER_59_260 ();
 sg13g2_fill_2 FILLER_59_307 ();
 sg13g2_fill_1 FILLER_59_309 ();
 sg13g2_decap_8 FILLER_59_315 ();
 sg13g2_decap_8 FILLER_59_322 ();
 sg13g2_decap_4 FILLER_59_329 ();
 sg13g2_fill_1 FILLER_59_333 ();
 sg13g2_decap_8 FILLER_59_339 ();
 sg13g2_decap_4 FILLER_59_346 ();
 sg13g2_fill_2 FILLER_59_350 ();
 sg13g2_fill_1 FILLER_59_380 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_56 ();
 sg13g2_fill_1 FILLER_60_60 ();
 sg13g2_fill_2 FILLER_60_87 ();
 sg13g2_fill_2 FILLER_60_93 ();
 sg13g2_fill_1 FILLER_60_108 ();
 sg13g2_fill_2 FILLER_60_123 ();
 sg13g2_fill_2 FILLER_60_155 ();
 sg13g2_fill_1 FILLER_60_157 ();
 sg13g2_fill_1 FILLER_60_233 ();
 sg13g2_decap_8 FILLER_60_260 ();
 sg13g2_decap_8 FILLER_60_267 ();
 sg13g2_decap_8 FILLER_60_274 ();
 sg13g2_decap_4 FILLER_60_281 ();
 sg13g2_fill_2 FILLER_60_285 ();
 sg13g2_decap_4 FILLER_60_305 ();
 sg13g2_fill_2 FILLER_60_309 ();
 sg13g2_decap_8 FILLER_60_314 ();
 sg13g2_decap_4 FILLER_60_325 ();
 sg13g2_fill_2 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_339 ();
 sg13g2_decap_8 FILLER_60_351 ();
 sg13g2_decap_8 FILLER_60_358 ();
 sg13g2_decap_8 FILLER_60_365 ();
 sg13g2_decap_4 FILLER_60_372 ();
 sg13g2_fill_2 FILLER_60_376 ();
 sg13g2_fill_1 FILLER_60_388 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_14 ();
 sg13g2_decap_4 FILLER_61_21 ();
 sg13g2_fill_1 FILLER_61_25 ();
 sg13g2_decap_4 FILLER_61_60 ();
 sg13g2_fill_2 FILLER_61_64 ();
 sg13g2_fill_2 FILLER_61_74 ();
 sg13g2_fill_2 FILLER_61_80 ();
 sg13g2_decap_8 FILLER_61_86 ();
 sg13g2_fill_1 FILLER_61_93 ();
 sg13g2_fill_1 FILLER_61_124 ();
 sg13g2_fill_2 FILLER_61_143 ();
 sg13g2_fill_1 FILLER_61_145 ();
 sg13g2_fill_2 FILLER_61_173 ();
 sg13g2_fill_2 FILLER_61_235 ();
 sg13g2_decap_8 FILLER_61_258 ();
 sg13g2_decap_8 FILLER_61_265 ();
 sg13g2_decap_8 FILLER_61_272 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_decap_8 FILLER_61_294 ();
 sg13g2_fill_1 FILLER_61_301 ();
 sg13g2_fill_1 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_334 ();
 sg13g2_fill_1 FILLER_61_362 ();
 sg13g2_fill_2 FILLER_61_368 ();
 sg13g2_decap_4 FILLER_61_374 ();
 sg13g2_fill_2 FILLER_61_378 ();
 sg13g2_decap_4 FILLER_61_388 ();
 sg13g2_fill_2 FILLER_61_392 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_fill_1 FILLER_62_31 ();
 sg13g2_fill_1 FILLER_62_41 ();
 sg13g2_fill_2 FILLER_62_47 ();
 sg13g2_fill_1 FILLER_62_49 ();
 sg13g2_fill_2 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_65 ();
 sg13g2_decap_8 FILLER_62_71 ();
 sg13g2_decap_8 FILLER_62_78 ();
 sg13g2_fill_1 FILLER_62_85 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_fill_2 FILLER_62_153 ();
 sg13g2_fill_1 FILLER_62_169 ();
 sg13g2_fill_1 FILLER_62_175 ();
 sg13g2_fill_1 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_226 ();
 sg13g2_decap_4 FILLER_62_262 ();
 sg13g2_fill_2 FILLER_62_266 ();
 sg13g2_decap_4 FILLER_62_405 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_31 ();
 sg13g2_decap_4 FILLER_63_43 ();
 sg13g2_fill_2 FILLER_63_69 ();
 sg13g2_fill_1 FILLER_63_71 ();
 sg13g2_fill_1 FILLER_63_98 ();
 sg13g2_fill_2 FILLER_63_114 ();
 sg13g2_fill_1 FILLER_63_208 ();
 sg13g2_fill_2 FILLER_63_227 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_fill_1 FILLER_63_304 ();
 sg13g2_fill_2 FILLER_63_341 ();
 sg13g2_fill_1 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_369 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_decap_4 FILLER_63_390 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_24 ();
 sg13g2_fill_2 FILLER_64_31 ();
 sg13g2_decap_4 FILLER_64_54 ();
 sg13g2_decap_4 FILLER_64_63 ();
 sg13g2_fill_1 FILLER_64_67 ();
 sg13g2_fill_1 FILLER_64_121 ();
 sg13g2_fill_1 FILLER_64_126 ();
 sg13g2_fill_2 FILLER_64_143 ();
 sg13g2_fill_1 FILLER_64_145 ();
 sg13g2_fill_2 FILLER_64_191 ();
 sg13g2_fill_2 FILLER_64_202 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_263 ();
 sg13g2_decap_8 FILLER_64_290 ();
 sg13g2_decap_4 FILLER_64_297 ();
 sg13g2_decap_8 FILLER_64_304 ();
 sg13g2_decap_8 FILLER_64_311 ();
 sg13g2_fill_2 FILLER_64_318 ();
 sg13g2_fill_1 FILLER_64_320 ();
 sg13g2_decap_8 FILLER_64_325 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_fill_2 FILLER_64_347 ();
 sg13g2_decap_8 FILLER_64_352 ();
 sg13g2_decap_8 FILLER_64_359 ();
 sg13g2_decap_8 FILLER_64_366 ();
 sg13g2_decap_8 FILLER_64_373 ();
 sg13g2_decap_4 FILLER_64_380 ();
 sg13g2_fill_1 FILLER_64_384 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_23 ();
 sg13g2_decap_4 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_32 ();
 sg13g2_fill_2 FILLER_65_54 ();
 sg13g2_fill_2 FILLER_65_64 ();
 sg13g2_fill_1 FILLER_65_66 ();
 sg13g2_fill_2 FILLER_65_87 ();
 sg13g2_fill_1 FILLER_65_103 ();
 sg13g2_fill_2 FILLER_65_142 ();
 sg13g2_fill_1 FILLER_65_144 ();
 sg13g2_fill_2 FILLER_65_189 ();
 sg13g2_fill_1 FILLER_65_191 ();
 sg13g2_fill_2 FILLER_65_201 ();
 sg13g2_fill_1 FILLER_65_203 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_decap_4 FILLER_65_222 ();
 sg13g2_decap_4 FILLER_65_239 ();
 sg13g2_fill_1 FILLER_65_243 ();
 sg13g2_decap_8 FILLER_65_255 ();
 sg13g2_fill_1 FILLER_65_262 ();
 sg13g2_decap_4 FILLER_65_267 ();
 sg13g2_fill_1 FILLER_65_284 ();
 sg13g2_decap_4 FILLER_65_302 ();
 sg13g2_fill_2 FILLER_65_306 ();
 sg13g2_fill_1 FILLER_65_321 ();
 sg13g2_decap_8 FILLER_65_330 ();
 sg13g2_fill_2 FILLER_65_337 ();
 sg13g2_decap_8 FILLER_65_344 ();
 sg13g2_decap_4 FILLER_65_351 ();
 sg13g2_decap_4 FILLER_65_363 ();
 sg13g2_decap_4 FILLER_65_375 ();
 sg13g2_decap_4 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_47 ();
 sg13g2_fill_1 FILLER_66_51 ();
 sg13g2_fill_2 FILLER_66_60 ();
 sg13g2_decap_8 FILLER_66_75 ();
 sg13g2_fill_2 FILLER_66_82 ();
 sg13g2_fill_1 FILLER_66_119 ();
 sg13g2_fill_1 FILLER_66_129 ();
 sg13g2_fill_2 FILLER_66_142 ();
 sg13g2_fill_2 FILLER_66_180 ();
 sg13g2_decap_4 FILLER_66_217 ();
 sg13g2_fill_1 FILLER_66_221 ();
 sg13g2_decap_8 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_242 ();
 sg13g2_fill_2 FILLER_66_287 ();
 sg13g2_decap_4 FILLER_66_307 ();
 sg13g2_fill_1 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_353 ();
 sg13g2_fill_2 FILLER_66_364 ();
 sg13g2_decap_4 FILLER_66_382 ();
 sg13g2_fill_2 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_402 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_11 ();
 sg13g2_fill_1 FILLER_67_45 ();
 sg13g2_fill_2 FILLER_67_59 ();
 sg13g2_fill_1 FILLER_67_61 ();
 sg13g2_fill_2 FILLER_67_72 ();
 sg13g2_fill_2 FILLER_67_83 ();
 sg13g2_fill_1 FILLER_67_85 ();
 sg13g2_fill_2 FILLER_67_93 ();
 sg13g2_fill_2 FILLER_67_113 ();
 sg13g2_fill_1 FILLER_67_154 ();
 sg13g2_fill_2 FILLER_67_173 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_decap_4 FILLER_67_233 ();
 sg13g2_decap_8 FILLER_67_246 ();
 sg13g2_decap_8 FILLER_67_253 ();
 sg13g2_decap_8 FILLER_67_260 ();
 sg13g2_decap_8 FILLER_67_267 ();
 sg13g2_fill_1 FILLER_67_274 ();
 sg13g2_fill_1 FILLER_67_306 ();
 sg13g2_decap_4 FILLER_67_350 ();
 sg13g2_fill_2 FILLER_67_354 ();
 sg13g2_fill_1 FILLER_67_364 ();
 sg13g2_fill_2 FILLER_67_374 ();
 sg13g2_fill_1 FILLER_67_376 ();
 sg13g2_fill_1 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_4 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_decap_8 FILLER_68_50 ();
 sg13g2_fill_1 FILLER_68_57 ();
 sg13g2_decap_4 FILLER_68_62 ();
 sg13g2_fill_1 FILLER_68_66 ();
 sg13g2_fill_2 FILLER_68_105 ();
 sg13g2_fill_1 FILLER_68_107 ();
 sg13g2_fill_2 FILLER_68_120 ();
 sg13g2_fill_1 FILLER_68_164 ();
 sg13g2_fill_1 FILLER_68_177 ();
 sg13g2_fill_2 FILLER_68_187 ();
 sg13g2_fill_2 FILLER_68_227 ();
 sg13g2_fill_1 FILLER_68_343 ();
 sg13g2_fill_1 FILLER_68_348 ();
 sg13g2_fill_2 FILLER_68_383 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_29 ();
 sg13g2_fill_1 FILLER_69_31 ();
 sg13g2_fill_2 FILLER_69_38 ();
 sg13g2_decap_4 FILLER_69_50 ();
 sg13g2_decap_4 FILLER_69_75 ();
 sg13g2_fill_1 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_120 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_fill_2 FILLER_69_216 ();
 sg13g2_fill_1 FILLER_69_226 ();
 sg13g2_decap_4 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_306 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_21 ();
 sg13g2_fill_1 FILLER_70_23 ();
 sg13g2_fill_1 FILLER_70_36 ();
 sg13g2_fill_2 FILLER_70_50 ();
 sg13g2_fill_1 FILLER_70_52 ();
 sg13g2_fill_2 FILLER_70_58 ();
 sg13g2_fill_1 FILLER_70_60 ();
 sg13g2_fill_2 FILLER_70_74 ();
 sg13g2_fill_1 FILLER_70_76 ();
 sg13g2_decap_8 FILLER_70_82 ();
 sg13g2_decap_8 FILLER_70_89 ();
 sg13g2_decap_4 FILLER_70_100 ();
 sg13g2_fill_1 FILLER_70_104 ();
 sg13g2_fill_1 FILLER_70_150 ();
 sg13g2_fill_2 FILLER_70_177 ();
 sg13g2_fill_2 FILLER_70_188 ();
 sg13g2_fill_2 FILLER_70_222 ();
 sg13g2_fill_1 FILLER_70_246 ();
 sg13g2_decap_4 FILLER_70_259 ();
 sg13g2_fill_1 FILLER_70_263 ();
 sg13g2_decap_8 FILLER_70_269 ();
 sg13g2_fill_2 FILLER_70_276 ();
 sg13g2_fill_2 FILLER_70_308 ();
 sg13g2_fill_2 FILLER_70_315 ();
 sg13g2_fill_2 FILLER_70_381 ();
 sg13g2_fill_1 FILLER_70_383 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_fill_2 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_16 ();
 sg13g2_fill_2 FILLER_71_61 ();
 sg13g2_fill_1 FILLER_71_63 ();
 sg13g2_decap_4 FILLER_71_96 ();
 sg13g2_fill_2 FILLER_71_126 ();
 sg13g2_fill_1 FILLER_71_151 ();
 sg13g2_decap_8 FILLER_71_219 ();
 sg13g2_fill_2 FILLER_71_226 ();
 sg13g2_fill_1 FILLER_71_228 ();
 sg13g2_decap_4 FILLER_71_233 ();
 sg13g2_fill_1 FILLER_71_253 ();
 sg13g2_fill_1 FILLER_71_311 ();
 sg13g2_fill_2 FILLER_71_321 ();
 sg13g2_fill_2 FILLER_71_328 ();
 sg13g2_fill_2 FILLER_71_335 ();
 sg13g2_fill_2 FILLER_71_342 ();
 sg13g2_fill_2 FILLER_71_348 ();
 sg13g2_fill_1 FILLER_71_350 ();
 sg13g2_fill_2 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_fill_2 FILLER_71_389 ();
 sg13g2_fill_1 FILLER_71_391 ();
 sg13g2_decap_8 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_52 ();
 sg13g2_fill_2 FILLER_72_74 ();
 sg13g2_fill_1 FILLER_72_76 ();
 sg13g2_fill_2 FILLER_72_103 ();
 sg13g2_fill_1 FILLER_72_136 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_fill_1 FILLER_72_173 ();
 sg13g2_fill_1 FILLER_72_189 ();
 sg13g2_decap_4 FILLER_72_217 ();
 sg13g2_fill_2 FILLER_72_256 ();
 sg13g2_fill_1 FILLER_72_258 ();
 sg13g2_fill_1 FILLER_72_288 ();
 sg13g2_fill_2 FILLER_72_319 ();
 sg13g2_fill_1 FILLER_72_321 ();
 sg13g2_decap_4 FILLER_72_327 ();
 sg13g2_decap_8 FILLER_72_346 ();
 sg13g2_fill_2 FILLER_72_353 ();
 sg13g2_decap_8 FILLER_72_373 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_fill_2 FILLER_73_28 ();
 sg13g2_fill_1 FILLER_73_30 ();
 sg13g2_fill_1 FILLER_73_54 ();
 sg13g2_decap_4 FILLER_73_68 ();
 sg13g2_fill_1 FILLER_73_124 ();
 sg13g2_fill_1 FILLER_73_146 ();
 sg13g2_fill_1 FILLER_73_174 ();
 sg13g2_fill_2 FILLER_73_218 ();
 sg13g2_fill_1 FILLER_73_263 ();
 sg13g2_fill_1 FILLER_73_288 ();
 sg13g2_fill_2 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_41 ();
 sg13g2_fill_1 FILLER_74_43 ();
 sg13g2_decap_8 FILLER_74_48 ();
 sg13g2_fill_2 FILLER_74_55 ();
 sg13g2_fill_1 FILLER_74_57 ();
 sg13g2_decap_8 FILLER_74_62 ();
 sg13g2_decap_8 FILLER_74_69 ();
 sg13g2_decap_8 FILLER_74_76 ();
 sg13g2_decap_8 FILLER_74_87 ();
 sg13g2_decap_8 FILLER_74_94 ();
 sg13g2_fill_1 FILLER_74_101 ();
 sg13g2_fill_1 FILLER_74_135 ();
 sg13g2_fill_1 FILLER_74_197 ();
 sg13g2_fill_1 FILLER_74_247 ();
 sg13g2_fill_2 FILLER_74_258 ();
 sg13g2_fill_1 FILLER_74_386 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_4 FILLER_75_98 ();
 sg13g2_fill_2 FILLER_75_102 ();
 sg13g2_fill_2 FILLER_75_150 ();
 sg13g2_decap_4 FILLER_75_243 ();
 sg13g2_fill_2 FILLER_75_260 ();
 sg13g2_fill_1 FILLER_75_262 ();
 sg13g2_fill_2 FILLER_75_279 ();
 sg13g2_fill_2 FILLER_75_291 ();
 sg13g2_fill_1 FILLER_75_302 ();
 sg13g2_fill_2 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_367 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_fill_2 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_2 FILLER_76_142 ();
 sg13g2_fill_2 FILLER_76_196 ();
 sg13g2_fill_1 FILLER_76_216 ();
 sg13g2_decap_8 FILLER_76_243 ();
 sg13g2_fill_1 FILLER_76_250 ();
 sg13g2_fill_1 FILLER_76_296 ();
 sg13g2_fill_2 FILLER_76_316 ();
 sg13g2_fill_2 FILLER_76_326 ();
 sg13g2_fill_2 FILLER_76_350 ();
 sg13g2_fill_2 FILLER_76_361 ();
 sg13g2_fill_2 FILLER_76_372 ();
 sg13g2_fill_2 FILLER_76_397 ();
 sg13g2_fill_1 FILLER_76_399 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_fill_2 FILLER_77_119 ();
 sg13g2_fill_1 FILLER_77_209 ();
 sg13g2_fill_1 FILLER_77_250 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_fill_2 FILLER_77_329 ();
 sg13g2_fill_2 FILLER_77_366 ();
 sg13g2_fill_1 FILLER_77_368 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_fill_2 FILLER_78_119 ();
 sg13g2_fill_1 FILLER_78_178 ();
 sg13g2_fill_2 FILLER_78_224 ();
 sg13g2_fill_1 FILLER_78_256 ();
 sg13g2_fill_1 FILLER_78_265 ();
 sg13g2_fill_1 FILLER_78_301 ();
 sg13g2_fill_2 FILLER_78_380 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_206 ();
 sg13g2_fill_2 FILLER_79_238 ();
 sg13g2_fill_1 FILLER_79_240 ();
 sg13g2_fill_2 FILLER_79_272 ();
 sg13g2_fill_2 FILLER_79_300 ();
 sg13g2_fill_1 FILLER_79_320 ();
 sg13g2_fill_2 FILLER_79_348 ();
 sg13g2_fill_2 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_fill_2 FILLER_80_108 ();
 sg13g2_fill_2 FILLER_80_164 ();
 sg13g2_fill_1 FILLER_80_166 ();
 sg13g2_fill_2 FILLER_80_172 ();
 sg13g2_fill_1 FILLER_80_174 ();
 sg13g2_fill_2 FILLER_80_194 ();
 sg13g2_fill_2 FILLER_80_204 ();
 sg13g2_fill_1 FILLER_80_206 ();
 sg13g2_fill_1 FILLER_80_216 ();
 sg13g2_fill_1 FILLER_80_257 ();
 sg13g2_fill_1 FILLER_80_267 ();
 sg13g2_decap_4 FILLER_80_277 ();
 sg13g2_fill_2 FILLER_80_300 ();
 sg13g2_fill_1 FILLER_80_302 ();
 sg13g2_decap_4 FILLER_80_321 ();
 sg13g2_fill_1 FILLER_80_325 ();
 sg13g2_fill_1 FILLER_80_344 ();
 sg13g2_fill_2 FILLER_80_358 ();
 sg13g2_fill_1 FILLER_80_360 ();
 sg13g2_fill_2 FILLER_80_374 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
 assign uo_out[2] = net21;
 assign uo_out[3] = net22;
 assign uo_out[4] = net23;
 assign uo_out[5] = net24;
 assign uo_out[6] = net25;
 assign uo_out[7] = net26;
endmodule

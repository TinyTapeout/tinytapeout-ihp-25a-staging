module tt_um_tommythorn_maxbw (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire \tokenflow_inst.i1.c.maj.C ;
 wire \tokenflow_inst.i10.cg.b ;
 wire \tokenflow_inst.i10.cg.maj.C ;
 wire \tokenflow_inst.i10.d0.inv_chain[0] ;
 wire \tokenflow_inst.i10.d0.inv_chain[1] ;
 wire \tokenflow_inst.i11.i.cg.maj.C ;
 wire \tokenflow_inst.i11.i.d0.inv_chain[0] ;
 wire \tokenflow_inst.i11.i.d0.inv_chain[1] ;
 wire \tokenflow_inst.i2.cg1.maj.C ;
 wire \tokenflow_inst.i2.cg2.a ;
 wire \tokenflow_inst.i2.cg2.maj.C ;
 wire \tokenflow_inst.i2.cg3.maj.C ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i3.ydata[0] ;
 wire \tokenflow_inst.i3.ydata[10] ;
 wire \tokenflow_inst.i3.ydata[11] ;
 wire \tokenflow_inst.i3.ydata[12] ;
 wire \tokenflow_inst.i3.ydata[13] ;
 wire \tokenflow_inst.i3.ydata[14] ;
 wire \tokenflow_inst.i3.ydata[15] ;
 wire \tokenflow_inst.i3.ydata[16] ;
 wire \tokenflow_inst.i3.ydata[17] ;
 wire \tokenflow_inst.i3.ydata[18] ;
 wire \tokenflow_inst.i3.ydata[19] ;
 wire \tokenflow_inst.i3.ydata[1] ;
 wire \tokenflow_inst.i3.ydata[20] ;
 wire \tokenflow_inst.i3.ydata[21] ;
 wire \tokenflow_inst.i3.ydata[22] ;
 wire \tokenflow_inst.i3.ydata[23] ;
 wire \tokenflow_inst.i3.ydata[24] ;
 wire \tokenflow_inst.i3.ydata[25] ;
 wire \tokenflow_inst.i3.ydata[26] ;
 wire \tokenflow_inst.i3.ydata[27] ;
 wire \tokenflow_inst.i3.ydata[28] ;
 wire \tokenflow_inst.i3.ydata[29] ;
 wire \tokenflow_inst.i3.ydata[2] ;
 wire \tokenflow_inst.i3.ydata[30] ;
 wire \tokenflow_inst.i3.ydata[31] ;
 wire \tokenflow_inst.i3.ydata[32] ;
 wire \tokenflow_inst.i3.ydata[33] ;
 wire \tokenflow_inst.i3.ydata[34] ;
 wire \tokenflow_inst.i3.ydata[35] ;
 wire \tokenflow_inst.i3.ydata[36] ;
 wire \tokenflow_inst.i3.ydata[37] ;
 wire \tokenflow_inst.i3.ydata[38] ;
 wire \tokenflow_inst.i3.ydata[39] ;
 wire \tokenflow_inst.i3.ydata[3] ;
 wire \tokenflow_inst.i3.ydata[40] ;
 wire \tokenflow_inst.i3.ydata[41] ;
 wire \tokenflow_inst.i3.ydata[42] ;
 wire \tokenflow_inst.i3.ydata[43] ;
 wire \tokenflow_inst.i3.ydata[44] ;
 wire \tokenflow_inst.i3.ydata[45] ;
 wire \tokenflow_inst.i3.ydata[46] ;
 wire \tokenflow_inst.i3.ydata[47] ;
 wire \tokenflow_inst.i3.ydata[48] ;
 wire \tokenflow_inst.i3.ydata[49] ;
 wire \tokenflow_inst.i3.ydata[4] ;
 wire \tokenflow_inst.i3.ydata[50] ;
 wire \tokenflow_inst.i3.ydata[51] ;
 wire \tokenflow_inst.i3.ydata[52] ;
 wire \tokenflow_inst.i3.ydata[53] ;
 wire \tokenflow_inst.i3.ydata[54] ;
 wire \tokenflow_inst.i3.ydata[55] ;
 wire \tokenflow_inst.i3.ydata[56] ;
 wire \tokenflow_inst.i3.ydata[57] ;
 wire \tokenflow_inst.i3.ydata[58] ;
 wire \tokenflow_inst.i3.ydata[59] ;
 wire \tokenflow_inst.i3.ydata[5] ;
 wire \tokenflow_inst.i3.ydata[60] ;
 wire \tokenflow_inst.i3.ydata[61] ;
 wire \tokenflow_inst.i3.ydata[62] ;
 wire \tokenflow_inst.i3.ydata[63] ;
 wire \tokenflow_inst.i3.ydata[64] ;
 wire \tokenflow_inst.i3.ydata[65] ;
 wire \tokenflow_inst.i3.ydata[66] ;
 wire \tokenflow_inst.i3.ydata[67] ;
 wire \tokenflow_inst.i3.ydata[68] ;
 wire \tokenflow_inst.i3.ydata[69] ;
 wire \tokenflow_inst.i3.ydata[6] ;
 wire \tokenflow_inst.i3.ydata[70] ;
 wire \tokenflow_inst.i3.ydata[71] ;
 wire \tokenflow_inst.i3.ydata[72] ;
 wire \tokenflow_inst.i3.ydata[73] ;
 wire \tokenflow_inst.i3.ydata[74] ;
 wire \tokenflow_inst.i3.ydata[75] ;
 wire \tokenflow_inst.i3.ydata[76] ;
 wire \tokenflow_inst.i3.ydata[77] ;
 wire \tokenflow_inst.i3.ydata[7] ;
 wire \tokenflow_inst.i3.ydata[8] ;
 wire \tokenflow_inst.i3.ydata[9] ;
 wire \tokenflow_inst.i6.cg_elem.maj.C ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[10] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[11] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[12] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[13] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[14] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[15] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[16] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[17] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[18] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[19] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[20] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[21] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[22] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[23] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[24] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[25] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[26] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[27] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[28] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[29] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[30] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[31] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[32] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[33] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[34] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[35] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[36] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[37] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[38] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[39] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[40] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[41] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[42] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[43] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[44] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[45] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[46] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[47] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[48] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[49] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[4] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[50] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[51] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[52] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[5] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[6] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[7] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[8] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[9] ;
 wire \tokenflow_inst.i6.ydata[0] ;
 wire \tokenflow_inst.i6.ydata[10] ;
 wire \tokenflow_inst.i6.ydata[11] ;
 wire \tokenflow_inst.i6.ydata[12] ;
 wire \tokenflow_inst.i6.ydata[13] ;
 wire \tokenflow_inst.i6.ydata[14] ;
 wire \tokenflow_inst.i6.ydata[15] ;
 wire \tokenflow_inst.i6.ydata[16] ;
 wire \tokenflow_inst.i6.ydata[17] ;
 wire \tokenflow_inst.i6.ydata[18] ;
 wire \tokenflow_inst.i6.ydata[19] ;
 wire \tokenflow_inst.i6.ydata[1] ;
 wire \tokenflow_inst.i6.ydata[20] ;
 wire \tokenflow_inst.i6.ydata[21] ;
 wire \tokenflow_inst.i6.ydata[22] ;
 wire \tokenflow_inst.i6.ydata[23] ;
 wire \tokenflow_inst.i6.ydata[24] ;
 wire \tokenflow_inst.i6.ydata[25] ;
 wire \tokenflow_inst.i6.ydata[26] ;
 wire \tokenflow_inst.i6.ydata[27] ;
 wire \tokenflow_inst.i6.ydata[28] ;
 wire \tokenflow_inst.i6.ydata[29] ;
 wire \tokenflow_inst.i6.ydata[2] ;
 wire \tokenflow_inst.i6.ydata[30] ;
 wire \tokenflow_inst.i6.ydata[31] ;
 wire \tokenflow_inst.i6.ydata[32] ;
 wire \tokenflow_inst.i6.ydata[33] ;
 wire \tokenflow_inst.i6.ydata[34] ;
 wire \tokenflow_inst.i6.ydata[35] ;
 wire \tokenflow_inst.i6.ydata[36] ;
 wire \tokenflow_inst.i6.ydata[37] ;
 wire \tokenflow_inst.i6.ydata[38] ;
 wire \tokenflow_inst.i6.ydata[39] ;
 wire \tokenflow_inst.i6.ydata[3] ;
 wire \tokenflow_inst.i6.ydata[40] ;
 wire \tokenflow_inst.i6.ydata[41] ;
 wire \tokenflow_inst.i6.ydata[42] ;
 wire \tokenflow_inst.i6.ydata[43] ;
 wire \tokenflow_inst.i6.ydata[44] ;
 wire \tokenflow_inst.i6.ydata[45] ;
 wire \tokenflow_inst.i6.ydata[46] ;
 wire \tokenflow_inst.i6.ydata[47] ;
 wire \tokenflow_inst.i6.ydata[48] ;
 wire \tokenflow_inst.i6.ydata[49] ;
 wire \tokenflow_inst.i6.ydata[4] ;
 wire \tokenflow_inst.i6.ydata[50] ;
 wire \tokenflow_inst.i6.ydata[51] ;
 wire \tokenflow_inst.i6.ydata[52] ;
 wire \tokenflow_inst.i6.ydata[53] ;
 wire \tokenflow_inst.i6.ydata[54] ;
 wire \tokenflow_inst.i6.ydata[55] ;
 wire \tokenflow_inst.i6.ydata[56] ;
 wire \tokenflow_inst.i6.ydata[57] ;
 wire \tokenflow_inst.i6.ydata[58] ;
 wire \tokenflow_inst.i6.ydata[59] ;
 wire \tokenflow_inst.i6.ydata[5] ;
 wire \tokenflow_inst.i6.ydata[60] ;
 wire \tokenflow_inst.i6.ydata[61] ;
 wire \tokenflow_inst.i6.ydata[62] ;
 wire \tokenflow_inst.i6.ydata[63] ;
 wire \tokenflow_inst.i6.ydata[64] ;
 wire \tokenflow_inst.i6.ydata[65] ;
 wire \tokenflow_inst.i6.ydata[66] ;
 wire \tokenflow_inst.i6.ydata[67] ;
 wire \tokenflow_inst.i6.ydata[68] ;
 wire \tokenflow_inst.i6.ydata[69] ;
 wire \tokenflow_inst.i6.ydata[6] ;
 wire \tokenflow_inst.i6.ydata[70] ;
 wire \tokenflow_inst.i6.ydata[71] ;
 wire \tokenflow_inst.i6.ydata[72] ;
 wire \tokenflow_inst.i6.ydata[73] ;
 wire \tokenflow_inst.i6.ydata[74] ;
 wire \tokenflow_inst.i6.ydata[75] ;
 wire \tokenflow_inst.i6.ydata[76] ;
 wire \tokenflow_inst.i6.ydata[77] ;
 wire \tokenflow_inst.i6.ydata[7] ;
 wire \tokenflow_inst.i6.ydata[8] ;
 wire \tokenflow_inst.i6.ydata[9] ;
 wire \tokenflow_inst.i78.cg_elem.maj.C ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i78.ydata[0] ;
 wire \tokenflow_inst.i78.ydata[10] ;
 wire \tokenflow_inst.i78.ydata[11] ;
 wire \tokenflow_inst.i78.ydata[12] ;
 wire \tokenflow_inst.i78.ydata[13] ;
 wire \tokenflow_inst.i78.ydata[14] ;
 wire \tokenflow_inst.i78.ydata[15] ;
 wire \tokenflow_inst.i78.ydata[16] ;
 wire \tokenflow_inst.i78.ydata[17] ;
 wire \tokenflow_inst.i78.ydata[18] ;
 wire \tokenflow_inst.i78.ydata[19] ;
 wire \tokenflow_inst.i78.ydata[1] ;
 wire \tokenflow_inst.i78.ydata[20] ;
 wire \tokenflow_inst.i78.ydata[21] ;
 wire \tokenflow_inst.i78.ydata[22] ;
 wire \tokenflow_inst.i78.ydata[23] ;
 wire \tokenflow_inst.i78.ydata[24] ;
 wire \tokenflow_inst.i78.ydata[25] ;
 wire \tokenflow_inst.i78.ydata[26] ;
 wire \tokenflow_inst.i78.ydata[27] ;
 wire \tokenflow_inst.i78.ydata[28] ;
 wire \tokenflow_inst.i78.ydata[29] ;
 wire \tokenflow_inst.i78.ydata[2] ;
 wire \tokenflow_inst.i78.ydata[30] ;
 wire \tokenflow_inst.i78.ydata[31] ;
 wire \tokenflow_inst.i78.ydata[32] ;
 wire \tokenflow_inst.i78.ydata[33] ;
 wire \tokenflow_inst.i78.ydata[34] ;
 wire \tokenflow_inst.i78.ydata[35] ;
 wire \tokenflow_inst.i78.ydata[36] ;
 wire \tokenflow_inst.i78.ydata[37] ;
 wire \tokenflow_inst.i78.ydata[38] ;
 wire \tokenflow_inst.i78.ydata[39] ;
 wire \tokenflow_inst.i78.ydata[3] ;
 wire \tokenflow_inst.i78.ydata[40] ;
 wire \tokenflow_inst.i78.ydata[41] ;
 wire \tokenflow_inst.i78.ydata[42] ;
 wire \tokenflow_inst.i78.ydata[43] ;
 wire \tokenflow_inst.i78.ydata[44] ;
 wire \tokenflow_inst.i78.ydata[45] ;
 wire \tokenflow_inst.i78.ydata[46] ;
 wire \tokenflow_inst.i78.ydata[47] ;
 wire \tokenflow_inst.i78.ydata[48] ;
 wire \tokenflow_inst.i78.ydata[49] ;
 wire \tokenflow_inst.i78.ydata[4] ;
 wire \tokenflow_inst.i78.ydata[54] ;
 wire \tokenflow_inst.i78.ydata[55] ;
 wire \tokenflow_inst.i78.ydata[56] ;
 wire \tokenflow_inst.i78.ydata[57] ;
 wire \tokenflow_inst.i78.ydata[58] ;
 wire \tokenflow_inst.i78.ydata[59] ;
 wire \tokenflow_inst.i78.ydata[5] ;
 wire \tokenflow_inst.i78.ydata[60] ;
 wire \tokenflow_inst.i78.ydata[61] ;
 wire \tokenflow_inst.i78.ydata[62] ;
 wire \tokenflow_inst.i78.ydata[63] ;
 wire \tokenflow_inst.i78.ydata[64] ;
 wire \tokenflow_inst.i78.ydata[65] ;
 wire \tokenflow_inst.i78.ydata[66] ;
 wire \tokenflow_inst.i78.ydata[67] ;
 wire \tokenflow_inst.i78.ydata[68] ;
 wire \tokenflow_inst.i78.ydata[69] ;
 wire \tokenflow_inst.i78.ydata[6] ;
 wire \tokenflow_inst.i78.ydata[70] ;
 wire \tokenflow_inst.i78.ydata[71] ;
 wire \tokenflow_inst.i78.ydata[72] ;
 wire \tokenflow_inst.i78.ydata[73] ;
 wire \tokenflow_inst.i78.ydata[74] ;
 wire \tokenflow_inst.i78.ydata[75] ;
 wire \tokenflow_inst.i78.ydata[76] ;
 wire \tokenflow_inst.i78.ydata[77] ;
 wire \tokenflow_inst.i78.ydata[7] ;
 wire \tokenflow_inst.i78.ydata[8] ;
 wire \tokenflow_inst.i78.ydata[9] ;
 wire \tokenflow_inst.i8.cg_elem.maj.C ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[10] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[11] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[12] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[13] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[14] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[15] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[16] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[17] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[18] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[19] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[20] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[21] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[22] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[23] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[24] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[25] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[26] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[27] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[28] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[29] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[30] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[31] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[32] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[33] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[34] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[35] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[36] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[37] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[38] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[39] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[40] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[41] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[42] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[43] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[44] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[45] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[46] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[47] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[48] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[49] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[4] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[50] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[51] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[52] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[5] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[6] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[7] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[8] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[9] ;
 wire \tokenflow_inst.i8.ydata[0] ;
 wire \tokenflow_inst.i8.ydata[10] ;
 wire \tokenflow_inst.i8.ydata[11] ;
 wire \tokenflow_inst.i8.ydata[12] ;
 wire \tokenflow_inst.i8.ydata[13] ;
 wire \tokenflow_inst.i8.ydata[14] ;
 wire \tokenflow_inst.i8.ydata[15] ;
 wire \tokenflow_inst.i8.ydata[16] ;
 wire \tokenflow_inst.i8.ydata[17] ;
 wire \tokenflow_inst.i8.ydata[18] ;
 wire \tokenflow_inst.i8.ydata[19] ;
 wire \tokenflow_inst.i8.ydata[1] ;
 wire \tokenflow_inst.i8.ydata[20] ;
 wire \tokenflow_inst.i8.ydata[21] ;
 wire \tokenflow_inst.i8.ydata[22] ;
 wire \tokenflow_inst.i8.ydata[23] ;
 wire \tokenflow_inst.i8.ydata[24] ;
 wire \tokenflow_inst.i8.ydata[25] ;
 wire \tokenflow_inst.i8.ydata[26] ;
 wire \tokenflow_inst.i8.ydata[27] ;
 wire \tokenflow_inst.i8.ydata[28] ;
 wire \tokenflow_inst.i8.ydata[29] ;
 wire \tokenflow_inst.i8.ydata[2] ;
 wire \tokenflow_inst.i8.ydata[30] ;
 wire \tokenflow_inst.i8.ydata[31] ;
 wire \tokenflow_inst.i8.ydata[32] ;
 wire \tokenflow_inst.i8.ydata[33] ;
 wire \tokenflow_inst.i8.ydata[34] ;
 wire \tokenflow_inst.i8.ydata[35] ;
 wire \tokenflow_inst.i8.ydata[36] ;
 wire \tokenflow_inst.i8.ydata[37] ;
 wire \tokenflow_inst.i8.ydata[38] ;
 wire \tokenflow_inst.i8.ydata[39] ;
 wire \tokenflow_inst.i8.ydata[3] ;
 wire \tokenflow_inst.i8.ydata[40] ;
 wire \tokenflow_inst.i8.ydata[41] ;
 wire \tokenflow_inst.i8.ydata[42] ;
 wire \tokenflow_inst.i8.ydata[43] ;
 wire \tokenflow_inst.i8.ydata[44] ;
 wire \tokenflow_inst.i8.ydata[45] ;
 wire \tokenflow_inst.i8.ydata[46] ;
 wire \tokenflow_inst.i8.ydata[47] ;
 wire \tokenflow_inst.i8.ydata[48] ;
 wire \tokenflow_inst.i8.ydata[49] ;
 wire \tokenflow_inst.i8.ydata[4] ;
 wire \tokenflow_inst.i8.ydata[50] ;
 wire net2;
 wire \tokenflow_inst.i8.ydata[53] ;
 wire \tokenflow_inst.i8.ydata[54] ;
 wire \tokenflow_inst.i8.ydata[55] ;
 wire \tokenflow_inst.i8.ydata[56] ;
 wire \tokenflow_inst.i8.ydata[57] ;
 wire \tokenflow_inst.i8.ydata[58] ;
 wire \tokenflow_inst.i8.ydata[59] ;
 wire \tokenflow_inst.i8.ydata[5] ;
 wire \tokenflow_inst.i8.ydata[60] ;
 wire \tokenflow_inst.i8.ydata[61] ;
 wire \tokenflow_inst.i8.ydata[62] ;
 wire \tokenflow_inst.i8.ydata[63] ;
 wire \tokenflow_inst.i8.ydata[64] ;
 wire \tokenflow_inst.i8.ydata[65] ;
 wire \tokenflow_inst.i8.ydata[66] ;
 wire \tokenflow_inst.i8.ydata[67] ;
 wire \tokenflow_inst.i8.ydata[68] ;
 wire \tokenflow_inst.i8.ydata[69] ;
 wire \tokenflow_inst.i8.ydata[6] ;
 wire \tokenflow_inst.i8.ydata[70] ;
 wire \tokenflow_inst.i8.ydata[71] ;
 wire \tokenflow_inst.i8.ydata[72] ;
 wire \tokenflow_inst.i8.ydata[73] ;
 wire \tokenflow_inst.i8.ydata[74] ;
 wire \tokenflow_inst.i8.ydata[75] ;
 wire \tokenflow_inst.i8.ydata[76] ;
 wire \tokenflow_inst.i8.ydata[77] ;
 wire \tokenflow_inst.i8.ydata[7] ;
 wire \tokenflow_inst.i8.ydata[8] ;
 wire \tokenflow_inst.i8.ydata[9] ;
 wire \tokenflow_inst.i9.c.maj.C ;
 wire \tokenflow_inst.ii1.cg_elem.maj.C ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.ii1.ydata[0] ;
 wire \tokenflow_inst.ii1.ydata[10] ;
 wire \tokenflow_inst.ii1.ydata[11] ;
 wire \tokenflow_inst.ii1.ydata[12] ;
 wire \tokenflow_inst.ii1.ydata[13] ;
 wire \tokenflow_inst.ii1.ydata[14] ;
 wire \tokenflow_inst.ii1.ydata[15] ;
 wire \tokenflow_inst.ii1.ydata[16] ;
 wire \tokenflow_inst.ii1.ydata[17] ;
 wire \tokenflow_inst.ii1.ydata[18] ;
 wire \tokenflow_inst.ii1.ydata[19] ;
 wire \tokenflow_inst.ii1.ydata[1] ;
 wire \tokenflow_inst.ii1.ydata[20] ;
 wire \tokenflow_inst.ii1.ydata[21] ;
 wire \tokenflow_inst.ii1.ydata[22] ;
 wire \tokenflow_inst.ii1.ydata[23] ;
 wire \tokenflow_inst.ii1.ydata[24] ;
 wire \tokenflow_inst.ii1.ydata[25] ;
 wire \tokenflow_inst.ii1.ydata[2] ;
 wire \tokenflow_inst.ii1.ydata[3] ;
 wire \tokenflow_inst.ii1.ydata[4] ;
 wire \tokenflow_inst.ii1.ydata[5] ;
 wire \tokenflow_inst.ii1.ydata[6] ;
 wire \tokenflow_inst.ii1.ydata[7] ;
 wire \tokenflow_inst.ii1.ydata[8] ;
 wire \tokenflow_inst.ii1.ydata[9] ;
 wire \tokenflow_inst.ii2.cg_elem.maj.C ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.ii2.ydata[0] ;
 wire \tokenflow_inst.ii2.ydata[10] ;
 wire \tokenflow_inst.ii2.ydata[11] ;
 wire \tokenflow_inst.ii2.ydata[12] ;
 wire \tokenflow_inst.ii2.ydata[13] ;
 wire \tokenflow_inst.ii2.ydata[14] ;
 wire \tokenflow_inst.ii2.ydata[15] ;
 wire \tokenflow_inst.ii2.ydata[16] ;
 wire \tokenflow_inst.ii2.ydata[17] ;
 wire \tokenflow_inst.ii2.ydata[18] ;
 wire \tokenflow_inst.ii2.ydata[19] ;
 wire \tokenflow_inst.ii2.ydata[1] ;
 wire \tokenflow_inst.ii2.ydata[20] ;
 wire \tokenflow_inst.ii2.ydata[21] ;
 wire \tokenflow_inst.ii2.ydata[22] ;
 wire \tokenflow_inst.ii2.ydata[23] ;
 wire \tokenflow_inst.ii2.ydata[24] ;
 wire \tokenflow_inst.ii2.ydata[25] ;
 wire \tokenflow_inst.ii2.ydata[2] ;
 wire \tokenflow_inst.ii2.ydata[3] ;
 wire \tokenflow_inst.ii2.ydata[4] ;
 wire \tokenflow_inst.ii2.ydata[5] ;
 wire \tokenflow_inst.ii2.ydata[6] ;
 wire \tokenflow_inst.ii2.ydata[7] ;
 wire \tokenflow_inst.ii2.ydata[8] ;
 wire \tokenflow_inst.ii2.ydata[9] ;
 wire \tokenflow_inst.ii3.i.cg_elem.maj.C ;
 wire \tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii3.i.ydata[0] ;
 wire \tokenflow_inst.ii3.i.ydata[10] ;
 wire \tokenflow_inst.ii3.i.ydata[11] ;
 wire \tokenflow_inst.ii3.i.ydata[12] ;
 wire \tokenflow_inst.ii3.i.ydata[13] ;
 wire \tokenflow_inst.ii3.i.ydata[14] ;
 wire \tokenflow_inst.ii3.i.ydata[15] ;
 wire \tokenflow_inst.ii3.i.ydata[16] ;
 wire \tokenflow_inst.ii3.i.ydata[17] ;
 wire \tokenflow_inst.ii3.i.ydata[18] ;
 wire \tokenflow_inst.ii3.i.ydata[19] ;
 wire \tokenflow_inst.ii3.i.ydata[1] ;
 wire \tokenflow_inst.ii3.i.ydata[20] ;
 wire \tokenflow_inst.ii3.i.ydata[21] ;
 wire \tokenflow_inst.ii3.i.ydata[22] ;
 wire \tokenflow_inst.ii3.i.ydata[23] ;
 wire \tokenflow_inst.ii3.i.ydata[24] ;
 wire \tokenflow_inst.ii3.i.ydata[25] ;
 wire \tokenflow_inst.ii3.i.ydata[2] ;
 wire \tokenflow_inst.ii3.i.ydata[3] ;
 wire \tokenflow_inst.ii3.i.ydata[4] ;
 wire \tokenflow_inst.ii3.i.ydata[5] ;
 wire \tokenflow_inst.ii3.i.ydata[6] ;
 wire \tokenflow_inst.ii3.i.ydata[7] ;
 wire \tokenflow_inst.ii3.i.ydata[8] ;
 wire \tokenflow_inst.ii3.i.ydata[9] ;
 wire \tokenflow_inst.ii4.c.maj.C ;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net1;

 sg13g2_inv_1 _1253_ (.Y(_0738_),
    .A(net686));
 sg13g2_inv_1 _1254_ (.Y(_0739_),
    .A(\tokenflow_inst.i6.ydata[21] ));
 sg13g2_inv_2 _1255_ (.Y(_0740_),
    .A(\tokenflow_inst.ii3.i.ydata[7] ));
 sg13g2_inv_1 _1256_ (.Y(_0741_),
    .A(\tokenflow_inst.ii3.i.ydata[8] ));
 sg13g2_inv_1 _1257_ (.Y(_0742_),
    .A(\tokenflow_inst.ii3.i.ydata[10] ));
 sg13g2_inv_2 _1258_ (.Y(_0743_),
    .A(\tokenflow_inst.ii3.i.ydata[13] ));
 sg13g2_inv_1 _1259_ (.Y(_0744_),
    .A(\tokenflow_inst.ii3.i.ydata[19] ));
 sg13g2_inv_1 _1260_ (.Y(_0745_),
    .A(\tokenflow_inst.ii3.i.ydata[25] ));
 sg13g2_inv_1 _1261_ (.Y(_0746_),
    .A(\tokenflow_inst.i8.ydata[22] ));
 sg13g2_inv_1 _1262_ (.Y(_0747_),
    .A(\tokenflow_inst.i1.c.maj.C ));
 sg13g2_inv_1 _1263_ (.Y(_0748_),
    .A(\tokenflow_inst.i10.cg.maj.C ));
 sg13g2_inv_1 _1264_ (.Y(_0749_),
    .A(\tokenflow_inst.ii4.c.maj.C ));
 sg13g2_a21oi_1 _1265_ (.A1(\tokenflow_inst.i10.cg.maj.C ),
    .A2(\tokenflow_inst.i9.c.maj.C ),
    .Y(_0750_),
    .B1(net1));
 sg13g2_o21ai_1 _1266_ (.B1(net692),
    .Y(_0751_),
    .A1(\tokenflow_inst.i10.cg.maj.C ),
    .A2(\tokenflow_inst.i9.c.maj.C ));
 sg13g2_nor2_1 _1267_ (.A(_0750_),
    .B(_0751_),
    .Y(\tokenflow_inst.i9.c.maj.C ));
 sg13g2_nor2_1 _1268_ (.A(net653),
    .B(\tokenflow_inst.i11.i.cg.maj.C ),
    .Y(_0752_));
 sg13g2_nor4_2 _1269_ (.A(\tokenflow_inst.i3.ydata[49] ),
    .B(\tokenflow_inst.i3.ydata[48] ),
    .C(\tokenflow_inst.i3.ydata[51] ),
    .Y(_0753_),
    .D(\tokenflow_inst.i3.ydata[50] ));
 sg13g2_nor4_1 _1270_ (.A(\tokenflow_inst.i3.ydata[45] ),
    .B(\tokenflow_inst.i3.ydata[44] ),
    .C(\tokenflow_inst.i3.ydata[47] ),
    .D(\tokenflow_inst.i3.ydata[46] ),
    .Y(_0754_));
 sg13g2_nor4_1 _1271_ (.A(\tokenflow_inst.i3.ydata[41] ),
    .B(\tokenflow_inst.i3.ydata[40] ),
    .C(\tokenflow_inst.i3.ydata[43] ),
    .D(\tokenflow_inst.i3.ydata[42] ),
    .Y(_0755_));
 sg13g2_nand3_1 _1272_ (.B(_0754_),
    .C(_0755_),
    .A(_0753_),
    .Y(_0756_));
 sg13g2_nor2_1 _1273_ (.A(\tokenflow_inst.i3.ydata[27] ),
    .B(\tokenflow_inst.i3.ydata[26] ),
    .Y(_0757_));
 sg13g2_nor4_1 _1274_ (.A(\tokenflow_inst.i3.ydata[29] ),
    .B(\tokenflow_inst.i3.ydata[28] ),
    .C(\tokenflow_inst.i3.ydata[31] ),
    .D(\tokenflow_inst.i3.ydata[30] ),
    .Y(_0758_));
 sg13g2_nor4_2 _1275_ (.A(\tokenflow_inst.i3.ydata[37] ),
    .B(\tokenflow_inst.i3.ydata[36] ),
    .C(\tokenflow_inst.i3.ydata[39] ),
    .Y(_0759_),
    .D(\tokenflow_inst.i3.ydata[38] ));
 sg13g2_nor4_1 _1276_ (.A(\tokenflow_inst.i3.ydata[33] ),
    .B(\tokenflow_inst.i3.ydata[32] ),
    .C(\tokenflow_inst.i3.ydata[35] ),
    .D(\tokenflow_inst.i3.ydata[34] ),
    .Y(_0760_));
 sg13g2_nand4_1 _1277_ (.B(_0758_),
    .C(_0759_),
    .A(_0757_),
    .Y(_0761_),
    .D(_0760_));
 sg13g2_nor2_1 _1278_ (.A(_0756_),
    .B(_0761_),
    .Y(_0762_));
 sg13g2_and2_1 _1279_ (.A(net692),
    .B(\tokenflow_inst.i2.cg2.a ),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[0] ));
 sg13g2_and2_1 _1280_ (.A(_0762_),
    .B(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i10.cg.b ));
 sg13g2_a21oi_1 _1281_ (.A1(\tokenflow_inst.i10.cg.maj.C ),
    .A2(_0752_),
    .Y(_0763_),
    .B1(\tokenflow_inst.i10.cg.b ));
 sg13g2_a21oi_2 _1282_ (.B1(_0763_),
    .Y(\tokenflow_inst.i10.cg.maj.C ),
    .A2(_0748_),
    .A1(\tokenflow_inst.i11.i.cg.maj.C ));
 sg13g2_nor2_1 _1283_ (.A(net653),
    .B(_0748_),
    .Y(\tokenflow_inst.i10.d0.inv_chain[0] ));
 sg13g2_nand2_1 _1284_ (.Y(_0764_),
    .A(net686),
    .B(\tokenflow_inst.i2.cg3.maj.C ));
 sg13g2_nand2_1 _1285_ (.Y(_0765_),
    .A(net685),
    .B(\tokenflow_inst.ii1.cg_elem.maj.C ));
 sg13g2_inv_1 _1286_ (.Y(\tokenflow_inst.ii1.d0_elem.inv_chain[0] ),
    .A(_0765_));
 sg13g2_o21ai_1 _1287_ (.B1(\tokenflow_inst.ii1.d0_elem.inv_chain[0] ),
    .Y(_0766_),
    .A1(\tokenflow_inst.i2.cg3.maj.C ),
    .A2(\tokenflow_inst.ii4.c.maj.C ));
 sg13g2_o21ai_1 _1288_ (.B1(_0766_),
    .Y(\tokenflow_inst.ii4.c.maj.C ),
    .A1(_0749_),
    .A2(_0764_));
 sg13g2_nor2_1 _1289_ (.A(net654),
    .B(\tokenflow_inst.ii2.cg_elem.maj.C ),
    .Y(_0363_));
 sg13g2_nor2_1 _1290_ (.A(net652),
    .B(\tokenflow_inst.ii3.i.cg_elem.maj.C ),
    .Y(_0390_));
 sg13g2_nand2b_1 _1291_ (.Y(_0767_),
    .B(\tokenflow_inst.ii2.cg_elem.maj.C ),
    .A_N(\tokenflow_inst.ii4.c.maj.C ));
 sg13g2_a22oi_1 _1292_ (.Y(\tokenflow_inst.ii3.i.cg_elem.maj.C ),
    .B1(net631),
    .B2(_0767_),
    .A2(net613),
    .A1(\tokenflow_inst.ii4.c.maj.C ));
 sg13g2_nand2_1 _1293_ (.Y(_0768_),
    .A(\tokenflow_inst.ii2.cg_elem.maj.C ),
    .B(net630));
 sg13g2_nor2b_1 _1294_ (.A(\tokenflow_inst.ii2.cg_elem.maj.C ),
    .B_N(\tokenflow_inst.ii3.i.cg_elem.maj.C ),
    .Y(_0769_));
 sg13g2_and2_1 _1295_ (.A(net686),
    .B(\tokenflow_inst.ii2.cg_elem.maj.C ),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[0] ));
 sg13g2_o21ai_1 _1296_ (.B1(_0768_),
    .Y(\tokenflow_inst.ii2.cg_elem.maj.C ),
    .A1(_0765_),
    .A2(_0769_));
 sg13g2_nand2_1 _1297_ (.Y(_0770_),
    .A(\tokenflow_inst.ii3.i.cg_elem.maj.C ),
    .B(net613));
 sg13g2_nor2b_1 _1298_ (.A(\tokenflow_inst.ii3.i.cg_elem.maj.C ),
    .B_N(\tokenflow_inst.ii2.cg_elem.maj.C ),
    .Y(_0771_));
 sg13g2_and2_1 _1299_ (.A(net686),
    .B(\tokenflow_inst.ii3.i.cg_elem.maj.C ),
    .X(\tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ));
 sg13g2_o21ai_1 _1300_ (.B1(_0770_),
    .Y(\tokenflow_inst.ii1.cg_elem.maj.C ),
    .A1(_0765_),
    .A2(_0771_));
 sg13g2_o21ai_1 _1301_ (.B1(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .Y(_0772_),
    .A1(\tokenflow_inst.i1.c.maj.C ),
    .A2(\tokenflow_inst.i2.cg3.maj.C ));
 sg13g2_o21ai_1 _1302_ (.B1(_0772_),
    .Y(\tokenflow_inst.i2.cg3.maj.C ),
    .A1(_0747_),
    .A2(_0764_));
 sg13g2_and2_1 _1303_ (.A(net686),
    .B(\tokenflow_inst.i11.i.cg.maj.C ),
    .X(\tokenflow_inst.i11.i.d0.inv_chain[0] ));
 sg13g2_nand2_1 _1304_ (.Y(_0773_),
    .A(\tokenflow_inst.i1.c.maj.C ),
    .B(\tokenflow_inst.i11.i.d0.inv_chain[0] ));
 sg13g2_o21ai_1 _1305_ (.B1(\tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ),
    .Y(_0774_),
    .A1(\tokenflow_inst.i11.i.cg.maj.C ),
    .A2(\tokenflow_inst.i1.c.maj.C ));
 sg13g2_nand2_2 _1306_ (.Y(\tokenflow_inst.i1.c.maj.C ),
    .A(_0773_),
    .B(_0774_));
 sg13g2_a21oi_1 _1307_ (.A1(\tokenflow_inst.i11.i.cg.maj.C ),
    .A2(\tokenflow_inst.i10.cg.maj.C ),
    .Y(_0775_),
    .B1(_0764_));
 sg13g2_a21oi_2 _1308_ (.B1(_0775_),
    .Y(\tokenflow_inst.i11.i.cg.maj.C ),
    .A2(_0752_),
    .A1(_0748_));
 sg13g2_nor2_1 _1309_ (.A(net653),
    .B(\tokenflow_inst.i6.cg_elem.maj.C ),
    .Y(_0157_));
 sg13g2_nor3_1 _1310_ (.A(net653),
    .B(\tokenflow_inst.i6.cg_elem.maj.C ),
    .C(\tokenflow_inst.i9.c.maj.C ),
    .Y(_0776_));
 sg13g2_nor2_1 _1311_ (.A(\tokenflow_inst.i2.cg2.a ),
    .B(_0776_),
    .Y(_0777_));
 sg13g2_nand2_1 _1312_ (.Y(_0778_),
    .A(\tokenflow_inst.i2.cg2.a ),
    .B(_0776_));
 sg13g2_nor2_1 _1313_ (.A(net650),
    .B(net649),
    .Y(_0779_));
 sg13g2_and2_1 _1314_ (.A(net660),
    .B(net649),
    .X(_0780_));
 sg13g2_a22oi_1 _1315_ (.Y(_0781_),
    .B1(net641),
    .B2(\tokenflow_inst.i78.cg_elem.maj.C ),
    .A2(net648),
    .A1(\tokenflow_inst.i1.c.maj.C ));
 sg13g2_o21ai_1 _1316_ (.B1(_0778_),
    .Y(\tokenflow_inst.i2.cg2.a ),
    .A1(_0777_),
    .A2(_0781_));
 sg13g2_a21oi_1 _1317_ (.A1(net649),
    .A2(\tokenflow_inst.i78.cg_elem.maj.C ),
    .Y(_0782_),
    .B1(_0747_));
 sg13g2_and2_1 _1318_ (.A(net691),
    .B(\tokenflow_inst.i78.cg_elem.maj.C ),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[0] ));
 sg13g2_nor2_1 _1319_ (.A(net640),
    .B(\tokenflow_inst.i78.d0_elem.inv_chain[0] ),
    .Y(_0783_));
 sg13g2_nor2_1 _1320_ (.A(_0782_),
    .B(_0783_),
    .Y(\tokenflow_inst.i2.cg1.maj.C ));
 sg13g2_nand2_1 _1321_ (.Y(_0784_),
    .A(\tokenflow_inst.i78.cg_elem.maj.C ),
    .B(\tokenflow_inst.i8.cg_elem.maj.C ));
 sg13g2_and2_1 _1322_ (.A(net690),
    .B(\tokenflow_inst.i8.cg_elem.maj.C ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[0] ));
 sg13g2_nor2_1 _1323_ (.A(\tokenflow_inst.i78.d0_elem.inv_chain[0] ),
    .B(net592),
    .Y(_0785_));
 sg13g2_a21oi_2 _1324_ (.B1(_0785_),
    .Y(\tokenflow_inst.i78.cg_elem.maj.C ),
    .A2(_0784_),
    .A1(\tokenflow_inst.i2.cg2.maj.C ));
 sg13g2_nor2_1 _1325_ (.A(\tokenflow_inst.i2.cg2.a ),
    .B(\tokenflow_inst.i2.cg2.maj.C ),
    .Y(_0786_));
 sg13g2_a21oi_1 _1326_ (.A1(\tokenflow_inst.i2.cg2.maj.C ),
    .A2(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .Y(_0787_),
    .B1(\tokenflow_inst.i78.d0_elem.inv_chain[0] ));
 sg13g2_nor2_1 _1327_ (.A(_0786_),
    .B(_0787_),
    .Y(\tokenflow_inst.i2.cg2.maj.C ));
 sg13g2_nor2_2 _1328_ (.A(net653),
    .B(\tokenflow_inst.i8.cg_elem.maj.C ),
    .Y(_0309_));
 sg13g2_and2_1 _1329_ (.A(net692),
    .B(\tokenflow_inst.i6.cg_elem.maj.C ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[0] ));
 sg13g2_o21ai_1 _1330_ (.B1(\tokenflow_inst.i2.cg2.a ),
    .Y(_0788_),
    .A1(net577),
    .A2(\tokenflow_inst.i6.d0_elem.inv_chain[0] ));
 sg13g2_nand2_1 _1331_ (.Y(_0789_),
    .A(\tokenflow_inst.i6.cg_elem.maj.C ),
    .B(net577));
 sg13g2_o21ai_1 _1332_ (.B1(_0789_),
    .Y(\tokenflow_inst.i6.cg_elem.maj.C ),
    .A1(_0762_),
    .A2(_0788_));
 sg13g2_nor2_1 _1333_ (.A(net652),
    .B(\tokenflow_inst.i78.cg_elem.maj.C ),
    .Y(_0232_));
 sg13g2_nand2b_1 _1334_ (.Y(_0790_),
    .B(\tokenflow_inst.i78.cg_elem.maj.C ),
    .A_N(\tokenflow_inst.i8.cg_elem.maj.C ));
 sg13g2_a22oi_1 _1335_ (.Y(_0791_),
    .B1(_0790_),
    .B2(\tokenflow_inst.i6.d0_elem.inv_chain[0] ),
    .A2(net606),
    .A1(\tokenflow_inst.i8.cg_elem.maj.C ));
 sg13g2_inv_2 _1336_ (.Y(\tokenflow_inst.i8.cg_elem.maj.C ),
    .A(_0791_));
 sg13g2_a21oi_1 _1337_ (.A1(net534),
    .A2(\tokenflow_inst.i6.ydata[52] ),
    .Y(_0792_),
    .B1(\tokenflow_inst.i6.ydata[0] ));
 sg13g2_nand3_1 _1338_ (.B(\tokenflow_inst.i6.ydata[52] ),
    .C(\tokenflow_inst.i6.ydata[0] ),
    .A(net535),
    .Y(_0793_));
 sg13g2_nand2_1 _1339_ (.Y(_0794_),
    .A(net704),
    .B(_0793_));
 sg13g2_nor2_1 _1340_ (.A(_0792_),
    .B(_0794_),
    .Y(_0233_));
 sg13g2_nand3_1 _1341_ (.B(\tokenflow_inst.i6.ydata[53] ),
    .C(\tokenflow_inst.i6.ydata[1] ),
    .A(net534),
    .Y(_0795_));
 sg13g2_a21oi_1 _1342_ (.A1(net535),
    .A2(\tokenflow_inst.i6.ydata[53] ),
    .Y(_0796_),
    .B1(\tokenflow_inst.i6.ydata[1] ));
 sg13g2_a21o_1 _1343_ (.A2(\tokenflow_inst.i6.ydata[53] ),
    .A1(net535),
    .B1(\tokenflow_inst.i6.ydata[1] ),
    .X(_0797_));
 sg13g2_nand2_1 _1344_ (.Y(_0798_),
    .A(_0795_),
    .B(_0797_));
 sg13g2_o21ai_1 _1345_ (.B1(net704),
    .Y(_0799_),
    .A1(_0793_),
    .A2(_0798_));
 sg13g2_a21oi_1 _1346_ (.A1(_0793_),
    .A2(_0798_),
    .Y(_0244_),
    .B1(_0799_));
 sg13g2_a21oi_1 _1347_ (.A1(net534),
    .A2(\tokenflow_inst.i6.ydata[54] ),
    .Y(_0800_),
    .B1(\tokenflow_inst.i6.ydata[2] ));
 sg13g2_and3_1 _1348_ (.X(_0801_),
    .A(net534),
    .B(\tokenflow_inst.i6.ydata[54] ),
    .C(\tokenflow_inst.i6.ydata[2] ));
 sg13g2_nand3_1 _1349_ (.B(\tokenflow_inst.i6.ydata[54] ),
    .C(\tokenflow_inst.i6.ydata[2] ),
    .A(net534),
    .Y(_0802_));
 sg13g2_nor2_1 _1350_ (.A(_0800_),
    .B(_0801_),
    .Y(_0803_));
 sg13g2_o21ai_1 _1351_ (.B1(_0795_),
    .Y(_0804_),
    .A1(_0793_),
    .A2(_0796_));
 sg13g2_nand2_1 _1352_ (.Y(_0805_),
    .A(_0803_),
    .B(_0804_));
 sg13g2_o21ai_1 _1353_ (.B1(net705),
    .Y(_0806_),
    .A1(_0803_),
    .A2(_0804_));
 sg13g2_nor2b_1 _1354_ (.A(_0806_),
    .B_N(_0805_),
    .Y(_0255_));
 sg13g2_and3_1 _1355_ (.X(_0807_),
    .A(net534),
    .B(\tokenflow_inst.i6.ydata[55] ),
    .C(\tokenflow_inst.i6.ydata[3] ));
 sg13g2_nand3_1 _1356_ (.B(\tokenflow_inst.i6.ydata[55] ),
    .C(\tokenflow_inst.i6.ydata[3] ),
    .A(net534),
    .Y(_0808_));
 sg13g2_a21oi_1 _1357_ (.A1(net534),
    .A2(\tokenflow_inst.i6.ydata[55] ),
    .Y(_0809_),
    .B1(\tokenflow_inst.i6.ydata[3] ));
 sg13g2_or2_1 _1358_ (.X(_0810_),
    .B(_0809_),
    .A(_0807_));
 sg13g2_and2_1 _1359_ (.A(_0802_),
    .B(_0810_),
    .X(_0811_));
 sg13g2_nor4_2 _1360_ (.A(_0800_),
    .B(_0801_),
    .C(_0807_),
    .Y(_0812_),
    .D(_0809_));
 sg13g2_o21ai_1 _1361_ (.B1(net705),
    .Y(_0813_),
    .A1(_0802_),
    .A2(_0810_));
 sg13g2_a221oi_1 _1362_ (.B2(_0804_),
    .C1(_0813_),
    .B1(_0812_),
    .A1(_0805_),
    .Y(_0266_),
    .A2(_0811_));
 sg13g2_a21oi_1 _1363_ (.A1(net536),
    .A2(\tokenflow_inst.i6.ydata[56] ),
    .Y(_0814_),
    .B1(\tokenflow_inst.i6.ydata[4] ));
 sg13g2_nand3_1 _1364_ (.B(\tokenflow_inst.i6.ydata[56] ),
    .C(\tokenflow_inst.i6.ydata[4] ),
    .A(net536),
    .Y(_0815_));
 sg13g2_nand2b_2 _1365_ (.Y(_0816_),
    .B(_0815_),
    .A_N(_0814_));
 sg13g2_o21ai_1 _1366_ (.B1(_0808_),
    .Y(_0817_),
    .A1(_0802_),
    .A2(_0809_));
 sg13g2_a21oi_1 _1367_ (.A1(_0804_),
    .A2(_0812_),
    .Y(_0818_),
    .B1(_0817_));
 sg13g2_a21o_1 _1368_ (.A2(_0812_),
    .A1(_0804_),
    .B1(_0817_),
    .X(_0819_));
 sg13g2_nand2b_1 _1369_ (.Y(_0820_),
    .B(_0819_),
    .A_N(_0816_));
 sg13g2_a21oi_1 _1370_ (.A1(_0816_),
    .A2(_0818_),
    .Y(_0821_),
    .B1(net655));
 sg13g2_and2_1 _1371_ (.A(_0820_),
    .B(_0821_),
    .X(_0277_));
 sg13g2_nand3_1 _1372_ (.B(\tokenflow_inst.i6.ydata[57] ),
    .C(\tokenflow_inst.i6.ydata[5] ),
    .A(net536),
    .Y(_0822_));
 sg13g2_a21oi_1 _1373_ (.A1(net533),
    .A2(\tokenflow_inst.i6.ydata[57] ),
    .Y(_0823_),
    .B1(\tokenflow_inst.i6.ydata[5] ));
 sg13g2_a21o_1 _1374_ (.A2(\tokenflow_inst.i6.ydata[57] ),
    .A1(net533),
    .B1(\tokenflow_inst.i6.ydata[5] ),
    .X(_0824_));
 sg13g2_nand2_1 _1375_ (.Y(_0825_),
    .A(_0822_),
    .B(_0824_));
 sg13g2_and2_1 _1376_ (.A(_0815_),
    .B(_0820_),
    .X(_0826_));
 sg13g2_o21ai_1 _1377_ (.B1(_0815_),
    .Y(_0827_),
    .A1(_0816_),
    .A2(_0818_));
 sg13g2_nand2b_1 _1378_ (.Y(_0828_),
    .B(_0827_),
    .A_N(_0825_));
 sg13g2_nand2_1 _1379_ (.Y(_0829_),
    .A(net702),
    .B(_0828_));
 sg13g2_a21oi_1 _1380_ (.A1(_0825_),
    .A2(_0826_),
    .Y(_0286_),
    .B1(_0829_));
 sg13g2_a21oi_1 _1381_ (.A1(net533),
    .A2(\tokenflow_inst.i6.ydata[58] ),
    .Y(_0830_),
    .B1(\tokenflow_inst.i6.ydata[6] ));
 sg13g2_and3_1 _1382_ (.X(_0831_),
    .A(net533),
    .B(\tokenflow_inst.i6.ydata[6] ),
    .C(\tokenflow_inst.i6.ydata[58] ));
 sg13g2_nand3_1 _1383_ (.B(\tokenflow_inst.i6.ydata[6] ),
    .C(\tokenflow_inst.i6.ydata[58] ),
    .A(net533),
    .Y(_0832_));
 sg13g2_nand2b_1 _1384_ (.Y(_0833_),
    .B(_0832_),
    .A_N(_0830_));
 sg13g2_and2_1 _1385_ (.A(_0822_),
    .B(_0828_),
    .X(_0834_));
 sg13g2_or2_1 _1386_ (.X(_0835_),
    .B(_0834_),
    .A(_0833_));
 sg13g2_nand2_1 _1387_ (.Y(_0836_),
    .A(net702),
    .B(_0835_));
 sg13g2_a21oi_1 _1388_ (.A1(_0833_),
    .A2(_0834_),
    .Y(_0297_),
    .B1(_0836_));
 sg13g2_and3_1 _1389_ (.X(_0837_),
    .A(net533),
    .B(\tokenflow_inst.i6.ydata[59] ),
    .C(\tokenflow_inst.i6.ydata[7] ));
 sg13g2_nand3_1 _1390_ (.B(\tokenflow_inst.i6.ydata[59] ),
    .C(\tokenflow_inst.i6.ydata[7] ),
    .A(net533),
    .Y(_0838_));
 sg13g2_a21oi_1 _1391_ (.A1(net533),
    .A2(\tokenflow_inst.i6.ydata[59] ),
    .Y(_0839_),
    .B1(\tokenflow_inst.i6.ydata[7] ));
 sg13g2_or2_1 _1392_ (.X(_0840_),
    .B(_0839_),
    .A(_0837_));
 sg13g2_nand3_1 _1393_ (.B(_0835_),
    .C(_0840_),
    .A(_0832_),
    .Y(_0841_));
 sg13g2_a21oi_1 _1394_ (.A1(_0832_),
    .A2(_0835_),
    .Y(_0842_),
    .B1(_0840_));
 sg13g2_nor2_1 _1395_ (.A(net655),
    .B(_0842_),
    .Y(_0843_));
 sg13g2_and2_1 _1396_ (.A(_0841_),
    .B(_0843_),
    .X(_0306_));
 sg13g2_nor4_1 _1397_ (.A(_0830_),
    .B(_0831_),
    .C(_0837_),
    .D(_0839_),
    .Y(_0844_));
 sg13g2_nor4_2 _1398_ (.A(_0816_),
    .B(_0825_),
    .C(_0833_),
    .Y(_0845_),
    .D(_0840_));
 sg13g2_o21ai_1 _1399_ (.B1(_0822_),
    .Y(_0846_),
    .A1(_0815_),
    .A2(_0823_));
 sg13g2_o21ai_1 _1400_ (.B1(_0838_),
    .Y(_0847_),
    .A1(_0832_),
    .A2(_0839_));
 sg13g2_a21o_1 _1401_ (.A2(_0846_),
    .A1(_0844_),
    .B1(_0847_),
    .X(_0848_));
 sg13g2_a21oi_1 _1402_ (.A1(_0819_),
    .A2(_0845_),
    .Y(_0849_),
    .B1(_0848_));
 sg13g2_a21o_1 _1403_ (.A2(_0845_),
    .A1(_0819_),
    .B1(_0848_),
    .X(_0850_));
 sg13g2_a21oi_1 _1404_ (.A1(net530),
    .A2(\tokenflow_inst.i6.ydata[60] ),
    .Y(_0851_),
    .B1(\tokenflow_inst.i6.ydata[8] ));
 sg13g2_nand3_1 _1405_ (.B(\tokenflow_inst.i6.ydata[8] ),
    .C(\tokenflow_inst.i6.ydata[60] ),
    .A(net530),
    .Y(_0852_));
 sg13g2_nand2b_1 _1406_ (.Y(_0853_),
    .B(_0852_),
    .A_N(_0851_));
 sg13g2_nand2b_1 _1407_ (.Y(_0854_),
    .B(_0850_),
    .A_N(_0853_));
 sg13g2_nand2_1 _1408_ (.Y(_0855_),
    .A(net678),
    .B(_0854_));
 sg13g2_a21oi_1 _1409_ (.A1(_0849_),
    .A2(_0853_),
    .Y(_0307_),
    .B1(_0855_));
 sg13g2_nand3_1 _1410_ (.B(\tokenflow_inst.i6.ydata[61] ),
    .C(\tokenflow_inst.i6.ydata[9] ),
    .A(net530),
    .Y(_0856_));
 sg13g2_a21oi_1 _1411_ (.A1(net530),
    .A2(\tokenflow_inst.i6.ydata[61] ),
    .Y(_0857_),
    .B1(\tokenflow_inst.i6.ydata[9] ));
 sg13g2_a21o_1 _1412_ (.A2(\tokenflow_inst.i6.ydata[61] ),
    .A1(net530),
    .B1(\tokenflow_inst.i6.ydata[9] ),
    .X(_0858_));
 sg13g2_nand2_1 _1413_ (.Y(_0859_),
    .A(_0856_),
    .B(_0858_));
 sg13g2_xnor2_1 _1414_ (.Y(_0860_),
    .A(_0852_),
    .B(_0859_));
 sg13g2_nor2_1 _1415_ (.A(_0853_),
    .B(_0859_),
    .Y(_0861_));
 sg13g2_nor2_1 _1416_ (.A(_0854_),
    .B(_0859_),
    .Y(_0862_));
 sg13g2_a221oi_1 _1417_ (.B2(_0850_),
    .C1(net656),
    .B1(_0861_),
    .A1(_0854_),
    .Y(_0308_),
    .A2(_0860_));
 sg13g2_a21oi_1 _1418_ (.A1(net529),
    .A2(\tokenflow_inst.i6.ydata[62] ),
    .Y(_0863_),
    .B1(\tokenflow_inst.i6.ydata[10] ));
 sg13g2_and3_1 _1419_ (.X(_0864_),
    .A(net529),
    .B(\tokenflow_inst.i6.ydata[10] ),
    .C(\tokenflow_inst.i6.ydata[62] ));
 sg13g2_nand3_1 _1420_ (.B(\tokenflow_inst.i6.ydata[10] ),
    .C(\tokenflow_inst.i6.ydata[62] ),
    .A(net528),
    .Y(_0865_));
 sg13g2_nor2_1 _1421_ (.A(_0863_),
    .B(_0864_),
    .Y(_0866_));
 sg13g2_o21ai_1 _1422_ (.B1(_0856_),
    .Y(_0867_),
    .A1(_0852_),
    .A2(_0857_));
 sg13g2_or3_1 _1423_ (.A(_0862_),
    .B(_0866_),
    .C(_0867_),
    .X(_0868_));
 sg13g2_o21ai_1 _1424_ (.B1(_0866_),
    .Y(_0391_),
    .A1(_0862_),
    .A2(_0867_));
 sg13g2_and3_1 _1425_ (.X(_0234_),
    .A(net679),
    .B(_0868_),
    .C(_0391_));
 sg13g2_and3_1 _1426_ (.X(_0392_),
    .A(net528),
    .B(\tokenflow_inst.i6.ydata[63] ),
    .C(\tokenflow_inst.i6.ydata[11] ));
 sg13g2_nand3_1 _1427_ (.B(\tokenflow_inst.i6.ydata[63] ),
    .C(\tokenflow_inst.i6.ydata[11] ),
    .A(net528),
    .Y(_0393_));
 sg13g2_a21oi_2 _1428_ (.B1(\tokenflow_inst.i6.ydata[11] ),
    .Y(_0394_),
    .A2(\tokenflow_inst.i6.ydata[63] ),
    .A1(net528));
 sg13g2_nor2_1 _1429_ (.A(_0392_),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_nand2_1 _1430_ (.Y(_0396_),
    .A(_0865_),
    .B(_0391_));
 sg13g2_o21ai_1 _1431_ (.B1(net672),
    .Y(_0397_),
    .A1(_0395_),
    .A2(_0396_));
 sg13g2_a21oi_1 _1432_ (.A1(_0395_),
    .A2(_0396_),
    .Y(_0235_),
    .B1(_0397_));
 sg13g2_a21oi_1 _1433_ (.A1(net528),
    .A2(\tokenflow_inst.i6.ydata[64] ),
    .Y(_0398_),
    .B1(\tokenflow_inst.i6.ydata[12] ));
 sg13g2_nand3_1 _1434_ (.B(\tokenflow_inst.i6.ydata[12] ),
    .C(\tokenflow_inst.i6.ydata[64] ),
    .A(net528),
    .Y(_0399_));
 sg13g2_nand2b_2 _1435_ (.Y(_0400_),
    .B(_0399_),
    .A_N(_0398_));
 sg13g2_o21ai_1 _1436_ (.B1(_0393_),
    .Y(_0401_),
    .A1(_0865_),
    .A2(_0394_));
 sg13g2_nor4_2 _1437_ (.A(_0863_),
    .B(_0864_),
    .C(_0392_),
    .Y(_0402_),
    .D(_0394_));
 sg13g2_a21oi_1 _1438_ (.A1(_0867_),
    .A2(_0402_),
    .Y(_0403_),
    .B1(_0401_));
 sg13g2_a21o_1 _1439_ (.A2(_0402_),
    .A1(_0867_),
    .B1(_0401_),
    .X(_0404_));
 sg13g2_nand3_1 _1440_ (.B(_0861_),
    .C(_0402_),
    .A(_0850_),
    .Y(_0405_));
 sg13g2_and3_1 _1441_ (.X(_0406_),
    .A(_0400_),
    .B(_0403_),
    .C(_0405_));
 sg13g2_a21oi_2 _1442_ (.B1(_0400_),
    .Y(_0407_),
    .A2(_0405_),
    .A1(_0403_));
 sg13g2_nor3_1 _1443_ (.A(net656),
    .B(_0406_),
    .C(_0407_),
    .Y(_0236_));
 sg13g2_nand3_1 _1444_ (.B(\tokenflow_inst.i6.ydata[65] ),
    .C(\tokenflow_inst.i6.ydata[13] ),
    .A(net528),
    .Y(_0408_));
 sg13g2_a21o_1 _1445_ (.A2(\tokenflow_inst.i6.ydata[65] ),
    .A1(net528),
    .B1(\tokenflow_inst.i6.ydata[13] ),
    .X(_0409_));
 sg13g2_nand2_2 _1446_ (.Y(_0410_),
    .A(_0408_),
    .B(_0409_));
 sg13g2_nand2_1 _1447_ (.Y(_0411_),
    .A(_0399_),
    .B(_0410_));
 sg13g2_nor2_1 _1448_ (.A(_0407_),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_and3_1 _1449_ (.X(_0413_),
    .A(_0407_),
    .B(_0408_),
    .C(_0409_));
 sg13g2_o21ai_1 _1450_ (.B1(net672),
    .Y(_0414_),
    .A1(_0399_),
    .A2(_0410_));
 sg13g2_nor3_1 _1451_ (.A(_0412_),
    .B(_0413_),
    .C(_0414_),
    .Y(_0237_));
 sg13g2_a21oi_1 _1452_ (.A1(net530),
    .A2(\tokenflow_inst.i6.ydata[66] ),
    .Y(_0415_),
    .B1(\tokenflow_inst.i6.ydata[14] ));
 sg13g2_nand3_1 _1453_ (.B(\tokenflow_inst.i6.ydata[14] ),
    .C(\tokenflow_inst.i6.ydata[66] ),
    .A(net530),
    .Y(_0416_));
 sg13g2_nand2b_1 _1454_ (.Y(_0417_),
    .B(_0416_),
    .A_N(_0415_));
 sg13g2_inv_1 _1455_ (.Y(_0418_),
    .A(_0417_));
 sg13g2_o21ai_1 _1456_ (.B1(_0408_),
    .Y(_0419_),
    .A1(_0399_),
    .A2(_0410_));
 sg13g2_nor3_1 _1457_ (.A(_0413_),
    .B(_0418_),
    .C(_0419_),
    .Y(_0420_));
 sg13g2_o21ai_1 _1458_ (.B1(_0418_),
    .Y(_0421_),
    .A1(_0413_),
    .A2(_0419_));
 sg13g2_nand2_1 _1459_ (.Y(_0422_),
    .A(net672),
    .B(_0421_));
 sg13g2_nor2_1 _1460_ (.A(_0420_),
    .B(_0422_),
    .Y(_0238_));
 sg13g2_a21oi_1 _1461_ (.A1(net530),
    .A2(\tokenflow_inst.i6.ydata[67] ),
    .Y(_0423_),
    .B1(\tokenflow_inst.i6.ydata[15] ));
 sg13g2_nand3_1 _1462_ (.B(\tokenflow_inst.i6.ydata[67] ),
    .C(\tokenflow_inst.i6.ydata[15] ),
    .A(net531),
    .Y(_0424_));
 sg13g2_nand2b_1 _1463_ (.Y(_0425_),
    .B(_0424_),
    .A_N(_0423_));
 sg13g2_and3_1 _1464_ (.X(_0426_),
    .A(_0416_),
    .B(_0421_),
    .C(_0425_));
 sg13g2_a21oi_1 _1465_ (.A1(_0416_),
    .A2(_0421_),
    .Y(_0427_),
    .B1(_0425_));
 sg13g2_nor3_1 _1466_ (.A(net651),
    .B(_0426_),
    .C(_0427_),
    .Y(_0239_));
 sg13g2_a21oi_1 _1467_ (.A1(net537),
    .A2(\tokenflow_inst.i6.ydata[68] ),
    .Y(_0428_),
    .B1(\tokenflow_inst.i6.ydata[16] ));
 sg13g2_nand3_1 _1468_ (.B(\tokenflow_inst.i6.ydata[16] ),
    .C(\tokenflow_inst.i6.ydata[68] ),
    .A(net537),
    .Y(_0429_));
 sg13g2_nor2b_1 _1469_ (.A(_0428_),
    .B_N(_0429_),
    .Y(_0430_));
 sg13g2_nand2b_1 _1470_ (.Y(_0431_),
    .B(_0429_),
    .A_N(_0428_));
 sg13g2_nor2_1 _1471_ (.A(_0417_),
    .B(_0425_),
    .Y(_0432_));
 sg13g2_nor4_2 _1472_ (.A(_0400_),
    .B(_0410_),
    .C(_0417_),
    .Y(_0433_),
    .D(_0425_));
 sg13g2_o21ai_1 _1473_ (.B1(_0424_),
    .Y(_0434_),
    .A1(_0416_),
    .A2(_0423_));
 sg13g2_a221oi_1 _1474_ (.B2(_0404_),
    .C1(_0434_),
    .B1(_0433_),
    .A1(_0419_),
    .Y(_0435_),
    .A2(_0432_));
 sg13g2_nand3_1 _1475_ (.B(_0402_),
    .C(_0433_),
    .A(_0861_),
    .Y(_0436_));
 sg13g2_o21ai_1 _1476_ (.B1(_0435_),
    .Y(_0437_),
    .A1(_0849_),
    .A2(_0436_));
 sg13g2_or2_1 _1477_ (.X(_0438_),
    .B(_0437_),
    .A(_0430_));
 sg13g2_nand2_1 _1478_ (.Y(_0439_),
    .A(_0430_),
    .B(_0437_));
 sg13g2_and3_1 _1479_ (.X(_0240_),
    .A(net681),
    .B(_0438_),
    .C(_0439_));
 sg13g2_a21oi_1 _1480_ (.A1(net537),
    .A2(\tokenflow_inst.i6.ydata[69] ),
    .Y(_0440_),
    .B1(\tokenflow_inst.i6.ydata[17] ));
 sg13g2_nand3_1 _1481_ (.B(\tokenflow_inst.i6.ydata[17] ),
    .C(\tokenflow_inst.i6.ydata[69] ),
    .A(net537),
    .Y(_0441_));
 sg13g2_nand2b_1 _1482_ (.Y(_0442_),
    .B(_0441_),
    .A_N(_0440_));
 sg13g2_nand3_1 _1483_ (.B(_0439_),
    .C(_0442_),
    .A(_0429_),
    .Y(_0443_));
 sg13g2_a21o_1 _1484_ (.A2(_0439_),
    .A1(_0429_),
    .B1(_0442_),
    .X(_0444_));
 sg13g2_and3_1 _1485_ (.X(_0241_),
    .A(net699),
    .B(_0443_),
    .C(_0444_));
 sg13g2_a21oi_1 _1486_ (.A1(net537),
    .A2(\tokenflow_inst.i6.ydata[70] ),
    .Y(_0445_),
    .B1(\tokenflow_inst.i6.ydata[18] ));
 sg13g2_nand3_1 _1487_ (.B(\tokenflow_inst.i6.ydata[18] ),
    .C(\tokenflow_inst.i6.ydata[70] ),
    .A(net537),
    .Y(_0446_));
 sg13g2_nand2b_2 _1488_ (.Y(_0447_),
    .B(_0446_),
    .A_N(_0445_));
 sg13g2_nand3_1 _1489_ (.B(_0444_),
    .C(_0447_),
    .A(_0441_),
    .Y(_0448_));
 sg13g2_a21o_1 _1490_ (.A2(_0444_),
    .A1(_0441_),
    .B1(_0447_),
    .X(_0449_));
 sg13g2_and3_1 _1491_ (.X(_0242_),
    .A(net699),
    .B(_0448_),
    .C(_0449_));
 sg13g2_and2_1 _1492_ (.A(net537),
    .B(\tokenflow_inst.i6.ydata[71] ),
    .X(_0450_));
 sg13g2_nor2_1 _1493_ (.A(\tokenflow_inst.i6.ydata[19] ),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_xnor2_1 _1494_ (.Y(_0452_),
    .A(\tokenflow_inst.i6.ydata[19] ),
    .B(_0450_));
 sg13g2_nand3_1 _1495_ (.B(_0449_),
    .C(_0452_),
    .A(_0446_),
    .Y(_0453_));
 sg13g2_a21o_1 _1496_ (.A2(_0449_),
    .A1(_0446_),
    .B1(_0452_),
    .X(_0454_));
 sg13g2_and3_1 _1497_ (.X(_0243_),
    .A(net700),
    .B(_0453_),
    .C(_0454_));
 sg13g2_nor2_1 _1498_ (.A(_0447_),
    .B(_0452_),
    .Y(_0455_));
 sg13g2_nor4_2 _1499_ (.A(_0431_),
    .B(_0442_),
    .C(_0447_),
    .Y(_0456_),
    .D(_0452_));
 sg13g2_o21ai_1 _1500_ (.B1(_0441_),
    .Y(_0457_),
    .A1(_0429_),
    .A2(_0440_));
 sg13g2_a22oi_1 _1501_ (.Y(_0458_),
    .B1(_0455_),
    .B2(_0457_),
    .A2(_0450_),
    .A1(\tokenflow_inst.i6.ydata[19] ));
 sg13g2_o21ai_1 _1502_ (.B1(_0458_),
    .Y(_0459_),
    .A1(_0446_),
    .A2(_0451_));
 sg13g2_a21oi_2 _1503_ (.B1(_0459_),
    .Y(_0460_),
    .A2(_0456_),
    .A1(_0437_));
 sg13g2_a21o_1 _1504_ (.A2(_0456_),
    .A1(_0437_),
    .B1(_0459_),
    .X(_0461_));
 sg13g2_a21oi_1 _1505_ (.A1(net531),
    .A2(\tokenflow_inst.i6.ydata[72] ),
    .Y(_0462_),
    .B1(\tokenflow_inst.i6.ydata[20] ));
 sg13g2_nand3_1 _1506_ (.B(\tokenflow_inst.i6.ydata[20] ),
    .C(\tokenflow_inst.i6.ydata[72] ),
    .A(net531),
    .Y(_0463_));
 sg13g2_nand2b_1 _1507_ (.Y(_0464_),
    .B(_0463_),
    .A_N(_0462_));
 sg13g2_o21ai_1 _1508_ (.B1(net681),
    .Y(_0465_),
    .A1(_0460_),
    .A2(_0464_));
 sg13g2_a21oi_1 _1509_ (.A1(_0460_),
    .A2(_0464_),
    .Y(_0245_),
    .B1(_0465_));
 sg13g2_nand2_1 _1510_ (.Y(_0466_),
    .A(net531),
    .B(\tokenflow_inst.i6.ydata[73] ));
 sg13g2_xnor2_1 _1511_ (.Y(_0467_),
    .A(_0739_),
    .B(_0466_));
 sg13g2_and2_1 _1512_ (.A(_0463_),
    .B(_0467_),
    .X(_0468_));
 sg13g2_o21ai_1 _1513_ (.B1(_0468_),
    .Y(_0469_),
    .A1(_0460_),
    .A2(_0464_));
 sg13g2_nor2_1 _1514_ (.A(_0464_),
    .B(_0467_),
    .Y(_0470_));
 sg13g2_nand2_1 _1515_ (.Y(_0471_),
    .A(_0461_),
    .B(_0470_));
 sg13g2_or2_1 _1516_ (.X(_0472_),
    .B(_0467_),
    .A(_0463_));
 sg13g2_and4_1 _1517_ (.A(net680),
    .B(_0469_),
    .C(_0471_),
    .D(_0472_),
    .X(_0246_));
 sg13g2_a21oi_1 _1518_ (.A1(net529),
    .A2(\tokenflow_inst.i6.ydata[74] ),
    .Y(_0473_),
    .B1(\tokenflow_inst.i6.ydata[22] ));
 sg13g2_nand3_1 _1519_ (.B(\tokenflow_inst.i6.ydata[22] ),
    .C(\tokenflow_inst.i6.ydata[74] ),
    .A(net529),
    .Y(_0474_));
 sg13g2_nand2b_1 _1520_ (.Y(_0475_),
    .B(_0474_),
    .A_N(_0473_));
 sg13g2_o21ai_1 _1521_ (.B1(_0472_),
    .Y(_0476_),
    .A1(_0739_),
    .A2(_0466_));
 sg13g2_a21oi_2 _1522_ (.B1(_0476_),
    .Y(_0477_),
    .A2(_0470_),
    .A1(_0461_));
 sg13g2_o21ai_1 _1523_ (.B1(net680),
    .Y(_0478_),
    .A1(_0475_),
    .A2(_0477_));
 sg13g2_a21oi_1 _1524_ (.A1(_0475_),
    .A2(_0477_),
    .Y(_0247_),
    .B1(_0478_));
 sg13g2_nand3_1 _1525_ (.B(\tokenflow_inst.i6.ydata[23] ),
    .C(\tokenflow_inst.i6.ydata[75] ),
    .A(net532),
    .Y(_0479_));
 sg13g2_a21oi_1 _1526_ (.A1(net532),
    .A2(\tokenflow_inst.i6.ydata[75] ),
    .Y(_0480_),
    .B1(\tokenflow_inst.i6.ydata[23] ));
 sg13g2_a21o_1 _1527_ (.A2(\tokenflow_inst.i6.ydata[75] ),
    .A1(net532),
    .B1(\tokenflow_inst.i6.ydata[23] ),
    .X(_0481_));
 sg13g2_nand2_1 _1528_ (.Y(_0482_),
    .A(_0479_),
    .B(_0481_));
 sg13g2_inv_1 _1529_ (.Y(_0483_),
    .A(_0482_));
 sg13g2_o21ai_1 _1530_ (.B1(_0474_),
    .Y(_0484_),
    .A1(_0475_),
    .A2(_0477_));
 sg13g2_o21ai_1 _1531_ (.B1(net675),
    .Y(_0485_),
    .A1(_0483_),
    .A2(_0484_));
 sg13g2_a21oi_1 _1532_ (.A1(_0483_),
    .A2(_0484_),
    .Y(_0248_),
    .B1(_0485_));
 sg13g2_nor2_1 _1533_ (.A(_0475_),
    .B(_0482_),
    .Y(_0486_));
 sg13g2_nand2_1 _1534_ (.Y(_0487_),
    .A(_0470_),
    .B(_0486_));
 sg13g2_o21ai_1 _1535_ (.B1(_0479_),
    .Y(_0488_),
    .A1(_0474_),
    .A2(_0480_));
 sg13g2_a21oi_1 _1536_ (.A1(_0476_),
    .A2(_0486_),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_o21ai_1 _1537_ (.B1(_0489_),
    .Y(_0490_),
    .A1(_0460_),
    .A2(_0487_));
 sg13g2_and3_1 _1538_ (.X(_0491_),
    .A(net529),
    .B(\tokenflow_inst.i6.ydata[76] ),
    .C(\tokenflow_inst.i6.ydata[24] ));
 sg13g2_a21o_1 _1539_ (.A2(\tokenflow_inst.i6.ydata[76] ),
    .A1(net529),
    .B1(\tokenflow_inst.i6.ydata[24] ),
    .X(_0492_));
 sg13g2_nand2b_1 _1540_ (.Y(_0493_),
    .B(_0492_),
    .A_N(_0491_));
 sg13g2_nor2b_1 _1541_ (.A(_0490_),
    .B_N(_0493_),
    .Y(_0494_));
 sg13g2_nor2b_1 _1542_ (.A(_0493_),
    .B_N(_0490_),
    .Y(_0495_));
 sg13g2_nor3_1 _1543_ (.A(net651),
    .B(_0494_),
    .C(_0495_),
    .Y(_0249_));
 sg13g2_nand2_1 _1544_ (.Y(_0496_),
    .A(net529),
    .B(\tokenflow_inst.i6.ydata[77] ));
 sg13g2_xor2_1 _1545_ (.B(_0496_),
    .A(\tokenflow_inst.i6.ydata[25] ),
    .X(_0497_));
 sg13g2_a21oi_1 _1546_ (.A1(_0490_),
    .A2(_0492_),
    .Y(_0498_),
    .B1(_0491_));
 sg13g2_o21ai_1 _1547_ (.B1(net674),
    .Y(_0499_),
    .A1(_0497_),
    .A2(_0498_));
 sg13g2_a21oi_1 _1548_ (.A1(_0497_),
    .A2(_0498_),
    .Y(_0250_),
    .B1(_0499_));
 sg13g2_and2_1 _1549_ (.A(net703),
    .B(\tokenflow_inst.i6.ydata[27] ),
    .X(_0251_));
 sg13g2_and2_1 _1550_ (.A(net694),
    .B(\tokenflow_inst.i6.ydata[28] ),
    .X(_0252_));
 sg13g2_and2_1 _1551_ (.A(net694),
    .B(\tokenflow_inst.i6.ydata[29] ),
    .X(_0253_));
 sg13g2_and2_1 _1552_ (.A(net693),
    .B(\tokenflow_inst.i6.ydata[30] ),
    .X(_0254_));
 sg13g2_and2_1 _1553_ (.A(net693),
    .B(\tokenflow_inst.i6.ydata[31] ),
    .X(_0256_));
 sg13g2_and2_1 _1554_ (.A(net692),
    .B(\tokenflow_inst.i6.ydata[32] ),
    .X(_0257_));
 sg13g2_and2_1 _1555_ (.A(net695),
    .B(\tokenflow_inst.i6.ydata[33] ),
    .X(_0258_));
 sg13g2_and2_1 _1556_ (.A(net689),
    .B(\tokenflow_inst.i6.ydata[34] ),
    .X(_0259_));
 sg13g2_and2_1 _1557_ (.A(net696),
    .B(\tokenflow_inst.i6.ydata[35] ),
    .X(_0260_));
 sg13g2_and2_1 _1558_ (.A(net669),
    .B(\tokenflow_inst.i6.ydata[36] ),
    .X(_0261_));
 sg13g2_and2_1 _1559_ (.A(net666),
    .B(\tokenflow_inst.i6.ydata[37] ),
    .X(_0262_));
 sg13g2_and2_1 _1560_ (.A(net660),
    .B(\tokenflow_inst.i6.ydata[38] ),
    .X(_0263_));
 sg13g2_and2_1 _1561_ (.A(net658),
    .B(\tokenflow_inst.i6.ydata[39] ),
    .X(_0264_));
 sg13g2_and2_1 _1562_ (.A(net661),
    .B(\tokenflow_inst.i6.ydata[40] ),
    .X(_0265_));
 sg13g2_and2_1 _1563_ (.A(net661),
    .B(\tokenflow_inst.i6.ydata[41] ),
    .X(_0267_));
 sg13g2_and2_1 _1564_ (.A(net669),
    .B(\tokenflow_inst.i6.ydata[42] ),
    .X(_0268_));
 sg13g2_and2_1 _1565_ (.A(net668),
    .B(\tokenflow_inst.i6.ydata[43] ),
    .X(_0269_));
 sg13g2_and2_1 _1566_ (.A(net689),
    .B(\tokenflow_inst.i6.ydata[44] ),
    .X(_0270_));
 sg13g2_and2_1 _1567_ (.A(net684),
    .B(\tokenflow_inst.i6.ydata[45] ),
    .X(_0271_));
 sg13g2_and2_1 _1568_ (.A(net689),
    .B(\tokenflow_inst.i6.ydata[46] ),
    .X(_0272_));
 sg13g2_and2_1 _1569_ (.A(net688),
    .B(\tokenflow_inst.i6.ydata[47] ),
    .X(_0273_));
 sg13g2_and2_1 _1570_ (.A(net663),
    .B(\tokenflow_inst.i6.ydata[48] ),
    .X(_0274_));
 sg13g2_and2_1 _1571_ (.A(net663),
    .B(\tokenflow_inst.i6.ydata[49] ),
    .X(_0275_));
 sg13g2_and2_1 _1572_ (.A(net661),
    .B(\tokenflow_inst.i6.ydata[50] ),
    .X(_0276_));
 sg13g2_and2_1 _1573_ (.A(net662),
    .B(\tokenflow_inst.i6.ydata[51] ),
    .X(_0278_));
 sg13g2_and2_1 _1574_ (.A(net704),
    .B(\tokenflow_inst.i6.ydata[52] ),
    .X(_0279_));
 sg13g2_and2_1 _1575_ (.A(net704),
    .B(\tokenflow_inst.i6.ydata[53] ),
    .X(_0280_));
 sg13g2_and2_1 _1576_ (.A(net705),
    .B(\tokenflow_inst.i6.ydata[54] ),
    .X(_0281_));
 sg13g2_and2_1 _1577_ (.A(net702),
    .B(\tokenflow_inst.i6.ydata[55] ),
    .X(_0282_));
 sg13g2_and2_1 _1578_ (.A(net703),
    .B(\tokenflow_inst.i6.ydata[56] ),
    .X(_0283_));
 sg13g2_and2_1 _1579_ (.A(net703),
    .B(\tokenflow_inst.i6.ydata[57] ),
    .X(_0284_));
 sg13g2_and2_1 _1580_ (.A(net697),
    .B(\tokenflow_inst.i6.ydata[58] ),
    .X(_0285_));
 sg13g2_and2_1 _1581_ (.A(net698),
    .B(\tokenflow_inst.i6.ydata[59] ),
    .X(_0287_));
 sg13g2_and2_1 _1582_ (.A(net678),
    .B(\tokenflow_inst.i6.ydata[60] ),
    .X(_0288_));
 sg13g2_and2_1 _1583_ (.A(net670),
    .B(\tokenflow_inst.i6.ydata[61] ),
    .X(_0289_));
 sg13g2_and2_1 _1584_ (.A(net663),
    .B(\tokenflow_inst.i6.ydata[62] ),
    .X(_0290_));
 sg13g2_and2_1 _1585_ (.A(net673),
    .B(\tokenflow_inst.i6.ydata[63] ),
    .X(_0291_));
 sg13g2_and2_1 _1586_ (.A(net673),
    .B(\tokenflow_inst.i6.ydata[64] ),
    .X(_0292_));
 sg13g2_and2_1 _1587_ (.A(net672),
    .B(\tokenflow_inst.i6.ydata[65] ),
    .X(_0293_));
 sg13g2_and2_1 _1588_ (.A(net679),
    .B(\tokenflow_inst.i6.ydata[66] ),
    .X(_0294_));
 sg13g2_and2_1 _1589_ (.A(net678),
    .B(\tokenflow_inst.i6.ydata[67] ),
    .X(_0295_));
 sg13g2_and2_1 _1590_ (.A(net699),
    .B(\tokenflow_inst.i6.ydata[68] ),
    .X(_0296_));
 sg13g2_and2_1 _1591_ (.A(net697),
    .B(\tokenflow_inst.i6.ydata[69] ),
    .X(_0298_));
 sg13g2_and2_1 _1592_ (.A(net699),
    .B(\tokenflow_inst.i6.ydata[70] ),
    .X(_0299_));
 sg13g2_and2_1 _1593_ (.A(net700),
    .B(\tokenflow_inst.i6.ydata[71] ),
    .X(_0300_));
 sg13g2_and2_1 _1594_ (.A(net680),
    .B(\tokenflow_inst.i6.ydata[72] ),
    .X(_0301_));
 sg13g2_and2_1 _1595_ (.A(net680),
    .B(\tokenflow_inst.i6.ydata[73] ),
    .X(_0302_));
 sg13g2_and2_1 _1596_ (.A(net676),
    .B(\tokenflow_inst.i6.ydata[74] ),
    .X(_0303_));
 sg13g2_and2_1 _1597_ (.A(net675),
    .B(\tokenflow_inst.i6.ydata[75] ),
    .X(_0304_));
 sg13g2_and2_1 _1598_ (.A(net676),
    .B(\tokenflow_inst.i6.ydata[76] ),
    .X(_0305_));
 sg13g2_and2_1 _1599_ (.A(net706),
    .B(\tokenflow_inst.i3.ydata[0] ),
    .X(_0079_));
 sg13g2_and2_1 _1600_ (.A(net704),
    .B(\tokenflow_inst.i3.ydata[1] ),
    .X(_0090_));
 sg13g2_and2_1 _1601_ (.A(net706),
    .B(\tokenflow_inst.i3.ydata[2] ),
    .X(_0101_));
 sg13g2_and2_1 _1602_ (.A(net706),
    .B(\tokenflow_inst.i3.ydata[3] ),
    .X(_0112_));
 sg13g2_and2_1 _1603_ (.A(net706),
    .B(\tokenflow_inst.i3.ydata[4] ),
    .X(_0123_));
 sg13g2_and2_1 _1604_ (.A(net702),
    .B(\tokenflow_inst.i3.ydata[5] ),
    .X(_0134_));
 sg13g2_and2_1 _1605_ (.A(net697),
    .B(\tokenflow_inst.i3.ydata[6] ),
    .X(_0145_));
 sg13g2_and2_1 _1606_ (.A(net698),
    .B(\tokenflow_inst.i3.ydata[7] ),
    .X(_0154_));
 sg13g2_and2_1 _1607_ (.A(net678),
    .B(\tokenflow_inst.i3.ydata[8] ),
    .X(_0155_));
 sg13g2_and2_1 _1608_ (.A(net678),
    .B(\tokenflow_inst.i3.ydata[9] ),
    .X(_0156_));
 sg13g2_and2_1 _1609_ (.A(net670),
    .B(\tokenflow_inst.i3.ydata[10] ),
    .X(_0080_));
 sg13g2_and2_1 _1610_ (.A(net672),
    .B(\tokenflow_inst.i3.ydata[11] ),
    .X(_0081_));
 sg13g2_and2_1 _1611_ (.A(net673),
    .B(\tokenflow_inst.i3.ydata[12] ),
    .X(_0082_));
 sg13g2_and2_1 _1612_ (.A(net672),
    .B(\tokenflow_inst.i3.ydata[13] ),
    .X(_0083_));
 sg13g2_and2_1 _1613_ (.A(net680),
    .B(\tokenflow_inst.i3.ydata[14] ),
    .X(_0084_));
 sg13g2_and2_1 _1614_ (.A(net678),
    .B(\tokenflow_inst.i3.ydata[15] ),
    .X(_0085_));
 sg13g2_and2_1 _1615_ (.A(net699),
    .B(\tokenflow_inst.i3.ydata[16] ),
    .X(_0086_));
 sg13g2_and2_1 _1616_ (.A(net699),
    .B(\tokenflow_inst.i3.ydata[17] ),
    .X(_0087_));
 sg13g2_and2_1 _1617_ (.A(net700),
    .B(\tokenflow_inst.i3.ydata[18] ),
    .X(_0088_));
 sg13g2_and2_1 _1618_ (.A(net701),
    .B(\tokenflow_inst.i3.ydata[19] ),
    .X(_0089_));
 sg13g2_and2_1 _1619_ (.A(net681),
    .B(\tokenflow_inst.i3.ydata[20] ),
    .X(_0091_));
 sg13g2_and2_1 _1620_ (.A(net681),
    .B(\tokenflow_inst.i3.ydata[21] ),
    .X(_0092_));
 sg13g2_and2_1 _1621_ (.A(net680),
    .B(\tokenflow_inst.i3.ydata[22] ),
    .X(_0093_));
 sg13g2_and2_1 _1622_ (.A(net675),
    .B(\tokenflow_inst.i3.ydata[23] ),
    .X(_0094_));
 sg13g2_and2_1 _1623_ (.A(net674),
    .B(\tokenflow_inst.i3.ydata[24] ),
    .X(_0095_));
 sg13g2_and2_1 _1624_ (.A(net674),
    .B(\tokenflow_inst.i3.ydata[25] ),
    .X(_0096_));
 sg13g2_and2_1 _1625_ (.A(net694),
    .B(\tokenflow_inst.i3.ydata[26] ),
    .X(_0097_));
 sg13g2_and2_1 _1626_ (.A(net694),
    .B(\tokenflow_inst.i3.ydata[27] ),
    .X(_0098_));
 sg13g2_and2_1 _1627_ (.A(net694),
    .B(\tokenflow_inst.i3.ydata[28] ),
    .X(_0099_));
 sg13g2_and2_1 _1628_ (.A(net693),
    .B(\tokenflow_inst.i3.ydata[29] ),
    .X(_0100_));
 sg13g2_and2_1 _1629_ (.A(net693),
    .B(\tokenflow_inst.i3.ydata[30] ),
    .X(_0102_));
 sg13g2_and2_1 _1630_ (.A(net693),
    .B(\tokenflow_inst.i3.ydata[31] ),
    .X(_0103_));
 sg13g2_and2_1 _1631_ (.A(net692),
    .B(\tokenflow_inst.i3.ydata[32] ),
    .X(_0104_));
 sg13g2_and2_1 _1632_ (.A(net692),
    .B(\tokenflow_inst.i3.ydata[33] ),
    .X(_0105_));
 sg13g2_and2_1 _1633_ (.A(net689),
    .B(\tokenflow_inst.i3.ydata[34] ),
    .X(_0106_));
 sg13g2_and2_1 _1634_ (.A(net688),
    .B(\tokenflow_inst.i3.ydata[35] ),
    .X(_0107_));
 sg13g2_and2_1 _1635_ (.A(net669),
    .B(\tokenflow_inst.i3.ydata[36] ),
    .X(_0108_));
 sg13g2_and2_1 _1636_ (.A(net660),
    .B(\tokenflow_inst.i3.ydata[37] ),
    .X(_0109_));
 sg13g2_and2_1 _1637_ (.A(net663),
    .B(\tokenflow_inst.i3.ydata[38] ),
    .X(_0110_));
 sg13g2_and2_1 _1638_ (.A(net658),
    .B(\tokenflow_inst.i3.ydata[39] ),
    .X(_0111_));
 sg13g2_and2_1 _1639_ (.A(net661),
    .B(\tokenflow_inst.i3.ydata[40] ),
    .X(_0113_));
 sg13g2_and2_1 _1640_ (.A(net669),
    .B(\tokenflow_inst.i3.ydata[41] ),
    .X(_0114_));
 sg13g2_and2_1 _1641_ (.A(net671),
    .B(\tokenflow_inst.i3.ydata[42] ),
    .X(_0115_));
 sg13g2_and2_1 _1642_ (.A(net670),
    .B(\tokenflow_inst.i3.ydata[43] ),
    .X(_0116_));
 sg13g2_and2_1 _1643_ (.A(net688),
    .B(\tokenflow_inst.i3.ydata[44] ),
    .X(_0117_));
 sg13g2_and2_1 _1644_ (.A(net688),
    .B(\tokenflow_inst.i3.ydata[45] ),
    .X(_0118_));
 sg13g2_and2_1 _1645_ (.A(net670),
    .B(\tokenflow_inst.i3.ydata[46] ),
    .X(_0119_));
 sg13g2_and2_1 _1646_ (.A(net688),
    .B(\tokenflow_inst.i3.ydata[47] ),
    .X(_0120_));
 sg13g2_and2_1 _1647_ (.A(net663),
    .B(\tokenflow_inst.i3.ydata[48] ),
    .X(_0121_));
 sg13g2_and2_1 _1648_ (.A(net663),
    .B(\tokenflow_inst.i3.ydata[49] ),
    .X(_0122_));
 sg13g2_and2_1 _1649_ (.A(net661),
    .B(\tokenflow_inst.i3.ydata[50] ),
    .X(_0124_));
 sg13g2_and2_1 _1650_ (.A(net662),
    .B(\tokenflow_inst.i3.ydata[51] ),
    .X(_0125_));
 sg13g2_and2_1 _1651_ (.A(net704),
    .B(\tokenflow_inst.i3.ydata[52] ),
    .X(_0126_));
 sg13g2_and2_1 _1652_ (.A(net704),
    .B(\tokenflow_inst.i3.ydata[53] ),
    .X(_0127_));
 sg13g2_and2_1 _1653_ (.A(net705),
    .B(\tokenflow_inst.i3.ydata[54] ),
    .X(_0128_));
 sg13g2_and2_1 _1654_ (.A(net705),
    .B(\tokenflow_inst.i3.ydata[55] ),
    .X(_0129_));
 sg13g2_and2_1 _1655_ (.A(net703),
    .B(\tokenflow_inst.i3.ydata[56] ),
    .X(_0130_));
 sg13g2_and2_1 _1656_ (.A(net703),
    .B(\tokenflow_inst.i3.ydata[57] ),
    .X(_0131_));
 sg13g2_and2_1 _1657_ (.A(net692),
    .B(\tokenflow_inst.i3.ydata[58] ),
    .X(_0132_));
 sg13g2_and2_1 _1658_ (.A(net689),
    .B(\tokenflow_inst.i3.ydata[59] ),
    .X(_0133_));
 sg13g2_and2_1 _1659_ (.A(net697),
    .B(\tokenflow_inst.i3.ydata[60] ),
    .X(_0135_));
 sg13g2_and2_1 _1660_ (.A(net670),
    .B(\tokenflow_inst.i3.ydata[61] ),
    .X(_0136_));
 sg13g2_and2_1 _1661_ (.A(net663),
    .B(\tokenflow_inst.i3.ydata[62] ),
    .X(_0137_));
 sg13g2_and2_1 _1662_ (.A(net661),
    .B(\tokenflow_inst.i3.ydata[63] ),
    .X(_0138_));
 sg13g2_and2_1 _1663_ (.A(net673),
    .B(\tokenflow_inst.i3.ydata[64] ),
    .X(_0139_));
 sg13g2_and2_1 _1664_ (.A(net673),
    .B(\tokenflow_inst.i3.ydata[65] ),
    .X(_0140_));
 sg13g2_and2_1 _1665_ (.A(net675),
    .B(\tokenflow_inst.i3.ydata[66] ),
    .X(_0141_));
 sg13g2_and2_1 _1666_ (.A(net678),
    .B(\tokenflow_inst.i3.ydata[67] ),
    .X(_0142_));
 sg13g2_and2_1 _1667_ (.A(net697),
    .B(\tokenflow_inst.i3.ydata[68] ),
    .X(_0143_));
 sg13g2_and2_1 _1668_ (.A(net697),
    .B(\tokenflow_inst.i3.ydata[69] ),
    .X(_0144_));
 sg13g2_and2_1 _1669_ (.A(net700),
    .B(\tokenflow_inst.i3.ydata[70] ),
    .X(_0146_));
 sg13g2_and2_1 _1670_ (.A(net700),
    .B(\tokenflow_inst.i3.ydata[71] ),
    .X(_0147_));
 sg13g2_and2_1 _1671_ (.A(net680),
    .B(\tokenflow_inst.i3.ydata[72] ),
    .X(_0148_));
 sg13g2_and2_1 _1672_ (.A(net681),
    .B(\tokenflow_inst.i3.ydata[73] ),
    .X(_0149_));
 sg13g2_and2_1 _1673_ (.A(net675),
    .B(\tokenflow_inst.i3.ydata[74] ),
    .X(_0150_));
 sg13g2_and2_1 _1674_ (.A(net675),
    .B(\tokenflow_inst.i3.ydata[75] ),
    .X(_0151_));
 sg13g2_and2_1 _1675_ (.A(net674),
    .B(\tokenflow_inst.i3.ydata[76] ),
    .X(_0152_));
 sg13g2_and2_1 _1676_ (.A(net673),
    .B(\tokenflow_inst.i3.ydata[77] ),
    .X(_0153_));
 sg13g2_and2_2 _1677_ (.A(\tokenflow_inst.ii3.i.ydata[0] ),
    .B(net648),
    .X(_0047_));
 sg13g2_a21o_1 _1678_ (.A2(net643),
    .A1(\tokenflow_inst.i78.ydata[0] ),
    .B1(_0047_),
    .X(_0000_));
 sg13g2_and2_2 _1679_ (.A(\tokenflow_inst.ii3.i.ydata[1] ),
    .B(net647),
    .X(_0048_));
 sg13g2_a21o_1 _1680_ (.A2(net645),
    .A1(\tokenflow_inst.i78.ydata[1] ),
    .B1(_0048_),
    .X(_0011_));
 sg13g2_and2_2 _1681_ (.A(\tokenflow_inst.ii3.i.ydata[2] ),
    .B(net647),
    .X(_0500_));
 sg13g2_a21o_1 _1682_ (.A2(net643),
    .A1(\tokenflow_inst.i78.ydata[2] ),
    .B1(_0500_),
    .X(_0022_));
 sg13g2_and2_2 _1683_ (.A(\tokenflow_inst.ii3.i.ydata[3] ),
    .B(net647),
    .X(_0501_));
 sg13g2_a21o_1 _1684_ (.A2(net643),
    .A1(\tokenflow_inst.i78.ydata[3] ),
    .B1(_0501_),
    .X(_0033_));
 sg13g2_and2_2 _1685_ (.A(\tokenflow_inst.ii3.i.ydata[4] ),
    .B(net647),
    .X(_0502_));
 sg13g2_a21o_1 _1686_ (.A2(net643),
    .A1(\tokenflow_inst.i78.ydata[4] ),
    .B1(_0502_),
    .X(_0044_));
 sg13g2_and2_1 _1687_ (.A(\tokenflow_inst.ii3.i.ydata[5] ),
    .B(net647),
    .X(_0503_));
 sg13g2_a21o_1 _1688_ (.A2(net643),
    .A1(\tokenflow_inst.i78.ydata[5] ),
    .B1(_0503_),
    .X(_0055_));
 sg13g2_and2_1 _1689_ (.A(\tokenflow_inst.ii3.i.ydata[6] ),
    .B(net647),
    .X(_0504_));
 sg13g2_a21o_1 _1690_ (.A2(net642),
    .A1(\tokenflow_inst.i78.ydata[6] ),
    .B1(_0504_),
    .X(_0066_));
 sg13g2_nor3_2 _1691_ (.A(net652),
    .B(_0740_),
    .C(\tokenflow_inst.i2.cg1.maj.C ),
    .Y(_0505_));
 sg13g2_a21o_1 _1692_ (.A2(net642),
    .A1(\tokenflow_inst.i78.ydata[7] ),
    .B1(_0505_),
    .X(_0075_));
 sg13g2_nor3_2 _1693_ (.A(net654),
    .B(_0741_),
    .C(net649),
    .Y(_0506_));
 sg13g2_a21o_1 _1694_ (.A2(net640),
    .A1(\tokenflow_inst.i78.ydata[8] ),
    .B1(_0506_),
    .X(_0076_));
 sg13g2_and2_1 _1695_ (.A(\tokenflow_inst.ii3.i.ydata[9] ),
    .B(net648),
    .X(_0507_));
 sg13g2_a21o_1 _1696_ (.A2(net634),
    .A1(\tokenflow_inst.i78.ydata[9] ),
    .B1(_0507_),
    .X(_0077_));
 sg13g2_nor3_2 _1697_ (.A(net651),
    .B(_0742_),
    .C(net649),
    .Y(_0508_));
 sg13g2_a21o_1 _1698_ (.A2(net635),
    .A1(\tokenflow_inst.i78.ydata[10] ),
    .B1(_0508_),
    .X(_0001_));
 sg13g2_and2_1 _1699_ (.A(\tokenflow_inst.ii3.i.ydata[11] ),
    .B(net646),
    .X(_0509_));
 sg13g2_a21o_1 _1700_ (.A2(net635),
    .A1(\tokenflow_inst.i78.ydata[11] ),
    .B1(_0509_),
    .X(_0002_));
 sg13g2_and2_1 _1701_ (.A(\tokenflow_inst.ii3.i.ydata[12] ),
    .B(net646),
    .X(_0510_));
 sg13g2_a21o_1 _1702_ (.A2(net633),
    .A1(\tokenflow_inst.i78.ydata[12] ),
    .B1(_0510_),
    .X(_0003_));
 sg13g2_nor3_2 _1703_ (.A(net650),
    .B(_0743_),
    .C(net649),
    .Y(_0511_));
 sg13g2_a21o_1 _1704_ (.A2(net636),
    .A1(\tokenflow_inst.i78.ydata[13] ),
    .B1(_0511_),
    .X(_0004_));
 sg13g2_and2_2 _1705_ (.A(\tokenflow_inst.ii3.i.ydata[14] ),
    .B(net646),
    .X(_0512_));
 sg13g2_a21o_1 _1706_ (.A2(net636),
    .A1(\tokenflow_inst.i78.ydata[14] ),
    .B1(_0512_),
    .X(_0005_));
 sg13g2_and2_2 _1707_ (.A(\tokenflow_inst.ii3.i.ydata[15] ),
    .B(net648),
    .X(_0513_));
 sg13g2_a21o_1 _1708_ (.A2(net638),
    .A1(\tokenflow_inst.i78.ydata[15] ),
    .B1(_0513_),
    .X(_0006_));
 sg13g2_and2_2 _1709_ (.A(\tokenflow_inst.ii3.i.ydata[16] ),
    .B(net648),
    .X(_0514_));
 sg13g2_a21o_1 _1710_ (.A2(net638),
    .A1(\tokenflow_inst.i78.ydata[16] ),
    .B1(_0514_),
    .X(_0007_));
 sg13g2_and2_2 _1711_ (.A(\tokenflow_inst.ii3.i.ydata[17] ),
    .B(net647),
    .X(_0515_));
 sg13g2_a21o_1 _1712_ (.A2(net644),
    .A1(\tokenflow_inst.i78.ydata[17] ),
    .B1(_0515_),
    .X(_0008_));
 sg13g2_and2_2 _1713_ (.A(\tokenflow_inst.ii3.i.ydata[18] ),
    .B(net647),
    .X(_0516_));
 sg13g2_a21o_1 _1714_ (.A2(net644),
    .A1(\tokenflow_inst.i78.ydata[18] ),
    .B1(_0516_),
    .X(_0009_));
 sg13g2_nor3_2 _1715_ (.A(net654),
    .B(_0744_),
    .C(net649),
    .Y(_0517_));
 sg13g2_a21o_1 _1716_ (.A2(net644),
    .A1(\tokenflow_inst.i78.ydata[19] ),
    .B1(_0517_),
    .X(_0010_));
 sg13g2_and2_2 _1717_ (.A(\tokenflow_inst.ii3.i.ydata[20] ),
    .B(net646),
    .X(_0518_));
 sg13g2_a21o_1 _1718_ (.A2(net638),
    .A1(\tokenflow_inst.i78.ydata[20] ),
    .B1(_0518_),
    .X(_0012_));
 sg13g2_and2_2 _1719_ (.A(\tokenflow_inst.ii3.i.ydata[21] ),
    .B(net646),
    .X(_0519_));
 sg13g2_a21o_1 _1720_ (.A2(net638),
    .A1(\tokenflow_inst.i78.ydata[21] ),
    .B1(_0519_),
    .X(_0013_));
 sg13g2_and2_2 _1721_ (.A(\tokenflow_inst.ii3.i.ydata[22] ),
    .B(net646),
    .X(_0520_));
 sg13g2_a21o_1 _1722_ (.A2(net636),
    .A1(\tokenflow_inst.i78.ydata[22] ),
    .B1(_0520_),
    .X(_0014_));
 sg13g2_and2_2 _1723_ (.A(\tokenflow_inst.ii3.i.ydata[23] ),
    .B(net646),
    .X(_0521_));
 sg13g2_a21o_1 _1724_ (.A2(net637),
    .A1(\tokenflow_inst.i78.ydata[23] ),
    .B1(_0521_),
    .X(_0015_));
 sg13g2_and2_2 _1725_ (.A(\tokenflow_inst.ii3.i.ydata[24] ),
    .B(net646),
    .X(_0045_));
 sg13g2_a21o_1 _1726_ (.A2(net637),
    .A1(\tokenflow_inst.i78.ydata[24] ),
    .B1(_0045_),
    .X(_0016_));
 sg13g2_nor3_2 _1727_ (.A(net650),
    .B(_0745_),
    .C(net649),
    .Y(_0046_));
 sg13g2_a21o_1 _1728_ (.A2(net636),
    .A1(\tokenflow_inst.i78.ydata[25] ),
    .B1(_0046_),
    .X(_0017_));
 sg13g2_a21o_1 _1729_ (.A2(net641),
    .A1(\tokenflow_inst.i78.ydata[26] ),
    .B1(_0047_),
    .X(_0018_));
 sg13g2_a21o_1 _1730_ (.A2(net642),
    .A1(\tokenflow_inst.i78.ydata[27] ),
    .B1(_0048_),
    .X(_0019_));
 sg13g2_a21o_1 _1731_ (.A2(net641),
    .A1(\tokenflow_inst.i78.ydata[28] ),
    .B1(_0500_),
    .X(_0020_));
 sg13g2_a21o_1 _1732_ (.A2(net641),
    .A1(\tokenflow_inst.i78.ydata[29] ),
    .B1(_0501_),
    .X(_0021_));
 sg13g2_a21o_1 _1733_ (.A2(net641),
    .A1(\tokenflow_inst.i78.ydata[30] ),
    .B1(_0502_),
    .X(_0023_));
 sg13g2_a21o_1 _1734_ (.A2(net641),
    .A1(\tokenflow_inst.i78.ydata[31] ),
    .B1(_0503_),
    .X(_0024_));
 sg13g2_a21o_1 _1735_ (.A2(net641),
    .A1(\tokenflow_inst.i78.ydata[32] ),
    .B1(_0504_),
    .X(_0025_));
 sg13g2_a21o_1 _1736_ (.A2(net640),
    .A1(\tokenflow_inst.i78.ydata[33] ),
    .B1(_0505_),
    .X(_0026_));
 sg13g2_a21o_1 _1737_ (.A2(net640),
    .A1(\tokenflow_inst.i78.ydata[34] ),
    .B1(_0506_),
    .X(_0027_));
 sg13g2_a21o_1 _1738_ (.A2(net634),
    .A1(\tokenflow_inst.i78.ydata[35] ),
    .B1(_0507_),
    .X(_0028_));
 sg13g2_a21o_1 _1739_ (.A2(net634),
    .A1(\tokenflow_inst.i78.ydata[36] ),
    .B1(_0508_),
    .X(_0029_));
 sg13g2_a21o_1 _1740_ (.A2(net633),
    .A1(\tokenflow_inst.i78.ydata[37] ),
    .B1(_0509_),
    .X(_0030_));
 sg13g2_a21o_1 _1741_ (.A2(net633),
    .A1(\tokenflow_inst.i78.ydata[38] ),
    .B1(_0510_),
    .X(_0031_));
 sg13g2_a21o_1 _1742_ (.A2(net633),
    .A1(\tokenflow_inst.i78.ydata[39] ),
    .B1(_0511_),
    .X(_0032_));
 sg13g2_a21o_1 _1743_ (.A2(net633),
    .A1(\tokenflow_inst.i78.ydata[40] ),
    .B1(_0512_),
    .X(_0034_));
 sg13g2_a21o_1 _1744_ (.A2(net634),
    .A1(\tokenflow_inst.i78.ydata[41] ),
    .B1(_0513_),
    .X(_0035_));
 sg13g2_a21o_1 _1745_ (.A2(net634),
    .A1(\tokenflow_inst.i78.ydata[42] ),
    .B1(_0514_),
    .X(_0036_));
 sg13g2_a21o_1 _1746_ (.A2(net640),
    .A1(\tokenflow_inst.i78.ydata[43] ),
    .B1(_0515_),
    .X(_0037_));
 sg13g2_a21o_1 _1747_ (.A2(net640),
    .A1(\tokenflow_inst.i78.ydata[44] ),
    .B1(_0516_),
    .X(_0038_));
 sg13g2_a21o_1 _1748_ (.A2(net640),
    .A1(\tokenflow_inst.i78.ydata[45] ),
    .B1(_0517_),
    .X(_0039_));
 sg13g2_a21o_1 _1749_ (.A2(net634),
    .A1(\tokenflow_inst.i78.ydata[46] ),
    .B1(_0518_),
    .X(_0040_));
 sg13g2_a21o_1 _1750_ (.A2(net634),
    .A1(\tokenflow_inst.i78.ydata[47] ),
    .B1(_0519_),
    .X(_0041_));
 sg13g2_a21o_1 _1751_ (.A2(net633),
    .A1(\tokenflow_inst.i78.ydata[48] ),
    .B1(_0520_),
    .X(_0042_));
 sg13g2_a21o_1 _1752_ (.A2(net633),
    .A1(\tokenflow_inst.i78.ydata[49] ),
    .B1(_0521_),
    .X(_0043_));
 sg13g2_a21o_1 _1753_ (.A2(net643),
    .A1(\tokenflow_inst.i78.ydata[54] ),
    .B1(_0500_),
    .X(_0049_));
 sg13g2_a21o_1 _1754_ (.A2(net644),
    .A1(\tokenflow_inst.i78.ydata[55] ),
    .B1(_0501_),
    .X(_0050_));
 sg13g2_a21o_1 _1755_ (.A2(net643),
    .A1(\tokenflow_inst.i78.ydata[56] ),
    .B1(_0502_),
    .X(_0051_));
 sg13g2_a21o_1 _1756_ (.A2(net643),
    .A1(\tokenflow_inst.i78.ydata[57] ),
    .B1(_0503_),
    .X(_0052_));
 sg13g2_a21o_1 _1757_ (.A2(net641),
    .A1(\tokenflow_inst.i78.ydata[58] ),
    .B1(_0504_),
    .X(_0053_));
 sg13g2_a21o_1 _1758_ (.A2(net642),
    .A1(\tokenflow_inst.i78.ydata[59] ),
    .B1(_0505_),
    .X(_0054_));
 sg13g2_a21o_1 _1759_ (.A2(net640),
    .A1(\tokenflow_inst.i78.ydata[60] ),
    .B1(_0506_),
    .X(_0056_));
 sg13g2_a21o_1 _1760_ (.A2(net642),
    .A1(\tokenflow_inst.i78.ydata[61] ),
    .B1(_0507_),
    .X(_0057_));
 sg13g2_a21o_1 _1761_ (.A2(net634),
    .A1(\tokenflow_inst.i78.ydata[62] ),
    .B1(_0508_),
    .X(_0058_));
 sg13g2_a21o_1 _1762_ (.A2(net633),
    .A1(\tokenflow_inst.i78.ydata[63] ),
    .B1(_0509_),
    .X(_0059_));
 sg13g2_a21o_1 _1763_ (.A2(net635),
    .A1(\tokenflow_inst.i78.ydata[64] ),
    .B1(_0510_),
    .X(_0060_));
 sg13g2_a21o_1 _1764_ (.A2(net636),
    .A1(\tokenflow_inst.i78.ydata[65] ),
    .B1(_0511_),
    .X(_0061_));
 sg13g2_a21o_1 _1765_ (.A2(net636),
    .A1(\tokenflow_inst.i78.ydata[66] ),
    .B1(_0512_),
    .X(_0062_));
 sg13g2_a21o_1 _1766_ (.A2(net639),
    .A1(\tokenflow_inst.i78.ydata[67] ),
    .B1(_0513_),
    .X(_0063_));
 sg13g2_a21o_1 _1767_ (.A2(net638),
    .A1(\tokenflow_inst.i78.ydata[68] ),
    .B1(_0514_),
    .X(_0064_));
 sg13g2_a21o_1 _1768_ (.A2(net644),
    .A1(\tokenflow_inst.i78.ydata[69] ),
    .B1(_0515_),
    .X(_0065_));
 sg13g2_a21o_1 _1769_ (.A2(net644),
    .A1(\tokenflow_inst.i78.ydata[70] ),
    .B1(_0516_),
    .X(_0067_));
 sg13g2_a21o_1 _1770_ (.A2(net644),
    .A1(\tokenflow_inst.i78.ydata[71] ),
    .B1(_0517_),
    .X(_0068_));
 sg13g2_a21o_1 _1771_ (.A2(net638),
    .A1(\tokenflow_inst.i78.ydata[72] ),
    .B1(_0518_),
    .X(_0069_));
 sg13g2_a21o_1 _1772_ (.A2(net639),
    .A1(\tokenflow_inst.i78.ydata[73] ),
    .B1(_0519_),
    .X(_0070_));
 sg13g2_a21o_1 _1773_ (.A2(net636),
    .A1(\tokenflow_inst.i78.ydata[74] ),
    .B1(_0520_),
    .X(_0071_));
 sg13g2_a21o_1 _1774_ (.A2(net637),
    .A1(\tokenflow_inst.i78.ydata[75] ),
    .B1(_0521_),
    .X(_0072_));
 sg13g2_a21o_1 _1775_ (.A2(net637),
    .A1(\tokenflow_inst.i78.ydata[76] ),
    .B1(_0045_),
    .X(_0073_));
 sg13g2_a21o_1 _1776_ (.A2(net636),
    .A1(\tokenflow_inst.i78.ydata[77] ),
    .B1(_0046_),
    .X(_0074_));
 sg13g2_and2_1 _1777_ (.A(net690),
    .B(\tokenflow_inst.ii2.ydata[0] ),
    .X(_0364_));
 sg13g2_and2_1 _1778_ (.A(net691),
    .B(\tokenflow_inst.ii2.ydata[1] ),
    .X(_0375_));
 sg13g2_and2_1 _1779_ (.A(net691),
    .B(\tokenflow_inst.ii2.ydata[2] ),
    .X(_0382_));
 sg13g2_and2_1 _1780_ (.A(net696),
    .B(\tokenflow_inst.ii2.ydata[3] ),
    .X(_0383_));
 sg13g2_and2_1 _1781_ (.A(net690),
    .B(\tokenflow_inst.ii2.ydata[4] ),
    .X(_0384_));
 sg13g2_and2_1 _1782_ (.A(net690),
    .B(\tokenflow_inst.ii2.ydata[5] ),
    .X(_0385_));
 sg13g2_and2_1 _1783_ (.A(net685),
    .B(\tokenflow_inst.ii2.ydata[6] ),
    .X(_0386_));
 sg13g2_and2_1 _1784_ (.A(net685),
    .B(\tokenflow_inst.ii2.ydata[7] ),
    .X(_0387_));
 sg13g2_and2_1 _1785_ (.A(net683),
    .B(\tokenflow_inst.ii2.ydata[8] ),
    .X(_0388_));
 sg13g2_and2_1 _1786_ (.A(net667),
    .B(\tokenflow_inst.ii2.ydata[9] ),
    .X(_0389_));
 sg13g2_and2_1 _1787_ (.A(net666),
    .B(\tokenflow_inst.ii2.ydata[10] ),
    .X(_0365_));
 sg13g2_and2_1 _1788_ (.A(net666),
    .B(\tokenflow_inst.ii2.ydata[11] ),
    .X(_0366_));
 sg13g2_and2_1 _1789_ (.A(net659),
    .B(\tokenflow_inst.ii2.ydata[12] ),
    .X(_0367_));
 sg13g2_and2_1 _1790_ (.A(net659),
    .B(\tokenflow_inst.ii2.ydata[13] ),
    .X(_0368_));
 sg13g2_and2_1 _1791_ (.A(net659),
    .B(\tokenflow_inst.ii2.ydata[14] ),
    .X(_0369_));
 sg13g2_and2_1 _1792_ (.A(net668),
    .B(\tokenflow_inst.ii2.ydata[15] ),
    .X(_0370_));
 sg13g2_and2_1 _1793_ (.A(net667),
    .B(\tokenflow_inst.ii2.ydata[16] ),
    .X(_0371_));
 sg13g2_and2_1 _1794_ (.A(net683),
    .B(\tokenflow_inst.ii2.ydata[17] ),
    .X(_0372_));
 sg13g2_and2_1 _1795_ (.A(net683),
    .B(\tokenflow_inst.ii2.ydata[18] ),
    .X(_0373_));
 sg13g2_and2_1 _1796_ (.A(net684),
    .B(\tokenflow_inst.ii2.ydata[19] ),
    .X(_0374_));
 sg13g2_and2_1 _1797_ (.A(net667),
    .B(\tokenflow_inst.ii2.ydata[20] ),
    .X(_0376_));
 sg13g2_and2_1 _1798_ (.A(net668),
    .B(\tokenflow_inst.ii2.ydata[21] ),
    .X(_0377_));
 sg13g2_and2_1 _1799_ (.A(net657),
    .B(\tokenflow_inst.ii2.ydata[22] ),
    .X(_0378_));
 sg13g2_and2_1 _1800_ (.A(net657),
    .B(\tokenflow_inst.ii2.ydata[23] ),
    .X(_0379_));
 sg13g2_and2_1 _1801_ (.A(net658),
    .B(\tokenflow_inst.ii2.ydata[24] ),
    .X(_0380_));
 sg13g2_and2_1 _1802_ (.A(net657),
    .B(\tokenflow_inst.ii2.ydata[25] ),
    .X(_0381_));
 sg13g2_and2_1 _1803_ (.A(net690),
    .B(\tokenflow_inst.ii1.ydata[0] ),
    .X(_0337_));
 sg13g2_and2_1 _1804_ (.A(net691),
    .B(\tokenflow_inst.ii1.ydata[1] ),
    .X(_0348_));
 sg13g2_and2_1 _1805_ (.A(net691),
    .B(\tokenflow_inst.ii1.ydata[2] ),
    .X(_0355_));
 sg13g2_and2_1 _1806_ (.A(net691),
    .B(\tokenflow_inst.ii1.ydata[3] ),
    .X(_0356_));
 sg13g2_and2_1 _1807_ (.A(net690),
    .B(\tokenflow_inst.ii1.ydata[4] ),
    .X(_0357_));
 sg13g2_and2_1 _1808_ (.A(net690),
    .B(\tokenflow_inst.ii1.ydata[5] ),
    .X(_0358_));
 sg13g2_and2_1 _1809_ (.A(net685),
    .B(\tokenflow_inst.ii1.ydata[6] ),
    .X(_0359_));
 sg13g2_and2_1 _1810_ (.A(net685),
    .B(\tokenflow_inst.ii1.ydata[7] ),
    .X(_0360_));
 sg13g2_and2_1 _1811_ (.A(net683),
    .B(\tokenflow_inst.ii1.ydata[8] ),
    .X(_0361_));
 sg13g2_and2_1 _1812_ (.A(net667),
    .B(\tokenflow_inst.ii1.ydata[9] ),
    .X(_0362_));
 sg13g2_and2_1 _1813_ (.A(net666),
    .B(\tokenflow_inst.ii1.ydata[10] ),
    .X(_0338_));
 sg13g2_and2_1 _1814_ (.A(net666),
    .B(\tokenflow_inst.ii1.ydata[11] ),
    .X(_0339_));
 sg13g2_and2_1 _1815_ (.A(net659),
    .B(\tokenflow_inst.ii1.ydata[12] ),
    .X(_0340_));
 sg13g2_and2_1 _1816_ (.A(net659),
    .B(\tokenflow_inst.ii1.ydata[13] ),
    .X(_0341_));
 sg13g2_and2_1 _1817_ (.A(net659),
    .B(\tokenflow_inst.ii1.ydata[14] ),
    .X(_0342_));
 sg13g2_and2_1 _1818_ (.A(net660),
    .B(\tokenflow_inst.ii1.ydata[15] ),
    .X(_0343_));
 sg13g2_and2_1 _1819_ (.A(net667),
    .B(\tokenflow_inst.ii1.ydata[16] ),
    .X(_0344_));
 sg13g2_and2_1 _1820_ (.A(net683),
    .B(\tokenflow_inst.ii1.ydata[17] ),
    .X(_0345_));
 sg13g2_and2_1 _1821_ (.A(net683),
    .B(\tokenflow_inst.ii1.ydata[18] ),
    .X(_0346_));
 sg13g2_and2_1 _1822_ (.A(net684),
    .B(\tokenflow_inst.ii1.ydata[19] ),
    .X(_0347_));
 sg13g2_and2_1 _1823_ (.A(net667),
    .B(\tokenflow_inst.ii1.ydata[20] ),
    .X(_0349_));
 sg13g2_and2_1 _1824_ (.A(net666),
    .B(\tokenflow_inst.ii1.ydata[21] ),
    .X(_0350_));
 sg13g2_and2_1 _1825_ (.A(net657),
    .B(\tokenflow_inst.ii1.ydata[22] ),
    .X(_0351_));
 sg13g2_and2_1 _1826_ (.A(net657),
    .B(\tokenflow_inst.ii1.ydata[23] ),
    .X(_0352_));
 sg13g2_and2_1 _1827_ (.A(net658),
    .B(\tokenflow_inst.ii1.ydata[24] ),
    .X(_0353_));
 sg13g2_and2_1 _1828_ (.A(net657),
    .B(\tokenflow_inst.ii1.ydata[25] ),
    .X(_0354_));
 sg13g2_nor2_1 _1829_ (.A(net652),
    .B(\tokenflow_inst.ii3.i.ydata[0] ),
    .Y(_0310_));
 sg13g2_xnor2_1 _1830_ (.Y(_0522_),
    .A(\tokenflow_inst.ii3.i.ydata[0] ),
    .B(\tokenflow_inst.ii3.i.ydata[1] ));
 sg13g2_nor2_1 _1831_ (.A(net652),
    .B(_0522_),
    .Y(_0321_));
 sg13g2_a21oi_1 _1832_ (.A1(\tokenflow_inst.ii3.i.ydata[0] ),
    .A2(\tokenflow_inst.ii3.i.ydata[1] ),
    .Y(_0523_),
    .B1(\tokenflow_inst.ii3.i.ydata[2] ));
 sg13g2_nand3_1 _1833_ (.B(\tokenflow_inst.ii3.i.ydata[1] ),
    .C(\tokenflow_inst.ii3.i.ydata[2] ),
    .A(\tokenflow_inst.ii3.i.ydata[0] ),
    .Y(_0524_));
 sg13g2_nand2_1 _1834_ (.Y(_0525_),
    .A(net691),
    .B(_0524_));
 sg13g2_nor2_1 _1835_ (.A(_0523_),
    .B(_0525_),
    .Y(_0328_));
 sg13g2_nor2b_1 _1836_ (.A(\tokenflow_inst.ii3.i.ydata[3] ),
    .B_N(_0524_),
    .Y(_0526_));
 sg13g2_and4_1 _1837_ (.A(\tokenflow_inst.ii3.i.ydata[0] ),
    .B(\tokenflow_inst.ii3.i.ydata[1] ),
    .C(\tokenflow_inst.ii3.i.ydata[2] ),
    .D(\tokenflow_inst.ii3.i.ydata[3] ),
    .X(_0527_));
 sg13g2_nor3_1 _1838_ (.A(net652),
    .B(_0526_),
    .C(_0527_),
    .Y(_0329_));
 sg13g2_nor2_1 _1839_ (.A(\tokenflow_inst.ii3.i.ydata[4] ),
    .B(_0527_),
    .Y(_0528_));
 sg13g2_and2_1 _1840_ (.A(\tokenflow_inst.ii3.i.ydata[4] ),
    .B(_0527_),
    .X(_0529_));
 sg13g2_nor3_1 _1841_ (.A(net652),
    .B(_0528_),
    .C(_0529_),
    .Y(_0330_));
 sg13g2_o21ai_1 _1842_ (.B1(net690),
    .Y(_0530_),
    .A1(\tokenflow_inst.ii3.i.ydata[5] ),
    .A2(_0529_));
 sg13g2_a21oi_1 _1843_ (.A1(\tokenflow_inst.ii3.i.ydata[5] ),
    .A2(_0529_),
    .Y(_0331_),
    .B1(_0530_));
 sg13g2_a21oi_1 _1844_ (.A1(\tokenflow_inst.ii3.i.ydata[5] ),
    .A2(_0529_),
    .Y(_0531_),
    .B1(\tokenflow_inst.ii3.i.ydata[6] ));
 sg13g2_nand4_1 _1845_ (.B(\tokenflow_inst.ii3.i.ydata[5] ),
    .C(\tokenflow_inst.ii3.i.ydata[6] ),
    .A(\tokenflow_inst.ii3.i.ydata[4] ),
    .Y(_0532_),
    .D(_0527_));
 sg13g2_nand2_1 _1846_ (.Y(_0533_),
    .A(net685),
    .B(_0532_));
 sg13g2_nor2_1 _1847_ (.A(_0531_),
    .B(_0533_),
    .Y(_0332_));
 sg13g2_o21ai_1 _1848_ (.B1(net685),
    .Y(_0534_),
    .A1(_0740_),
    .A2(_0532_));
 sg13g2_a21oi_1 _1849_ (.A1(_0740_),
    .A2(_0532_),
    .Y(_0333_),
    .B1(_0534_));
 sg13g2_o21ai_1 _1850_ (.B1(_0741_),
    .Y(_0535_),
    .A1(_0740_),
    .A2(_0532_));
 sg13g2_nor3_2 _1851_ (.A(_0740_),
    .B(_0741_),
    .C(_0532_),
    .Y(_0536_));
 sg13g2_nand2_1 _1852_ (.Y(_0537_),
    .A(net685),
    .B(_0535_));
 sg13g2_nor2_1 _1853_ (.A(_0536_),
    .B(_0537_),
    .Y(_0334_));
 sg13g2_or2_1 _1854_ (.X(_0538_),
    .B(_0536_),
    .A(\tokenflow_inst.ii3.i.ydata[9] ));
 sg13g2_nand2_1 _1855_ (.Y(_0539_),
    .A(\tokenflow_inst.ii3.i.ydata[9] ),
    .B(_0536_));
 sg13g2_and3_1 _1856_ (.X(_0335_),
    .A(net666),
    .B(_0538_),
    .C(_0539_));
 sg13g2_nand3_1 _1857_ (.B(\tokenflow_inst.ii3.i.ydata[10] ),
    .C(_0536_),
    .A(\tokenflow_inst.ii3.i.ydata[9] ),
    .Y(_0540_));
 sg13g2_nand2_1 _1858_ (.Y(_0541_),
    .A(net666),
    .B(_0540_));
 sg13g2_a21oi_1 _1859_ (.A1(_0742_),
    .A2(_0539_),
    .Y(_0311_),
    .B1(_0541_));
 sg13g2_nor2b_1 _1860_ (.A(\tokenflow_inst.ii3.i.ydata[11] ),
    .B_N(_0540_),
    .Y(_0542_));
 sg13g2_and4_1 _1861_ (.A(\tokenflow_inst.ii3.i.ydata[9] ),
    .B(\tokenflow_inst.ii3.i.ydata[10] ),
    .C(\tokenflow_inst.ii3.i.ydata[11] ),
    .D(_0536_),
    .X(_0543_));
 sg13g2_nor3_1 _1862_ (.A(net650),
    .B(_0542_),
    .C(_0543_),
    .Y(_0312_));
 sg13g2_or2_1 _1863_ (.X(_0544_),
    .B(_0543_),
    .A(\tokenflow_inst.ii3.i.ydata[12] ));
 sg13g2_nand2_2 _1864_ (.Y(_0545_),
    .A(\tokenflow_inst.ii3.i.ydata[12] ),
    .B(_0543_));
 sg13g2_and3_1 _1865_ (.X(_0313_),
    .A(net659),
    .B(_0544_),
    .C(_0545_));
 sg13g2_nor2_2 _1866_ (.A(_0743_),
    .B(_0545_),
    .Y(_0546_));
 sg13g2_a21oi_1 _1867_ (.A1(_0743_),
    .A2(_0545_),
    .Y(_0547_),
    .B1(net650));
 sg13g2_nor2b_1 _1868_ (.A(_0546_),
    .B_N(_0547_),
    .Y(_0314_));
 sg13g2_o21ai_1 _1869_ (.B1(net659),
    .Y(_0548_),
    .A1(\tokenflow_inst.ii3.i.ydata[14] ),
    .A2(_0546_));
 sg13g2_a21oi_1 _1870_ (.A1(\tokenflow_inst.ii3.i.ydata[14] ),
    .A2(_0546_),
    .Y(_0315_),
    .B1(_0548_));
 sg13g2_a21oi_1 _1871_ (.A1(\tokenflow_inst.ii3.i.ydata[14] ),
    .A2(_0546_),
    .Y(_0549_),
    .B1(\tokenflow_inst.ii3.i.ydata[15] ));
 sg13g2_nand2_1 _1872_ (.Y(_0550_),
    .A(\tokenflow_inst.ii3.i.ydata[14] ),
    .B(\tokenflow_inst.ii3.i.ydata[15] ));
 sg13g2_nor3_2 _1873_ (.A(_0743_),
    .B(_0545_),
    .C(_0550_),
    .Y(_0551_));
 sg13g2_nor3_1 _1874_ (.A(net650),
    .B(_0549_),
    .C(_0551_),
    .Y(_0316_));
 sg13g2_xnor2_1 _1875_ (.Y(_0552_),
    .A(\tokenflow_inst.ii3.i.ydata[16] ),
    .B(_0551_));
 sg13g2_nor2_1 _1876_ (.A(net650),
    .B(_0552_),
    .Y(_0317_));
 sg13g2_a21oi_1 _1877_ (.A1(\tokenflow_inst.ii3.i.ydata[16] ),
    .A2(_0551_),
    .Y(_0553_),
    .B1(\tokenflow_inst.ii3.i.ydata[17] ));
 sg13g2_nand3_1 _1878_ (.B(\tokenflow_inst.ii3.i.ydata[17] ),
    .C(_0551_),
    .A(\tokenflow_inst.ii3.i.ydata[16] ),
    .Y(_0554_));
 sg13g2_nand2_1 _1879_ (.Y(_0555_),
    .A(net683),
    .B(_0554_));
 sg13g2_nor2_1 _1880_ (.A(_0553_),
    .B(_0555_),
    .Y(_0318_));
 sg13g2_nand2b_1 _1881_ (.Y(_0556_),
    .B(_0554_),
    .A_N(\tokenflow_inst.ii3.i.ydata[18] ));
 sg13g2_nand4_1 _1882_ (.B(\tokenflow_inst.ii3.i.ydata[17] ),
    .C(\tokenflow_inst.ii3.i.ydata[18] ),
    .A(\tokenflow_inst.ii3.i.ydata[16] ),
    .Y(_0557_),
    .D(_0551_));
 sg13g2_and3_1 _1883_ (.X(_0319_),
    .A(net683),
    .B(_0556_),
    .C(_0557_));
 sg13g2_nand4_1 _1884_ (.B(\tokenflow_inst.ii3.i.ydata[17] ),
    .C(\tokenflow_inst.ii3.i.ydata[18] ),
    .A(\tokenflow_inst.ii3.i.ydata[16] ),
    .Y(_0558_),
    .D(\tokenflow_inst.ii3.i.ydata[19] ));
 sg13g2_nor4_2 _1885_ (.A(_0743_),
    .B(_0545_),
    .C(_0550_),
    .Y(_0559_),
    .D(_0558_));
 sg13g2_nand2b_1 _1886_ (.Y(_0560_),
    .B(net667),
    .A_N(_0559_));
 sg13g2_a21oi_1 _1887_ (.A1(_0744_),
    .A2(_0557_),
    .Y(_0320_),
    .B1(_0560_));
 sg13g2_o21ai_1 _1888_ (.B1(net668),
    .Y(_0561_),
    .A1(\tokenflow_inst.ii3.i.ydata[20] ),
    .A2(_0559_));
 sg13g2_a21oi_1 _1889_ (.A1(\tokenflow_inst.ii3.i.ydata[20] ),
    .A2(_0559_),
    .Y(_0322_),
    .B1(_0561_));
 sg13g2_a21oi_1 _1890_ (.A1(\tokenflow_inst.ii3.i.ydata[20] ),
    .A2(_0559_),
    .Y(_0562_),
    .B1(\tokenflow_inst.ii3.i.ydata[21] ));
 sg13g2_and3_2 _1891_ (.X(_0563_),
    .A(\tokenflow_inst.ii3.i.ydata[20] ),
    .B(\tokenflow_inst.ii3.i.ydata[21] ),
    .C(_0559_));
 sg13g2_nor3_1 _1892_ (.A(net651),
    .B(_0562_),
    .C(_0563_),
    .Y(_0323_));
 sg13g2_o21ai_1 _1893_ (.B1(net657),
    .Y(_0564_),
    .A1(\tokenflow_inst.ii3.i.ydata[22] ),
    .A2(_0563_));
 sg13g2_a21oi_1 _1894_ (.A1(\tokenflow_inst.ii3.i.ydata[22] ),
    .A2(_0563_),
    .Y(_0324_),
    .B1(_0564_));
 sg13g2_a21oi_1 _1895_ (.A1(\tokenflow_inst.ii3.i.ydata[22] ),
    .A2(_0563_),
    .Y(_0565_),
    .B1(\tokenflow_inst.ii3.i.ydata[23] ));
 sg13g2_and3_1 _1896_ (.X(_0566_),
    .A(\tokenflow_inst.ii3.i.ydata[22] ),
    .B(\tokenflow_inst.ii3.i.ydata[23] ),
    .C(_0563_));
 sg13g2_nor3_1 _1897_ (.A(net650),
    .B(_0565_),
    .C(_0566_),
    .Y(_0325_));
 sg13g2_or2_1 _1898_ (.X(_0567_),
    .B(_0566_),
    .A(\tokenflow_inst.ii3.i.ydata[24] ));
 sg13g2_nand4_1 _1899_ (.B(\tokenflow_inst.ii3.i.ydata[23] ),
    .C(\tokenflow_inst.ii3.i.ydata[24] ),
    .A(\tokenflow_inst.ii3.i.ydata[22] ),
    .Y(_0568_),
    .D(_0563_));
 sg13g2_and3_1 _1900_ (.X(_0326_),
    .A(net657),
    .B(_0567_),
    .C(_0568_));
 sg13g2_o21ai_1 _1901_ (.B1(net658),
    .Y(_0569_),
    .A1(_0745_),
    .A2(_0568_));
 sg13g2_a21oi_1 _1902_ (.A1(_0745_),
    .A2(_0568_),
    .Y(_0327_),
    .B1(_0569_));
 sg13g2_and2_1 _1903_ (.A(net706),
    .B(\tokenflow_inst.i8.ydata[0] ),
    .X(_0158_));
 sg13g2_a21oi_1 _1904_ (.A1(net566),
    .A2(\tokenflow_inst.i8.ydata[53] ),
    .Y(_0570_),
    .B1(\tokenflow_inst.i8.ydata[1] ));
 sg13g2_nand3_1 _1905_ (.B(\tokenflow_inst.i8.ydata[53] ),
    .C(\tokenflow_inst.i8.ydata[1] ),
    .A(net567),
    .Y(_0571_));
 sg13g2_nand2_1 _1906_ (.Y(_0572_),
    .A(net704),
    .B(_0571_));
 sg13g2_nor2_1 _1907_ (.A(_0570_),
    .B(_0572_),
    .Y(_0169_));
 sg13g2_nand3_1 _1908_ (.B(\tokenflow_inst.i8.ydata[54] ),
    .C(\tokenflow_inst.i8.ydata[2] ),
    .A(net567),
    .Y(_0573_));
 sg13g2_a21oi_1 _1909_ (.A1(net567),
    .A2(\tokenflow_inst.i8.ydata[54] ),
    .Y(_0574_),
    .B1(\tokenflow_inst.i8.ydata[2] ));
 sg13g2_a21o_1 _1910_ (.A2(\tokenflow_inst.i8.ydata[54] ),
    .A1(net567),
    .B1(\tokenflow_inst.i8.ydata[2] ),
    .X(_0575_));
 sg13g2_nand2_1 _1911_ (.Y(_0576_),
    .A(_0573_),
    .B(_0575_));
 sg13g2_o21ai_1 _1912_ (.B1(net706),
    .Y(_0577_),
    .A1(_0571_),
    .A2(_0576_));
 sg13g2_a21oi_1 _1913_ (.A1(_0571_),
    .A2(_0576_),
    .Y(_0180_),
    .B1(_0577_));
 sg13g2_a21oi_1 _1914_ (.A1(net567),
    .A2(\tokenflow_inst.i8.ydata[55] ),
    .Y(_0578_),
    .B1(\tokenflow_inst.i8.ydata[3] ));
 sg13g2_and3_1 _1915_ (.X(_0579_),
    .A(net567),
    .B(\tokenflow_inst.i8.ydata[55] ),
    .C(\tokenflow_inst.i8.ydata[3] ));
 sg13g2_or2_1 _1916_ (.X(_0580_),
    .B(_0579_),
    .A(_0578_));
 sg13g2_o21ai_1 _1917_ (.B1(_0573_),
    .Y(_0581_),
    .A1(_0571_),
    .A2(_0574_));
 sg13g2_nand2b_1 _1918_ (.Y(_0582_),
    .B(_0580_),
    .A_N(_0581_));
 sg13g2_nand2b_1 _1919_ (.Y(_0583_),
    .B(_0581_),
    .A_N(_0580_));
 sg13g2_and3_1 _1920_ (.X(_0191_),
    .A(net705),
    .B(_0582_),
    .C(_0583_));
 sg13g2_and3_1 _1921_ (.X(_0584_),
    .A(net566),
    .B(\tokenflow_inst.i8.ydata[56] ),
    .C(\tokenflow_inst.i8.ydata[4] ));
 sg13g2_a21oi_1 _1922_ (.A1(net566),
    .A2(\tokenflow_inst.i8.ydata[56] ),
    .Y(_0585_),
    .B1(\tokenflow_inst.i8.ydata[4] ));
 sg13g2_nor2_1 _1923_ (.A(_0584_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_nor2_1 _1924_ (.A(_0579_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_nor4_1 _1925_ (.A(_0578_),
    .B(_0579_),
    .C(_0584_),
    .D(_0585_),
    .Y(_0588_));
 sg13g2_a21o_1 _1926_ (.A2(_0586_),
    .A1(_0579_),
    .B1(net655),
    .X(_0589_));
 sg13g2_a221oi_1 _1927_ (.B2(_0581_),
    .C1(_0589_),
    .B1(_0588_),
    .A1(_0583_),
    .Y(_0202_),
    .A2(_0587_));
 sg13g2_a21oi_1 _1928_ (.A1(net566),
    .A2(\tokenflow_inst.i8.ydata[57] ),
    .Y(_0590_),
    .B1(\tokenflow_inst.i8.ydata[5] ));
 sg13g2_nand3_1 _1929_ (.B(\tokenflow_inst.i8.ydata[57] ),
    .C(\tokenflow_inst.i8.ydata[5] ),
    .A(net566),
    .Y(_0591_));
 sg13g2_nand2b_1 _1930_ (.Y(_0592_),
    .B(_0591_),
    .A_N(_0590_));
 sg13g2_a221oi_1 _1931_ (.B2(_0581_),
    .C1(_0584_),
    .B1(_0588_),
    .A1(_0579_),
    .Y(_0593_),
    .A2(_0586_));
 sg13g2_nor2_1 _1932_ (.A(_0592_),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_or2_1 _1933_ (.X(_0595_),
    .B(_0593_),
    .A(_0592_));
 sg13g2_nand2_1 _1934_ (.Y(_0596_),
    .A(net702),
    .B(_0595_));
 sg13g2_a21oi_1 _1935_ (.A1(_0592_),
    .A2(_0593_),
    .Y(_0209_),
    .B1(_0596_));
 sg13g2_and3_1 _1936_ (.X(_0597_),
    .A(net566),
    .B(\tokenflow_inst.i8.ydata[58] ),
    .C(\tokenflow_inst.i8.ydata[6] ));
 sg13g2_nand3_1 _1937_ (.B(\tokenflow_inst.i8.ydata[58] ),
    .C(\tokenflow_inst.i8.ydata[6] ),
    .A(net566),
    .Y(_0598_));
 sg13g2_a21oi_1 _1938_ (.A1(net566),
    .A2(\tokenflow_inst.i8.ydata[58] ),
    .Y(_0599_),
    .B1(\tokenflow_inst.i8.ydata[6] ));
 sg13g2_nor2_2 _1939_ (.A(_0597_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_inv_1 _1940_ (.Y(_0601_),
    .A(_0600_));
 sg13g2_nand3_1 _1941_ (.B(_0595_),
    .C(_0601_),
    .A(_0591_),
    .Y(_0602_));
 sg13g2_o21ai_1 _1942_ (.B1(net702),
    .Y(_0603_),
    .A1(_0591_),
    .A2(_0601_));
 sg13g2_a21oi_1 _1943_ (.A1(_0594_),
    .A2(_0600_),
    .Y(_0604_),
    .B1(_0603_));
 sg13g2_and2_1 _1944_ (.A(_0602_),
    .B(_0604_),
    .X(_0220_));
 sg13g2_a21oi_1 _1945_ (.A1(net564),
    .A2(\tokenflow_inst.i8.ydata[59] ),
    .Y(_0605_),
    .B1(\tokenflow_inst.i8.ydata[7] ));
 sg13g2_and3_1 _1946_ (.X(_0606_),
    .A(net564),
    .B(\tokenflow_inst.i8.ydata[7] ),
    .C(\tokenflow_inst.i8.ydata[59] ));
 sg13g2_nand3_1 _1947_ (.B(\tokenflow_inst.i8.ydata[7] ),
    .C(\tokenflow_inst.i8.ydata[59] ),
    .A(net564),
    .Y(_0607_));
 sg13g2_nand2b_1 _1948_ (.Y(_0608_),
    .B(_0607_),
    .A_N(_0605_));
 sg13g2_o21ai_1 _1949_ (.B1(_0598_),
    .Y(_0609_),
    .A1(_0591_),
    .A2(_0599_));
 sg13g2_a21oi_1 _1950_ (.A1(_0594_),
    .A2(_0600_),
    .Y(_0610_),
    .B1(_0609_));
 sg13g2_or2_1 _1951_ (.X(_0611_),
    .B(_0610_),
    .A(_0608_));
 sg13g2_nand2_1 _1952_ (.Y(_0612_),
    .A(net698),
    .B(_0611_));
 sg13g2_a21oi_1 _1953_ (.A1(_0608_),
    .A2(_0610_),
    .Y(_0229_),
    .B1(_0612_));
 sg13g2_and3_1 _1954_ (.X(_0613_),
    .A(net564),
    .B(\tokenflow_inst.i8.ydata[60] ),
    .C(\tokenflow_inst.i8.ydata[8] ));
 sg13g2_a21oi_1 _1955_ (.A1(net564),
    .A2(\tokenflow_inst.i8.ydata[60] ),
    .Y(_0614_),
    .B1(\tokenflow_inst.i8.ydata[8] ));
 sg13g2_nor2_1 _1956_ (.A(_0613_),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_nand2_1 _1957_ (.Y(_0616_),
    .A(_0607_),
    .B(_0611_));
 sg13g2_o21ai_1 _1958_ (.B1(net697),
    .Y(_0617_),
    .A1(_0615_),
    .A2(_0616_));
 sg13g2_a21oi_1 _1959_ (.A1(_0615_),
    .A2(_0616_),
    .Y(_0230_),
    .B1(_0617_));
 sg13g2_nor4_1 _1960_ (.A(_0605_),
    .B(_0606_),
    .C(_0613_),
    .D(_0614_),
    .Y(_0618_));
 sg13g2_nand3b_1 _1961_ (.B(_0600_),
    .C(_0618_),
    .Y(_0619_),
    .A_N(_0592_));
 sg13g2_a221oi_1 _1962_ (.B2(_0609_),
    .C1(_0613_),
    .B1(_0618_),
    .A1(_0606_),
    .Y(_0620_),
    .A2(_0615_));
 sg13g2_o21ai_1 _1963_ (.B1(_0620_),
    .Y(_0621_),
    .A1(_0593_),
    .A2(_0619_));
 sg13g2_a21oi_1 _1964_ (.A1(net562),
    .A2(\tokenflow_inst.i8.ydata[61] ),
    .Y(_0622_),
    .B1(\tokenflow_inst.i8.ydata[9] ));
 sg13g2_nand3_1 _1965_ (.B(\tokenflow_inst.i8.ydata[9] ),
    .C(\tokenflow_inst.i8.ydata[61] ),
    .A(net562),
    .Y(_0623_));
 sg13g2_nand2b_1 _1966_ (.Y(_0624_),
    .B(_0623_),
    .A_N(_0622_));
 sg13g2_nand2b_1 _1967_ (.Y(_0625_),
    .B(_0624_),
    .A_N(_0621_));
 sg13g2_nand2b_1 _1968_ (.Y(_0626_),
    .B(_0621_),
    .A_N(_0624_));
 sg13g2_and3_1 _1969_ (.X(_0231_),
    .A(net669),
    .B(_0625_),
    .C(_0626_));
 sg13g2_nand3_1 _1970_ (.B(\tokenflow_inst.i8.ydata[62] ),
    .C(\tokenflow_inst.i8.ydata[10] ),
    .A(net562),
    .Y(_0627_));
 sg13g2_a21oi_1 _1971_ (.A1(net562),
    .A2(\tokenflow_inst.i8.ydata[62] ),
    .Y(_0628_),
    .B1(\tokenflow_inst.i8.ydata[10] ));
 sg13g2_a21o_1 _1972_ (.A2(\tokenflow_inst.i8.ydata[62] ),
    .A1(net562),
    .B1(\tokenflow_inst.i8.ydata[10] ),
    .X(_0629_));
 sg13g2_nand2_1 _1973_ (.Y(_0630_),
    .A(_0627_),
    .B(_0629_));
 sg13g2_xnor2_1 _1974_ (.Y(_0631_),
    .A(_0623_),
    .B(_0630_));
 sg13g2_nor2_1 _1975_ (.A(_0624_),
    .B(_0630_),
    .Y(_0632_));
 sg13g2_a221oi_1 _1976_ (.B2(_0621_),
    .C1(net656),
    .B1(_0632_),
    .A1(_0626_),
    .Y(_0159_),
    .A2(_0631_));
 sg13g2_a21oi_1 _1977_ (.A1(net560),
    .A2(\tokenflow_inst.i8.ydata[63] ),
    .Y(_0633_),
    .B1(\tokenflow_inst.i8.ydata[11] ));
 sg13g2_and3_1 _1978_ (.X(_0634_),
    .A(net560),
    .B(\tokenflow_inst.i8.ydata[11] ),
    .C(\tokenflow_inst.i8.ydata[63] ));
 sg13g2_nand3_1 _1979_ (.B(\tokenflow_inst.i8.ydata[11] ),
    .C(\tokenflow_inst.i8.ydata[63] ),
    .A(net560),
    .Y(_0635_));
 sg13g2_nor2_1 _1980_ (.A(_0633_),
    .B(_0634_),
    .Y(_0636_));
 sg13g2_o21ai_1 _1981_ (.B1(_0627_),
    .Y(_0637_),
    .A1(_0623_),
    .A2(_0628_));
 sg13g2_a21o_1 _1982_ (.A2(_0632_),
    .A1(_0621_),
    .B1(_0637_),
    .X(_0638_));
 sg13g2_or2_1 _1983_ (.X(_0639_),
    .B(_0638_),
    .A(_0636_));
 sg13g2_nand2_1 _1984_ (.Y(_0640_),
    .A(_0636_),
    .B(_0638_));
 sg13g2_and3_1 _1985_ (.X(_0160_),
    .A(net664),
    .B(_0639_),
    .C(_0640_));
 sg13g2_and3_1 _1986_ (.X(_0641_),
    .A(net560),
    .B(\tokenflow_inst.i8.ydata[64] ),
    .C(\tokenflow_inst.i8.ydata[12] ));
 sg13g2_nand3_1 _1987_ (.B(\tokenflow_inst.i8.ydata[64] ),
    .C(\tokenflow_inst.i8.ydata[12] ),
    .A(net560),
    .Y(_0642_));
 sg13g2_a21oi_2 _1988_ (.B1(\tokenflow_inst.i8.ydata[12] ),
    .Y(_0643_),
    .A2(\tokenflow_inst.i8.ydata[64] ),
    .A1(net560));
 sg13g2_nor2_1 _1989_ (.A(_0641_),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_nand2_1 _1990_ (.Y(_0645_),
    .A(_0635_),
    .B(_0640_));
 sg13g2_o21ai_1 _1991_ (.B1(net673),
    .Y(_0646_),
    .A1(_0644_),
    .A2(_0645_));
 sg13g2_a21oi_1 _1992_ (.A1(_0644_),
    .A2(_0645_),
    .Y(_0161_),
    .B1(_0646_));
 sg13g2_a21oi_1 _1993_ (.A1(net561),
    .A2(\tokenflow_inst.i8.ydata[65] ),
    .Y(_0647_),
    .B1(\tokenflow_inst.i8.ydata[13] ));
 sg13g2_nand3_1 _1994_ (.B(\tokenflow_inst.i8.ydata[13] ),
    .C(\tokenflow_inst.i8.ydata[65] ),
    .A(net561),
    .Y(_0648_));
 sg13g2_nand2b_2 _1995_ (.Y(_0649_),
    .B(_0648_),
    .A_N(_0647_));
 sg13g2_o21ai_1 _1996_ (.B1(_0642_),
    .Y(_0650_),
    .A1(_0635_),
    .A2(_0643_));
 sg13g2_nor4_2 _1997_ (.A(_0633_),
    .B(_0634_),
    .C(_0641_),
    .Y(_0651_),
    .D(_0643_));
 sg13g2_a21o_1 _1998_ (.A2(_0651_),
    .A1(_0637_),
    .B1(_0650_),
    .X(_0652_));
 sg13g2_a21oi_2 _1999_ (.B1(_0650_),
    .Y(_0653_),
    .A2(_0651_),
    .A1(_0638_));
 sg13g2_or2_1 _2000_ (.X(_0654_),
    .B(_0653_),
    .A(_0649_));
 sg13g2_nand2_1 _2001_ (.Y(_0655_),
    .A(net672),
    .B(_0654_));
 sg13g2_a21oi_1 _2002_ (.A1(_0649_),
    .A2(_0653_),
    .Y(_0162_),
    .B1(_0655_));
 sg13g2_nand3_1 _2003_ (.B(\tokenflow_inst.i8.ydata[66] ),
    .C(\tokenflow_inst.i8.ydata[14] ),
    .A(net560),
    .Y(_0656_));
 sg13g2_a21o_1 _2004_ (.A2(\tokenflow_inst.i8.ydata[66] ),
    .A1(net560),
    .B1(\tokenflow_inst.i8.ydata[14] ),
    .X(_0657_));
 sg13g2_nand2_2 _2005_ (.Y(_0658_),
    .A(_0656_),
    .B(_0657_));
 sg13g2_nor3_2 _2006_ (.A(_0649_),
    .B(_0653_),
    .C(_0658_),
    .Y(_0659_));
 sg13g2_and3_1 _2007_ (.X(_0660_),
    .A(_0648_),
    .B(_0654_),
    .C(_0658_));
 sg13g2_o21ai_1 _2008_ (.B1(net672),
    .Y(_0661_),
    .A1(_0648_),
    .A2(_0658_));
 sg13g2_nor3_1 _2009_ (.A(_0659_),
    .B(_0660_),
    .C(_0661_),
    .Y(_0163_));
 sg13g2_a21oi_1 _2010_ (.A1(net562),
    .A2(\tokenflow_inst.i8.ydata[67] ),
    .Y(_0662_),
    .B1(\tokenflow_inst.i8.ydata[15] ));
 sg13g2_nand3_1 _2011_ (.B(\tokenflow_inst.i8.ydata[15] ),
    .C(\tokenflow_inst.i8.ydata[67] ),
    .A(net562),
    .Y(_0663_));
 sg13g2_nand2b_1 _2012_ (.Y(_0664_),
    .B(_0663_),
    .A_N(_0662_));
 sg13g2_inv_1 _2013_ (.Y(_0665_),
    .A(_0664_));
 sg13g2_o21ai_1 _2014_ (.B1(_0656_),
    .Y(_0666_),
    .A1(_0648_),
    .A2(_0658_));
 sg13g2_nor3_1 _2015_ (.A(_0659_),
    .B(_0665_),
    .C(_0666_),
    .Y(_0667_));
 sg13g2_o21ai_1 _2016_ (.B1(_0665_),
    .Y(_0668_),
    .A1(_0659_),
    .A2(_0666_));
 sg13g2_nand2_1 _2017_ (.Y(_0669_),
    .A(net679),
    .B(_0668_));
 sg13g2_nor2_1 _2018_ (.A(_0667_),
    .B(_0669_),
    .Y(_0164_));
 sg13g2_a21oi_1 _2019_ (.A1(net563),
    .A2(\tokenflow_inst.i8.ydata[68] ),
    .Y(_0670_),
    .B1(\tokenflow_inst.i8.ydata[16] ));
 sg13g2_nand3_1 _2020_ (.B(\tokenflow_inst.i8.ydata[68] ),
    .C(\tokenflow_inst.i8.ydata[16] ),
    .A(net562),
    .Y(_0671_));
 sg13g2_nand2b_1 _2021_ (.Y(_0672_),
    .B(_0671_),
    .A_N(_0670_));
 sg13g2_and3_1 _2022_ (.X(_0673_),
    .A(_0663_),
    .B(_0668_),
    .C(_0672_));
 sg13g2_a21oi_1 _2023_ (.A1(_0663_),
    .A2(_0668_),
    .Y(_0674_),
    .B1(_0672_));
 sg13g2_nor3_1 _2024_ (.A(net651),
    .B(_0673_),
    .C(_0674_),
    .Y(_0165_));
 sg13g2_a21oi_1 _2025_ (.A1(net565),
    .A2(\tokenflow_inst.i8.ydata[69] ),
    .Y(_0675_),
    .B1(\tokenflow_inst.i8.ydata[17] ));
 sg13g2_nand3_1 _2026_ (.B(\tokenflow_inst.i8.ydata[17] ),
    .C(\tokenflow_inst.i8.ydata[69] ),
    .A(net565),
    .Y(_0676_));
 sg13g2_nand2b_1 _2027_ (.Y(_0677_),
    .B(_0676_),
    .A_N(_0675_));
 sg13g2_nor2_1 _2028_ (.A(_0664_),
    .B(_0672_),
    .Y(_0678_));
 sg13g2_nor4_1 _2029_ (.A(_0649_),
    .B(_0658_),
    .C(_0664_),
    .D(_0672_),
    .Y(_0679_));
 sg13g2_o21ai_1 _2030_ (.B1(_0671_),
    .Y(_0680_),
    .A1(_0663_),
    .A2(_0670_));
 sg13g2_and3_1 _2031_ (.X(_0681_),
    .A(_0632_),
    .B(_0651_),
    .C(_0679_));
 sg13g2_a21o_1 _2032_ (.A2(_0679_),
    .A1(_0652_),
    .B1(_0680_),
    .X(_0682_));
 sg13g2_a221oi_1 _2033_ (.B2(_0621_),
    .C1(_0682_),
    .B1(_0681_),
    .A1(_0666_),
    .Y(_0683_),
    .A2(_0678_));
 sg13g2_or2_1 _2034_ (.X(_0684_),
    .B(_0683_),
    .A(_0677_));
 sg13g2_nand2_1 _2035_ (.Y(_0685_),
    .A(net699),
    .B(_0684_));
 sg13g2_a21oi_1 _2036_ (.A1(_0677_),
    .A2(_0683_),
    .Y(_0166_),
    .B1(_0685_));
 sg13g2_nand3_1 _2037_ (.B(\tokenflow_inst.i8.ydata[18] ),
    .C(\tokenflow_inst.i8.ydata[70] ),
    .A(net564),
    .Y(_0686_));
 sg13g2_a21o_1 _2038_ (.A2(\tokenflow_inst.i8.ydata[70] ),
    .A1(net564),
    .B1(\tokenflow_inst.i8.ydata[18] ),
    .X(_0687_));
 sg13g2_nand2_1 _2039_ (.Y(_0688_),
    .A(_0686_),
    .B(_0687_));
 sg13g2_nand3_1 _2040_ (.B(_0684_),
    .C(_0688_),
    .A(_0676_),
    .Y(_0689_));
 sg13g2_a21o_1 _2041_ (.A2(_0684_),
    .A1(_0676_),
    .B1(_0688_),
    .X(_0690_));
 sg13g2_and3_1 _2042_ (.X(_0167_),
    .A(net701),
    .B(_0689_),
    .C(_0690_));
 sg13g2_a21oi_1 _2043_ (.A1(net565),
    .A2(\tokenflow_inst.i8.ydata[71] ),
    .Y(_0691_),
    .B1(\tokenflow_inst.i8.ydata[19] ));
 sg13g2_nand3_1 _2044_ (.B(\tokenflow_inst.i8.ydata[19] ),
    .C(\tokenflow_inst.i8.ydata[71] ),
    .A(net565),
    .Y(_0692_));
 sg13g2_nand2b_1 _2045_ (.Y(_0693_),
    .B(_0692_),
    .A_N(_0691_));
 sg13g2_nand3_1 _2046_ (.B(_0690_),
    .C(_0693_),
    .A(_0686_),
    .Y(_0694_));
 sg13g2_a21o_1 _2047_ (.A2(_0690_),
    .A1(_0686_),
    .B1(_0693_),
    .X(_0695_));
 sg13g2_and3_1 _2048_ (.X(_0168_),
    .A(net699),
    .B(_0694_),
    .C(_0695_));
 sg13g2_and3_1 _2049_ (.X(_0696_),
    .A(net565),
    .B(\tokenflow_inst.i8.ydata[72] ),
    .C(\tokenflow_inst.i8.ydata[20] ));
 sg13g2_a21oi_1 _2050_ (.A1(net564),
    .A2(\tokenflow_inst.i8.ydata[72] ),
    .Y(_0697_),
    .B1(\tokenflow_inst.i8.ydata[20] ));
 sg13g2_or2_1 _2051_ (.X(_0698_),
    .B(_0697_),
    .A(_0696_));
 sg13g2_and3_1 _2052_ (.X(_0699_),
    .A(_0692_),
    .B(_0695_),
    .C(_0698_));
 sg13g2_a21oi_1 _2053_ (.A1(_0692_),
    .A2(_0695_),
    .Y(_0700_),
    .B1(_0698_));
 sg13g2_nor3_1 _2054_ (.A(net655),
    .B(_0699_),
    .C(_0700_),
    .Y(_0170_));
 sg13g2_nor2_1 _2055_ (.A(_0693_),
    .B(_0698_),
    .Y(_0701_));
 sg13g2_or4_1 _2056_ (.A(_0677_),
    .B(_0688_),
    .C(_0693_),
    .D(_0698_),
    .X(_0702_));
 sg13g2_nand2_1 _2057_ (.Y(_0703_),
    .A(_0676_),
    .B(_0686_));
 sg13g2_and2_1 _2058_ (.A(_0687_),
    .B(_0703_),
    .X(_0704_));
 sg13g2_nor2_1 _2059_ (.A(_0692_),
    .B(_0697_),
    .Y(_0705_));
 sg13g2_a21oi_1 _2060_ (.A1(_0701_),
    .A2(_0704_),
    .Y(_0706_),
    .B1(_0696_));
 sg13g2_nor2b_1 _2061_ (.A(_0705_),
    .B_N(_0706_),
    .Y(_0707_));
 sg13g2_o21ai_1 _2062_ (.B1(_0707_),
    .Y(_0708_),
    .A1(_0683_),
    .A2(_0702_));
 sg13g2_a21oi_1 _2063_ (.A1(net563),
    .A2(\tokenflow_inst.i8.ydata[73] ),
    .Y(_0709_),
    .B1(\tokenflow_inst.i8.ydata[21] ));
 sg13g2_nand3_1 _2064_ (.B(\tokenflow_inst.i8.ydata[21] ),
    .C(\tokenflow_inst.i8.ydata[73] ),
    .A(net563),
    .Y(_0710_));
 sg13g2_nand2b_1 _2065_ (.Y(_0711_),
    .B(_0710_),
    .A_N(_0709_));
 sg13g2_nand2b_1 _2066_ (.Y(_0712_),
    .B(_0711_),
    .A_N(_0708_));
 sg13g2_nand2b_1 _2067_ (.Y(_0713_),
    .B(_0708_),
    .A_N(_0711_));
 sg13g2_and3_1 _2068_ (.X(_0171_),
    .A(net680),
    .B(_0712_),
    .C(_0713_));
 sg13g2_nand2_1 _2069_ (.Y(_0714_),
    .A(net561),
    .B(\tokenflow_inst.i8.ydata[74] ));
 sg13g2_xnor2_1 _2070_ (.Y(_0715_),
    .A(_0746_),
    .B(_0714_));
 sg13g2_nand3_1 _2071_ (.B(_0713_),
    .C(_0715_),
    .A(_0710_),
    .Y(_0716_));
 sg13g2_nor2_1 _2072_ (.A(_0711_),
    .B(_0715_),
    .Y(_0717_));
 sg13g2_or2_1 _2073_ (.X(_0718_),
    .B(_0715_),
    .A(_0710_));
 sg13g2_a21oi_1 _2074_ (.A1(_0708_),
    .A2(_0717_),
    .Y(_0719_),
    .B1(net651));
 sg13g2_and3_1 _2075_ (.X(_0172_),
    .A(_0716_),
    .B(_0718_),
    .C(_0719_));
 sg13g2_o21ai_1 _2076_ (.B1(_0718_),
    .Y(_0720_),
    .A1(_0746_),
    .A2(_0714_));
 sg13g2_a21oi_2 _2077_ (.B1(_0720_),
    .Y(_0721_),
    .A2(_0717_),
    .A1(_0708_));
 sg13g2_a21oi_1 _2078_ (.A1(net569),
    .A2(\tokenflow_inst.i8.ydata[75] ),
    .Y(_0722_),
    .B1(\tokenflow_inst.i8.ydata[23] ));
 sg13g2_nand3_1 _2079_ (.B(\tokenflow_inst.i8.ydata[23] ),
    .C(\tokenflow_inst.i8.ydata[75] ),
    .A(net561),
    .Y(_0723_));
 sg13g2_nand2b_1 _2080_ (.Y(_0724_),
    .B(_0723_),
    .A_N(_0722_));
 sg13g2_or2_1 _2081_ (.X(_0725_),
    .B(_0724_),
    .A(_0721_));
 sg13g2_nand2_1 _2082_ (.Y(_0726_),
    .A(net674),
    .B(_0725_));
 sg13g2_a21oi_1 _2083_ (.A1(_0721_),
    .A2(_0724_),
    .Y(_0173_),
    .B1(_0726_));
 sg13g2_nand3_1 _2084_ (.B(\tokenflow_inst.i8.ydata[24] ),
    .C(\tokenflow_inst.i8.ydata[76] ),
    .A(net561),
    .Y(_0727_));
 sg13g2_a21o_1 _2085_ (.A2(\tokenflow_inst.i8.ydata[76] ),
    .A1(net561),
    .B1(\tokenflow_inst.i8.ydata[24] ),
    .X(_0728_));
 sg13g2_nand2_1 _2086_ (.Y(_0729_),
    .A(_0727_),
    .B(_0728_));
 sg13g2_nand3_1 _2087_ (.B(_0725_),
    .C(_0729_),
    .A(_0723_),
    .Y(_0730_));
 sg13g2_or3_1 _2088_ (.A(_0721_),
    .B(_0724_),
    .C(_0729_),
    .X(_0731_));
 sg13g2_or2_1 _2089_ (.X(_0732_),
    .B(_0729_),
    .A(_0723_));
 sg13g2_and4_1 _2090_ (.A(net674),
    .B(_0730_),
    .C(_0731_),
    .D(_0732_),
    .X(_0174_));
 sg13g2_nand2_1 _2091_ (.Y(_0733_),
    .A(net561),
    .B(\tokenflow_inst.i8.ydata[77] ));
 sg13g2_xor2_1 _2092_ (.B(_0733_),
    .A(\tokenflow_inst.i8.ydata[25] ),
    .X(_0734_));
 sg13g2_and2_1 _2093_ (.A(_0727_),
    .B(_0732_),
    .X(_0735_));
 sg13g2_and3_1 _2094_ (.X(_0736_),
    .A(_0731_),
    .B(_0734_),
    .C(_0735_));
 sg13g2_a21oi_1 _2095_ (.A1(_0731_),
    .A2(_0735_),
    .Y(_0737_),
    .B1(_0734_));
 sg13g2_nor3_1 _2096_ (.A(net651),
    .B(_0736_),
    .C(_0737_),
    .Y(_0175_));
 sg13g2_and2_1 _2097_ (.A(net693),
    .B(\tokenflow_inst.i8.ydata[27] ),
    .X(_0176_));
 sg13g2_and2_1 _2098_ (.A(net694),
    .B(\tokenflow_inst.i8.ydata[28] ),
    .X(_0177_));
 sg13g2_and2_1 _2099_ (.A(net693),
    .B(\tokenflow_inst.i8.ydata[29] ),
    .X(_0178_));
 sg13g2_and2_1 _2100_ (.A(net693),
    .B(\tokenflow_inst.i8.ydata[30] ),
    .X(_0179_));
 sg13g2_and2_1 _2101_ (.A(net692),
    .B(\tokenflow_inst.i8.ydata[31] ),
    .X(_0181_));
 sg13g2_and2_1 _2102_ (.A(net695),
    .B(\tokenflow_inst.i8.ydata[32] ),
    .X(_0182_));
 sg13g2_and2_1 _2103_ (.A(net689),
    .B(\tokenflow_inst.i8.ydata[33] ),
    .X(_0183_));
 sg13g2_and2_1 _2104_ (.A(net689),
    .B(\tokenflow_inst.i8.ydata[34] ),
    .X(_0184_));
 sg13g2_and2_1 _2105_ (.A(net670),
    .B(\tokenflow_inst.i8.ydata[35] ),
    .X(_0185_));
 sg13g2_and2_1 _2106_ (.A(net667),
    .B(\tokenflow_inst.i8.ydata[36] ),
    .X(_0186_));
 sg13g2_and2_1 _2107_ (.A(net668),
    .B(\tokenflow_inst.i8.ydata[37] ),
    .X(_0187_));
 sg13g2_and2_1 _2108_ (.A(net658),
    .B(\tokenflow_inst.i8.ydata[38] ),
    .X(_0188_));
 sg13g2_and2_1 _2109_ (.A(net661),
    .B(\tokenflow_inst.i8.ydata[39] ),
    .X(_0189_));
 sg13g2_and2_1 _2110_ (.A(net658),
    .B(\tokenflow_inst.i8.ydata[40] ),
    .X(_0190_));
 sg13g2_and2_1 _2111_ (.A(net669),
    .B(\tokenflow_inst.i8.ydata[41] ),
    .X(_0192_));
 sg13g2_and2_1 _2112_ (.A(net668),
    .B(\tokenflow_inst.i8.ydata[42] ),
    .X(_0193_));
 sg13g2_and2_1 _2113_ (.A(net688),
    .B(\tokenflow_inst.i8.ydata[43] ),
    .X(_0194_));
 sg13g2_and2_1 _2114_ (.A(net684),
    .B(\tokenflow_inst.i8.ydata[44] ),
    .X(_0195_));
 sg13g2_and2_1 _2115_ (.A(net688),
    .B(\tokenflow_inst.i8.ydata[45] ),
    .X(_0196_));
 sg13g2_and2_1 _2116_ (.A(net688),
    .B(\tokenflow_inst.i8.ydata[46] ),
    .X(_0197_));
 sg13g2_and2_1 _2117_ (.A(net669),
    .B(\tokenflow_inst.i8.ydata[47] ),
    .X(_0198_));
 sg13g2_and2_1 _2118_ (.A(net669),
    .B(\tokenflow_inst.i8.ydata[48] ),
    .X(_0199_));
 sg13g2_and2_1 _2119_ (.A(net661),
    .B(\tokenflow_inst.i8.ydata[49] ),
    .X(_0200_));
 sg13g2_and2_1 _2120_ (.A(net662),
    .B(\tokenflow_inst.i8.ydata[50] ),
    .X(_0201_));
 sg13g2_and2_1 _2121_ (.A(net706),
    .B(\tokenflow_inst.i8.ydata[53] ),
    .X(_0203_));
 sg13g2_and2_1 _2122_ (.A(net705),
    .B(\tokenflow_inst.i8.ydata[54] ),
    .X(_0204_));
 sg13g2_and2_1 _2123_ (.A(net703),
    .B(\tokenflow_inst.i8.ydata[55] ),
    .X(_0205_));
 sg13g2_and2_1 _2124_ (.A(net703),
    .B(\tokenflow_inst.i8.ydata[56] ),
    .X(_0206_));
 sg13g2_and2_1 _2125_ (.A(net702),
    .B(\tokenflow_inst.i8.ydata[57] ),
    .X(_0207_));
 sg13g2_and2_1 _2126_ (.A(net702),
    .B(\tokenflow_inst.i8.ydata[58] ),
    .X(_0208_));
 sg13g2_and2_1 _2127_ (.A(net698),
    .B(\tokenflow_inst.i8.ydata[59] ),
    .X(_0210_));
 sg13g2_and2_1 _2128_ (.A(net697),
    .B(\tokenflow_inst.i8.ydata[60] ),
    .X(_0211_));
 sg13g2_and2_1 _2129_ (.A(net670),
    .B(\tokenflow_inst.i8.ydata[61] ),
    .X(_0212_));
 sg13g2_and2_1 _2130_ (.A(net663),
    .B(\tokenflow_inst.i8.ydata[62] ),
    .X(_0213_));
 sg13g2_and2_1 _2131_ (.A(net662),
    .B(\tokenflow_inst.i8.ydata[63] ),
    .X(_0214_));
 sg13g2_and2_1 _2132_ (.A(net673),
    .B(\tokenflow_inst.i8.ydata[64] ),
    .X(_0215_));
 sg13g2_and2_1 _2133_ (.A(net677),
    .B(\tokenflow_inst.i8.ydata[65] ),
    .X(_0216_));
 sg13g2_and2_1 _2134_ (.A(net679),
    .B(\tokenflow_inst.i8.ydata[66] ),
    .X(_0217_));
 sg13g2_and2_1 _2135_ (.A(net679),
    .B(\tokenflow_inst.i8.ydata[67] ),
    .X(_0218_));
 sg13g2_and2_1 _2136_ (.A(net678),
    .B(\tokenflow_inst.i8.ydata[68] ),
    .X(_0219_));
 sg13g2_and2_1 _2137_ (.A(net700),
    .B(\tokenflow_inst.i8.ydata[69] ),
    .X(_0221_));
 sg13g2_and2_1 _2138_ (.A(net701),
    .B(\tokenflow_inst.i8.ydata[70] ),
    .X(_0222_));
 sg13g2_and2_1 _2139_ (.A(net700),
    .B(\tokenflow_inst.i8.ydata[71] ),
    .X(_0223_));
 sg13g2_and2_1 _2140_ (.A(net681),
    .B(\tokenflow_inst.i8.ydata[72] ),
    .X(_0224_));
 sg13g2_and2_1 _2141_ (.A(net675),
    .B(\tokenflow_inst.i8.ydata[73] ),
    .X(_0225_));
 sg13g2_and2_1 _2142_ (.A(net675),
    .B(\tokenflow_inst.i8.ydata[74] ),
    .X(_0226_));
 sg13g2_and2_1 _2143_ (.A(net674),
    .B(\tokenflow_inst.i8.ydata[75] ),
    .X(_0227_));
 sg13g2_and2_1 _2144_ (.A(net674),
    .B(\tokenflow_inst.i8.ydata[76] ),
    .X(_0228_));
 sg13g2_nor2_1 _2145_ (.A(net653),
    .B(\tokenflow_inst.i2.cg2.a ),
    .Y(_0078_));
 sg13g2_nor2_1 _2146_ (.A(net652),
    .B(\tokenflow_inst.ii1.cg_elem.maj.C ),
    .Y(_0336_));
 sg13g2_xor2_1 _2147_ (.B(\tokenflow_inst.i3.ydata[15] ),
    .A(\tokenflow_inst.i3.ydata[0] ),
    .X(uo_out[1]));
 sg13g2_xor2_1 _2148_ (.B(\tokenflow_inst.i3.ydata[16] ),
    .A(\tokenflow_inst.i3.ydata[1] ),
    .X(uo_out[2]));
 sg13g2_xor2_1 _2149_ (.B(\tokenflow_inst.i3.ydata[17] ),
    .A(\tokenflow_inst.i3.ydata[2] ),
    .X(uo_out[3]));
 sg13g2_xor2_1 _2150_ (.B(\tokenflow_inst.i3.ydata[18] ),
    .A(\tokenflow_inst.i3.ydata[3] ),
    .X(uo_out[4]));
 sg13g2_xor2_1 _2151_ (.B(\tokenflow_inst.i3.ydata[19] ),
    .A(\tokenflow_inst.i3.ydata[4] ),
    .X(uo_out[5]));
 sg13g2_xor2_1 _2152_ (.B(\tokenflow_inst.i3.ydata[20] ),
    .A(\tokenflow_inst.i3.ydata[5] ),
    .X(uo_out[6]));
 sg13g2_xor2_1 _2153_ (.B(\tokenflow_inst.i3.ydata[21] ),
    .A(\tokenflow_inst.i3.ydata[6] ),
    .X(uo_out[7]));
 sg13g2_xor2_1 _2154_ (.B(\tokenflow_inst.i3.ydata[22] ),
    .A(\tokenflow_inst.i3.ydata[7] ),
    .X(uio_out[0]));
 sg13g2_xor2_1 _2155_ (.B(\tokenflow_inst.i3.ydata[23] ),
    .A(\tokenflow_inst.i3.ydata[8] ),
    .X(uio_out[1]));
 sg13g2_xor2_1 _2156_ (.B(\tokenflow_inst.i3.ydata[24] ),
    .A(\tokenflow_inst.i3.ydata[9] ),
    .X(uio_out[2]));
 sg13g2_xor2_1 _2157_ (.B(\tokenflow_inst.i3.ydata[25] ),
    .A(\tokenflow_inst.i3.ydata[10] ),
    .X(uio_out[3]));
 sg13g2_dllrq_1 _2158_ (.D(_0228_),
    .GATE_N(net601),
    .RESET_B(net2),
    .Q(\tokenflow_inst.i78.ydata[77] ));
 sg13g2_dllrq_1 _2159_ (.D(_0079_),
    .GATE_N(net557),
    .RESET_B(net3),
    .Q(\tokenflow_inst.i6.ydata[0] ));
 sg13g2_dllrq_1 _2160_ (.D(_0090_),
    .GATE_N(net557),
    .RESET_B(net4),
    .Q(\tokenflow_inst.i6.ydata[1] ));
 sg13g2_dllrq_1 _2161_ (.D(_0101_),
    .GATE_N(net557),
    .RESET_B(net5),
    .Q(\tokenflow_inst.i6.ydata[2] ));
 sg13g2_dllrq_1 _2162_ (.D(_0112_),
    .GATE_N(net558),
    .RESET_B(net6),
    .Q(\tokenflow_inst.i6.ydata[3] ));
 sg13g2_dllrq_1 _2163_ (.D(_0123_),
    .GATE_N(net557),
    .RESET_B(net7),
    .Q(\tokenflow_inst.i6.ydata[4] ));
 sg13g2_dllrq_1 _2164_ (.D(_0134_),
    .GATE_N(net557),
    .RESET_B(net8),
    .Q(\tokenflow_inst.i6.ydata[5] ));
 sg13g2_dllrq_1 _2165_ (.D(_0145_),
    .GATE_N(net556),
    .RESET_B(net9),
    .Q(\tokenflow_inst.i6.ydata[6] ));
 sg13g2_dllrq_1 _2166_ (.D(_0154_),
    .GATE_N(net556),
    .RESET_B(net10),
    .Q(\tokenflow_inst.i6.ydata[7] ));
 sg13g2_dllrq_1 _2167_ (.D(_0155_),
    .GATE_N(net549),
    .RESET_B(net11),
    .Q(\tokenflow_inst.i6.ydata[8] ));
 sg13g2_dllrq_1 _2168_ (.D(_0156_),
    .GATE_N(net549),
    .RESET_B(net12),
    .Q(\tokenflow_inst.i6.ydata[9] ));
 sg13g2_dllrq_1 _2169_ (.D(_0080_),
    .GATE_N(net549),
    .RESET_B(net13),
    .Q(\tokenflow_inst.i6.ydata[10] ));
 sg13g2_dllrq_1 _2170_ (.D(_0081_),
    .GATE_N(net548),
    .RESET_B(net14),
    .Q(\tokenflow_inst.i6.ydata[11] ));
 sg13g2_dllrq_1 _2171_ (.D(_0082_),
    .GATE_N(net548),
    .RESET_B(net15),
    .Q(\tokenflow_inst.i6.ydata[12] ));
 sg13g2_dllrq_1 _2172_ (.D(_0083_),
    .GATE_N(net550),
    .RESET_B(net16),
    .Q(\tokenflow_inst.i6.ydata[13] ));
 sg13g2_dllrq_1 _2173_ (.D(_0084_),
    .GATE_N(net551),
    .RESET_B(net17),
    .Q(\tokenflow_inst.i6.ydata[14] ));
 sg13g2_dllrq_1 _2174_ (.D(_0085_),
    .GATE_N(net551),
    .RESET_B(net18),
    .Q(\tokenflow_inst.i6.ydata[15] ));
 sg13g2_dllrq_1 _2175_ (.D(_0086_),
    .GATE_N(net558),
    .RESET_B(net19),
    .Q(\tokenflow_inst.i6.ydata[16] ));
 sg13g2_dllrq_1 _2176_ (.D(_0087_),
    .GATE_N(net556),
    .RESET_B(net20),
    .Q(\tokenflow_inst.i6.ydata[17] ));
 sg13g2_dllrq_1 _2177_ (.D(_0088_),
    .GATE_N(net556),
    .RESET_B(net21),
    .Q(\tokenflow_inst.i6.ydata[18] ));
 sg13g2_dllrq_1 _2178_ (.D(_0089_),
    .GATE_N(net558),
    .RESET_B(net22),
    .Q(\tokenflow_inst.i6.ydata[19] ));
 sg13g2_dllrq_1 _2179_ (.D(_0091_),
    .GATE_N(net551),
    .RESET_B(net23),
    .Q(\tokenflow_inst.i6.ydata[20] ));
 sg13g2_dllrq_1 _2180_ (.D(_0092_),
    .GATE_N(net551),
    .RESET_B(net24),
    .Q(\tokenflow_inst.i6.ydata[21] ));
 sg13g2_dllrq_1 _2181_ (.D(_0093_),
    .GATE_N(net552),
    .RESET_B(net25),
    .Q(\tokenflow_inst.i6.ydata[22] ));
 sg13g2_dllrq_1 _2182_ (.D(_0094_),
    .GATE_N(net550),
    .RESET_B(net26),
    .Q(\tokenflow_inst.i6.ydata[23] ));
 sg13g2_dllrq_1 _2183_ (.D(_0095_),
    .GATE_N(net550),
    .RESET_B(net27),
    .Q(\tokenflow_inst.i6.ydata[24] ));
 sg13g2_dllrq_1 _2184_ (.D(_0096_),
    .GATE_N(net550),
    .RESET_B(net28),
    .Q(\tokenflow_inst.i6.ydata[25] ));
 sg13g2_dllrq_1 _2185_ (.D(_0097_),
    .GATE_N(net554),
    .RESET_B(net29),
    .Q(\tokenflow_inst.i6.ydata[26] ));
 sg13g2_dllrq_1 _2186_ (.D(_0098_),
    .GATE_N(net559),
    .RESET_B(net30),
    .Q(\tokenflow_inst.i6.ydata[27] ));
 sg13g2_dllrq_1 _2187_ (.D(_0099_),
    .GATE_N(net554),
    .RESET_B(net31),
    .Q(\tokenflow_inst.i6.ydata[28] ));
 sg13g2_dllrq_1 _2188_ (.D(_0100_),
    .GATE_N(net554),
    .RESET_B(net32),
    .Q(\tokenflow_inst.i6.ydata[29] ));
 sg13g2_dllrq_1 _2189_ (.D(_0102_),
    .GATE_N(net554),
    .RESET_B(net33),
    .Q(\tokenflow_inst.i6.ydata[30] ));
 sg13g2_dllrq_1 _2190_ (.D(_0103_),
    .GATE_N(net554),
    .RESET_B(net34),
    .Q(\tokenflow_inst.i6.ydata[31] ));
 sg13g2_dllrq_1 _2191_ (.D(_0104_),
    .GATE_N(net554),
    .RESET_B(net35),
    .Q(\tokenflow_inst.i6.ydata[32] ));
 sg13g2_dllrq_1 _2192_ (.D(_0105_),
    .GATE_N(net554),
    .RESET_B(net36),
    .Q(\tokenflow_inst.i6.ydata[33] ));
 sg13g2_dllrq_1 _2193_ (.D(_0106_),
    .GATE_N(net555),
    .RESET_B(net37),
    .Q(\tokenflow_inst.i6.ydata[34] ));
 sg13g2_dllrq_1 _2194_ (.D(_0107_),
    .GATE_N(net555),
    .RESET_B(net38),
    .Q(\tokenflow_inst.i6.ydata[35] ));
 sg13g2_dllrq_1 _2195_ (.D(_0108_),
    .GATE_N(net553),
    .RESET_B(net39),
    .Q(\tokenflow_inst.i6.ydata[36] ));
 sg13g2_dllrq_1 _2196_ (.D(_0109_),
    .GATE_N(net549),
    .RESET_B(net40),
    .Q(\tokenflow_inst.i6.ydata[37] ));
 sg13g2_dllrq_1 _2197_ (.D(_0110_),
    .GATE_N(net547),
    .RESET_B(net41),
    .Q(\tokenflow_inst.i6.ydata[38] ));
 sg13g2_dllrq_1 _2198_ (.D(_0111_),
    .GATE_N(net547),
    .RESET_B(net42),
    .Q(\tokenflow_inst.i6.ydata[39] ));
 sg13g2_dllrq_1 _2199_ (.D(_0113_),
    .GATE_N(net547),
    .RESET_B(net43),
    .Q(\tokenflow_inst.i6.ydata[40] ));
 sg13g2_dllrq_1 _2200_ (.D(_0114_),
    .GATE_N(net547),
    .RESET_B(net44),
    .Q(\tokenflow_inst.i6.ydata[41] ));
 sg13g2_dllrq_1 _2201_ (.D(_0115_),
    .GATE_N(net553),
    .RESET_B(net45),
    .Q(\tokenflow_inst.i6.ydata[42] ));
 sg13g2_dllrq_1 _2202_ (.D(_0116_),
    .GATE_N(net549),
    .RESET_B(net46),
    .Q(\tokenflow_inst.i6.ydata[43] ));
 sg13g2_dllrq_1 _2203_ (.D(_0117_),
    .GATE_N(net555),
    .RESET_B(net47),
    .Q(\tokenflow_inst.i6.ydata[44] ));
 sg13g2_dllrq_1 _2204_ (.D(_0118_),
    .GATE_N(net555),
    .RESET_B(net48),
    .Q(\tokenflow_inst.i6.ydata[45] ));
 sg13g2_dllrq_1 _2205_ (.D(_0119_),
    .GATE_N(net555),
    .RESET_B(net49),
    .Q(\tokenflow_inst.i6.ydata[46] ));
 sg13g2_dllrq_1 _2206_ (.D(_0120_),
    .GATE_N(net555),
    .RESET_B(net50),
    .Q(\tokenflow_inst.i6.ydata[47] ));
 sg13g2_dllrq_1 _2207_ (.D(_0121_),
    .GATE_N(net547),
    .RESET_B(net51),
    .Q(\tokenflow_inst.i6.ydata[48] ));
 sg13g2_dllrq_1 _2208_ (.D(_0122_),
    .GATE_N(net547),
    .RESET_B(net52),
    .Q(\tokenflow_inst.i6.ydata[49] ));
 sg13g2_dllrq_1 _2209_ (.D(_0124_),
    .GATE_N(net547),
    .RESET_B(net53),
    .Q(\tokenflow_inst.i6.ydata[50] ));
 sg13g2_dllrq_1 _2210_ (.D(_0125_),
    .GATE_N(net547),
    .RESET_B(net54),
    .Q(\tokenflow_inst.i6.ydata[51] ));
 sg13g2_dllrq_1 _2211_ (.D(_0126_),
    .GATE_N(net557),
    .RESET_B(net55),
    .Q(\tokenflow_inst.i6.ydata[52] ));
 sg13g2_dllrq_1 _2212_ (.D(_0127_),
    .GATE_N(net558),
    .RESET_B(net56),
    .Q(\tokenflow_inst.i6.ydata[53] ));
 sg13g2_dllrq_1 _2213_ (.D(_0128_),
    .GATE_N(net558),
    .RESET_B(net57),
    .Q(\tokenflow_inst.i6.ydata[54] ));
 sg13g2_dllrq_1 _2214_ (.D(_0129_),
    .GATE_N(net557),
    .RESET_B(net58),
    .Q(\tokenflow_inst.i6.ydata[55] ));
 sg13g2_dllrq_1 _2215_ (.D(_0130_),
    .GATE_N(net557),
    .RESET_B(net59),
    .Q(\tokenflow_inst.i6.ydata[56] ));
 sg13g2_dllrq_1 _2216_ (.D(_0131_),
    .GATE_N(net559),
    .RESET_B(net60),
    .Q(\tokenflow_inst.i6.ydata[57] ));
 sg13g2_dllrq_1 _2217_ (.D(_0132_),
    .GATE_N(net559),
    .RESET_B(net61),
    .Q(\tokenflow_inst.i6.ydata[58] ));
 sg13g2_dllrq_1 _2218_ (.D(_0133_),
    .GATE_N(net554),
    .RESET_B(net62),
    .Q(\tokenflow_inst.i6.ydata[59] ));
 sg13g2_dllrq_1 _2219_ (.D(_0135_),
    .GATE_N(net555),
    .RESET_B(net63),
    .Q(\tokenflow_inst.i6.ydata[60] ));
 sg13g2_dllrq_1 _2220_ (.D(_0136_),
    .GATE_N(net549),
    .RESET_B(net64),
    .Q(\tokenflow_inst.i6.ydata[61] ));
 sg13g2_dllrq_1 _2221_ (.D(_0137_),
    .GATE_N(net548),
    .RESET_B(net65),
    .Q(\tokenflow_inst.i6.ydata[62] ));
 sg13g2_dllrq_1 _2222_ (.D(_0138_),
    .GATE_N(net548),
    .RESET_B(net66),
    .Q(\tokenflow_inst.i6.ydata[63] ));
 sg13g2_dllrq_1 _2223_ (.D(_0139_),
    .GATE_N(net548),
    .RESET_B(net67),
    .Q(\tokenflow_inst.i6.ydata[64] ));
 sg13g2_dllrq_1 _2224_ (.D(_0140_),
    .GATE_N(net550),
    .RESET_B(net68),
    .Q(\tokenflow_inst.i6.ydata[65] ));
 sg13g2_dllrq_1 _2225_ (.D(_0141_),
    .GATE_N(net551),
    .RESET_B(net69),
    .Q(\tokenflow_inst.i6.ydata[66] ));
 sg13g2_dllrq_1 _2226_ (.D(_0142_),
    .GATE_N(net551),
    .RESET_B(net70),
    .Q(\tokenflow_inst.i6.ydata[67] ));
 sg13g2_dllrq_1 _2227_ (.D(_0143_),
    .GATE_N(net556),
    .RESET_B(net71),
    .Q(\tokenflow_inst.i6.ydata[68] ));
 sg13g2_dllrq_1 _2228_ (.D(_0144_),
    .GATE_N(net556),
    .RESET_B(net72),
    .Q(\tokenflow_inst.i6.ydata[69] ));
 sg13g2_dllrq_1 _2229_ (.D(_0146_),
    .GATE_N(net556),
    .RESET_B(net73),
    .Q(\tokenflow_inst.i6.ydata[70] ));
 sg13g2_dllrq_1 _2230_ (.D(_0147_),
    .GATE_N(net556),
    .RESET_B(net74),
    .Q(\tokenflow_inst.i6.ydata[71] ));
 sg13g2_dllrq_1 _2231_ (.D(_0148_),
    .GATE_N(net551),
    .RESET_B(net75),
    .Q(\tokenflow_inst.i6.ydata[72] ));
 sg13g2_dllrq_1 _2232_ (.D(_0149_),
    .GATE_N(net551),
    .RESET_B(net76),
    .Q(\tokenflow_inst.i6.ydata[73] ));
 sg13g2_dllrq_1 _2233_ (.D(_0150_),
    .GATE_N(net550),
    .RESET_B(net77),
    .Q(\tokenflow_inst.i6.ydata[74] ));
 sg13g2_dllrq_1 _2234_ (.D(_0151_),
    .GATE_N(net552),
    .RESET_B(net78),
    .Q(\tokenflow_inst.i6.ydata[75] ));
 sg13g2_dllrq_1 _2235_ (.D(_0152_),
    .GATE_N(net550),
    .RESET_B(net79),
    .Q(\tokenflow_inst.i6.ydata[76] ));
 sg13g2_dllrq_1 _2236_ (.D(_0153_),
    .GATE_N(net550),
    .RESET_B(net80),
    .Q(\tokenflow_inst.i6.ydata[77] ));
 sg13g2_dllrq_1 _2237_ (.D(_0000_),
    .GATE_N(net624),
    .RESET_B(net81),
    .Q(\tokenflow_inst.i3.ydata[0] ));
 sg13g2_dllrq_1 _2238_ (.D(_0011_),
    .GATE_N(net624),
    .RESET_B(net82),
    .Q(\tokenflow_inst.i3.ydata[1] ));
 sg13g2_dllrq_1 _2239_ (.D(_0022_),
    .GATE_N(net624),
    .RESET_B(net83),
    .Q(\tokenflow_inst.i3.ydata[2] ));
 sg13g2_dllrq_1 _2240_ (.D(_0033_),
    .GATE_N(net626),
    .RESET_B(net84),
    .Q(\tokenflow_inst.i3.ydata[3] ));
 sg13g2_dllrq_1 _2241_ (.D(_0044_),
    .GATE_N(net624),
    .RESET_B(net85),
    .Q(\tokenflow_inst.i3.ydata[4] ));
 sg13g2_dllrq_1 _2242_ (.D(_0055_),
    .GATE_N(net624),
    .RESET_B(net86),
    .Q(\tokenflow_inst.i3.ydata[5] ));
 sg13g2_dllrq_1 _2243_ (.D(_0066_),
    .GATE_N(net625),
    .RESET_B(net87),
    .Q(\tokenflow_inst.i3.ydata[6] ));
 sg13g2_dllrq_1 _2244_ (.D(_0075_),
    .GATE_N(net621),
    .RESET_B(net88),
    .Q(\tokenflow_inst.i3.ydata[7] ));
 sg13g2_dllrq_1 _2245_ (.D(_0076_),
    .GATE_N(net621),
    .RESET_B(net89),
    .Q(\tokenflow_inst.i3.ydata[8] ));
 sg13g2_dllrq_1 _2246_ (.D(_0077_),
    .GATE_N(net617),
    .RESET_B(net90),
    .Q(\tokenflow_inst.i3.ydata[9] ));
 sg13g2_dllrq_1 _2247_ (.D(_0001_),
    .GATE_N(net617),
    .RESET_B(net91),
    .Q(\tokenflow_inst.i3.ydata[10] ));
 sg13g2_dllrq_1 _2248_ (.D(_0002_),
    .GATE_N(net617),
    .RESET_B(net92),
    .Q(\tokenflow_inst.i3.ydata[11] ));
 sg13g2_dllrq_1 _2249_ (.D(_0003_),
    .GATE_N(net617),
    .RESET_B(net93),
    .Q(\tokenflow_inst.i3.ydata[12] ));
 sg13g2_dllrq_1 _2250_ (.D(_0004_),
    .GATE_N(net618),
    .RESET_B(net94),
    .Q(\tokenflow_inst.i3.ydata[13] ));
 sg13g2_dllrq_1 _2251_ (.D(_0005_),
    .GATE_N(net618),
    .RESET_B(net95),
    .Q(\tokenflow_inst.i3.ydata[14] ));
 sg13g2_dllrq_1 _2252_ (.D(_0006_),
    .GATE_N(net620),
    .RESET_B(net96),
    .Q(\tokenflow_inst.i3.ydata[15] ));
 sg13g2_dllrq_1 _2253_ (.D(_0007_),
    .GATE_N(net625),
    .RESET_B(net97),
    .Q(\tokenflow_inst.i3.ydata[16] ));
 sg13g2_dllrq_1 _2254_ (.D(_0008_),
    .GATE_N(net625),
    .RESET_B(net98),
    .Q(\tokenflow_inst.i3.ydata[17] ));
 sg13g2_dllrq_1 _2255_ (.D(_0009_),
    .GATE_N(net625),
    .RESET_B(net99),
    .Q(\tokenflow_inst.i3.ydata[18] ));
 sg13g2_dllrq_1 _2256_ (.D(_0010_),
    .GATE_N(net625),
    .RESET_B(net100),
    .Q(\tokenflow_inst.i3.ydata[19] ));
 sg13g2_dllrq_1 _2257_ (.D(_0012_),
    .GATE_N(net619),
    .RESET_B(net101),
    .Q(\tokenflow_inst.i3.ydata[20] ));
 sg13g2_dllrq_1 _2258_ (.D(_0013_),
    .GATE_N(net619),
    .RESET_B(net102),
    .Q(\tokenflow_inst.i3.ydata[21] ));
 sg13g2_dllrq_1 _2259_ (.D(_0014_),
    .GATE_N(net620),
    .RESET_B(net103),
    .Q(\tokenflow_inst.i3.ydata[22] ));
 sg13g2_dllrq_1 _2260_ (.D(_0015_),
    .GATE_N(net618),
    .RESET_B(net104),
    .Q(\tokenflow_inst.i3.ydata[23] ));
 sg13g2_dllrq_1 _2261_ (.D(_0016_),
    .GATE_N(net619),
    .RESET_B(net105),
    .Q(\tokenflow_inst.i3.ydata[24] ));
 sg13g2_dllrq_1 _2262_ (.D(_0017_),
    .GATE_N(net618),
    .RESET_B(net106),
    .Q(\tokenflow_inst.i3.ydata[25] ));
 sg13g2_dllrq_1 _2263_ (.D(_0018_),
    .GATE_N(net623),
    .RESET_B(net107),
    .Q(\tokenflow_inst.i3.ydata[26] ));
 sg13g2_dllrq_1 _2264_ (.D(_0019_),
    .GATE_N(net622),
    .RESET_B(net108),
    .Q(\tokenflow_inst.i3.ydata[27] ));
 sg13g2_dllrq_1 _2265_ (.D(_0020_),
    .GATE_N(net622),
    .RESET_B(net109),
    .Q(\tokenflow_inst.i3.ydata[28] ));
 sg13g2_dllrq_1 _2266_ (.D(_0021_),
    .GATE_N(net622),
    .RESET_B(net110),
    .Q(\tokenflow_inst.i3.ydata[29] ));
 sg13g2_dllrq_1 _2267_ (.D(_0023_),
    .GATE_N(net622),
    .RESET_B(net111),
    .Q(\tokenflow_inst.i3.ydata[30] ));
 sg13g2_dllrq_1 _2268_ (.D(_0024_),
    .GATE_N(net622),
    .RESET_B(net112),
    .Q(\tokenflow_inst.i3.ydata[31] ));
 sg13g2_dllrq_1 _2269_ (.D(_0025_),
    .GATE_N(net622),
    .RESET_B(net113),
    .Q(\tokenflow_inst.i3.ydata[32] ));
 sg13g2_dllrq_1 _2270_ (.D(_0026_),
    .GATE_N(net621),
    .RESET_B(net114),
    .Q(\tokenflow_inst.i3.ydata[33] ));
 sg13g2_dllrq_1 _2271_ (.D(_0027_),
    .GATE_N(net621),
    .RESET_B(net115),
    .Q(\tokenflow_inst.i3.ydata[34] ));
 sg13g2_dllrq_1 _2272_ (.D(_0028_),
    .GATE_N(net621),
    .RESET_B(net116),
    .Q(\tokenflow_inst.i3.ydata[35] ));
 sg13g2_dllrq_1 _2273_ (.D(_0029_),
    .GATE_N(net616),
    .RESET_B(net117),
    .Q(\tokenflow_inst.i3.ydata[36] ));
 sg13g2_dllrq_1 _2274_ (.D(_0030_),
    .GATE_N(net615),
    .RESET_B(net118),
    .Q(\tokenflow_inst.i3.ydata[37] ));
 sg13g2_dllrq_1 _2275_ (.D(_0031_),
    .GATE_N(net615),
    .RESET_B(net119),
    .Q(\tokenflow_inst.i3.ydata[38] ));
 sg13g2_dllrq_1 _2276_ (.D(_0032_),
    .GATE_N(net615),
    .RESET_B(net120),
    .Q(\tokenflow_inst.i3.ydata[39] ));
 sg13g2_dllrq_1 _2277_ (.D(_0034_),
    .GATE_N(net616),
    .RESET_B(net121),
    .Q(\tokenflow_inst.i3.ydata[40] ));
 sg13g2_dllrq_1 _2278_ (.D(_0035_),
    .GATE_N(net616),
    .RESET_B(net122),
    .Q(\tokenflow_inst.i3.ydata[41] ));
 sg13g2_dllrq_1 _2279_ (.D(_0036_),
    .GATE_N(net616),
    .RESET_B(net123),
    .Q(\tokenflow_inst.i3.ydata[42] ));
 sg13g2_dllrq_1 _2280_ (.D(_0037_),
    .GATE_N(net616),
    .RESET_B(net124),
    .Q(\tokenflow_inst.i3.ydata[43] ));
 sg13g2_dllrq_1 _2281_ (.D(_0038_),
    .GATE_N(net621),
    .RESET_B(net125),
    .Q(\tokenflow_inst.i3.ydata[44] ));
 sg13g2_dllrq_1 _2282_ (.D(_0039_),
    .GATE_N(net621),
    .RESET_B(net126),
    .Q(\tokenflow_inst.i3.ydata[45] ));
 sg13g2_dllrq_1 _2283_ (.D(_0040_),
    .GATE_N(net616),
    .RESET_B(net127),
    .Q(\tokenflow_inst.i3.ydata[46] ));
 sg13g2_dllrq_1 _2284_ (.D(_0041_),
    .GATE_N(net616),
    .RESET_B(net128),
    .Q(\tokenflow_inst.i3.ydata[47] ));
 sg13g2_dllrq_1 _2285_ (.D(_0042_),
    .GATE_N(net615),
    .RESET_B(net129),
    .Q(\tokenflow_inst.i3.ydata[48] ));
 sg13g2_dllrq_1 _2286_ (.D(_0043_),
    .GATE_N(net615),
    .RESET_B(net130),
    .Q(\tokenflow_inst.i3.ydata[49] ));
 sg13g2_dllrq_1 _2287_ (.D(_0045_),
    .GATE_N(net615),
    .RESET_B(net131),
    .Q(\tokenflow_inst.i3.ydata[50] ));
 sg13g2_dllrq_1 _2288_ (.D(_0046_),
    .GATE_N(net615),
    .RESET_B(net132),
    .Q(\tokenflow_inst.i3.ydata[51] ));
 sg13g2_dllrq_1 _2289_ (.D(_0047_),
    .GATE_N(net624),
    .RESET_B(net133),
    .Q(\tokenflow_inst.i3.ydata[52] ));
 sg13g2_dllrq_1 _2290_ (.D(_0048_),
    .GATE_N(net626),
    .RESET_B(net134),
    .Q(\tokenflow_inst.i3.ydata[53] ));
 sg13g2_dllrq_1 _2291_ (.D(_0049_),
    .GATE_N(net624),
    .RESET_B(net135),
    .Q(\tokenflow_inst.i3.ydata[54] ));
 sg13g2_dllrq_1 _2292_ (.D(_0050_),
    .GATE_N(net626),
    .RESET_B(net136),
    .Q(\tokenflow_inst.i3.ydata[55] ));
 sg13g2_dllrq_1 _2293_ (.D(_0051_),
    .GATE_N(net624),
    .RESET_B(net137),
    .Q(\tokenflow_inst.i3.ydata[56] ));
 sg13g2_dllrq_1 _2294_ (.D(_0052_),
    .GATE_N(net622),
    .RESET_B(net138),
    .Q(\tokenflow_inst.i3.ydata[57] ));
 sg13g2_dllrq_1 _2295_ (.D(_0053_),
    .GATE_N(net622),
    .RESET_B(net139),
    .Q(\tokenflow_inst.i3.ydata[58] ));
 sg13g2_dllrq_1 _2296_ (.D(_0054_),
    .GATE_N(net621),
    .RESET_B(net140),
    .Q(\tokenflow_inst.i3.ydata[59] ));
 sg13g2_dllrq_1 _2297_ (.D(_0056_),
    .GATE_N(net623),
    .RESET_B(net141),
    .Q(\tokenflow_inst.i3.ydata[60] ));
 sg13g2_dllrq_1 _2298_ (.D(_0057_),
    .GATE_N(net623),
    .RESET_B(net142),
    .Q(\tokenflow_inst.i3.ydata[61] ));
 sg13g2_dllrq_1 _2299_ (.D(_0058_),
    .GATE_N(net616),
    .RESET_B(net143),
    .Q(\tokenflow_inst.i3.ydata[62] ));
 sg13g2_dllrq_1 _2300_ (.D(_0059_),
    .GATE_N(net615),
    .RESET_B(net144),
    .Q(\tokenflow_inst.i3.ydata[63] ));
 sg13g2_dllrq_1 _2301_ (.D(_0060_),
    .GATE_N(net617),
    .RESET_B(net145),
    .Q(\tokenflow_inst.i3.ydata[64] ));
 sg13g2_dllrq_1 _2302_ (.D(_0061_),
    .GATE_N(net618),
    .RESET_B(net146),
    .Q(\tokenflow_inst.i3.ydata[65] ));
 sg13g2_dllrq_1 _2303_ (.D(_0062_),
    .GATE_N(net618),
    .RESET_B(net147),
    .Q(\tokenflow_inst.i3.ydata[66] ));
 sg13g2_dllrq_1 _2304_ (.D(_0063_),
    .GATE_N(net617),
    .RESET_B(net148),
    .Q(\tokenflow_inst.i3.ydata[67] ));
 sg13g2_dllrq_1 _2305_ (.D(_0064_),
    .GATE_N(net620),
    .RESET_B(net149),
    .Q(\tokenflow_inst.i3.ydata[68] ));
 sg13g2_dllrq_1 _2306_ (.D(_0065_),
    .GATE_N(net625),
    .RESET_B(net150),
    .Q(\tokenflow_inst.i3.ydata[69] ));
 sg13g2_dllrq_1 _2307_ (.D(_0067_),
    .GATE_N(net625),
    .RESET_B(net151),
    .Q(\tokenflow_inst.i3.ydata[70] ));
 sg13g2_dllrq_1 _2308_ (.D(_0068_),
    .GATE_N(net625),
    .RESET_B(net152),
    .Q(\tokenflow_inst.i3.ydata[71] ));
 sg13g2_dllrq_1 _2309_ (.D(_0069_),
    .GATE_N(net619),
    .RESET_B(net153),
    .Q(\tokenflow_inst.i3.ydata[72] ));
 sg13g2_dllrq_1 _2310_ (.D(_0070_),
    .GATE_N(net619),
    .RESET_B(net154),
    .Q(\tokenflow_inst.i3.ydata[73] ));
 sg13g2_dllrq_1 _2311_ (.D(_0071_),
    .GATE_N(net618),
    .RESET_B(net155),
    .Q(\tokenflow_inst.i3.ydata[74] ));
 sg13g2_dllrq_1 _2312_ (.D(_0072_),
    .GATE_N(net619),
    .RESET_B(net156),
    .Q(\tokenflow_inst.i3.ydata[75] ));
 sg13g2_dllrq_1 _2313_ (.D(_0073_),
    .GATE_N(net619),
    .RESET_B(net157),
    .Q(\tokenflow_inst.i3.ydata[76] ));
 sg13g2_dllrq_1 _2314_ (.D(_0074_),
    .GATE_N(net618),
    .RESET_B(net158),
    .Q(\tokenflow_inst.i3.ydata[77] ));
 sg13g2_dllrq_1 _2315_ (.D(_0364_),
    .GATE_N(net631),
    .RESET_B(net159),
    .Q(\tokenflow_inst.ii3.i.ydata[0] ));
 sg13g2_dllrq_1 _2316_ (.D(_0375_),
    .GATE_N(net631),
    .RESET_B(net160),
    .Q(\tokenflow_inst.ii3.i.ydata[1] ));
 sg13g2_dllrq_1 _2317_ (.D(_0382_),
    .GATE_N(net631),
    .RESET_B(net161),
    .Q(\tokenflow_inst.ii3.i.ydata[2] ));
 sg13g2_dllrq_1 _2318_ (.D(_0383_),
    .GATE_N(net630),
    .RESET_B(net162),
    .Q(\tokenflow_inst.ii3.i.ydata[3] ));
 sg13g2_dllrq_1 _2319_ (.D(_0384_),
    .GATE_N(net631),
    .RESET_B(net163),
    .Q(\tokenflow_inst.ii3.i.ydata[4] ));
 sg13g2_dllrq_1 _2320_ (.D(_0385_),
    .GATE_N(net631),
    .RESET_B(net164),
    .Q(\tokenflow_inst.ii3.i.ydata[5] ));
 sg13g2_dllrq_1 _2321_ (.D(_0386_),
    .GATE_N(net631),
    .RESET_B(net165),
    .Q(\tokenflow_inst.ii3.i.ydata[6] ));
 sg13g2_dllrq_1 _2322_ (.D(_0387_),
    .GATE_N(net630),
    .RESET_B(net166),
    .Q(\tokenflow_inst.ii3.i.ydata[7] ));
 sg13g2_dllrq_1 _2323_ (.D(_0388_),
    .GATE_N(net630),
    .RESET_B(net167),
    .Q(\tokenflow_inst.ii3.i.ydata[8] ));
 sg13g2_dllrq_1 _2324_ (.D(_0389_),
    .GATE_N(net628),
    .RESET_B(net168),
    .Q(\tokenflow_inst.ii3.i.ydata[9] ));
 sg13g2_dllrq_1 _2325_ (.D(_0365_),
    .GATE_N(net629),
    .RESET_B(net169),
    .Q(\tokenflow_inst.ii3.i.ydata[10] ));
 sg13g2_dllrq_1 _2326_ (.D(_0366_),
    .GATE_N(net629),
    .RESET_B(net170),
    .Q(\tokenflow_inst.ii3.i.ydata[11] ));
 sg13g2_dllrq_1 _2327_ (.D(_0367_),
    .GATE_N(net628),
    .RESET_B(net171),
    .Q(\tokenflow_inst.ii3.i.ydata[12] ));
 sg13g2_dllrq_1 _2328_ (.D(_0368_),
    .GATE_N(net628),
    .RESET_B(net172),
    .Q(\tokenflow_inst.ii3.i.ydata[13] ));
 sg13g2_dllrq_1 _2329_ (.D(_0369_),
    .GATE_N(net628),
    .RESET_B(net173),
    .Q(\tokenflow_inst.ii3.i.ydata[14] ));
 sg13g2_dllrq_1 _2330_ (.D(_0370_),
    .GATE_N(net629),
    .RESET_B(net174),
    .Q(\tokenflow_inst.ii3.i.ydata[15] ));
 sg13g2_dllrq_1 _2331_ (.D(_0371_),
    .GATE_N(net630),
    .RESET_B(net175),
    .Q(\tokenflow_inst.ii3.i.ydata[16] ));
 sg13g2_dllrq_1 _2332_ (.D(_0372_),
    .GATE_N(net630),
    .RESET_B(net176),
    .Q(\tokenflow_inst.ii3.i.ydata[17] ));
 sg13g2_dllrq_1 _2333_ (.D(_0373_),
    .GATE_N(net630),
    .RESET_B(net177),
    .Q(\tokenflow_inst.ii3.i.ydata[18] ));
 sg13g2_dllrq_1 _2334_ (.D(_0374_),
    .GATE_N(net630),
    .RESET_B(net178),
    .Q(\tokenflow_inst.ii3.i.ydata[19] ));
 sg13g2_dllrq_1 _2335_ (.D(_0376_),
    .GATE_N(net629),
    .RESET_B(net179),
    .Q(\tokenflow_inst.ii3.i.ydata[20] ));
 sg13g2_dllrq_1 _2336_ (.D(_0377_),
    .GATE_N(net629),
    .RESET_B(net180),
    .Q(\tokenflow_inst.ii3.i.ydata[21] ));
 sg13g2_dllrq_1 _2337_ (.D(_0378_),
    .GATE_N(net628),
    .RESET_B(net181),
    .Q(\tokenflow_inst.ii3.i.ydata[22] ));
 sg13g2_dllrq_1 _2338_ (.D(_0379_),
    .GATE_N(net628),
    .RESET_B(net182),
    .Q(\tokenflow_inst.ii3.i.ydata[23] ));
 sg13g2_dllrq_1 _2339_ (.D(_0380_),
    .GATE_N(net628),
    .RESET_B(net183),
    .Q(\tokenflow_inst.ii3.i.ydata[24] ));
 sg13g2_dllrq_1 _2340_ (.D(_0381_),
    .GATE_N(net628),
    .RESET_B(net184),
    .Q(\tokenflow_inst.ii3.i.ydata[25] ));
 sg13g2_dllrq_1 _2341_ (.D(_0337_),
    .GATE_N(net613),
    .RESET_B(net185),
    .Q(\tokenflow_inst.ii2.ydata[0] ));
 sg13g2_dllrq_1 _2342_ (.D(_0348_),
    .GATE_N(net614),
    .RESET_B(net186),
    .Q(\tokenflow_inst.ii2.ydata[1] ));
 sg13g2_dllrq_1 _2343_ (.D(_0355_),
    .GATE_N(net613),
    .RESET_B(net187),
    .Q(\tokenflow_inst.ii2.ydata[2] ));
 sg13g2_dllrq_1 _2344_ (.D(_0356_),
    .GATE_N(net613),
    .RESET_B(net188),
    .Q(\tokenflow_inst.ii2.ydata[3] ));
 sg13g2_dllrq_1 _2345_ (.D(_0357_),
    .GATE_N(net613),
    .RESET_B(net189),
    .Q(\tokenflow_inst.ii2.ydata[4] ));
 sg13g2_dllrq_1 _2346_ (.D(_0358_),
    .GATE_N(net613),
    .RESET_B(net190),
    .Q(\tokenflow_inst.ii2.ydata[5] ));
 sg13g2_dllrq_1 _2347_ (.D(_0359_),
    .GATE_N(net613),
    .RESET_B(net191),
    .Q(\tokenflow_inst.ii2.ydata[6] ));
 sg13g2_dllrq_1 _2348_ (.D(_0360_),
    .GATE_N(net614),
    .RESET_B(net192),
    .Q(\tokenflow_inst.ii2.ydata[7] ));
 sg13g2_dllrq_1 _2349_ (.D(_0361_),
    .GATE_N(net614),
    .RESET_B(net193),
    .Q(\tokenflow_inst.ii2.ydata[8] ));
 sg13g2_dllrq_1 _2350_ (.D(_0362_),
    .GATE_N(net611),
    .RESET_B(net194),
    .Q(\tokenflow_inst.ii2.ydata[9] ));
 sg13g2_dllrq_1 _2351_ (.D(_0338_),
    .GATE_N(net612),
    .RESET_B(net195),
    .Q(\tokenflow_inst.ii2.ydata[10] ));
 sg13g2_dllrq_1 _2352_ (.D(_0339_),
    .GATE_N(net612),
    .RESET_B(net196),
    .Q(\tokenflow_inst.ii2.ydata[11] ));
 sg13g2_dllrq_1 _2353_ (.D(_0340_),
    .GATE_N(net611),
    .RESET_B(net197),
    .Q(\tokenflow_inst.ii2.ydata[12] ));
 sg13g2_dllrq_1 _2354_ (.D(_0341_),
    .GATE_N(net611),
    .RESET_B(net198),
    .Q(\tokenflow_inst.ii2.ydata[13] ));
 sg13g2_dllrq_1 _2355_ (.D(_0342_),
    .GATE_N(net611),
    .RESET_B(net199),
    .Q(\tokenflow_inst.ii2.ydata[14] ));
 sg13g2_dllrq_1 _2356_ (.D(_0343_),
    .GATE_N(net612),
    .RESET_B(net200),
    .Q(\tokenflow_inst.ii2.ydata[15] ));
 sg13g2_dllrq_1 _2357_ (.D(_0344_),
    .GATE_N(net614),
    .RESET_B(net201),
    .Q(\tokenflow_inst.ii2.ydata[16] ));
 sg13g2_dllrq_1 _2358_ (.D(_0345_),
    .GATE_N(net614),
    .RESET_B(net202),
    .Q(\tokenflow_inst.ii2.ydata[17] ));
 sg13g2_dllrq_1 _2359_ (.D(_0346_),
    .GATE_N(net614),
    .RESET_B(net203),
    .Q(\tokenflow_inst.ii2.ydata[18] ));
 sg13g2_dllrq_1 _2360_ (.D(_0347_),
    .GATE_N(net614),
    .RESET_B(net204),
    .Q(\tokenflow_inst.ii2.ydata[19] ));
 sg13g2_dllrq_1 _2361_ (.D(_0349_),
    .GATE_N(net612),
    .RESET_B(net205),
    .Q(\tokenflow_inst.ii2.ydata[20] ));
 sg13g2_dllrq_1 _2362_ (.D(_0350_),
    .GATE_N(net612),
    .RESET_B(net206),
    .Q(\tokenflow_inst.ii2.ydata[21] ));
 sg13g2_dllrq_1 _2363_ (.D(_0351_),
    .GATE_N(net611),
    .RESET_B(net207),
    .Q(\tokenflow_inst.ii2.ydata[22] ));
 sg13g2_dllrq_1 _2364_ (.D(_0352_),
    .GATE_N(net611),
    .RESET_B(net208),
    .Q(\tokenflow_inst.ii2.ydata[23] ));
 sg13g2_dllrq_1 _2365_ (.D(_0353_),
    .GATE_N(net611),
    .RESET_B(net209),
    .Q(\tokenflow_inst.ii2.ydata[24] ));
 sg13g2_dllrq_1 _2366_ (.D(_0354_),
    .GATE_N(net611),
    .RESET_B(net210),
    .Q(\tokenflow_inst.ii2.ydata[25] ));
 sg13g2_dllrq_1 _2367_ (.D(_0310_),
    .GATE_N(net596),
    .RESET_B(net211),
    .Q(\tokenflow_inst.ii1.ydata[0] ));
 sg13g2_dllrq_1 _2368_ (.D(_0321_),
    .GATE_N(net596),
    .RESET_B(net212),
    .Q(\tokenflow_inst.ii1.ydata[1] ));
 sg13g2_dllrq_1 _2369_ (.D(_0328_),
    .GATE_N(net596),
    .RESET_B(net213),
    .Q(\tokenflow_inst.ii1.ydata[2] ));
 sg13g2_dllrq_1 _2370_ (.D(_0329_),
    .GATE_N(net596),
    .RESET_B(net214),
    .Q(\tokenflow_inst.ii1.ydata[3] ));
 sg13g2_dllrq_1 _2371_ (.D(_0330_),
    .GATE_N(net595),
    .RESET_B(net215),
    .Q(\tokenflow_inst.ii1.ydata[4] ));
 sg13g2_dllrq_1 _2372_ (.D(_0331_),
    .GATE_N(net595),
    .RESET_B(net216),
    .Q(\tokenflow_inst.ii1.ydata[5] ));
 sg13g2_dllrq_1 _2373_ (.D(_0332_),
    .GATE_N(net595),
    .RESET_B(net217),
    .Q(\tokenflow_inst.ii1.ydata[6] ));
 sg13g2_dllrq_1 _2374_ (.D(_0333_),
    .GATE_N(net596),
    .RESET_B(net218),
    .Q(\tokenflow_inst.ii1.ydata[7] ));
 sg13g2_dllrq_1 _2375_ (.D(_0334_),
    .GATE_N(net595),
    .RESET_B(net219),
    .Q(\tokenflow_inst.ii1.ydata[8] ));
 sg13g2_dllrq_1 _2376_ (.D(_0335_),
    .GATE_N(net593),
    .RESET_B(net220),
    .Q(\tokenflow_inst.ii1.ydata[9] ));
 sg13g2_dllrq_1 _2377_ (.D(_0311_),
    .GATE_N(net594),
    .RESET_B(net221),
    .Q(\tokenflow_inst.ii1.ydata[10] ));
 sg13g2_dllrq_1 _2378_ (.D(_0312_),
    .GATE_N(net594),
    .RESET_B(net222),
    .Q(\tokenflow_inst.ii1.ydata[11] ));
 sg13g2_dllrq_1 _2379_ (.D(_0313_),
    .GATE_N(net593),
    .RESET_B(net223),
    .Q(\tokenflow_inst.ii1.ydata[12] ));
 sg13g2_dllrq_1 _2380_ (.D(_0314_),
    .GATE_N(net593),
    .RESET_B(net224),
    .Q(\tokenflow_inst.ii1.ydata[13] ));
 sg13g2_dllrq_1 _2381_ (.D(_0315_),
    .GATE_N(net593),
    .RESET_B(net225),
    .Q(\tokenflow_inst.ii1.ydata[14] ));
 sg13g2_dllrq_1 _2382_ (.D(_0316_),
    .GATE_N(net594),
    .RESET_B(net226),
    .Q(\tokenflow_inst.ii1.ydata[15] ));
 sg13g2_dllrq_1 _2383_ (.D(_0317_),
    .GATE_N(net595),
    .RESET_B(net227),
    .Q(\tokenflow_inst.ii1.ydata[16] ));
 sg13g2_dllrq_1 _2384_ (.D(_0318_),
    .GATE_N(net595),
    .RESET_B(net228),
    .Q(\tokenflow_inst.ii1.ydata[17] ));
 sg13g2_dllrq_1 _2385_ (.D(_0319_),
    .GATE_N(net595),
    .RESET_B(net229),
    .Q(\tokenflow_inst.ii1.ydata[18] ));
 sg13g2_dllrq_1 _2386_ (.D(_0320_),
    .GATE_N(net595),
    .RESET_B(net230),
    .Q(\tokenflow_inst.ii1.ydata[19] ));
 sg13g2_dllrq_1 _2387_ (.D(_0322_),
    .GATE_N(net594),
    .RESET_B(net231),
    .Q(\tokenflow_inst.ii1.ydata[20] ));
 sg13g2_dllrq_1 _2388_ (.D(_0323_),
    .GATE_N(net594),
    .RESET_B(net232),
    .Q(\tokenflow_inst.ii1.ydata[21] ));
 sg13g2_dllrq_1 _2389_ (.D(_0324_),
    .GATE_N(net593),
    .RESET_B(net233),
    .Q(\tokenflow_inst.ii1.ydata[22] ));
 sg13g2_dllrq_1 _2390_ (.D(_0325_),
    .GATE_N(net593),
    .RESET_B(net234),
    .Q(\tokenflow_inst.ii1.ydata[23] ));
 sg13g2_dllrq_1 _2391_ (.D(_0326_),
    .GATE_N(net593),
    .RESET_B(net235),
    .Q(\tokenflow_inst.ii1.ydata[24] ));
 sg13g2_dllrq_1 _2392_ (.D(_0327_),
    .GATE_N(net593),
    .RESET_B(net236),
    .Q(\tokenflow_inst.ii1.ydata[25] ));
 sg13g2_dllrq_1 _2393_ (.D(_0233_),
    .GATE_N(net580),
    .RESET_B(net237),
    .Q(\tokenflow_inst.i8.ydata[0] ));
 sg13g2_dllrq_1 _2394_ (.D(_0244_),
    .GATE_N(net582),
    .RESET_B(net238),
    .Q(\tokenflow_inst.i8.ydata[1] ));
 sg13g2_dllrq_1 _2395_ (.D(_0255_),
    .GATE_N(net582),
    .RESET_B(net239),
    .Q(\tokenflow_inst.i8.ydata[2] ));
 sg13g2_dllrq_1 _2396_ (.D(_0266_),
    .GATE_N(net580),
    .RESET_B(net240),
    .Q(\tokenflow_inst.i8.ydata[3] ));
 sg13g2_dllrq_1 _2397_ (.D(_0277_),
    .GATE_N(net580),
    .RESET_B(net241),
    .Q(\tokenflow_inst.i8.ydata[4] ));
 sg13g2_dllrq_1 _2398_ (.D(_0286_),
    .GATE_N(net580),
    .RESET_B(net242),
    .Q(\tokenflow_inst.i8.ydata[5] ));
 sg13g2_dllrq_1 _2399_ (.D(_0297_),
    .GATE_N(net577),
    .RESET_B(net243),
    .Q(\tokenflow_inst.i8.ydata[6] ));
 sg13g2_dllrq_1 _2400_ (.D(_0306_),
    .GATE_N(net581),
    .RESET_B(net244),
    .Q(\tokenflow_inst.i8.ydata[7] ));
 sg13g2_dllrq_1 _2401_ (.D(_0307_),
    .GATE_N(net579),
    .RESET_B(net245),
    .Q(\tokenflow_inst.i8.ydata[8] ));
 sg13g2_dllrq_1 _2402_ (.D(_0308_),
    .GATE_N(net571),
    .RESET_B(net246),
    .Q(\tokenflow_inst.i8.ydata[9] ));
 sg13g2_dllrq_1 _2403_ (.D(_0234_),
    .GATE_N(net572),
    .RESET_B(net247),
    .Q(\tokenflow_inst.i8.ydata[10] ));
 sg13g2_dllrq_1 _2404_ (.D(_0235_),
    .GATE_N(net572),
    .RESET_B(net248),
    .Q(\tokenflow_inst.i8.ydata[11] ));
 sg13g2_dllrq_1 _2405_ (.D(_0236_),
    .GATE_N(net570),
    .RESET_B(net249),
    .Q(\tokenflow_inst.i8.ydata[12] ));
 sg13g2_dllrq_1 _2406_ (.D(_0237_),
    .GATE_N(net573),
    .RESET_B(net250),
    .Q(\tokenflow_inst.i8.ydata[13] ));
 sg13g2_dllrq_1 _2407_ (.D(_0238_),
    .GATE_N(net573),
    .RESET_B(net251),
    .Q(\tokenflow_inst.i8.ydata[14] ));
 sg13g2_dllrq_1 _2408_ (.D(_0239_),
    .GATE_N(net574),
    .RESET_B(net252),
    .Q(\tokenflow_inst.i8.ydata[15] ));
 sg13g2_dllrq_1 _2409_ (.D(_0240_),
    .GATE_N(net574),
    .RESET_B(net253),
    .Q(\tokenflow_inst.i8.ydata[16] ));
 sg13g2_dllrq_1 _2410_ (.D(_0241_),
    .GATE_N(net581),
    .RESET_B(net254),
    .Q(\tokenflow_inst.i8.ydata[17] ));
 sg13g2_dllrq_1 _2411_ (.D(_0242_),
    .GATE_N(net581),
    .RESET_B(net255),
    .Q(\tokenflow_inst.i8.ydata[18] ));
 sg13g2_dllrq_1 _2412_ (.D(_0243_),
    .GATE_N(net581),
    .RESET_B(net256),
    .Q(\tokenflow_inst.i8.ydata[19] ));
 sg13g2_dllrq_1 _2413_ (.D(_0245_),
    .GATE_N(net574),
    .RESET_B(net257),
    .Q(\tokenflow_inst.i8.ydata[20] ));
 sg13g2_dllrq_1 _2414_ (.D(_0246_),
    .GATE_N(net575),
    .RESET_B(net258),
    .Q(\tokenflow_inst.i8.ydata[21] ));
 sg13g2_dllrq_1 _2415_ (.D(_0247_),
    .GATE_N(net574),
    .RESET_B(net259),
    .Q(\tokenflow_inst.i8.ydata[22] ));
 sg13g2_dllrq_1 _2416_ (.D(_0248_),
    .GATE_N(net575),
    .RESET_B(net260),
    .Q(\tokenflow_inst.i8.ydata[23] ));
 sg13g2_dllrq_1 _2417_ (.D(_0249_),
    .GATE_N(net575),
    .RESET_B(net261),
    .Q(\tokenflow_inst.i8.ydata[24] ));
 sg13g2_dllrq_1 _2418_ (.D(_0250_),
    .GATE_N(net573),
    .RESET_B(net262),
    .Q(\tokenflow_inst.i8.ydata[25] ));
 sg13g2_dllrq_1 _2419_ (.D(_0251_),
    .GATE_N(net578),
    .RESET_B(net263),
    .Q(\tokenflow_inst.i8.ydata[26] ));
 sg13g2_dllrq_1 _2420_ (.D(_0252_),
    .GATE_N(net578),
    .RESET_B(net264),
    .Q(\tokenflow_inst.i8.ydata[27] ));
 sg13g2_dllrq_1 _2421_ (.D(_0253_),
    .GATE_N(net578),
    .RESET_B(net265),
    .Q(\tokenflow_inst.i8.ydata[28] ));
 sg13g2_dllrq_1 _2422_ (.D(_0254_),
    .GATE_N(net577),
    .RESET_B(net266),
    .Q(\tokenflow_inst.i8.ydata[29] ));
 sg13g2_dllrq_1 _2423_ (.D(_0256_),
    .GATE_N(net577),
    .RESET_B(net267),
    .Q(\tokenflow_inst.i8.ydata[30] ));
 sg13g2_dllrq_1 _2424_ (.D(_0257_),
    .GATE_N(net577),
    .RESET_B(net268),
    .Q(\tokenflow_inst.i8.ydata[31] ));
 sg13g2_dllrq_1 _2425_ (.D(_0258_),
    .GATE_N(net577),
    .RESET_B(net269),
    .Q(\tokenflow_inst.i8.ydata[32] ));
 sg13g2_dllrq_1 _2426_ (.D(_0259_),
    .GATE_N(net576),
    .RESET_B(net270),
    .Q(\tokenflow_inst.i8.ydata[33] ));
 sg13g2_dllrq_1 _2427_ (.D(_0260_),
    .GATE_N(net576),
    .RESET_B(net271),
    .Q(\tokenflow_inst.i8.ydata[34] ));
 sg13g2_dllrq_1 _2428_ (.D(_0261_),
    .GATE_N(net571),
    .RESET_B(net272),
    .Q(\tokenflow_inst.i8.ydata[35] ));
 sg13g2_dllrq_1 _2429_ (.D(_0262_),
    .GATE_N(net571),
    .RESET_B(net273),
    .Q(\tokenflow_inst.i8.ydata[36] ));
 sg13g2_dllrq_1 _2430_ (.D(_0263_),
    .GATE_N(net570),
    .RESET_B(net274),
    .Q(\tokenflow_inst.i8.ydata[37] ));
 sg13g2_dllrq_1 _2431_ (.D(_0264_),
    .GATE_N(net570),
    .RESET_B(net275),
    .Q(\tokenflow_inst.i8.ydata[38] ));
 sg13g2_dllrq_1 _2432_ (.D(_0265_),
    .GATE_N(net570),
    .RESET_B(net276),
    .Q(\tokenflow_inst.i8.ydata[39] ));
 sg13g2_dllrq_1 _2433_ (.D(_0267_),
    .GATE_N(net570),
    .RESET_B(net277),
    .Q(\tokenflow_inst.i8.ydata[40] ));
 sg13g2_dllrq_1 _2434_ (.D(_0268_),
    .GATE_N(net571),
    .RESET_B(net278),
    .Q(\tokenflow_inst.i8.ydata[41] ));
 sg13g2_dllrq_1 _2435_ (.D(_0269_),
    .GATE_N(net571),
    .RESET_B(net279),
    .Q(\tokenflow_inst.i8.ydata[42] ));
 sg13g2_dllrq_1 _2436_ (.D(_0270_),
    .GATE_N(net576),
    .RESET_B(net280),
    .Q(\tokenflow_inst.i8.ydata[43] ));
 sg13g2_dllrq_1 _2437_ (.D(_0271_),
    .GATE_N(net576),
    .RESET_B(net281),
    .Q(\tokenflow_inst.i8.ydata[44] ));
 sg13g2_dllrq_1 _2438_ (.D(_0272_),
    .GATE_N(net576),
    .RESET_B(net282),
    .Q(\tokenflow_inst.i8.ydata[45] ));
 sg13g2_dllrq_1 _2439_ (.D(_0273_),
    .GATE_N(net576),
    .RESET_B(net283),
    .Q(\tokenflow_inst.i8.ydata[46] ));
 sg13g2_dllrq_1 _2440_ (.D(_0274_),
    .GATE_N(net571),
    .RESET_B(net284),
    .Q(\tokenflow_inst.i8.ydata[47] ));
 sg13g2_dllrq_1 _2441_ (.D(_0275_),
    .GATE_N(net571),
    .RESET_B(net285),
    .Q(\tokenflow_inst.i8.ydata[48] ));
 sg13g2_dllrq_1 _2442_ (.D(_0276_),
    .GATE_N(net570),
    .RESET_B(net286),
    .Q(\tokenflow_inst.i8.ydata[49] ));
 sg13g2_dllrq_1 _2443_ (.D(_0278_),
    .GATE_N(net570),
    .RESET_B(net287),
    .Q(\tokenflow_inst.i8.ydata[50] ));
 sg13g2_dllrq_1 _2444_ (.D(_0279_),
    .GATE_N(net580),
    .RESET_B(net288),
    .Q(\tokenflow_inst.i8.ydata[53] ));
 sg13g2_dllrq_1 _2445_ (.D(_0280_),
    .GATE_N(net580),
    .RESET_B(net289),
    .Q(\tokenflow_inst.i8.ydata[54] ));
 sg13g2_dllrq_1 _2446_ (.D(_0281_),
    .GATE_N(net580),
    .RESET_B(net290),
    .Q(\tokenflow_inst.i8.ydata[55] ));
 sg13g2_dllrq_1 _2447_ (.D(_0282_),
    .GATE_N(net580),
    .RESET_B(net291),
    .Q(\tokenflow_inst.i8.ydata[56] ));
 sg13g2_dllrq_1 _2448_ (.D(_0283_),
    .GATE_N(net578),
    .RESET_B(net292),
    .Q(\tokenflow_inst.i8.ydata[57] ));
 sg13g2_dllrq_1 _2449_ (.D(_0284_),
    .GATE_N(net577),
    .RESET_B(net293),
    .Q(\tokenflow_inst.i8.ydata[58] ));
 sg13g2_dllrq_1 _2450_ (.D(_0285_),
    .GATE_N(net576),
    .RESET_B(net294),
    .Q(\tokenflow_inst.i8.ydata[59] ));
 sg13g2_dllrq_1 _2451_ (.D(_0287_),
    .GATE_N(net576),
    .RESET_B(net295),
    .Q(\tokenflow_inst.i8.ydata[60] ));
 sg13g2_dllrq_1 _2452_ (.D(_0288_),
    .GATE_N(net572),
    .RESET_B(net296),
    .Q(\tokenflow_inst.i8.ydata[61] ));
 sg13g2_dllrq_1 _2453_ (.D(_0289_),
    .GATE_N(net571),
    .RESET_B(net297),
    .Q(\tokenflow_inst.i8.ydata[62] ));
 sg13g2_dllrq_1 _2454_ (.D(_0290_),
    .GATE_N(net570),
    .RESET_B(net298),
    .Q(\tokenflow_inst.i8.ydata[63] ));
 sg13g2_dllrq_1 _2455_ (.D(_0291_),
    .GATE_N(net572),
    .RESET_B(net299),
    .Q(\tokenflow_inst.i8.ydata[64] ));
 sg13g2_dllrq_1 _2456_ (.D(_0292_),
    .GATE_N(net573),
    .RESET_B(net300),
    .Q(\tokenflow_inst.i8.ydata[65] ));
 sg13g2_dllrq_1 _2457_ (.D(_0293_),
    .GATE_N(net573),
    .RESET_B(net301),
    .Q(\tokenflow_inst.i8.ydata[66] ));
 sg13g2_dllrq_1 _2458_ (.D(_0294_),
    .GATE_N(net574),
    .RESET_B(net302),
    .Q(\tokenflow_inst.i8.ydata[67] ));
 sg13g2_dllrq_1 _2459_ (.D(_0295_),
    .GATE_N(net574),
    .RESET_B(net303),
    .Q(\tokenflow_inst.i8.ydata[68] ));
 sg13g2_dllrq_1 _2460_ (.D(_0296_),
    .GATE_N(net581),
    .RESET_B(net304),
    .Q(\tokenflow_inst.i8.ydata[69] ));
 sg13g2_dllrq_1 _2461_ (.D(_0298_),
    .GATE_N(net581),
    .RESET_B(net305),
    .Q(\tokenflow_inst.i8.ydata[70] ));
 sg13g2_dllrq_1 _2462_ (.D(_0299_),
    .GATE_N(net581),
    .RESET_B(net306),
    .Q(\tokenflow_inst.i8.ydata[71] ));
 sg13g2_dllrq_1 _2463_ (.D(_0300_),
    .GATE_N(net581),
    .RESET_B(net307),
    .Q(\tokenflow_inst.i8.ydata[72] ));
 sg13g2_dllrq_1 _2464_ (.D(_0301_),
    .GATE_N(net574),
    .RESET_B(net308),
    .Q(\tokenflow_inst.i8.ydata[73] ));
 sg13g2_dllrq_1 _2465_ (.D(_0302_),
    .GATE_N(net574),
    .RESET_B(net309),
    .Q(\tokenflow_inst.i8.ydata[74] ));
 sg13g2_dllrq_1 _2466_ (.D(_0303_),
    .GATE_N(net573),
    .RESET_B(net310),
    .Q(\tokenflow_inst.i8.ydata[75] ));
 sg13g2_dllrq_1 _2467_ (.D(_0304_),
    .GATE_N(net573),
    .RESET_B(net311),
    .Q(\tokenflow_inst.i8.ydata[76] ));
 sg13g2_dllrq_1 _2468_ (.D(_0305_),
    .GATE_N(net573),
    .RESET_B(net312),
    .Q(\tokenflow_inst.i8.ydata[77] ));
 sg13g2_dllrq_1 _2469_ (.D(_0158_),
    .GATE_N(net608),
    .RESET_B(net313),
    .Q(\tokenflow_inst.i78.ydata[0] ));
 sg13g2_dllrq_1 _2470_ (.D(_0169_),
    .GATE_N(net610),
    .RESET_B(net314),
    .Q(\tokenflow_inst.i78.ydata[1] ));
 sg13g2_dllrq_1 _2471_ (.D(_0180_),
    .GATE_N(net609),
    .RESET_B(net315),
    .Q(\tokenflow_inst.i78.ydata[2] ));
 sg13g2_dllrq_1 _2472_ (.D(_0191_),
    .GATE_N(net608),
    .RESET_B(net316),
    .Q(\tokenflow_inst.i78.ydata[3] ));
 sg13g2_dllrq_1 _2473_ (.D(_0202_),
    .GATE_N(net608),
    .RESET_B(net317),
    .Q(\tokenflow_inst.i78.ydata[4] ));
 sg13g2_dllrq_1 _2474_ (.D(_0209_),
    .GATE_N(net608),
    .RESET_B(net318),
    .Q(\tokenflow_inst.i78.ydata[5] ));
 sg13g2_dllrq_1 _2475_ (.D(_0220_),
    .GATE_N(net607),
    .RESET_B(net319),
    .Q(\tokenflow_inst.i78.ydata[6] ));
 sg13g2_dllrq_1 _2476_ (.D(_0229_),
    .GATE_N(net605),
    .RESET_B(net320),
    .Q(\tokenflow_inst.i78.ydata[7] ));
 sg13g2_dllrq_1 _2477_ (.D(_0230_),
    .GATE_N(net605),
    .RESET_B(net321),
    .Q(\tokenflow_inst.i78.ydata[8] ));
 sg13g2_dllrq_1 _2478_ (.D(_0231_),
    .GATE_N(net599),
    .RESET_B(net322),
    .Q(\tokenflow_inst.i78.ydata[9] ));
 sg13g2_dllrq_1 _2479_ (.D(_0159_),
    .GATE_N(net599),
    .RESET_B(net323),
    .Q(\tokenflow_inst.i78.ydata[10] ));
 sg13g2_dllrq_1 _2480_ (.D(_0160_),
    .GATE_N(net599),
    .RESET_B(net324),
    .Q(\tokenflow_inst.i78.ydata[11] ));
 sg13g2_dllrq_1 _2481_ (.D(_0161_),
    .GATE_N(net598),
    .RESET_B(net325),
    .Q(\tokenflow_inst.i78.ydata[12] ));
 sg13g2_dllrq_1 _2482_ (.D(_0162_),
    .GATE_N(net601),
    .RESET_B(net326),
    .Q(\tokenflow_inst.i78.ydata[13] ));
 sg13g2_dllrq_1 _2483_ (.D(_0163_),
    .GATE_N(net601),
    .RESET_B(net327),
    .Q(\tokenflow_inst.i78.ydata[14] ));
 sg13g2_dllrq_1 _2484_ (.D(_0164_),
    .GATE_N(net603),
    .RESET_B(net328),
    .Q(\tokenflow_inst.i78.ydata[15] ));
 sg13g2_dllrq_1 _2485_ (.D(_0165_),
    .GATE_N(net603),
    .RESET_B(net329),
    .Q(\tokenflow_inst.i78.ydata[16] ));
 sg13g2_dllrq_1 _2486_ (.D(_0166_),
    .GATE_N(net609),
    .RESET_B(net330),
    .Q(\tokenflow_inst.i78.ydata[17] ));
 sg13g2_dllrq_1 _2487_ (.D(_0167_),
    .GATE_N(net609),
    .RESET_B(net331),
    .Q(\tokenflow_inst.i78.ydata[18] ));
 sg13g2_dllrq_1 _2488_ (.D(_0168_),
    .GATE_N(net609),
    .RESET_B(net332),
    .Q(\tokenflow_inst.i78.ydata[19] ));
 sg13g2_dllrq_1 _2489_ (.D(_0170_),
    .GATE_N(net603),
    .RESET_B(net333),
    .Q(\tokenflow_inst.i78.ydata[20] ));
 sg13g2_dllrq_1 _2490_ (.D(_0171_),
    .GATE_N(net604),
    .RESET_B(net334),
    .Q(\tokenflow_inst.i78.ydata[21] ));
 sg13g2_dllrq_1 _2491_ (.D(_0172_),
    .GATE_N(net601),
    .RESET_B(net335),
    .Q(\tokenflow_inst.i78.ydata[22] ));
 sg13g2_dllrq_1 _2492_ (.D(_0173_),
    .GATE_N(net602),
    .RESET_B(net336),
    .Q(\tokenflow_inst.i78.ydata[23] ));
 sg13g2_dllrq_1 _2493_ (.D(_0174_),
    .GATE_N(net601),
    .RESET_B(net337),
    .Q(\tokenflow_inst.i78.ydata[24] ));
 sg13g2_dllrq_1 _2494_ (.D(_0175_),
    .GATE_N(net602),
    .RESET_B(net338),
    .Q(\tokenflow_inst.i78.ydata[25] ));
 sg13g2_dllrq_1 _2495_ (.D(_0176_),
    .GATE_N(net606),
    .RESET_B(net339),
    .Q(\tokenflow_inst.i78.ydata[26] ));
 sg13g2_dllrq_1 _2496_ (.D(_0177_),
    .GATE_N(net606),
    .RESET_B(net340),
    .Q(\tokenflow_inst.i78.ydata[27] ));
 sg13g2_dllrq_1 _2497_ (.D(_0178_),
    .GATE_N(net606),
    .RESET_B(net341),
    .Q(\tokenflow_inst.i78.ydata[28] ));
 sg13g2_dllrq_1 _2498_ (.D(_0179_),
    .GATE_N(net606),
    .RESET_B(net342),
    .Q(\tokenflow_inst.i78.ydata[29] ));
 sg13g2_dllrq_1 _2499_ (.D(_0181_),
    .GATE_N(net606),
    .RESET_B(net343),
    .Q(\tokenflow_inst.i78.ydata[30] ));
 sg13g2_dllrq_1 _2500_ (.D(_0182_),
    .GATE_N(net606),
    .RESET_B(net344),
    .Q(\tokenflow_inst.i78.ydata[31] ));
 sg13g2_dllrq_1 _2501_ (.D(_0183_),
    .GATE_N(net607),
    .RESET_B(net345),
    .Q(\tokenflow_inst.i78.ydata[32] ));
 sg13g2_dllrq_1 _2502_ (.D(_0184_),
    .GATE_N(net605),
    .RESET_B(net346),
    .Q(\tokenflow_inst.i78.ydata[33] ));
 sg13g2_dllrq_1 _2503_ (.D(_0185_),
    .GATE_N(net605),
    .RESET_B(net347),
    .Q(\tokenflow_inst.i78.ydata[34] ));
 sg13g2_dllrq_1 _2504_ (.D(_0186_),
    .GATE_N(net599),
    .RESET_B(net348),
    .Q(\tokenflow_inst.i78.ydata[35] ));
 sg13g2_dllrq_1 _2505_ (.D(_0187_),
    .GATE_N(net598),
    .RESET_B(net349),
    .Q(\tokenflow_inst.i78.ydata[36] ));
 sg13g2_dllrq_1 _2506_ (.D(_0188_),
    .GATE_N(net598),
    .RESET_B(net350),
    .Q(\tokenflow_inst.i78.ydata[37] ));
 sg13g2_dllrq_1 _2507_ (.D(_0189_),
    .GATE_N(net598),
    .RESET_B(net351),
    .Q(\tokenflow_inst.i78.ydata[38] ));
 sg13g2_dllrq_1 _2508_ (.D(_0190_),
    .GATE_N(net598),
    .RESET_B(net352),
    .Q(\tokenflow_inst.i78.ydata[39] ));
 sg13g2_dllrq_1 _2509_ (.D(_0192_),
    .GATE_N(net598),
    .RESET_B(net353),
    .Q(\tokenflow_inst.i78.ydata[40] ));
 sg13g2_dllrq_1 _2510_ (.D(_0193_),
    .GATE_N(net600),
    .RESET_B(net354),
    .Q(\tokenflow_inst.i78.ydata[41] ));
 sg13g2_dllrq_1 _2511_ (.D(_0194_),
    .GATE_N(net599),
    .RESET_B(net355),
    .Q(\tokenflow_inst.i78.ydata[42] ));
 sg13g2_dllrq_1 _2512_ (.D(_0195_),
    .GATE_N(net605),
    .RESET_B(net356),
    .Q(\tokenflow_inst.i78.ydata[43] ));
 sg13g2_dllrq_1 _2513_ (.D(_0196_),
    .GATE_N(net605),
    .RESET_B(net357),
    .Q(\tokenflow_inst.i78.ydata[44] ));
 sg13g2_dllrq_1 _2514_ (.D(_0197_),
    .GATE_N(net605),
    .RESET_B(net358),
    .Q(\tokenflow_inst.i78.ydata[45] ));
 sg13g2_dllrq_1 _2515_ (.D(_0198_),
    .GATE_N(net600),
    .RESET_B(net359),
    .Q(\tokenflow_inst.i78.ydata[46] ));
 sg13g2_dllrq_1 _2516_ (.D(_0199_),
    .GATE_N(net600),
    .RESET_B(net360),
    .Q(\tokenflow_inst.i78.ydata[47] ));
 sg13g2_dllrq_1 _2517_ (.D(_0200_),
    .GATE_N(net598),
    .RESET_B(net361),
    .Q(\tokenflow_inst.i78.ydata[48] ));
 sg13g2_dllrq_1 _2518_ (.D(_0201_),
    .GATE_N(net598),
    .RESET_B(net362),
    .Q(\tokenflow_inst.i78.ydata[49] ));
 sg13g2_dllrq_1 _2519_ (.D(_0203_),
    .GATE_N(net608),
    .RESET_B(net363),
    .Q(\tokenflow_inst.i78.ydata[54] ));
 sg13g2_dllrq_1 _2520_ (.D(_0204_),
    .GATE_N(net608),
    .RESET_B(net364),
    .Q(\tokenflow_inst.i78.ydata[55] ));
 sg13g2_dllrq_1 _2521_ (.D(_0205_),
    .GATE_N(net608),
    .RESET_B(net365),
    .Q(\tokenflow_inst.i78.ydata[56] ));
 sg13g2_dllrq_1 _2522_ (.D(_0206_),
    .GATE_N(net608),
    .RESET_B(net366),
    .Q(\tokenflow_inst.i78.ydata[57] ));
 sg13g2_dllrq_1 _2523_ (.D(_0207_),
    .GATE_N(net606),
    .RESET_B(net367),
    .Q(\tokenflow_inst.i78.ydata[58] ));
 sg13g2_dllrq_1 _2524_ (.D(_0208_),
    .GATE_N(net607),
    .RESET_B(net368),
    .Q(\tokenflow_inst.i78.ydata[59] ));
 sg13g2_dllrq_1 _2525_ (.D(_0210_),
    .GATE_N(net605),
    .RESET_B(net369),
    .Q(\tokenflow_inst.i78.ydata[60] ));
 sg13g2_dllrq_1 _2526_ (.D(_0211_),
    .GATE_N(net607),
    .RESET_B(net370),
    .Q(\tokenflow_inst.i78.ydata[61] ));
 sg13g2_dllrq_1 _2527_ (.D(_0212_),
    .GATE_N(net600),
    .RESET_B(net371),
    .Q(\tokenflow_inst.i78.ydata[62] ));
 sg13g2_dllrq_1 _2528_ (.D(_0213_),
    .GATE_N(net599),
    .RESET_B(net372),
    .Q(\tokenflow_inst.i78.ydata[63] ));
 sg13g2_dllrq_1 _2529_ (.D(_0214_),
    .GATE_N(net599),
    .RESET_B(net373),
    .Q(\tokenflow_inst.i78.ydata[64] ));
 sg13g2_dllrq_1 _2530_ (.D(_0215_),
    .GATE_N(net601),
    .RESET_B(net374),
    .Q(\tokenflow_inst.i78.ydata[65] ));
 sg13g2_dllrq_1 _2531_ (.D(_0216_),
    .GATE_N(net601),
    .RESET_B(net375),
    .Q(\tokenflow_inst.i78.ydata[66] ));
 sg13g2_dllrq_1 _2532_ (.D(_0217_),
    .GATE_N(net604),
    .RESET_B(net376),
    .Q(\tokenflow_inst.i78.ydata[67] ));
 sg13g2_dllrq_1 _2533_ (.D(_0218_),
    .GATE_N(net603),
    .RESET_B(net377),
    .Q(\tokenflow_inst.i78.ydata[68] ));
 sg13g2_dllrq_1 _2534_ (.D(_0219_),
    .GATE_N(net609),
    .RESET_B(net378),
    .Q(\tokenflow_inst.i78.ydata[69] ));
 sg13g2_dllrq_1 _2535_ (.D(_0221_),
    .GATE_N(net609),
    .RESET_B(net379),
    .Q(\tokenflow_inst.i78.ydata[70] ));
 sg13g2_dllrq_1 _2536_ (.D(_0222_),
    .GATE_N(net609),
    .RESET_B(net380),
    .Q(\tokenflow_inst.i78.ydata[71] ));
 sg13g2_dllrq_1 _2537_ (.D(_0223_),
    .GATE_N(net603),
    .RESET_B(net381),
    .Q(\tokenflow_inst.i78.ydata[72] ));
 sg13g2_dllrq_1 _2538_ (.D(_0224_),
    .GATE_N(net603),
    .RESET_B(net382),
    .Q(\tokenflow_inst.i78.ydata[73] ));
 sg13g2_dllrq_1 _2539_ (.D(_0225_),
    .GATE_N(net601),
    .RESET_B(net383),
    .Q(\tokenflow_inst.i78.ydata[74] ));
 sg13g2_dllrq_1 _2540_ (.D(_0226_),
    .GATE_N(net602),
    .RESET_B(net384),
    .Q(\tokenflow_inst.i78.ydata[75] ));
 sg13g2_dllrq_1 _2541_ (.D(_0227_),
    .GATE_N(net602),
    .RESET_B(net385),
    .Q(\tokenflow_inst.i78.ydata[76] ));
 sg13g2_tiehi _2159__3 (.L_HI(net3));
 sg13g2_tiehi _2160__4 (.L_HI(net4));
 sg13g2_tiehi _2161__5 (.L_HI(net5));
 sg13g2_tiehi _2162__6 (.L_HI(net6));
 sg13g2_tiehi _2163__7 (.L_HI(net7));
 sg13g2_tiehi _2164__8 (.L_HI(net8));
 sg13g2_tiehi _2165__9 (.L_HI(net9));
 sg13g2_tiehi _2166__10 (.L_HI(net10));
 sg13g2_tiehi _2167__11 (.L_HI(net11));
 sg13g2_tiehi _2168__12 (.L_HI(net12));
 sg13g2_tiehi _2169__13 (.L_HI(net13));
 sg13g2_tiehi _2170__14 (.L_HI(net14));
 sg13g2_tiehi _2171__15 (.L_HI(net15));
 sg13g2_tiehi _2172__16 (.L_HI(net16));
 sg13g2_tiehi _2173__17 (.L_HI(net17));
 sg13g2_tiehi _2174__18 (.L_HI(net18));
 sg13g2_tiehi _2175__19 (.L_HI(net19));
 sg13g2_tiehi _2176__20 (.L_HI(net20));
 sg13g2_tiehi _2177__21 (.L_HI(net21));
 sg13g2_tiehi _2178__22 (.L_HI(net22));
 sg13g2_tiehi _2179__23 (.L_HI(net23));
 sg13g2_tiehi _2180__24 (.L_HI(net24));
 sg13g2_tiehi _2181__25 (.L_HI(net25));
 sg13g2_tiehi _2182__26 (.L_HI(net26));
 sg13g2_tiehi _2183__27 (.L_HI(net27));
 sg13g2_tiehi _2184__28 (.L_HI(net28));
 sg13g2_tiehi _2185__29 (.L_HI(net29));
 sg13g2_tiehi _2186__30 (.L_HI(net30));
 sg13g2_tiehi _2187__31 (.L_HI(net31));
 sg13g2_tiehi _2188__32 (.L_HI(net32));
 sg13g2_tiehi _2189__33 (.L_HI(net33));
 sg13g2_tiehi _2190__34 (.L_HI(net34));
 sg13g2_tiehi _2191__35 (.L_HI(net35));
 sg13g2_tiehi _2192__36 (.L_HI(net36));
 sg13g2_tiehi _2193__37 (.L_HI(net37));
 sg13g2_tiehi _2194__38 (.L_HI(net38));
 sg13g2_tiehi _2195__39 (.L_HI(net39));
 sg13g2_tiehi _2196__40 (.L_HI(net40));
 sg13g2_tiehi _2197__41 (.L_HI(net41));
 sg13g2_tiehi _2198__42 (.L_HI(net42));
 sg13g2_tiehi _2199__43 (.L_HI(net43));
 sg13g2_tiehi _2200__44 (.L_HI(net44));
 sg13g2_tiehi _2201__45 (.L_HI(net45));
 sg13g2_tiehi _2202__46 (.L_HI(net46));
 sg13g2_tiehi _2203__47 (.L_HI(net47));
 sg13g2_tiehi _2204__48 (.L_HI(net48));
 sg13g2_tiehi _2205__49 (.L_HI(net49));
 sg13g2_tiehi _2206__50 (.L_HI(net50));
 sg13g2_tiehi _2207__51 (.L_HI(net51));
 sg13g2_tiehi _2208__52 (.L_HI(net52));
 sg13g2_tiehi _2209__53 (.L_HI(net53));
 sg13g2_tiehi _2210__54 (.L_HI(net54));
 sg13g2_tiehi _2211__55 (.L_HI(net55));
 sg13g2_tiehi _2212__56 (.L_HI(net56));
 sg13g2_tiehi _2213__57 (.L_HI(net57));
 sg13g2_tiehi _2214__58 (.L_HI(net58));
 sg13g2_tiehi _2215__59 (.L_HI(net59));
 sg13g2_tiehi _2216__60 (.L_HI(net60));
 sg13g2_tiehi _2217__61 (.L_HI(net61));
 sg13g2_tiehi _2218__62 (.L_HI(net62));
 sg13g2_tiehi _2219__63 (.L_HI(net63));
 sg13g2_tiehi _2220__64 (.L_HI(net64));
 sg13g2_tiehi _2221__65 (.L_HI(net65));
 sg13g2_tiehi _2222__66 (.L_HI(net66));
 sg13g2_tiehi _2223__67 (.L_HI(net67));
 sg13g2_tiehi _2224__68 (.L_HI(net68));
 sg13g2_tiehi _2225__69 (.L_HI(net69));
 sg13g2_tiehi _2226__70 (.L_HI(net70));
 sg13g2_tiehi _2227__71 (.L_HI(net71));
 sg13g2_tiehi _2228__72 (.L_HI(net72));
 sg13g2_tiehi _2229__73 (.L_HI(net73));
 sg13g2_tiehi _2230__74 (.L_HI(net74));
 sg13g2_tiehi _2231__75 (.L_HI(net75));
 sg13g2_tiehi _2232__76 (.L_HI(net76));
 sg13g2_tiehi _2233__77 (.L_HI(net77));
 sg13g2_tiehi _2234__78 (.L_HI(net78));
 sg13g2_tiehi _2235__79 (.L_HI(net79));
 sg13g2_tiehi _2236__80 (.L_HI(net80));
 sg13g2_tiehi _2237__81 (.L_HI(net81));
 sg13g2_tiehi _2238__82 (.L_HI(net82));
 sg13g2_tiehi _2239__83 (.L_HI(net83));
 sg13g2_tiehi _2240__84 (.L_HI(net84));
 sg13g2_tiehi _2241__85 (.L_HI(net85));
 sg13g2_tiehi _2242__86 (.L_HI(net86));
 sg13g2_tiehi _2243__87 (.L_HI(net87));
 sg13g2_tiehi _2244__88 (.L_HI(net88));
 sg13g2_tiehi _2245__89 (.L_HI(net89));
 sg13g2_tiehi _2246__90 (.L_HI(net90));
 sg13g2_tiehi _2247__91 (.L_HI(net91));
 sg13g2_tiehi _2248__92 (.L_HI(net92));
 sg13g2_tiehi _2249__93 (.L_HI(net93));
 sg13g2_tiehi _2250__94 (.L_HI(net94));
 sg13g2_tiehi _2251__95 (.L_HI(net95));
 sg13g2_tiehi _2252__96 (.L_HI(net96));
 sg13g2_tiehi _2253__97 (.L_HI(net97));
 sg13g2_tiehi _2254__98 (.L_HI(net98));
 sg13g2_tiehi _2255__99 (.L_HI(net99));
 sg13g2_tiehi _2256__100 (.L_HI(net100));
 sg13g2_tiehi _2257__101 (.L_HI(net101));
 sg13g2_tiehi _2258__102 (.L_HI(net102));
 sg13g2_tiehi _2259__103 (.L_HI(net103));
 sg13g2_tiehi _2260__104 (.L_HI(net104));
 sg13g2_tiehi _2261__105 (.L_HI(net105));
 sg13g2_tiehi _2262__106 (.L_HI(net106));
 sg13g2_tiehi _2263__107 (.L_HI(net107));
 sg13g2_tiehi _2264__108 (.L_HI(net108));
 sg13g2_tiehi _2265__109 (.L_HI(net109));
 sg13g2_tiehi _2266__110 (.L_HI(net110));
 sg13g2_tiehi _2267__111 (.L_HI(net111));
 sg13g2_tiehi _2268__112 (.L_HI(net112));
 sg13g2_tiehi _2269__113 (.L_HI(net113));
 sg13g2_tiehi _2270__114 (.L_HI(net114));
 sg13g2_tiehi _2271__115 (.L_HI(net115));
 sg13g2_tiehi _2272__116 (.L_HI(net116));
 sg13g2_tiehi _2273__117 (.L_HI(net117));
 sg13g2_tiehi _2274__118 (.L_HI(net118));
 sg13g2_tiehi _2275__119 (.L_HI(net119));
 sg13g2_tiehi _2276__120 (.L_HI(net120));
 sg13g2_tiehi _2277__121 (.L_HI(net121));
 sg13g2_tiehi _2278__122 (.L_HI(net122));
 sg13g2_tiehi _2279__123 (.L_HI(net123));
 sg13g2_tiehi _2280__124 (.L_HI(net124));
 sg13g2_tiehi _2281__125 (.L_HI(net125));
 sg13g2_tiehi _2282__126 (.L_HI(net126));
 sg13g2_tiehi _2283__127 (.L_HI(net127));
 sg13g2_tiehi _2284__128 (.L_HI(net128));
 sg13g2_tiehi _2285__129 (.L_HI(net129));
 sg13g2_tiehi _2286__130 (.L_HI(net130));
 sg13g2_tiehi _2287__131 (.L_HI(net131));
 sg13g2_tiehi _2288__132 (.L_HI(net132));
 sg13g2_tiehi _2289__133 (.L_HI(net133));
 sg13g2_tiehi _2290__134 (.L_HI(net134));
 sg13g2_tiehi _2291__135 (.L_HI(net135));
 sg13g2_tiehi _2292__136 (.L_HI(net136));
 sg13g2_tiehi _2293__137 (.L_HI(net137));
 sg13g2_tiehi _2294__138 (.L_HI(net138));
 sg13g2_tiehi _2295__139 (.L_HI(net139));
 sg13g2_tiehi _2296__140 (.L_HI(net140));
 sg13g2_tiehi _2297__141 (.L_HI(net141));
 sg13g2_tiehi _2298__142 (.L_HI(net142));
 sg13g2_tiehi _2299__143 (.L_HI(net143));
 sg13g2_tiehi _2300__144 (.L_HI(net144));
 sg13g2_tiehi _2301__145 (.L_HI(net145));
 sg13g2_tiehi _2302__146 (.L_HI(net146));
 sg13g2_tiehi _2303__147 (.L_HI(net147));
 sg13g2_tiehi _2304__148 (.L_HI(net148));
 sg13g2_tiehi _2305__149 (.L_HI(net149));
 sg13g2_tiehi _2306__150 (.L_HI(net150));
 sg13g2_tiehi _2307__151 (.L_HI(net151));
 sg13g2_tiehi _2308__152 (.L_HI(net152));
 sg13g2_tiehi _2309__153 (.L_HI(net153));
 sg13g2_tiehi _2310__154 (.L_HI(net154));
 sg13g2_tiehi _2311__155 (.L_HI(net155));
 sg13g2_tiehi _2312__156 (.L_HI(net156));
 sg13g2_tiehi _2313__157 (.L_HI(net157));
 sg13g2_tiehi _2314__158 (.L_HI(net158));
 sg13g2_tiehi _2315__159 (.L_HI(net159));
 sg13g2_tiehi _2316__160 (.L_HI(net160));
 sg13g2_tiehi _2317__161 (.L_HI(net161));
 sg13g2_tiehi _2318__162 (.L_HI(net162));
 sg13g2_tiehi _2319__163 (.L_HI(net163));
 sg13g2_tiehi _2320__164 (.L_HI(net164));
 sg13g2_tiehi _2321__165 (.L_HI(net165));
 sg13g2_tiehi _2322__166 (.L_HI(net166));
 sg13g2_tiehi _2323__167 (.L_HI(net167));
 sg13g2_tiehi _2324__168 (.L_HI(net168));
 sg13g2_tiehi _2325__169 (.L_HI(net169));
 sg13g2_tiehi _2326__170 (.L_HI(net170));
 sg13g2_tiehi _2327__171 (.L_HI(net171));
 sg13g2_tiehi _2328__172 (.L_HI(net172));
 sg13g2_tiehi _2329__173 (.L_HI(net173));
 sg13g2_tiehi _2330__174 (.L_HI(net174));
 sg13g2_tiehi _2331__175 (.L_HI(net175));
 sg13g2_tiehi _2332__176 (.L_HI(net176));
 sg13g2_tiehi _2333__177 (.L_HI(net177));
 sg13g2_tiehi _2334__178 (.L_HI(net178));
 sg13g2_tiehi _2335__179 (.L_HI(net179));
 sg13g2_tiehi _2336__180 (.L_HI(net180));
 sg13g2_tiehi _2337__181 (.L_HI(net181));
 sg13g2_tiehi _2338__182 (.L_HI(net182));
 sg13g2_tiehi _2339__183 (.L_HI(net183));
 sg13g2_tiehi _2340__184 (.L_HI(net184));
 sg13g2_tiehi _2341__185 (.L_HI(net185));
 sg13g2_tiehi _2342__186 (.L_HI(net186));
 sg13g2_tiehi _2343__187 (.L_HI(net187));
 sg13g2_tiehi _2344__188 (.L_HI(net188));
 sg13g2_tiehi _2345__189 (.L_HI(net189));
 sg13g2_tiehi _2346__190 (.L_HI(net190));
 sg13g2_tiehi _2347__191 (.L_HI(net191));
 sg13g2_tiehi _2348__192 (.L_HI(net192));
 sg13g2_tiehi _2349__193 (.L_HI(net193));
 sg13g2_tiehi _2350__194 (.L_HI(net194));
 sg13g2_tiehi _2351__195 (.L_HI(net195));
 sg13g2_tiehi _2352__196 (.L_HI(net196));
 sg13g2_tiehi _2353__197 (.L_HI(net197));
 sg13g2_tiehi _2354__198 (.L_HI(net198));
 sg13g2_tiehi _2355__199 (.L_HI(net199));
 sg13g2_tiehi _2356__200 (.L_HI(net200));
 sg13g2_tiehi _2357__201 (.L_HI(net201));
 sg13g2_tiehi _2358__202 (.L_HI(net202));
 sg13g2_tiehi _2359__203 (.L_HI(net203));
 sg13g2_tiehi _2360__204 (.L_HI(net204));
 sg13g2_tiehi _2361__205 (.L_HI(net205));
 sg13g2_tiehi _2362__206 (.L_HI(net206));
 sg13g2_tiehi _2363__207 (.L_HI(net207));
 sg13g2_tiehi _2364__208 (.L_HI(net208));
 sg13g2_tiehi _2365__209 (.L_HI(net209));
 sg13g2_tiehi _2366__210 (.L_HI(net210));
 sg13g2_tiehi _2367__211 (.L_HI(net211));
 sg13g2_tiehi _2368__212 (.L_HI(net212));
 sg13g2_tiehi _2369__213 (.L_HI(net213));
 sg13g2_tiehi _2370__214 (.L_HI(net214));
 sg13g2_tiehi _2371__215 (.L_HI(net215));
 sg13g2_tiehi _2372__216 (.L_HI(net216));
 sg13g2_tiehi _2373__217 (.L_HI(net217));
 sg13g2_tiehi _2374__218 (.L_HI(net218));
 sg13g2_tiehi _2375__219 (.L_HI(net219));
 sg13g2_tiehi _2376__220 (.L_HI(net220));
 sg13g2_tiehi _2377__221 (.L_HI(net221));
 sg13g2_tiehi _2378__222 (.L_HI(net222));
 sg13g2_tiehi _2379__223 (.L_HI(net223));
 sg13g2_tiehi _2380__224 (.L_HI(net224));
 sg13g2_tiehi _2381__225 (.L_HI(net225));
 sg13g2_tiehi _2382__226 (.L_HI(net226));
 sg13g2_tiehi _2383__227 (.L_HI(net227));
 sg13g2_tiehi _2384__228 (.L_HI(net228));
 sg13g2_tiehi _2385__229 (.L_HI(net229));
 sg13g2_tiehi _2386__230 (.L_HI(net230));
 sg13g2_tiehi _2387__231 (.L_HI(net231));
 sg13g2_tiehi _2388__232 (.L_HI(net232));
 sg13g2_tiehi _2389__233 (.L_HI(net233));
 sg13g2_tiehi _2390__234 (.L_HI(net234));
 sg13g2_tiehi _2391__235 (.L_HI(net235));
 sg13g2_tiehi _2392__236 (.L_HI(net236));
 sg13g2_tiehi _2393__237 (.L_HI(net237));
 sg13g2_tiehi _2394__238 (.L_HI(net238));
 sg13g2_tiehi _2395__239 (.L_HI(net239));
 sg13g2_tiehi _2396__240 (.L_HI(net240));
 sg13g2_tiehi _2397__241 (.L_HI(net241));
 sg13g2_tiehi _2398__242 (.L_HI(net242));
 sg13g2_tiehi _2399__243 (.L_HI(net243));
 sg13g2_tiehi _2400__244 (.L_HI(net244));
 sg13g2_tiehi _2401__245 (.L_HI(net245));
 sg13g2_tiehi _2402__246 (.L_HI(net246));
 sg13g2_tiehi _2403__247 (.L_HI(net247));
 sg13g2_tiehi _2404__248 (.L_HI(net248));
 sg13g2_tiehi _2405__249 (.L_HI(net249));
 sg13g2_tiehi _2406__250 (.L_HI(net250));
 sg13g2_tiehi _2407__251 (.L_HI(net251));
 sg13g2_tiehi _2408__252 (.L_HI(net252));
 sg13g2_tiehi _2409__253 (.L_HI(net253));
 sg13g2_tiehi _2410__254 (.L_HI(net254));
 sg13g2_tiehi _2411__255 (.L_HI(net255));
 sg13g2_tiehi _2412__256 (.L_HI(net256));
 sg13g2_tiehi _2413__257 (.L_HI(net257));
 sg13g2_tiehi _2414__258 (.L_HI(net258));
 sg13g2_tiehi _2415__259 (.L_HI(net259));
 sg13g2_tiehi _2416__260 (.L_HI(net260));
 sg13g2_tiehi _2417__261 (.L_HI(net261));
 sg13g2_tiehi _2418__262 (.L_HI(net262));
 sg13g2_tiehi _2419__263 (.L_HI(net263));
 sg13g2_tiehi _2420__264 (.L_HI(net264));
 sg13g2_tiehi _2421__265 (.L_HI(net265));
 sg13g2_tiehi _2422__266 (.L_HI(net266));
 sg13g2_tiehi _2423__267 (.L_HI(net267));
 sg13g2_tiehi _2424__268 (.L_HI(net268));
 sg13g2_tiehi _2425__269 (.L_HI(net269));
 sg13g2_tiehi _2426__270 (.L_HI(net270));
 sg13g2_tiehi _2427__271 (.L_HI(net271));
 sg13g2_tiehi _2428__272 (.L_HI(net272));
 sg13g2_tiehi _2429__273 (.L_HI(net273));
 sg13g2_tiehi _2430__274 (.L_HI(net274));
 sg13g2_tiehi _2431__275 (.L_HI(net275));
 sg13g2_tiehi _2432__276 (.L_HI(net276));
 sg13g2_tiehi _2433__277 (.L_HI(net277));
 sg13g2_tiehi _2434__278 (.L_HI(net278));
 sg13g2_tiehi _2435__279 (.L_HI(net279));
 sg13g2_tiehi _2436__280 (.L_HI(net280));
 sg13g2_tiehi _2437__281 (.L_HI(net281));
 sg13g2_tiehi _2438__282 (.L_HI(net282));
 sg13g2_tiehi _2439__283 (.L_HI(net283));
 sg13g2_tiehi _2440__284 (.L_HI(net284));
 sg13g2_tiehi _2441__285 (.L_HI(net285));
 sg13g2_tiehi _2442__286 (.L_HI(net286));
 sg13g2_tiehi _2443__287 (.L_HI(net287));
 sg13g2_tiehi _2444__288 (.L_HI(net288));
 sg13g2_tiehi _2445__289 (.L_HI(net289));
 sg13g2_tiehi _2446__290 (.L_HI(net290));
 sg13g2_tiehi _2447__291 (.L_HI(net291));
 sg13g2_tiehi _2448__292 (.L_HI(net292));
 sg13g2_tiehi _2449__293 (.L_HI(net293));
 sg13g2_tiehi _2450__294 (.L_HI(net294));
 sg13g2_tiehi _2451__295 (.L_HI(net295));
 sg13g2_tiehi _2452__296 (.L_HI(net296));
 sg13g2_tiehi _2453__297 (.L_HI(net297));
 sg13g2_tiehi _2454__298 (.L_HI(net298));
 sg13g2_tiehi _2455__299 (.L_HI(net299));
 sg13g2_tiehi _2456__300 (.L_HI(net300));
 sg13g2_tiehi _2457__301 (.L_HI(net301));
 sg13g2_tiehi _2458__302 (.L_HI(net302));
 sg13g2_tiehi _2459__303 (.L_HI(net303));
 sg13g2_tiehi _2460__304 (.L_HI(net304));
 sg13g2_tiehi _2461__305 (.L_HI(net305));
 sg13g2_tiehi _2462__306 (.L_HI(net306));
 sg13g2_tiehi _2463__307 (.L_HI(net307));
 sg13g2_tiehi _2464__308 (.L_HI(net308));
 sg13g2_tiehi _2465__309 (.L_HI(net309));
 sg13g2_tiehi _2466__310 (.L_HI(net310));
 sg13g2_tiehi _2467__311 (.L_HI(net311));
 sg13g2_tiehi _2468__312 (.L_HI(net312));
 sg13g2_tiehi _2469__313 (.L_HI(net313));
 sg13g2_tiehi _2470__314 (.L_HI(net314));
 sg13g2_tiehi _2471__315 (.L_HI(net315));
 sg13g2_tiehi _2472__316 (.L_HI(net316));
 sg13g2_tiehi _2473__317 (.L_HI(net317));
 sg13g2_tiehi _2474__318 (.L_HI(net318));
 sg13g2_tiehi _2475__319 (.L_HI(net319));
 sg13g2_tiehi _2476__320 (.L_HI(net320));
 sg13g2_tiehi _2477__321 (.L_HI(net321));
 sg13g2_tiehi _2478__322 (.L_HI(net322));
 sg13g2_tiehi _2479__323 (.L_HI(net323));
 sg13g2_tiehi _2480__324 (.L_HI(net324));
 sg13g2_tiehi _2481__325 (.L_HI(net325));
 sg13g2_tiehi _2482__326 (.L_HI(net326));
 sg13g2_tiehi _2483__327 (.L_HI(net327));
 sg13g2_tiehi _2484__328 (.L_HI(net328));
 sg13g2_tiehi _2485__329 (.L_HI(net329));
 sg13g2_tiehi _2486__330 (.L_HI(net330));
 sg13g2_tiehi _2487__331 (.L_HI(net331));
 sg13g2_tiehi _2488__332 (.L_HI(net332));
 sg13g2_tiehi _2489__333 (.L_HI(net333));
 sg13g2_tiehi _2490__334 (.L_HI(net334));
 sg13g2_tiehi _2491__335 (.L_HI(net335));
 sg13g2_tiehi _2492__336 (.L_HI(net336));
 sg13g2_tiehi _2493__337 (.L_HI(net337));
 sg13g2_tiehi _2494__338 (.L_HI(net338));
 sg13g2_tiehi _2495__339 (.L_HI(net339));
 sg13g2_tiehi _2496__340 (.L_HI(net340));
 sg13g2_tiehi _2497__341 (.L_HI(net341));
 sg13g2_tiehi _2498__342 (.L_HI(net342));
 sg13g2_tiehi _2499__343 (.L_HI(net343));
 sg13g2_tiehi _2500__344 (.L_HI(net344));
 sg13g2_tiehi _2501__345 (.L_HI(net345));
 sg13g2_tiehi _2502__346 (.L_HI(net346));
 sg13g2_tiehi _2503__347 (.L_HI(net347));
 sg13g2_tiehi _2504__348 (.L_HI(net348));
 sg13g2_tiehi _2505__349 (.L_HI(net349));
 sg13g2_tiehi _2506__350 (.L_HI(net350));
 sg13g2_tiehi _2507__351 (.L_HI(net351));
 sg13g2_tiehi _2508__352 (.L_HI(net352));
 sg13g2_tiehi _2509__353 (.L_HI(net353));
 sg13g2_tiehi _2510__354 (.L_HI(net354));
 sg13g2_tiehi _2511__355 (.L_HI(net355));
 sg13g2_tiehi _2512__356 (.L_HI(net356));
 sg13g2_tiehi _2513__357 (.L_HI(net357));
 sg13g2_tiehi _2514__358 (.L_HI(net358));
 sg13g2_tiehi _2515__359 (.L_HI(net359));
 sg13g2_tiehi _2516__360 (.L_HI(net360));
 sg13g2_tiehi _2517__361 (.L_HI(net361));
 sg13g2_tiehi _2518__362 (.L_HI(net362));
 sg13g2_tiehi _2519__363 (.L_HI(net363));
 sg13g2_tiehi _2520__364 (.L_HI(net364));
 sg13g2_tiehi _2521__365 (.L_HI(net365));
 sg13g2_tiehi _2522__366 (.L_HI(net366));
 sg13g2_tiehi _2523__367 (.L_HI(net367));
 sg13g2_tiehi _2524__368 (.L_HI(net368));
 sg13g2_tiehi _2525__369 (.L_HI(net369));
 sg13g2_tiehi _2526__370 (.L_HI(net370));
 sg13g2_tiehi _2527__371 (.L_HI(net371));
 sg13g2_tiehi _2528__372 (.L_HI(net372));
 sg13g2_tiehi _2529__373 (.L_HI(net373));
 sg13g2_tiehi _2530__374 (.L_HI(net374));
 sg13g2_tiehi _2531__375 (.L_HI(net375));
 sg13g2_tiehi _2532__376 (.L_HI(net376));
 sg13g2_tiehi _2533__377 (.L_HI(net377));
 sg13g2_tiehi _2534__378 (.L_HI(net378));
 sg13g2_tiehi _2535__379 (.L_HI(net379));
 sg13g2_tiehi _2536__380 (.L_HI(net380));
 sg13g2_tiehi _2537__381 (.L_HI(net381));
 sg13g2_tiehi _2538__382 (.L_HI(net382));
 sg13g2_tiehi _2539__383 (.L_HI(net383));
 sg13g2_tiehi _2540__384 (.L_HI(net384));
 sg13g2_tiehi _2541__385 (.L_HI(net385));
 sg13g2_tiehi tt_um_tommythorn_maxbw_386 (.L_HI(net386));
 sg13g2_tiehi tt_um_tommythorn_maxbw_387 (.L_HI(net387));
 sg13g2_tiehi tt_um_tommythorn_maxbw_388 (.L_HI(net388));
 sg13g2_tiehi tt_um_tommythorn_maxbw_389 (.L_HI(net389));
 sg13g2_tiehi tt_um_tommythorn_maxbw_390 (.L_HI(net390));
 sg13g2_tiehi tt_um_tommythorn_maxbw_391 (.L_HI(net391));
 sg13g2_tiehi tt_um_tommythorn_maxbw_392 (.L_HI(net392));
 sg13g2_tiehi tt_um_tommythorn_maxbw_393 (.L_HI(net393));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_4 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_43 ();
 sg13g2_fill_2 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_tiehi _2158__2 (.L_HI(net2));
 sg13g2_buf_1 _2940_ (.A(\tokenflow_inst.i11.i.d0.inv_chain[0] ),
    .X(\tokenflow_inst.i11.i.d0.inv_chain[1] ));
 sg13g2_buf_1 _2941_ (.A(\tokenflow_inst.i10.d0.inv_chain[0] ),
    .X(\tokenflow_inst.i10.d0.inv_chain[1] ));
 sg13g2_buf_1 _2942_ (.A(\tokenflow_inst.i78.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[1] ));
 sg13g2_buf_1 _2943_ (.A(\tokenflow_inst.i78.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[2] ));
 sg13g2_buf_1 _2944_ (.A(\tokenflow_inst.i78.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[3] ));
 sg13g2_buf_1 _2945_ (.A(net591),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[1] ));
 sg13g2_buf_1 _2946_ (.A(net586),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[2] ));
 sg13g2_buf_1 _2947_ (.A(net588),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[3] ));
 sg13g2_buf_1 _2948_ (.A(net584),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[4] ));
 sg13g2_buf_1 _2949_ (.A(net591),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[5] ));
 sg13g2_buf_1 _2950_ (.A(net584),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[6] ));
 sg13g2_buf_1 _2951_ (.A(net586),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[7] ));
 sg13g2_buf_1 _2952_ (.A(net586),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[8] ));
 sg13g2_buf_1 _2953_ (.A(net591),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[9] ));
 sg13g2_buf_1 _2954_ (.A(net586),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[10] ));
 sg13g2_buf_1 _2955_ (.A(net584),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[11] ));
 sg13g2_buf_1 _2956_ (.A(net586),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[12] ));
 sg13g2_buf_1 _2957_ (.A(net585),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[13] ));
 sg13g2_buf_1 _2958_ (.A(net589),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[14] ));
 sg13g2_buf_1 _2959_ (.A(net584),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[15] ));
 sg13g2_buf_1 _2960_ (.A(net590),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[16] ));
 sg13g2_buf_1 _2961_ (.A(net584),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[17] ));
 sg13g2_buf_1 _2962_ (.A(net585),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[18] ));
 sg13g2_buf_1 _2963_ (.A(net583),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[19] ));
 sg13g2_buf_1 _2964_ (.A(net583),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[20] ));
 sg13g2_buf_1 _2965_ (.A(net585),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[21] ));
 sg13g2_buf_1 _2966_ (.A(net591),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[22] ));
 sg13g2_buf_1 _2967_ (.A(net588),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[23] ));
 sg13g2_buf_1 _2968_ (.A(net585),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[24] ));
 sg13g2_buf_1 _2969_ (.A(net589),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[25] ));
 sg13g2_buf_1 _2970_ (.A(net583),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[26] ));
 sg13g2_buf_1 _2971_ (.A(net588),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[27] ));
 sg13g2_buf_1 _2972_ (.A(net583),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[28] ));
 sg13g2_buf_1 _2973_ (.A(net590),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[29] ));
 sg13g2_buf_1 _2974_ (.A(net591),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[30] ));
 sg13g2_buf_1 _2975_ (.A(net592),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[31] ));
 sg13g2_buf_1 _2976_ (.A(net585),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[32] ));
 sg13g2_buf_1 _2977_ (.A(net585),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[33] ));
 sg13g2_buf_1 _2978_ (.A(net583),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[34] ));
 sg13g2_buf_1 _2979_ (.A(net585),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[35] ));
 sg13g2_buf_1 _2980_ (.A(net587),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[36] ));
 sg13g2_buf_1 _2981_ (.A(net587),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[37] ));
 sg13g2_buf_1 _2982_ (.A(net583),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[38] ));
 sg13g2_buf_1 _2983_ (.A(net587),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[39] ));
 sg13g2_buf_1 _2984_ (.A(net588),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[40] ));
 sg13g2_buf_1 _2985_ (.A(net592),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[41] ));
 sg13g2_buf_1 _2986_ (.A(net588),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[42] ));
 sg13g2_buf_1 _2987_ (.A(net585),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[43] ));
 sg13g2_buf_1 _2988_ (.A(net588),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[44] ));
 sg13g2_buf_1 _2989_ (.A(net583),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[45] ));
 sg13g2_buf_1 _2990_ (.A(net583),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[46] ));
 sg13g2_buf_1 _2991_ (.A(net588),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[47] ));
 sg13g2_buf_1 _2992_ (.A(net584),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[48] ));
 sg13g2_buf_1 _2993_ (.A(net589),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[49] ));
 sg13g2_buf_1 _2994_ (.A(net588),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[50] ));
 sg13g2_buf_1 _2995_ (.A(net586),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[51] ));
 sg13g2_buf_1 _2996_ (.A(net584),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[52] ));
 sg13g2_buf_1 _2997_ (.A(net541),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[1] ));
 sg13g2_buf_1 _2998_ (.A(net545),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[2] ));
 sg13g2_buf_1 _2999_ (.A(net544),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[3] ));
 sg13g2_buf_1 _3000_ (.A(net538),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[4] ));
 sg13g2_buf_1 _3001_ (.A(net541),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[5] ));
 sg13g2_buf_1 _3002_ (.A(net545),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[6] ));
 sg13g2_buf_1 _3003_ (.A(net538),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[7] ));
 sg13g2_buf_1 _3004_ (.A(net542),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[8] ));
 sg13g2_buf_1 _3005_ (.A(net544),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[9] ));
 sg13g2_buf_1 _3006_ (.A(net542),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[10] ));
 sg13g2_buf_1 _3007_ (.A(net539),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[11] ));
 sg13g2_buf_1 _3008_ (.A(net543),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[12] ));
 sg13g2_buf_1 _3009_ (.A(net541),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[13] ));
 sg13g2_buf_1 _3010_ (.A(net542),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[14] ));
 sg13g2_buf_1 _3011_ (.A(net544),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[15] ));
 sg13g2_buf_1 _3012_ (.A(net542),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[16] ));
 sg13g2_buf_1 _3013_ (.A(net540),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[17] ));
 sg13g2_buf_1 _3014_ (.A(net541),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[18] ));
 sg13g2_buf_1 _3015_ (.A(net538),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[19] ));
 sg13g2_buf_1 _3016_ (.A(net540),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[20] ));
 sg13g2_buf_1 _3017_ (.A(net538),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[21] ));
 sg13g2_buf_1 _3018_ (.A(net539),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[22] ));
 sg13g2_buf_1 _3019_ (.A(net542),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[23] ));
 sg13g2_buf_1 _3020_ (.A(net542),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[24] ));
 sg13g2_buf_1 _3021_ (.A(net544),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[25] ));
 sg13g2_buf_1 _3022_ (.A(net543),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[26] ));
 sg13g2_buf_1 _3023_ (.A(net543),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[27] ));
 sg13g2_buf_1 _3024_ (.A(net543),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[28] ));
 sg13g2_buf_1 _3025_ (.A(net539),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[29] ));
 sg13g2_buf_1 _3026_ (.A(net546),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[30] ));
 sg13g2_buf_1 _3027_ (.A(net539),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[31] ));
 sg13g2_buf_1 _3028_ (.A(net538),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[32] ));
 sg13g2_buf_1 _3029_ (.A(net544),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[33] ));
 sg13g2_buf_1 _3030_ (.A(net542),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[34] ));
 sg13g2_buf_1 _3031_ (.A(net538),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[35] ));
 sg13g2_buf_1 _3032_ (.A(net538),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[36] ));
 sg13g2_buf_1 _3033_ (.A(net541),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[37] ));
 sg13g2_buf_1 _3034_ (.A(net541),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[38] ));
 sg13g2_buf_1 _3035_ (.A(net539),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[39] ));
 sg13g2_buf_1 _3036_ (.A(net544),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[40] ));
 sg13g2_buf_1 _3037_ (.A(net540),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[41] ));
 sg13g2_buf_1 _3038_ (.A(net543),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[42] ));
 sg13g2_buf_1 _3039_ (.A(net543),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[43] ));
 sg13g2_buf_1 _3040_ (.A(net539),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[44] ));
 sg13g2_buf_1 _3041_ (.A(net543),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[45] ));
 sg13g2_buf_1 _3042_ (.A(net541),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[46] ));
 sg13g2_buf_1 _3043_ (.A(net542),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[47] ));
 sg13g2_buf_1 _3044_ (.A(net539),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[48] ));
 sg13g2_buf_1 _3045_ (.A(net538),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[49] ));
 sg13g2_buf_1 _3046_ (.A(net541),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[50] ));
 sg13g2_buf_1 _3047_ (.A(net539),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[51] ));
 sg13g2_buf_1 _3048_ (.A(net543),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[52] ));
 sg13g2_buf_1 _3049_ (.A(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[1] ));
 sg13g2_buf_1 _3050_ (.A(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[2] ));
 sg13g2_buf_1 _3051_ (.A(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[3] ));
 sg13g2_buf_1 _3052_ (.A(\tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ));
 sg13g2_buf_1 _3053_ (.A(\tokenflow_inst.ii2.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[1] ));
 sg13g2_buf_1 _3054_ (.A(\tokenflow_inst.ii2.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[2] ));
 sg13g2_buf_1 _3055_ (.A(\tokenflow_inst.ii1.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.ii1.d0_elem.inv_chain[2] ));
 sg13g2_buf_1 _3056_ (.A(\tokenflow_inst.ii1.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.ii1.d0_elem.inv_chain[1] ));
 sg13g2_buf_2 _3057_ (.A(\tokenflow_inst.i3.ydata[11] ),
    .X(uio_out[4]));
 sg13g2_buf_2 _3058_ (.A(\tokenflow_inst.i3.ydata[12] ),
    .X(uio_out[5]));
 sg13g2_buf_1 _3059_ (.A(\tokenflow_inst.i3.ydata[13] ),
    .X(uio_out[6]));
 sg13g2_buf_1 _3060_ (.A(\tokenflow_inst.i3.ydata[14] ),
    .X(uio_out[7]));
 sg13g2_buf_2 _3061_ (.A(\tokenflow_inst.i10.cg.b ),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(net532));
 sg13g2_buf_2 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(\tokenflow_inst.i6.ydata[26] ),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net536),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_1 fanout535 (.A(net536),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(\tokenflow_inst.i6.ydata[26] ),
    .X(net537));
 sg13g2_buf_1 fanout538 (.A(net540),
    .X(net538));
 sg13g2_buf_1 fanout539 (.A(net540),
    .X(net539));
 sg13g2_buf_1 fanout540 (.A(net546),
    .X(net540));
 sg13g2_buf_1 fanout541 (.A(net546),
    .X(net541));
 sg13g2_buf_1 fanout542 (.A(net545),
    .X(net542));
 sg13g2_buf_1 fanout543 (.A(net545),
    .X(net543));
 sg13g2_buf_1 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_1 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_1 fanout546 (.A(\tokenflow_inst.i6.d0_elem.inv_chain[0] ),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net549),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(net553));
 sg13g2_buf_2 fanout550 (.A(net552),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_0157_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net559),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net558),
    .X(net556));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(net558));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(net559));
 sg13g2_buf_2 fanout559 (.A(_0157_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net569),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net563),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net569),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net568),
    .X(net564));
 sg13g2_buf_1 fanout565 (.A(net568),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net568),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(\tokenflow_inst.i8.ydata[26] ),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net572),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_0309_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net575),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net575),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_0309_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net579),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net579),
    .X(net577));
 sg13g2_buf_1 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net582),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net582),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_0309_),
    .X(net582));
 sg13g2_buf_1 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_1 fanout584 (.A(net592),
    .X(net584));
 sg13g2_buf_1 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_1 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_1 fanout587 (.A(net590),
    .X(net587));
 sg13g2_buf_1 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_1 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_1 fanout590 (.A(net591),
    .X(net590));
 sg13g2_buf_1 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_1 fanout592 (.A(\tokenflow_inst.i8.d0_elem.inv_chain[0] ),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(net597),
    .X(net593));
 sg13g2_buf_1 fanout594 (.A(net597),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net597),
    .X(net595));
 sg13g2_buf_1 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_1 fanout597 (.A(_0336_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(net604),
    .X(net599));
 sg13g2_buf_1 fanout600 (.A(net604),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(net603),
    .X(net601));
 sg13g2_buf_1 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(net610),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(net607),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net610),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_0232_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_0363_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_0363_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_0363_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net617),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(net620),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(net627),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(net623),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(net627),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(net626),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(net627),
    .X(net625));
 sg13g2_buf_1 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_0078_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(net632),
    .X(net628));
 sg13g2_buf_1 fanout629 (.A(net632),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(net632),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_1 fanout632 (.A(_0390_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(net635),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net639),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net638),
    .X(net636));
 sg13g2_buf_1 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net645),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(net642),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net645),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_0780_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(net648),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_0779_),
    .X(net648));
 sg13g2_buf_4 fanout649 (.X(net649),
    .A(\tokenflow_inst.i2.cg1.maj.C ));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(net651));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(net656));
 sg13g2_buf_2 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_4 fanout655 (.X(net655),
    .A(net656));
 sg13g2_buf_2 fanout656 (.A(_0738_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(net665),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net665),
    .X(net659));
 sg13g2_buf_1 fanout660 (.A(net665),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(net664),
    .X(net661));
 sg13g2_buf_1 fanout662 (.A(net664),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_1 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net671),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(net668),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(net671),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_1 fanout671 (.A(net708),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net677),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(net677),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(net676),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net676),
    .X(net675));
 sg13g2_buf_1 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_1 fanout677 (.A(net682),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(net682),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(net682),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(net708),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(net687),
    .X(net683));
 sg13g2_buf_1 fanout684 (.A(net687),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net687),
    .X(net685));
 sg13g2_buf_1 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_1 fanout687 (.A(net696),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net696),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net696),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net695),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(net695),
    .X(net693));
 sg13g2_buf_1 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_1 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(net708),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net701),
    .X(net697));
 sg13g2_buf_1 fanout698 (.A(net701),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(net707),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net707),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net707),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(net706),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(net707),
    .X(net706));
 sg13g2_buf_1 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(rst_n),
    .X(net708));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_fill_2 FILLER_0_60 ();
 sg13g2_decap_8 FILLER_0_66 ();
 sg13g2_fill_2 FILLER_0_73 ();
 sg13g2_fill_1 FILLER_0_75 ();
 sg13g2_fill_1 FILLER_0_90 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_4 FILLER_0_117 ();
 sg13g2_fill_1 FILLER_0_121 ();
 sg13g2_fill_1 FILLER_0_138 ();
 sg13g2_decap_4 FILLER_0_169 ();
 sg13g2_fill_1 FILLER_0_173 ();
 sg13g2_decap_4 FILLER_0_178 ();
 sg13g2_fill_1 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_fill_1 FILLER_0_224 ();
 sg13g2_decap_4 FILLER_0_249 ();
 sg13g2_fill_1 FILLER_0_253 ();
 sg13g2_fill_2 FILLER_0_258 ();
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_fill_2 FILLER_0_266 ();
 sg13g2_fill_2 FILLER_0_277 ();
 sg13g2_fill_2 FILLER_0_307 ();
 sg13g2_fill_1 FILLER_0_329 ();
 sg13g2_fill_1 FILLER_0_362 ();
 sg13g2_fill_2 FILLER_0_383 ();
 sg13g2_fill_1 FILLER_0_385 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_fill_1 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_17 ();
 sg13g2_fill_1 FILLER_1_24 ();
 sg13g2_fill_1 FILLER_1_113 ();
 sg13g2_fill_2 FILLER_1_143 ();
 sg13g2_fill_1 FILLER_1_145 ();
 sg13g2_fill_1 FILLER_1_207 ();
 sg13g2_fill_1 FILLER_1_240 ();
 sg13g2_fill_2 FILLER_1_257 ();
 sg13g2_fill_2 FILLER_1_303 ();
 sg13g2_fill_1 FILLER_1_322 ();
 sg13g2_fill_1 FILLER_1_327 ();
 sg13g2_fill_1 FILLER_1_345 ();
 sg13g2_fill_2 FILLER_1_390 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_7 ();
 sg13g2_fill_1 FILLER_2_40 ();
 sg13g2_fill_2 FILLER_2_59 ();
 sg13g2_fill_1 FILLER_2_74 ();
 sg13g2_fill_2 FILLER_2_98 ();
 sg13g2_fill_1 FILLER_2_104 ();
 sg13g2_fill_2 FILLER_2_159 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_fill_2 FILLER_2_182 ();
 sg13g2_fill_1 FILLER_2_184 ();
 sg13g2_decap_4 FILLER_2_214 ();
 sg13g2_fill_2 FILLER_2_218 ();
 sg13g2_fill_1 FILLER_2_229 ();
 sg13g2_fill_2 FILLER_2_235 ();
 sg13g2_fill_1 FILLER_2_237 ();
 sg13g2_fill_1 FILLER_2_264 ();
 sg13g2_fill_2 FILLER_2_281 ();
 sg13g2_fill_2 FILLER_2_301 ();
 sg13g2_fill_1 FILLER_2_303 ();
 sg13g2_fill_2 FILLER_2_333 ();
 sg13g2_fill_1 FILLER_2_335 ();
 sg13g2_fill_2 FILLER_2_352 ();
 sg13g2_fill_1 FILLER_2_359 ();
 sg13g2_fill_2 FILLER_2_396 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_21 ();
 sg13g2_fill_1 FILLER_3_23 ();
 sg13g2_fill_1 FILLER_3_54 ();
 sg13g2_fill_2 FILLER_3_87 ();
 sg13g2_fill_2 FILLER_3_105 ();
 sg13g2_fill_1 FILLER_3_107 ();
 sg13g2_fill_1 FILLER_3_132 ();
 sg13g2_fill_2 FILLER_3_138 ();
 sg13g2_fill_2 FILLER_3_189 ();
 sg13g2_fill_2 FILLER_3_200 ();
 sg13g2_fill_1 FILLER_3_202 ();
 sg13g2_fill_1 FILLER_3_212 ();
 sg13g2_fill_2 FILLER_3_218 ();
 sg13g2_fill_1 FILLER_3_220 ();
 sg13g2_fill_2 FILLER_3_241 ();
 sg13g2_fill_2 FILLER_3_337 ();
 sg13g2_fill_2 FILLER_3_344 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_4 ();
 sg13g2_fill_2 FILLER_4_31 ();
 sg13g2_fill_2 FILLER_4_73 ();
 sg13g2_fill_1 FILLER_4_75 ();
 sg13g2_fill_1 FILLER_4_93 ();
 sg13g2_fill_2 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_120 ();
 sg13g2_fill_2 FILLER_4_135 ();
 sg13g2_fill_2 FILLER_4_162 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_decap_8 FILLER_4_178 ();
 sg13g2_fill_2 FILLER_4_185 ();
 sg13g2_fill_1 FILLER_4_187 ();
 sg13g2_decap_4 FILLER_4_235 ();
 sg13g2_fill_1 FILLER_4_239 ();
 sg13g2_fill_2 FILLER_4_245 ();
 sg13g2_fill_1 FILLER_4_247 ();
 sg13g2_fill_2 FILLER_4_278 ();
 sg13g2_fill_1 FILLER_4_280 ();
 sg13g2_fill_2 FILLER_4_301 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_fill_2 FILLER_4_337 ();
 sg13g2_fill_2 FILLER_4_343 ();
 sg13g2_fill_1 FILLER_4_376 ();
 sg13g2_fill_2 FILLER_4_381 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_22 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_decap_4 FILLER_5_113 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_fill_2 FILLER_5_157 ();
 sg13g2_fill_1 FILLER_5_184 ();
 sg13g2_decap_4 FILLER_5_190 ();
 sg13g2_fill_1 FILLER_5_194 ();
 sg13g2_decap_4 FILLER_5_208 ();
 sg13g2_fill_2 FILLER_5_212 ();
 sg13g2_decap_4 FILLER_5_218 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_fill_2 FILLER_5_304 ();
 sg13g2_fill_1 FILLER_5_328 ();
 sg13g2_fill_2 FILLER_5_382 ();
 sg13g2_fill_1 FILLER_5_396 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_27 ();
 sg13g2_fill_2 FILLER_6_44 ();
 sg13g2_fill_1 FILLER_6_46 ();
 sg13g2_decap_4 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_67 ();
 sg13g2_fill_2 FILLER_6_94 ();
 sg13g2_fill_1 FILLER_6_96 ();
 sg13g2_fill_2 FILLER_6_137 ();
 sg13g2_fill_1 FILLER_6_155 ();
 sg13g2_fill_1 FILLER_6_161 ();
 sg13g2_decap_4 FILLER_6_178 ();
 sg13g2_decap_4 FILLER_6_219 ();
 sg13g2_fill_2 FILLER_6_223 ();
 sg13g2_fill_1 FILLER_6_251 ();
 sg13g2_fill_1 FILLER_6_267 ();
 sg13g2_decap_4 FILLER_6_280 ();
 sg13g2_fill_2 FILLER_6_284 ();
 sg13g2_fill_2 FILLER_6_323 ();
 sg13g2_fill_1 FILLER_6_325 ();
 sg13g2_fill_2 FILLER_6_342 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_fill_2 FILLER_6_375 ();
 sg13g2_fill_1 FILLER_6_377 ();
 sg13g2_fill_1 FILLER_6_386 ();
 sg13g2_fill_2 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_27 ();
 sg13g2_fill_1 FILLER_7_29 ();
 sg13g2_decap_4 FILLER_7_34 ();
 sg13g2_fill_1 FILLER_7_38 ();
 sg13g2_fill_2 FILLER_7_92 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_100 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_134 ();
 sg13g2_fill_1 FILLER_7_140 ();
 sg13g2_fill_1 FILLER_7_157 ();
 sg13g2_decap_8 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_194 ();
 sg13g2_fill_2 FILLER_7_233 ();
 sg13g2_fill_1 FILLER_7_235 ();
 sg13g2_fill_2 FILLER_7_241 ();
 sg13g2_fill_1 FILLER_7_243 ();
 sg13g2_decap_4 FILLER_7_286 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_fill_2 FILLER_7_316 ();
 sg13g2_fill_1 FILLER_7_318 ();
 sg13g2_fill_2 FILLER_7_347 ();
 sg13g2_fill_1 FILLER_7_349 ();
 sg13g2_fill_2 FILLER_7_386 ();
 sg13g2_fill_2 FILLER_7_396 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_33 ();
 sg13g2_fill_1 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_41 ();
 sg13g2_fill_1 FILLER_8_46 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_81 ();
 sg13g2_fill_1 FILLER_8_87 ();
 sg13g2_fill_1 FILLER_8_102 ();
 sg13g2_fill_2 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_118 ();
 sg13g2_decap_4 FILLER_8_137 ();
 sg13g2_decap_4 FILLER_8_146 ();
 sg13g2_fill_1 FILLER_8_150 ();
 sg13g2_decap_4 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_169 ();
 sg13g2_fill_2 FILLER_8_197 ();
 sg13g2_fill_1 FILLER_8_199 ();
 sg13g2_fill_2 FILLER_8_213 ();
 sg13g2_fill_1 FILLER_8_215 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_decap_4 FILLER_8_248 ();
 sg13g2_fill_1 FILLER_8_252 ();
 sg13g2_fill_1 FILLER_8_265 ();
 sg13g2_fill_2 FILLER_8_270 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_324 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_fill_2 FILLER_8_363 ();
 sg13g2_fill_1 FILLER_8_365 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_fill_2 FILLER_9_26 ();
 sg13g2_fill_1 FILLER_9_28 ();
 sg13g2_fill_1 FILLER_9_52 ();
 sg13g2_fill_1 FILLER_9_57 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_fill_1 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_187 ();
 sg13g2_fill_2 FILLER_9_204 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_decap_4 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_237 ();
 sg13g2_fill_2 FILLER_9_250 ();
 sg13g2_fill_1 FILLER_9_283 ();
 sg13g2_fill_2 FILLER_9_296 ();
 sg13g2_fill_1 FILLER_9_303 ();
 sg13g2_fill_2 FILLER_9_312 ();
 sg13g2_fill_1 FILLER_9_314 ();
 sg13g2_fill_2 FILLER_9_324 ();
 sg13g2_fill_1 FILLER_9_326 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_363 ();
 sg13g2_fill_1 FILLER_9_365 ();
 sg13g2_fill_2 FILLER_9_382 ();
 sg13g2_fill_2 FILLER_9_392 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_17 ();
 sg13g2_fill_1 FILLER_10_19 ();
 sg13g2_decap_4 FILLER_10_66 ();
 sg13g2_fill_1 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_80 ();
 sg13g2_fill_2 FILLER_10_127 ();
 sg13g2_fill_1 FILLER_10_129 ();
 sg13g2_decap_4 FILLER_10_135 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_1 FILLER_10_150 ();
 sg13g2_fill_2 FILLER_10_156 ();
 sg13g2_fill_2 FILLER_10_177 ();
 sg13g2_fill_2 FILLER_10_195 ();
 sg13g2_fill_1 FILLER_10_197 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_260 ();
 sg13g2_fill_2 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_284 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_fill_2 FILLER_10_295 ();
 sg13g2_fill_1 FILLER_10_297 ();
 sg13g2_fill_2 FILLER_10_303 ();
 sg13g2_decap_4 FILLER_10_329 ();
 sg13g2_fill_2 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_374 ();
 sg13g2_fill_2 FILLER_10_396 ();
 sg13g2_fill_1 FILLER_10_402 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_38 ();
 sg13g2_fill_1 FILLER_11_40 ();
 sg13g2_fill_2 FILLER_11_57 ();
 sg13g2_fill_2 FILLER_11_104 ();
 sg13g2_fill_1 FILLER_11_106 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_fill_2 FILLER_11_142 ();
 sg13g2_fill_1 FILLER_11_144 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_decap_8 FILLER_11_202 ();
 sg13g2_decap_4 FILLER_11_233 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_259 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_fill_2 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_317 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_fill_2 FILLER_11_370 ();
 sg13g2_fill_1 FILLER_11_372 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_2 FILLER_12_12 ();
 sg13g2_fill_2 FILLER_12_27 ();
 sg13g2_fill_1 FILLER_12_29 ();
 sg13g2_fill_2 FILLER_12_34 ();
 sg13g2_fill_1 FILLER_12_36 ();
 sg13g2_fill_2 FILLER_12_53 ();
 sg13g2_fill_1 FILLER_12_55 ();
 sg13g2_fill_2 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_fill_1 FILLER_12_155 ();
 sg13g2_fill_2 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_313 ();
 sg13g2_fill_2 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_38 ();
 sg13g2_fill_1 FILLER_13_40 ();
 sg13g2_fill_2 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_80 ();
 sg13g2_fill_2 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_145 ();
 sg13g2_fill_1 FILLER_13_151 ();
 sg13g2_fill_2 FILLER_13_168 ();
 sg13g2_fill_1 FILLER_13_170 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_decap_4 FILLER_13_231 ();
 sg13g2_fill_2 FILLER_13_235 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_256 ();
 sg13g2_fill_2 FILLER_13_274 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_343 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_1 FILLER_13_376 ();
 sg13g2_fill_2 FILLER_13_387 ();
 sg13g2_fill_1 FILLER_13_389 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_12 ();
 sg13g2_fill_1 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_43 ();
 sg13g2_fill_2 FILLER_14_48 ();
 sg13g2_fill_1 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_103 ();
 sg13g2_fill_2 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_137 ();
 sg13g2_fill_2 FILLER_14_162 ();
 sg13g2_fill_1 FILLER_14_164 ();
 sg13g2_fill_1 FILLER_14_173 ();
 sg13g2_fill_2 FILLER_14_199 ();
 sg13g2_fill_2 FILLER_14_222 ();
 sg13g2_fill_2 FILLER_14_288 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_36 ();
 sg13g2_fill_1 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_55 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_2 FILLER_15_86 ();
 sg13g2_fill_2 FILLER_15_97 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_fill_2 FILLER_15_159 ();
 sg13g2_fill_1 FILLER_15_161 ();
 sg13g2_decap_4 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_189 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_fill_2 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_fill_2 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_292 ();
 sg13g2_decap_4 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_decap_4 FILLER_15_312 ();
 sg13g2_fill_1 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_347 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_378 ();
 sg13g2_fill_2 FILLER_15_387 ();
 sg13g2_fill_1 FILLER_15_402 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_1 FILLER_16_34 ();
 sg13g2_fill_2 FILLER_16_48 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_93 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_116 ();
 sg13g2_fill_1 FILLER_16_137 ();
 sg13g2_fill_2 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_164 ();
 sg13g2_decap_4 FILLER_16_201 ();
 sg13g2_decap_4 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_fill_1 FILLER_16_269 ();
 sg13g2_fill_2 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_fill_1 FILLER_16_389 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_22 ();
 sg13g2_fill_1 FILLER_17_29 ();
 sg13g2_fill_1 FILLER_17_53 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_fill_1 FILLER_17_79 ();
 sg13g2_fill_1 FILLER_17_94 ();
 sg13g2_decap_8 FILLER_17_100 ();
 sg13g2_fill_2 FILLER_17_107 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_fill_2 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_decap_8 FILLER_17_241 ();
 sg13g2_decap_4 FILLER_17_265 ();
 sg13g2_decap_4 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_fill_1 FILLER_17_385 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_26 ();
 sg13g2_fill_1 FILLER_18_31 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_fill_2 FILLER_18_122 ();
 sg13g2_fill_1 FILLER_18_143 ();
 sg13g2_decap_4 FILLER_18_204 ();
 sg13g2_fill_2 FILLER_18_208 ();
 sg13g2_decap_4 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_decap_4 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_332 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_12 ();
 sg13g2_fill_2 FILLER_19_30 ();
 sg13g2_fill_1 FILLER_19_32 ();
 sg13g2_fill_2 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_decap_4 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_decap_4 FILLER_19_113 ();
 sg13g2_fill_2 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_128 ();
 sg13g2_fill_2 FILLER_19_164 ();
 sg13g2_fill_1 FILLER_19_166 ();
 sg13g2_decap_4 FILLER_19_171 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_253 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_decap_4 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_297 ();
 sg13g2_fill_1 FILLER_19_302 ();
 sg13g2_fill_2 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_34 ();
 sg13g2_fill_2 FILLER_20_46 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_2 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_143 ();
 sg13g2_fill_1 FILLER_20_145 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_decap_4 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_228 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_fill_2 FILLER_20_323 ();
 sg13g2_fill_1 FILLER_20_325 ();
 sg13g2_fill_1 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_375 ();
 sg13g2_fill_2 FILLER_20_382 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_1 FILLER_21_52 ();
 sg13g2_fill_2 FILLER_21_67 ();
 sg13g2_fill_1 FILLER_21_69 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_147 ();
 sg13g2_decap_4 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_220 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_fill_2 FILLER_21_297 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_30 ();
 sg13g2_fill_2 FILLER_22_48 ();
 sg13g2_fill_2 FILLER_22_55 ();
 sg13g2_fill_2 FILLER_22_81 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_fill_2 FILLER_22_131 ();
 sg13g2_fill_1 FILLER_22_133 ();
 sg13g2_decap_4 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_decap_4 FILLER_22_165 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_fill_1 FILLER_22_258 ();
 sg13g2_decap_4 FILLER_22_296 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_336 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_fill_2 FILLER_22_367 ();
 sg13g2_fill_2 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_388 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_12 ();
 sg13g2_fill_1 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_33 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_decap_4 FILLER_23_96 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_decap_4 FILLER_23_125 ();
 sg13g2_decap_4 FILLER_23_134 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_192 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_decap_4 FILLER_23_240 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_decap_4 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_fill_2 FILLER_23_348 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_402 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_29 ();
 sg13g2_fill_1 FILLER_24_33 ();
 sg13g2_fill_2 FILLER_24_59 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_107 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_157 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_199 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_216 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_fill_1 FILLER_24_241 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_decap_4 FILLER_24_384 ();
 sg13g2_fill_1 FILLER_24_388 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_2 FILLER_25_19 ();
 sg13g2_fill_2 FILLER_25_101 ();
 sg13g2_fill_2 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_142 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_227 ();
 sg13g2_fill_2 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_251 ();
 sg13g2_fill_1 FILLER_25_253 ();
 sg13g2_fill_2 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_265 ();
 sg13g2_fill_1 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_decap_4 FILLER_25_321 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_fill_1 FILLER_25_336 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_45 ();
 sg13g2_fill_1 FILLER_26_52 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_decap_4 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_299 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_fill_2 FILLER_26_355 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_383 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_25 ();
 sg13g2_fill_1 FILLER_27_27 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_fill_1 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_2 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_fill_2 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_decap_4 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_241 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_decap_8 FILLER_27_278 ();
 sg13g2_decap_4 FILLER_27_285 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_fill_2 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_27 ();
 sg13g2_fill_2 FILLER_28_40 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_53 ();
 sg13g2_fill_2 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_fill_2 FILLER_28_87 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_fill_2 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_166 ();
 sg13g2_decap_4 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_fill_2 FILLER_28_228 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_328 ();
 sg13g2_fill_2 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_367 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_54 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_61 ();
 sg13g2_decap_8 FILLER_29_73 ();
 sg13g2_fill_1 FILLER_29_80 ();
 sg13g2_decap_4 FILLER_29_94 ();
 sg13g2_decap_4 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_decap_4 FILLER_29_236 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_268 ();
 sg13g2_decap_4 FILLER_29_279 ();
 sg13g2_decap_4 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_decap_4 FILLER_30_30 ();
 sg13g2_fill_2 FILLER_30_34 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_248 ();
 sg13g2_fill_2 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_307 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_339 ();
 sg13g2_fill_2 FILLER_30_352 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_decap_4 FILLER_31_75 ();
 sg13g2_decap_4 FILLER_31_87 ();
 sg13g2_fill_1 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_29 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_2 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_fill_1 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_278 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_390 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_2 FILLER_33_24 ();
 sg13g2_fill_2 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_51 ();
 sg13g2_fill_2 FILLER_33_57 ();
 sg13g2_fill_1 FILLER_33_64 ();
 sg13g2_fill_2 FILLER_33_86 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_decap_4 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_decap_4 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_1 FILLER_34_38 ();
 sg13g2_fill_1 FILLER_34_68 ();
 sg13g2_fill_1 FILLER_34_74 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_99 ();
 sg13g2_fill_2 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_fill_2 FILLER_34_148 ();
 sg13g2_fill_2 FILLER_34_171 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_decap_4 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_332 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_367 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_fill_2 FILLER_34_385 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_1 FILLER_35_20 ();
 sg13g2_fill_2 FILLER_35_26 ();
 sg13g2_fill_1 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_2 FILLER_35_62 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_fill_2 FILLER_35_81 ();
 sg13g2_fill_1 FILLER_35_83 ();
 sg13g2_fill_1 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_decap_4 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_348 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_12 ();
 sg13g2_fill_2 FILLER_36_37 ();
 sg13g2_fill_1 FILLER_36_49 ();
 sg13g2_fill_1 FILLER_36_55 ();
 sg13g2_fill_2 FILLER_36_68 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_fill_2 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_decap_4 FILLER_36_130 ();
 sg13g2_fill_2 FILLER_36_157 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_165 ();
 sg13g2_fill_2 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_183 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_205 ();
 sg13g2_decap_4 FILLER_36_211 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_371 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_fill_2 FILLER_36_403 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_166 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_211 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_fill_2 FILLER_37_375 ();
 sg13g2_fill_1 FILLER_37_377 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_61 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_110 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_149 ();
 sg13g2_decap_8 FILLER_38_169 ();
 sg13g2_fill_2 FILLER_38_176 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_211 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_2 FILLER_38_298 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net386;
 assign uio_oe[1] = net387;
 assign uio_oe[2] = net388;
 assign uio_oe[3] = net389;
 assign uio_oe[4] = net390;
 assign uio_oe[5] = net391;
 assign uio_oe[6] = net392;
 assign uio_oe[7] = net393;
endmodule

module tt_um_cellular_alchemist (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire net17;
 wire net18;
 wire net19;
 wire \hopfield_inst.active_neuron[0] ;
 wire \hopfield_inst.active_neuron[1] ;
 wire \hopfield_inst.active_neuron[2] ;
 wire \hopfield_inst.currents[0] ;
 wire \hopfield_inst.currents[1] ;
 wire \hopfield_inst.currents[2] ;
 wire \hopfield_inst.currents[3] ;
 wire \hopfield_inst.currents[4] ;
 wire \hopfield_inst.currents[5] ;
 wire \hopfield_inst.currents[6] ;
 wire \hopfield_inst.currents[7] ;
 wire \hopfield_inst.learning_inst.counter[0] ;
 wire \hopfield_inst.learning_inst.counter[1] ;
 wire \hopfield_inst.learning_inst.counter[2] ;
 wire \hopfield_inst.learning_inst.state[0] ;
 wire \hopfield_inst.learning_inst.state[1] ;
 wire \hopfield_inst.learning_inst.state[2] ;
 wire \hopfield_inst.learning_inst.temp_weight[0] ;
 wire \hopfield_inst.learning_inst.temp_weight[1] ;
 wire \hopfield_inst.learning_inst.temp_weight[2] ;
 wire \hopfield_inst.learning_inst.temp_weight[3] ;
 wire \hopfield_inst.learning_inst.temp_weight[4] ;
 wire \hopfield_inst.learning_inst.temp_weight[5] ;
 wire \hopfield_inst.learning_inst.weights[17][0] ;
 wire \hopfield_inst.learning_inst.weights[17][1] ;
 wire \hopfield_inst.learning_inst.weights[17][2] ;
 wire \hopfield_inst.learning_inst.weights[17][3] ;
 wire \hopfield_inst.learning_inst.weights[1][0] ;
 wire \hopfield_inst.learning_inst.weights[1][1] ;
 wire \hopfield_inst.learning_inst.weights[1][2] ;
 wire \hopfield_inst.learning_inst.weights[1][3] ;
 wire \hopfield_inst.learning_inst.weights[25][0] ;
 wire \hopfield_inst.learning_inst.weights[25][1] ;
 wire \hopfield_inst.learning_inst.weights[25][2] ;
 wire \hopfield_inst.learning_inst.weights[25][3] ;
 wire \hopfield_inst.learning_inst.weights[33][0] ;
 wire \hopfield_inst.learning_inst.weights[33][1] ;
 wire \hopfield_inst.learning_inst.weights[33][2] ;
 wire \hopfield_inst.learning_inst.weights[33][3] ;
 wire \hopfield_inst.learning_inst.weights[41][0] ;
 wire \hopfield_inst.learning_inst.weights[41][1] ;
 wire \hopfield_inst.learning_inst.weights[41][2] ;
 wire \hopfield_inst.learning_inst.weights[41][3] ;
 wire \hopfield_inst.learning_inst.weights[9][0] ;
 wire \hopfield_inst.learning_inst.weights[9][1] ;
 wire \hopfield_inst.learning_inst.weights[9][2] ;
 wire \hopfield_inst.learning_inst.weights[9][3] ;
 wire \hopfield_inst.neuron_inst.u[0] ;
 wire \hopfield_inst.neuron_inst.u[1] ;
 wire \hopfield_inst.neuron_inst.u[2] ;
 wire \hopfield_inst.neuron_inst.u[3] ;
 wire \hopfield_inst.neuron_inst.u[4] ;
 wire \hopfield_inst.neuron_inst.u[5] ;
 wire \hopfield_inst.neuron_inst.u[6] ;
 wire \hopfield_inst.neuron_inst.u[7] ;
 wire \hopfield_inst.neuron_inst.v[0] ;
 wire \hopfield_inst.neuron_inst.v[1] ;
 wire \hopfield_inst.neuron_inst.v[2] ;
 wire \hopfield_inst.neuron_inst.v[3] ;
 wire \hopfield_inst.neuron_inst.v[4] ;
 wire \hopfield_inst.neuron_inst.v[5] ;
 wire \hopfield_inst.neuron_inst.v[6] ;
 wire \hopfield_inst.neuron_inst.v[7] ;
 wire \temp_activity_count[0] ;
 wire \temp_activity_count[1] ;
 wire \temp_activity_count[2] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_0_clk;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;

 sg13g2_inv_1 _436_ (.Y(_088_),
    .A(net78));
 sg13g2_inv_1 _437_ (.Y(_089_),
    .A(uio_out[7]));
 sg13g2_inv_1 _438_ (.Y(_090_),
    .A(net68));
 sg13g2_inv_1 _439_ (.Y(_091_),
    .A(\hopfield_inst.neuron_inst.u[1] ));
 sg13g2_inv_1 _440_ (.Y(_092_),
    .A(\hopfield_inst.neuron_inst.v[5] ));
 sg13g2_inv_1 _441_ (.Y(_093_),
    .A(\hopfield_inst.currents[3] ));
 sg13g2_inv_1 _442_ (.Y(_094_),
    .A(\hopfield_inst.neuron_inst.u[3] ));
 sg13g2_inv_1 _443_ (.Y(_095_),
    .A(\hopfield_inst.currents[5] ));
 sg13g2_inv_1 _444_ (.Y(_096_),
    .A(net75));
 sg13g2_inv_1 _445_ (.Y(_097_),
    .A(net114));
 sg13g2_inv_1 _446_ (.Y(_098_),
    .A(net31));
 sg13g2_inv_1 _447_ (.Y(_099_),
    .A(net33));
 sg13g2_inv_1 _448_ (.Y(_100_),
    .A(net37));
 sg13g2_inv_1 _449_ (.Y(_101_),
    .A(net35));
 sg13g2_inv_1 _450_ (.Y(_102_),
    .A(net129));
 sg13g2_nor2b_1 _451_ (.A(\hopfield_inst.neuron_inst.u[6] ),
    .B_N(\hopfield_inst.currents[6] ),
    .Y(_103_));
 sg13g2_nor2b_1 _452_ (.A(\hopfield_inst.neuron_inst.u[4] ),
    .B_N(\hopfield_inst.currents[4] ),
    .Y(_104_));
 sg13g2_nor2b_1 _453_ (.A(\hopfield_inst.neuron_inst.u[2] ),
    .B_N(\hopfield_inst.currents[2] ),
    .Y(_105_));
 sg13g2_nand2b_1 _454_ (.Y(_106_),
    .B(\hopfield_inst.neuron_inst.u[2] ),
    .A_N(\hopfield_inst.currents[2] ));
 sg13g2_nand2b_1 _455_ (.Y(_107_),
    .B(_106_),
    .A_N(_105_));
 sg13g2_nor2_1 _456_ (.A(\hopfield_inst.currents[1] ),
    .B(_091_),
    .Y(_108_));
 sg13g2_nand2_1 _457_ (.Y(_109_),
    .A(\hopfield_inst.currents[1] ),
    .B(_091_));
 sg13g2_nor2b_1 _458_ (.A(\hopfield_inst.currents[0] ),
    .B_N(\hopfield_inst.neuron_inst.u[0] ),
    .Y(_110_));
 sg13g2_a21oi_1 _459_ (.A1(_109_),
    .A2(_110_),
    .Y(_111_),
    .B1(_108_));
 sg13g2_a21oi_1 _460_ (.A1(_106_),
    .A2(_111_),
    .Y(_112_),
    .B1(_105_));
 sg13g2_xnor2_1 _461_ (.Y(_113_),
    .A(\hopfield_inst.currents[3] ),
    .B(\hopfield_inst.neuron_inst.u[3] ));
 sg13g2_nand2b_1 _462_ (.Y(_114_),
    .B(_113_),
    .A_N(_112_));
 sg13g2_o21ai_1 _463_ (.B1(_114_),
    .Y(_115_),
    .A1(_093_),
    .A2(\hopfield_inst.neuron_inst.u[3] ));
 sg13g2_xor2_1 _464_ (.B(\hopfield_inst.neuron_inst.u[4] ),
    .A(\hopfield_inst.currents[4] ),
    .X(_116_));
 sg13g2_nor2b_1 _465_ (.A(_116_),
    .B_N(_115_),
    .Y(_117_));
 sg13g2_xnor2_1 _466_ (.Y(_118_),
    .A(\hopfield_inst.currents[5] ),
    .B(\hopfield_inst.neuron_inst.u[5] ));
 sg13g2_o21ai_1 _467_ (.B1(_118_),
    .Y(_119_),
    .A1(_104_),
    .A2(_117_));
 sg13g2_o21ai_1 _468_ (.B1(_119_),
    .Y(_120_),
    .A1(_095_),
    .A2(\hopfield_inst.neuron_inst.u[5] ));
 sg13g2_nand2b_1 _469_ (.Y(_121_),
    .B(\hopfield_inst.neuron_inst.u[6] ),
    .A_N(\hopfield_inst.currents[6] ));
 sg13g2_nand2b_1 _470_ (.Y(_122_),
    .B(_121_),
    .A_N(_103_));
 sg13g2_a21oi_1 _471_ (.A1(_120_),
    .A2(_121_),
    .Y(_123_),
    .B1(_103_));
 sg13g2_xnor2_1 _472_ (.Y(_124_),
    .A(\hopfield_inst.currents[7] ),
    .B(\hopfield_inst.neuron_inst.u[7] ));
 sg13g2_xnor2_1 _473_ (.Y(_125_),
    .A(_123_),
    .B(_124_));
 sg13g2_nand2_1 _474_ (.Y(_126_),
    .A(net125),
    .B(_125_));
 sg13g2_xnor2_1 _475_ (.Y(_127_),
    .A(\hopfield_inst.neuron_inst.v[6] ),
    .B(_125_));
 sg13g2_xnor2_1 _476_ (.Y(_128_),
    .A(net138),
    .B(_125_));
 sg13g2_xnor2_1 _477_ (.Y(_129_),
    .A(_120_),
    .B(_122_));
 sg13g2_nand2_1 _478_ (.Y(_130_),
    .A(net76),
    .B(_129_));
 sg13g2_or3_1 _479_ (.A(_104_),
    .B(_117_),
    .C(_118_),
    .X(_131_));
 sg13g2_and2_1 _480_ (.A(_119_),
    .B(_131_),
    .X(_132_));
 sg13g2_xnor2_1 _481_ (.Y(_133_),
    .A(_115_),
    .B(_116_));
 sg13g2_nand2_1 _482_ (.Y(_134_),
    .A(\hopfield_inst.neuron_inst.v[2] ),
    .B(_133_));
 sg13g2_xnor2_1 _483_ (.Y(_135_),
    .A(_112_),
    .B(_113_));
 sg13g2_nand2_1 _484_ (.Y(_136_),
    .A(net128),
    .B(_135_));
 sg13g2_xnor2_1 _485_ (.Y(_137_),
    .A(_107_),
    .B(_111_));
 sg13g2_nand2_1 _486_ (.Y(_138_),
    .A(net118),
    .B(_137_));
 sg13g2_xnor2_1 _487_ (.Y(_139_),
    .A(net128),
    .B(_135_));
 sg13g2_o21ai_1 _488_ (.B1(_136_),
    .Y(_140_),
    .A1(_138_),
    .A2(_139_));
 sg13g2_xnor2_1 _489_ (.Y(_141_),
    .A(net132),
    .B(_133_));
 sg13g2_nand2b_1 _490_ (.Y(_142_),
    .B(_140_),
    .A_N(_141_));
 sg13g2_and2_1 _491_ (.A(_134_),
    .B(_142_),
    .X(_143_));
 sg13g2_xnor2_1 _492_ (.Y(_144_),
    .A(net77),
    .B(_132_));
 sg13g2_nor2_1 _493_ (.A(_143_),
    .B(_144_),
    .Y(_145_));
 sg13g2_a21oi_1 _494_ (.A1(net77),
    .A2(_132_),
    .Y(_146_),
    .B1(_145_));
 sg13g2_xnor2_1 _495_ (.Y(_147_),
    .A(net76),
    .B(_129_));
 sg13g2_or2_1 _496_ (.X(_148_),
    .B(_147_),
    .A(_146_));
 sg13g2_a21oi_1 _497_ (.A1(_130_),
    .A2(_148_),
    .Y(_149_),
    .B1(_128_));
 sg13g2_a21oi_1 _498_ (.A1(net138),
    .A2(_125_),
    .Y(_150_),
    .B1(_149_));
 sg13g2_o21ai_1 _499_ (.B1(_126_),
    .Y(_151_),
    .A1(_127_),
    .A2(_150_));
 sg13g2_xnor2_1 _500_ (.Y(_152_),
    .A(net105),
    .B(_125_));
 sg13g2_nor2_1 _501_ (.A(\hopfield_inst.neuron_inst.v[2] ),
    .B(\hopfield_inst.neuron_inst.v[3] ),
    .Y(_153_));
 sg13g2_o21ai_1 _502_ (.B1(net76),
    .Y(_154_),
    .A1(\hopfield_inst.neuron_inst.v[2] ),
    .A2(net77));
 sg13g2_nor2_1 _503_ (.A(\hopfield_inst.neuron_inst.v[6] ),
    .B(\hopfield_inst.neuron_inst.v[5] ),
    .Y(_155_));
 sg13g2_a21oi_1 _504_ (.A1(_154_),
    .A2(_155_),
    .Y(_156_),
    .B1(net105));
 sg13g2_inv_2 _505_ (.Y(_157_),
    .A(net74));
 sg13g2_o21ai_1 _506_ (.B1(_157_),
    .Y(_158_),
    .A1(_151_),
    .A2(_152_));
 sg13g2_a21oi_1 _507_ (.A1(_151_),
    .A2(_152_),
    .Y(_050_),
    .B1(_158_));
 sg13g2_xor2_1 _508_ (.B(_150_),
    .A(_127_),
    .X(_159_));
 sg13g2_nor2_1 _509_ (.A(net73),
    .B(_159_),
    .Y(_049_));
 sg13g2_nand2_1 _510_ (.Y(_160_),
    .A(_146_),
    .B(_147_));
 sg13g2_a21oi_1 _511_ (.A1(_148_),
    .A2(_160_),
    .Y(_048_),
    .B1(net73));
 sg13g2_nand2b_1 _512_ (.Y(_161_),
    .B(_141_),
    .A_N(_140_));
 sg13g2_a21oi_1 _513_ (.A1(_142_),
    .A2(_161_),
    .Y(_047_),
    .B1(net73));
 sg13g2_xor2_1 _514_ (.B(_139_),
    .A(_138_),
    .X(_162_));
 sg13g2_nor2_1 _515_ (.A(net74),
    .B(_162_),
    .Y(_046_));
 sg13g2_nand2b_1 _516_ (.Y(_163_),
    .B(net99),
    .A_N(net1));
 sg13g2_nor2b_1 _517_ (.A(net79),
    .B_N(\hopfield_inst.learning_inst.counter[1] ),
    .Y(_164_));
 sg13g2_nand2_1 _518_ (.Y(_165_),
    .A(net78),
    .B(_164_));
 sg13g2_nand4_1 _519_ (.B(net81),
    .C(net68),
    .A(net78),
    .Y(_166_),
    .D(_164_));
 sg13g2_and2_1 _520_ (.A(_163_),
    .B(_166_),
    .X(_045_));
 sg13g2_nand3_1 _521_ (.B(net68),
    .C(_165_),
    .A(net81),
    .Y(_167_));
 sg13g2_nand2b_1 _522_ (.Y(_168_),
    .B(net81),
    .A_N(net99));
 sg13g2_o21ai_1 _523_ (.B1(_168_),
    .Y(_169_),
    .A1(net81),
    .A2(net47));
 sg13g2_nand2_1 _524_ (.Y(_000_),
    .A(_167_),
    .B(_169_));
 sg13g2_o21ai_1 _525_ (.B1(_157_),
    .Y(_170_),
    .A1(net118),
    .A2(_137_));
 sg13g2_nor2b_1 _526_ (.A(_170_),
    .B_N(_138_),
    .Y(_019_));
 sg13g2_a21oi_1 _527_ (.A1(_143_),
    .A2(_144_),
    .Y(_171_),
    .B1(net74));
 sg13g2_nor2b_1 _528_ (.A(_145_),
    .B_N(_171_),
    .Y(_020_));
 sg13g2_and3_1 _529_ (.X(_172_),
    .A(_128_),
    .B(_130_),
    .C(_148_));
 sg13g2_nor3_1 _530_ (.A(_149_),
    .B(net73),
    .C(_172_),
    .Y(_021_));
 sg13g2_nor3_2 _531_ (.A(\hopfield_inst.active_neuron[0] ),
    .B(_096_),
    .C(_097_),
    .Y(_173_));
 sg13g2_nor2b_1 _532_ (.A(_173_),
    .B_N(net45),
    .Y(_008_));
 sg13g2_xnor2_1 _533_ (.Y(_174_),
    .A(net119),
    .B(net75));
 sg13g2_nor2_1 _534_ (.A(net120),
    .B(_174_),
    .Y(_009_));
 sg13g2_a21oi_1 _535_ (.A1(\hopfield_inst.active_neuron[0] ),
    .A2(net75),
    .Y(_175_),
    .B1(net114));
 sg13g2_a21oi_1 _536_ (.A1(net75),
    .A2(net114),
    .Y(_010_),
    .B1(_175_));
 sg13g2_mux4_1 _537_ (.S0(\hopfield_inst.active_neuron[0] ),
    .A0(net2),
    .A1(net3),
    .A2(net4),
    .A3(net5),
    .S1(\hopfield_inst.active_neuron[1] ),
    .X(_176_));
 sg13g2_and2_1 _538_ (.A(net27),
    .B(_176_),
    .X(_011_));
 sg13g2_and2_1 _539_ (.A(net29),
    .B(_176_),
    .X(_012_));
 sg13g2_and2_1 _540_ (.A(net31),
    .B(_176_),
    .X(_013_));
 sg13g2_and2_1 _541_ (.A(net33),
    .B(_176_),
    .X(_014_));
 sg13g2_and2_1 _542_ (.A(_100_),
    .B(_176_),
    .X(_015_));
 sg13g2_and2_1 _543_ (.A(net35),
    .B(_015_),
    .X(_017_));
 sg13g2_nand3_1 _544_ (.B(_101_),
    .C(_176_),
    .A(net37),
    .Y(_177_));
 sg13g2_nand2b_1 _545_ (.Y(_016_),
    .B(_177_),
    .A_N(_017_));
 sg13g2_nor3_1 _546_ (.A(\hopfield_inst.active_neuron[0] ),
    .B(net75),
    .C(\hopfield_inst.active_neuron[2] ),
    .Y(_178_));
 sg13g2_nand2_1 _547_ (.Y(_179_),
    .A(net45),
    .B(_178_));
 sg13g2_a22oi_1 _548_ (.Y(_180_),
    .B1(_179_),
    .B2(net59),
    .A2(_178_),
    .A1(net74));
 sg13g2_inv_1 _549_ (.Y(_001_),
    .A(net106));
 sg13g2_or2_1 _550_ (.X(_181_),
    .B(_174_),
    .A(net45));
 sg13g2_o21ai_1 _551_ (.B1(net139),
    .Y(_182_),
    .A1(\hopfield_inst.active_neuron[0] ),
    .A2(net75));
 sg13g2_nor2_1 _552_ (.A(_157_),
    .B(_178_),
    .Y(_183_));
 sg13g2_nand2_1 _553_ (.Y(_184_),
    .A(_182_),
    .B(_183_));
 sg13g2_o21ai_1 _554_ (.B1(net102),
    .Y(_185_),
    .A1(\hopfield_inst.active_neuron[2] ),
    .A2(_181_));
 sg13g2_o21ai_1 _555_ (.B1(net103),
    .Y(_002_),
    .A1(_181_),
    .A2(_184_));
 sg13g2_nand2b_1 _556_ (.Y(_186_),
    .B(net75),
    .A_N(\hopfield_inst.active_neuron[0] ));
 sg13g2_o21ai_1 _557_ (.B1(net110),
    .Y(_187_),
    .A1(\hopfield_inst.active_neuron[2] ),
    .A2(_186_));
 sg13g2_o21ai_1 _558_ (.B1(net111),
    .Y(_003_),
    .A1(_184_),
    .A2(_186_));
 sg13g2_nor2_1 _559_ (.A(net45),
    .B(_175_),
    .Y(_188_));
 sg13g2_nand2_1 _560_ (.Y(_189_),
    .A(_182_),
    .B(_188_));
 sg13g2_mux2_1 _561_ (.A0(_183_),
    .A1(net113),
    .S(_189_),
    .X(_004_));
 sg13g2_nor3_1 _562_ (.A(\hopfield_inst.active_neuron[0] ),
    .B(net75),
    .C(_097_),
    .Y(_190_));
 sg13g2_mux2_1 _563_ (.A0(net109),
    .A1(net74),
    .S(_190_),
    .X(_005_));
 sg13g2_nor2_1 _564_ (.A(_097_),
    .B(_181_),
    .Y(_191_));
 sg13g2_nor2_1 _565_ (.A(net107),
    .B(_191_),
    .Y(_192_));
 sg13g2_a21oi_1 _566_ (.A1(_157_),
    .A2(_191_),
    .Y(_006_),
    .B1(net108));
 sg13g2_nor2_1 _567_ (.A(net40),
    .B(net120),
    .Y(_193_));
 sg13g2_a21oi_1 _568_ (.A1(_157_),
    .A2(_173_),
    .Y(_007_),
    .B1(_193_));
 sg13g2_and2_1 _569_ (.A(\hopfield_inst.neuron_inst.v[2] ),
    .B(net77),
    .X(_194_));
 sg13g2_o21ai_1 _570_ (.B1(\hopfield_inst.neuron_inst.v[1] ),
    .Y(_195_),
    .A1(\hopfield_inst.neuron_inst.v[0] ),
    .A2(\hopfield_inst.neuron_inst.v[2] ));
 sg13g2_nor3_1 _571_ (.A(_153_),
    .B(_194_),
    .C(_195_),
    .Y(_196_));
 sg13g2_nand3b_1 _572_ (.B(\hopfield_inst.neuron_inst.v[2] ),
    .C(net77),
    .Y(_197_),
    .A_N(net76));
 sg13g2_nand2b_1 _573_ (.Y(_198_),
    .B(net76),
    .A_N(net77));
 sg13g2_xnor2_1 _574_ (.Y(_199_),
    .A(net76),
    .B(net77));
 sg13g2_nand2b_1 _575_ (.Y(_200_),
    .B(_199_),
    .A_N(_194_));
 sg13g2_nor4_2 _576_ (.A(_153_),
    .B(_194_),
    .C(_195_),
    .Y(_201_),
    .D(_199_));
 sg13g2_a21oi_1 _577_ (.A1(_197_),
    .A2(_200_),
    .Y(_202_),
    .B1(_196_));
 sg13g2_or2_1 _578_ (.X(_203_),
    .B(_202_),
    .A(_201_));
 sg13g2_nand3_1 _579_ (.B(_197_),
    .C(_198_),
    .A(_092_),
    .Y(_204_));
 sg13g2_a21o_1 _580_ (.A2(_198_),
    .A1(_197_),
    .B1(_092_),
    .X(_205_));
 sg13g2_and3_1 _581_ (.X(_206_),
    .A(_201_),
    .B(_204_),
    .C(_205_));
 sg13g2_a21oi_1 _582_ (.A1(_204_),
    .A2(_205_),
    .Y(_207_),
    .B1(_201_));
 sg13g2_nor2_2 _583_ (.A(_206_),
    .B(_207_),
    .Y(_208_));
 sg13g2_nand2_1 _584_ (.Y(_209_),
    .A(_028_),
    .B(_208_));
 sg13g2_nand2_1 _585_ (.Y(_210_),
    .A(_203_),
    .B(_209_));
 sg13g2_or2_1 _586_ (.X(_211_),
    .B(_197_),
    .A(_092_));
 sg13g2_and2_1 _587_ (.A(\hopfield_inst.neuron_inst.v[5] ),
    .B(net76),
    .X(_212_));
 sg13g2_a21oi_1 _588_ (.A1(net76),
    .A2(net77),
    .Y(_213_),
    .B1(\hopfield_inst.neuron_inst.v[5] ));
 sg13g2_or3_1 _589_ (.A(\hopfield_inst.neuron_inst.v[6] ),
    .B(_212_),
    .C(_213_),
    .X(_214_));
 sg13g2_o21ai_1 _590_ (.B1(\hopfield_inst.neuron_inst.v[6] ),
    .Y(_215_),
    .A1(_212_),
    .A2(_213_));
 sg13g2_a21oi_1 _591_ (.A1(_214_),
    .A2(_215_),
    .Y(_216_),
    .B1(_211_));
 sg13g2_nand3_1 _592_ (.B(_214_),
    .C(_215_),
    .A(_211_),
    .Y(_217_));
 sg13g2_nand2b_1 _593_ (.Y(_218_),
    .B(_217_),
    .A_N(_216_));
 sg13g2_a21oi_1 _594_ (.A1(_206_),
    .A2(_217_),
    .Y(_219_),
    .B1(_216_));
 sg13g2_mux2_1 _595_ (.A0(_212_),
    .A1(_092_),
    .S(\hopfield_inst.neuron_inst.v[6] ),
    .X(_220_));
 sg13g2_nand4_1 _596_ (.B(_092_),
    .C(\hopfield_inst.neuron_inst.v[4] ),
    .A(\hopfield_inst.neuron_inst.v[6] ),
    .Y(_221_),
    .D(\hopfield_inst.neuron_inst.v[3] ));
 sg13g2_xor2_1 _597_ (.B(\hopfield_inst.neuron_inst.v[7] ),
    .A(\hopfield_inst.neuron_inst.v[0] ),
    .X(_222_));
 sg13g2_xnor2_1 _598_ (.Y(_223_),
    .A(_221_),
    .B(_222_));
 sg13g2_xnor2_1 _599_ (.Y(_224_),
    .A(_220_),
    .B(_223_));
 sg13g2_xnor2_1 _600_ (.Y(_225_),
    .A(_219_),
    .B(_224_));
 sg13g2_inv_1 _601_ (.Y(_226_),
    .A(_225_));
 sg13g2_xor2_1 _602_ (.B(_225_),
    .A(_026_),
    .X(_227_));
 sg13g2_nor2b_1 _603_ (.A(_227_),
    .B_N(_208_),
    .Y(_228_));
 sg13g2_xnor2_1 _604_ (.Y(_229_),
    .A(_208_),
    .B(_227_));
 sg13g2_xor2_1 _605_ (.B(_227_),
    .A(_208_),
    .X(_230_));
 sg13g2_xnor2_1 _606_ (.Y(_231_),
    .A(_206_),
    .B(_218_));
 sg13g2_inv_1 _607_ (.Y(_232_),
    .A(_231_));
 sg13g2_nor2_1 _608_ (.A(_203_),
    .B(_231_),
    .Y(_233_));
 sg13g2_xnor2_1 _609_ (.Y(_234_),
    .A(_229_),
    .B(_233_));
 sg13g2_a21oi_1 _610_ (.A1(_024_),
    .A2(_229_),
    .Y(_235_),
    .B1(_210_));
 sg13g2_xnor2_1 _611_ (.Y(_236_),
    .A(_203_),
    .B(_231_));
 sg13g2_nand2_1 _612_ (.Y(_237_),
    .A(_027_),
    .B(_236_));
 sg13g2_xor2_1 _613_ (.B(_236_),
    .A(_027_),
    .X(_238_));
 sg13g2_o21ai_1 _614_ (.B1(_238_),
    .Y(_239_),
    .A1(_028_),
    .A2(_208_));
 sg13g2_or2_1 _615_ (.X(_240_),
    .B(_239_),
    .A(_235_));
 sg13g2_a21oi_1 _616_ (.A1(_210_),
    .A2(_234_),
    .Y(_241_),
    .B1(_240_));
 sg13g2_inv_1 _617_ (.Y(_242_),
    .A(_241_));
 sg13g2_nor2_1 _618_ (.A(_234_),
    .B(_237_),
    .Y(_243_));
 sg13g2_a21oi_1 _619_ (.A1(_094_),
    .A2(_226_),
    .Y(_244_),
    .B1(_228_));
 sg13g2_nand2_1 _620_ (.Y(_245_),
    .A(_025_),
    .B(_208_));
 sg13g2_xnor2_1 _621_ (.Y(_246_),
    .A(_025_),
    .B(_208_));
 sg13g2_nand2_1 _622_ (.Y(_247_),
    .A(_225_),
    .B(_231_));
 sg13g2_xor2_1 _623_ (.B(_231_),
    .A(_225_),
    .X(_248_));
 sg13g2_nor2_1 _624_ (.A(_246_),
    .B(_248_),
    .Y(_249_));
 sg13g2_xnor2_1 _625_ (.Y(_250_),
    .A(_246_),
    .B(_248_));
 sg13g2_a21oi_1 _626_ (.A1(_230_),
    .A2(_232_),
    .Y(_251_),
    .B1(_203_));
 sg13g2_nand2b_1 _627_ (.Y(_252_),
    .B(_251_),
    .A_N(_250_));
 sg13g2_xnor2_1 _628_ (.Y(_253_),
    .A(_250_),
    .B(_251_));
 sg13g2_nand2b_1 _629_ (.Y(_254_),
    .B(_253_),
    .A_N(_244_));
 sg13g2_xnor2_1 _630_ (.Y(_255_),
    .A(_244_),
    .B(_253_));
 sg13g2_nand2_1 _631_ (.Y(_256_),
    .A(_243_),
    .B(_255_));
 sg13g2_xnor2_1 _632_ (.Y(_257_),
    .A(_243_),
    .B(_255_));
 sg13g2_xnor2_1 _633_ (.Y(_258_),
    .A(_241_),
    .B(_257_));
 sg13g2_nor2_1 _634_ (.A(net73),
    .B(_258_),
    .Y(_259_));
 sg13g2_xor2_1 _635_ (.B(_259_),
    .A(net26),
    .X(_031_));
 sg13g2_o21ai_1 _636_ (.B1(net116),
    .Y(_260_),
    .A1(net73),
    .A2(_258_));
 sg13g2_o21ai_1 _637_ (.B1(_256_),
    .Y(_261_),
    .A1(_242_),
    .A2(_257_));
 sg13g2_xor2_1 _638_ (.B(_247_),
    .A(_029_),
    .X(_262_));
 sg13g2_nand2b_1 _639_ (.Y(_263_),
    .B(_249_),
    .A_N(_262_));
 sg13g2_xor2_1 _640_ (.B(_262_),
    .A(_249_),
    .X(_264_));
 sg13g2_or2_1 _641_ (.X(_265_),
    .B(_264_),
    .A(_245_));
 sg13g2_xnor2_1 _642_ (.Y(_266_),
    .A(_245_),
    .B(_264_));
 sg13g2_a21oi_1 _643_ (.A1(_252_),
    .A2(_254_),
    .Y(_267_),
    .B1(_266_));
 sg13g2_nand3_1 _644_ (.B(_254_),
    .C(_266_),
    .A(_252_),
    .Y(_268_));
 sg13g2_nor2b_1 _645_ (.A(_267_),
    .B_N(_268_),
    .Y(_269_));
 sg13g2_a21oi_1 _646_ (.A1(_261_),
    .A2(_269_),
    .Y(_270_),
    .B1(net73));
 sg13g2_o21ai_1 _647_ (.B1(_270_),
    .Y(_271_),
    .A1(_261_),
    .A2(_269_));
 sg13g2_xnor2_1 _648_ (.Y(_272_),
    .A(_028_),
    .B(_271_));
 sg13g2_xor2_1 _649_ (.B(_272_),
    .A(_260_),
    .X(_032_));
 sg13g2_or2_1 _650_ (.X(_273_),
    .B(_271_),
    .A(_091_));
 sg13g2_o21ai_1 _651_ (.B1(_273_),
    .Y(_274_),
    .A1(_260_),
    .A2(_272_));
 sg13g2_a21o_1 _652_ (.A2(_269_),
    .A1(_261_),
    .B1(_267_),
    .X(_275_));
 sg13g2_o21ai_1 _653_ (.B1(_231_),
    .Y(_276_),
    .A1(_029_),
    .A2(_226_));
 sg13g2_or2_1 _654_ (.X(_277_),
    .B(_276_),
    .A(_102_));
 sg13g2_xnor2_1 _655_ (.Y(_278_),
    .A(_102_),
    .B(_276_));
 sg13g2_and2_1 _656_ (.A(_263_),
    .B(_265_),
    .X(_279_));
 sg13g2_nor2_1 _657_ (.A(_278_),
    .B(_279_),
    .Y(_280_));
 sg13g2_xor2_1 _658_ (.B(_279_),
    .A(_278_),
    .X(_281_));
 sg13g2_xnor2_1 _659_ (.Y(_282_),
    .A(_275_),
    .B(_281_));
 sg13g2_nand2_1 _660_ (.Y(_283_),
    .A(_157_),
    .B(_282_));
 sg13g2_xor2_1 _661_ (.B(_283_),
    .A(net131),
    .X(_284_));
 sg13g2_nand2_1 _662_ (.Y(_285_),
    .A(_274_),
    .B(_284_));
 sg13g2_xor2_1 _663_ (.B(_284_),
    .A(_274_),
    .X(_033_));
 sg13g2_nand2b_1 _664_ (.Y(_286_),
    .B(_283_),
    .A_N(net136));
 sg13g2_a21oi_1 _665_ (.A1(_275_),
    .A2(_281_),
    .Y(_287_),
    .B1(_280_));
 sg13g2_xnor2_1 _666_ (.Y(_288_),
    .A(\hopfield_inst.neuron_inst.u[7] ),
    .B(_225_));
 sg13g2_xnor2_1 _667_ (.Y(_289_),
    .A(_277_),
    .B(_288_));
 sg13g2_a21oi_1 _668_ (.A1(_287_),
    .A2(_289_),
    .Y(_290_),
    .B1(net73));
 sg13g2_o21ai_1 _669_ (.B1(_290_),
    .Y(_291_),
    .A1(_287_),
    .A2(_289_));
 sg13g2_inv_1 _670_ (.Y(_292_),
    .A(_291_));
 sg13g2_xnor2_1 _671_ (.Y(_293_),
    .A(_026_),
    .B(_291_));
 sg13g2_nand3_1 _672_ (.B(_286_),
    .C(_293_),
    .A(_285_),
    .Y(_294_));
 sg13g2_a21o_1 _673_ (.A2(_286_),
    .A1(_285_),
    .B1(_293_),
    .X(_295_));
 sg13g2_and2_1 _674_ (.A(net137),
    .B(_295_),
    .X(_034_));
 sg13g2_nand2_1 _675_ (.Y(_296_),
    .A(net133),
    .B(_292_));
 sg13g2_xnor2_1 _676_ (.Y(_297_),
    .A(_025_),
    .B(_291_));
 sg13g2_a21oi_1 _677_ (.A1(_295_),
    .A2(_296_),
    .Y(_298_),
    .B1(_297_));
 sg13g2_nand3_1 _678_ (.B(_296_),
    .C(_297_),
    .A(_295_),
    .Y(_299_));
 sg13g2_nor2b_1 _679_ (.A(_298_),
    .B_N(net134),
    .Y(_035_));
 sg13g2_a21oi_1 _680_ (.A1(net126),
    .A2(_292_),
    .Y(_300_),
    .B1(_298_));
 sg13g2_xor2_1 _681_ (.B(_291_),
    .A(_029_),
    .X(_301_));
 sg13g2_xnor2_1 _682_ (.Y(_036_),
    .A(_300_),
    .B(_301_));
 sg13g2_a21oi_1 _683_ (.A1(\hopfield_inst.neuron_inst.u[4] ),
    .A2(_029_),
    .Y(_302_),
    .B1(\hopfield_inst.neuron_inst.u[5] ));
 sg13g2_nor2_1 _684_ (.A(_291_),
    .B(_302_),
    .Y(_303_));
 sg13g2_a21o_1 _685_ (.A2(_301_),
    .A1(_298_),
    .B1(_303_),
    .X(_304_));
 sg13g2_xnor2_1 _686_ (.Y(_305_),
    .A(_102_),
    .B(_291_));
 sg13g2_xor2_1 _687_ (.B(_305_),
    .A(_304_),
    .X(_037_));
 sg13g2_a22oi_1 _688_ (.Y(_306_),
    .B1(_304_),
    .B2(_305_),
    .A2(_292_),
    .A1(net123));
 sg13g2_xnor2_1 _689_ (.Y(_307_),
    .A(\hopfield_inst.neuron_inst.u[7] ),
    .B(_291_));
 sg13g2_xnor2_1 _690_ (.Y(_038_),
    .A(_306_),
    .B(_307_));
 sg13g2_nand3_1 _691_ (.B(net25),
    .C(net86),
    .A(net40),
    .Y(_308_));
 sg13g2_a21o_1 _692_ (.A2(net86),
    .A1(net40),
    .B1(net25),
    .X(_309_));
 sg13g2_and2_1 _693_ (.A(_308_),
    .B(_309_),
    .X(_051_));
 sg13g2_nand4_1 _694_ (.B(net25),
    .C(net24),
    .A(net40),
    .Y(_310_),
    .D(net86));
 sg13g2_xnor2_1 _695_ (.Y(_052_),
    .A(net24),
    .B(_308_));
 sg13g2_xnor2_1 _696_ (.Y(_053_),
    .A(net23),
    .B(_310_));
 sg13g2_a21oi_1 _697_ (.A1(net79),
    .A2(_089_),
    .Y(_311_),
    .B1(net78));
 sg13g2_o21ai_1 _698_ (.B1(_311_),
    .Y(_312_),
    .A1(net79),
    .A2(uio_out[6]));
 sg13g2_nand2_1 _699_ (.Y(_313_),
    .A(net81),
    .B(net47));
 sg13g2_nor3_2 _700_ (.A(net79),
    .B(\hopfield_inst.learning_inst.counter[1] ),
    .C(net78),
    .Y(_314_));
 sg13g2_nand2b_1 _701_ (.Y(_315_),
    .B(_314_),
    .A_N(uio_out[4]));
 sg13g2_nor2b_1 _702_ (.A(\hopfield_inst.learning_inst.counter[1] ),
    .B_N(net79),
    .Y(_316_));
 sg13g2_and2_2 _703_ (.A(_088_),
    .B(_316_),
    .X(_317_));
 sg13g2_nor2b_1 _704_ (.A(uio_out[5]),
    .B_N(_317_),
    .Y(_318_));
 sg13g2_nor2b_1 _705_ (.A(net80),
    .B_N(uo_out[0]),
    .Y(_319_));
 sg13g2_a21oi_1 _706_ (.A1(net80),
    .A2(uo_out[1]),
    .Y(_320_),
    .B1(_319_));
 sg13g2_a221oi_1 _707_ (.B2(\hopfield_inst.learning_inst.counter[2] ),
    .C1(_318_),
    .B1(_320_),
    .A1(\hopfield_inst.learning_inst.counter[1] ),
    .Y(_321_),
    .A2(_312_));
 sg13g2_nand4_1 _708_ (.B(net47),
    .C(_315_),
    .A(net81),
    .Y(_322_),
    .D(net49));
 sg13g2_and2_2 _709_ (.A(net78),
    .B(_316_),
    .X(_323_));
 sg13g2_and2_2 _710_ (.A(_088_),
    .B(_164_),
    .X(_324_));
 sg13g2_nor3_2 _711_ (.A(net79),
    .B(\hopfield_inst.learning_inst.counter[1] ),
    .C(_088_),
    .Y(_325_));
 sg13g2_nand2_1 _712_ (.Y(_326_),
    .A(net79),
    .B(\hopfield_inst.learning_inst.counter[1] ));
 sg13g2_nor2_2 _713_ (.A(net78),
    .B(_326_),
    .Y(_327_));
 sg13g2_a22oi_1 _714_ (.Y(_328_),
    .B1(_327_),
    .B2(\hopfield_inst.learning_inst.weights[25][3] ),
    .A2(_325_),
    .A1(\hopfield_inst.learning_inst.weights[33][3] ));
 sg13g2_a22oi_1 _715_ (.Y(_329_),
    .B1(_323_),
    .B2(\hopfield_inst.learning_inst.weights[41][3] ),
    .A2(_314_),
    .A1(\hopfield_inst.learning_inst.weights[1][3] ));
 sg13g2_a22oi_1 _716_ (.Y(_330_),
    .B1(_324_),
    .B2(\hopfield_inst.learning_inst.weights[17][3] ),
    .A2(_317_),
    .A1(\hopfield_inst.learning_inst.weights[9][3] ));
 sg13g2_nand3_1 _717_ (.B(_329_),
    .C(_330_),
    .A(_328_),
    .Y(_331_));
 sg13g2_a22oi_1 _718_ (.Y(_332_),
    .B1(_327_),
    .B2(\hopfield_inst.learning_inst.weights[25][2] ),
    .A2(_323_),
    .A1(\hopfield_inst.learning_inst.weights[41][2] ));
 sg13g2_a22oi_1 _719_ (.Y(_333_),
    .B1(_317_),
    .B2(\hopfield_inst.learning_inst.weights[9][2] ),
    .A2(_314_),
    .A1(\hopfield_inst.learning_inst.weights[1][2] ));
 sg13g2_nand2_1 _720_ (.Y(_334_),
    .A(_332_),
    .B(_333_));
 sg13g2_a221oi_1 _721_ (.B2(\hopfield_inst.learning_inst.weights[33][2] ),
    .C1(_334_),
    .B1(_325_),
    .A1(\hopfield_inst.learning_inst.weights[17][2] ),
    .Y(_335_),
    .A2(_324_));
 sg13g2_a22oi_1 _722_ (.Y(_336_),
    .B1(_324_),
    .B2(\hopfield_inst.learning_inst.weights[17][0] ),
    .A2(_323_),
    .A1(\hopfield_inst.learning_inst.weights[41][0] ));
 sg13g2_a22oi_1 _723_ (.Y(_337_),
    .B1(_325_),
    .B2(\hopfield_inst.learning_inst.weights[33][0] ),
    .A2(_314_),
    .A1(\hopfield_inst.learning_inst.weights[1][0] ));
 sg13g2_nand2_1 _724_ (.Y(_338_),
    .A(_336_),
    .B(_337_));
 sg13g2_a221oi_1 _725_ (.B2(\hopfield_inst.learning_inst.weights[25][0] ),
    .C1(_338_),
    .B1(_327_),
    .A1(net50),
    .Y(_339_),
    .A2(_317_));
 sg13g2_a22oi_1 _726_ (.Y(_340_),
    .B1(_323_),
    .B2(\hopfield_inst.learning_inst.weights[41][1] ),
    .A2(_314_),
    .A1(\hopfield_inst.learning_inst.weights[1][1] ));
 sg13g2_a22oi_1 _727_ (.Y(_341_),
    .B1(_325_),
    .B2(\hopfield_inst.learning_inst.weights[33][1] ),
    .A2(_317_),
    .A1(\hopfield_inst.learning_inst.weights[9][1] ));
 sg13g2_a22oi_1 _728_ (.Y(_342_),
    .B1(_327_),
    .B2(\hopfield_inst.learning_inst.weights[25][1] ),
    .A2(_324_),
    .A1(\hopfield_inst.learning_inst.weights[17][1] ));
 sg13g2_nand3_1 _729_ (.B(_341_),
    .C(_342_),
    .A(_340_),
    .Y(_343_));
 sg13g2_nand2b_1 _730_ (.Y(_344_),
    .B(_343_),
    .A_N(net72));
 sg13g2_or2_1 _731_ (.X(_345_),
    .B(_344_),
    .A(_335_));
 sg13g2_nor2_1 _732_ (.A(_331_),
    .B(_345_),
    .Y(_346_));
 sg13g2_nor2_1 _733_ (.A(_322_),
    .B(_346_),
    .Y(_347_));
 sg13g2_mux2_1 _734_ (.A0(net27),
    .A1(net72),
    .S(net71),
    .X(_054_));
 sg13g2_xnor2_1 _735_ (.Y(_348_),
    .A(net72),
    .B(_343_));
 sg13g2_mux2_1 _736_ (.A0(net29),
    .A1(_348_),
    .S(net71),
    .X(_055_));
 sg13g2_xor2_1 _737_ (.B(_344_),
    .A(_335_),
    .X(_349_));
 sg13g2_nand2b_1 _738_ (.Y(_350_),
    .B(_349_),
    .A_N(_322_));
 sg13g2_o21ai_1 _739_ (.B1(_350_),
    .Y(_056_),
    .A1(_098_),
    .A2(net71));
 sg13g2_nand3b_1 _740_ (.B(_331_),
    .C(_345_),
    .Y(_351_),
    .A_N(_322_));
 sg13g2_inv_2 _741_ (.Y(_352_),
    .A(_351_));
 sg13g2_o21ai_1 _742_ (.B1(_351_),
    .Y(_057_),
    .A1(_099_),
    .A2(net70));
 sg13g2_o21ai_1 _743_ (.B1(_351_),
    .Y(_058_),
    .A1(_100_),
    .A2(net70));
 sg13g2_o21ai_1 _744_ (.B1(_351_),
    .Y(_059_),
    .A1(_101_),
    .A2(net70));
 sg13g2_nand3_1 _745_ (.B(_090_),
    .C(net99),
    .A(net81),
    .Y(_353_));
 sg13g2_and2_1 _746_ (.A(_167_),
    .B(_353_),
    .X(_354_));
 sg13g2_nand2_1 _747_ (.Y(_355_),
    .A(net79),
    .B(_354_));
 sg13g2_o21ai_1 _748_ (.B1(_355_),
    .Y(_060_),
    .A1(net80),
    .A2(_167_));
 sg13g2_nand2_1 _749_ (.Y(_356_),
    .A(net61),
    .B(_354_));
 sg13g2_nor2_1 _750_ (.A(_164_),
    .B(_316_),
    .Y(_357_));
 sg13g2_o21ai_1 _751_ (.B1(_356_),
    .Y(_061_),
    .A1(_167_),
    .A2(_357_));
 sg13g2_nand2_1 _752_ (.Y(_358_),
    .A(net78),
    .B(_354_));
 sg13g2_xnor2_1 _753_ (.Y(_359_),
    .A(net54),
    .B(_326_));
 sg13g2_o21ai_1 _754_ (.B1(_358_),
    .Y(_062_),
    .A1(_167_),
    .A2(_359_));
 sg13g2_nand2_2 _755_ (.Y(_360_),
    .A(_314_),
    .B(net71));
 sg13g2_mux2_1 _756_ (.A0(net51),
    .A1(net64),
    .S(_360_),
    .X(_063_));
 sg13g2_mux2_1 _757_ (.A0(_348_),
    .A1(net53),
    .S(_360_),
    .X(_064_));
 sg13g2_mux2_1 _758_ (.A0(_349_),
    .A1(net56),
    .S(_360_),
    .X(_065_));
 sg13g2_xnor2_1 _759_ (.Y(_361_),
    .A(_331_),
    .B(_345_));
 sg13g2_mux2_1 _760_ (.A0(_361_),
    .A1(net58),
    .S(_360_),
    .X(_066_));
 sg13g2_nand2_2 _761_ (.Y(_362_),
    .A(_317_),
    .B(net70));
 sg13g2_mux2_1 _762_ (.A0(net72),
    .A1(net50),
    .S(_362_),
    .X(_067_));
 sg13g2_mux2_1 _763_ (.A0(_348_),
    .A1(net57),
    .S(_362_),
    .X(_068_));
 sg13g2_mux2_1 _764_ (.A0(_349_),
    .A1(net60),
    .S(_362_),
    .X(_069_));
 sg13g2_a22oi_1 _765_ (.Y(_363_),
    .B1(_362_),
    .B2(net44),
    .A2(_352_),
    .A1(_317_));
 sg13g2_inv_1 _766_ (.Y(_070_),
    .A(_363_));
 sg13g2_nand2_2 _767_ (.Y(_364_),
    .A(_323_),
    .B(net70));
 sg13g2_mux2_1 _768_ (.A0(net72),
    .A1(net98),
    .S(_364_),
    .X(_071_));
 sg13g2_mux2_1 _769_ (.A0(_348_),
    .A1(net52),
    .S(_364_),
    .X(_072_));
 sg13g2_mux2_1 _770_ (.A0(_349_),
    .A1(net100),
    .S(_364_),
    .X(_073_));
 sg13g2_a22oi_1 _771_ (.Y(_365_),
    .B1(_364_),
    .B2(net43),
    .A2(_352_),
    .A1(_323_));
 sg13g2_inv_1 _772_ (.Y(_074_),
    .A(_365_));
 sg13g2_nand2_2 _773_ (.Y(_366_),
    .A(_324_),
    .B(net70));
 sg13g2_mux2_1 _774_ (.A0(net72),
    .A1(net62),
    .S(_366_),
    .X(_075_));
 sg13g2_mux2_1 _775_ (.A0(_348_),
    .A1(net63),
    .S(_366_),
    .X(_076_));
 sg13g2_mux2_1 _776_ (.A0(_349_),
    .A1(net96),
    .S(_366_),
    .X(_077_));
 sg13g2_a22oi_1 _777_ (.Y(_367_),
    .B1(_366_),
    .B2(net42),
    .A2(_352_),
    .A1(_324_));
 sg13g2_inv_1 _778_ (.Y(_078_),
    .A(_367_));
 sg13g2_nand2_2 _779_ (.Y(_368_),
    .A(_327_),
    .B(net70));
 sg13g2_mux2_1 _780_ (.A0(net72),
    .A1(net101),
    .S(_368_),
    .X(_079_));
 sg13g2_mux2_1 _781_ (.A0(_348_),
    .A1(net69),
    .S(_368_),
    .X(_080_));
 sg13g2_mux2_1 _782_ (.A0(_349_),
    .A1(net66),
    .S(_368_),
    .X(_081_));
 sg13g2_a22oi_1 _783_ (.Y(_369_),
    .B1(_368_),
    .B2(net38),
    .A2(_352_),
    .A1(_327_));
 sg13g2_inv_1 _784_ (.Y(_082_),
    .A(_369_));
 sg13g2_nand2_2 _785_ (.Y(_370_),
    .A(_325_),
    .B(net70));
 sg13g2_mux2_1 _786_ (.A0(net72),
    .A1(net67),
    .S(_370_),
    .X(_083_));
 sg13g2_mux2_1 _787_ (.A0(_348_),
    .A1(net97),
    .S(_370_),
    .X(_084_));
 sg13g2_mux2_1 _788_ (.A0(_349_),
    .A1(net65),
    .S(_370_),
    .X(_085_));
 sg13g2_a22oi_1 _789_ (.Y(_371_),
    .B1(_370_),
    .B2(net39),
    .A2(_352_),
    .A1(_325_));
 sg13g2_inv_1 _790_ (.Y(_086_),
    .A(_371_));
 sg13g2_o21ai_1 _791_ (.B1(_313_),
    .Y(_087_),
    .A1(net81),
    .A2(_090_));
 sg13g2_and2_1 _792_ (.A(net35),
    .B(_015_),
    .X(_018_));
 sg13g2_dfrbp_1 _793_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net86),
    .D(net25),
    .Q_N(_414_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _794_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net86),
    .D(net24),
    .Q_N(_415_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _795_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net87),
    .D(net23),
    .Q_N(_413_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _796_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net88),
    .D(_045_),
    .Q_N(\hopfield_inst.learning_inst.state[0] ),
    .Q(_039_));
 sg13g2_dfrbp_1 _797_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net88),
    .D(_000_),
    .Q_N(_412_),
    .Q(\hopfield_inst.learning_inst.state[2] ));
 sg13g2_dfrbp_1 _798_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net18),
    .D(_051_),
    .Q_N(_411_),
    .Q(\temp_activity_count[0] ));
 sg13g2_dfrbp_1 _799_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net17),
    .D(_052_),
    .Q_N(_410_),
    .Q(\temp_activity_count[1] ));
 sg13g2_dfrbp_1 _800_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net16),
    .D(_053_),
    .Q_N(_409_),
    .Q(\temp_activity_count[2] ));
 sg13g2_dfrbp_1 _801_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net84),
    .D(_054_),
    .Q_N(_408_),
    .Q(\hopfield_inst.learning_inst.temp_weight[0] ));
 sg13g2_dfrbp_1 _802_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net90),
    .D(_055_),
    .Q_N(_407_),
    .Q(\hopfield_inst.learning_inst.temp_weight[1] ));
 sg13g2_dfrbp_1 _803_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net84),
    .D(_056_),
    .Q_N(_406_),
    .Q(\hopfield_inst.learning_inst.temp_weight[2] ));
 sg13g2_dfrbp_1 _804_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_057_),
    .Q_N(_405_),
    .Q(\hopfield_inst.learning_inst.temp_weight[3] ));
 sg13g2_dfrbp_1 _805_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_058_),
    .Q_N(_404_),
    .Q(\hopfield_inst.learning_inst.temp_weight[4] ));
 sg13g2_dfrbp_1 _806_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_059_),
    .Q_N(_403_),
    .Q(\hopfield_inst.learning_inst.temp_weight[5] ));
 sg13g2_dfrbp_1 _807_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net88),
    .D(_060_),
    .Q_N(_402_),
    .Q(\hopfield_inst.learning_inst.counter[0] ));
 sg13g2_dfrbp_1 _808_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net87),
    .D(_061_),
    .Q_N(_401_),
    .Q(\hopfield_inst.learning_inst.counter[1] ));
 sg13g2_dfrbp_1 _809_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net87),
    .D(net55),
    .Q_N(_022_),
    .Q(\hopfield_inst.learning_inst.counter[2] ));
 sg13g2_dfrbp_1 _810_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net84),
    .D(_063_),
    .Q_N(_400_),
    .Q(\hopfield_inst.learning_inst.weights[1][0] ));
 sg13g2_dfrbp_1 _811_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net85),
    .D(_064_),
    .Q_N(_399_),
    .Q(\hopfield_inst.learning_inst.weights[1][1] ));
 sg13g2_dfrbp_1 _812_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net84),
    .D(_065_),
    .Q_N(_398_),
    .Q(\hopfield_inst.learning_inst.weights[1][2] ));
 sg13g2_dfrbp_1 _813_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net85),
    .D(_066_),
    .Q_N(_397_),
    .Q(\hopfield_inst.learning_inst.weights[1][3] ));
 sg13g2_dfrbp_1 _814_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net83),
    .D(_067_),
    .Q_N(_396_),
    .Q(\hopfield_inst.learning_inst.weights[9][0] ));
 sg13g2_dfrbp_1 _815_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net83),
    .D(_068_),
    .Q_N(_395_),
    .Q(\hopfield_inst.learning_inst.weights[9][1] ));
 sg13g2_dfrbp_1 _816_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net83),
    .D(_069_),
    .Q_N(_394_),
    .Q(\hopfield_inst.learning_inst.weights[9][2] ));
 sg13g2_dfrbp_1 _817_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net83),
    .D(_070_),
    .Q_N(_393_),
    .Q(\hopfield_inst.learning_inst.weights[9][3] ));
 sg13g2_dfrbp_1 _818_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net84),
    .D(_071_),
    .Q_N(_392_),
    .Q(\hopfield_inst.learning_inst.weights[41][0] ));
 sg13g2_dfrbp_1 _819_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net84),
    .D(_072_),
    .Q_N(_391_),
    .Q(\hopfield_inst.learning_inst.weights[41][1] ));
 sg13g2_dfrbp_1 _820_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net84),
    .D(_073_),
    .Q_N(_390_),
    .Q(\hopfield_inst.learning_inst.weights[41][2] ));
 sg13g2_dfrbp_1 _821_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net84),
    .D(_074_),
    .Q_N(_389_),
    .Q(\hopfield_inst.learning_inst.weights[41][3] ));
 sg13g2_dfrbp_1 _822_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(_075_),
    .Q_N(_388_),
    .Q(\hopfield_inst.learning_inst.weights[17][0] ));
 sg13g2_dfrbp_1 _823_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(_076_),
    .Q_N(_387_),
    .Q(\hopfield_inst.learning_inst.weights[17][1] ));
 sg13g2_dfrbp_1 _824_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(_077_),
    .Q_N(_386_),
    .Q(\hopfield_inst.learning_inst.weights[17][2] ));
 sg13g2_dfrbp_1 _825_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net82),
    .D(_078_),
    .Q_N(_385_),
    .Q(\hopfield_inst.learning_inst.weights[17][3] ));
 sg13g2_dfrbp_1 _826_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net82),
    .D(_079_),
    .Q_N(_384_),
    .Q(\hopfield_inst.learning_inst.weights[25][0] ));
 sg13g2_dfrbp_1 _827_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net82),
    .D(_080_),
    .Q_N(_383_),
    .Q(\hopfield_inst.learning_inst.weights[25][1] ));
 sg13g2_dfrbp_1 _828_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net82),
    .D(_081_),
    .Q_N(_382_),
    .Q(\hopfield_inst.learning_inst.weights[25][2] ));
 sg13g2_dfrbp_1 _829_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net82),
    .D(_082_),
    .Q_N(_381_),
    .Q(\hopfield_inst.learning_inst.weights[25][3] ));
 sg13g2_dfrbp_1 _830_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net83),
    .D(_083_),
    .Q_N(_380_),
    .Q(\hopfield_inst.learning_inst.weights[33][0] ));
 sg13g2_dfrbp_1 _831_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net87),
    .D(_084_),
    .Q_N(_379_),
    .Q(\hopfield_inst.learning_inst.weights[33][1] ));
 sg13g2_dfrbp_1 _832_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net83),
    .D(_085_),
    .Q_N(_378_),
    .Q(\hopfield_inst.learning_inst.weights[33][2] ));
 sg13g2_dfrbp_1 _833_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net83),
    .D(_086_),
    .Q_N(_377_),
    .Q(\hopfield_inst.learning_inst.weights[33][3] ));
 sg13g2_dfrbp_1 _834_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net90),
    .D(_031_),
    .Q_N(_024_),
    .Q(\hopfield_inst.neuron_inst.u[0] ));
 sg13g2_dfrbp_1 _835_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net90),
    .D(net117),
    .Q_N(_028_),
    .Q(\hopfield_inst.neuron_inst.u[1] ));
 sg13g2_dfrbp_1 _836_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net90),
    .D(_033_),
    .Q_N(_027_),
    .Q(\hopfield_inst.neuron_inst.u[2] ));
 sg13g2_dfrbp_1 _837_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(_034_),
    .Q_N(_026_),
    .Q(\hopfield_inst.neuron_inst.u[3] ));
 sg13g2_dfrbp_1 _838_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(net135),
    .Q_N(_025_),
    .Q(\hopfield_inst.neuron_inst.u[4] ));
 sg13g2_dfrbp_1 _839_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(net127),
    .Q_N(_029_),
    .Q(\hopfield_inst.neuron_inst.u[5] ));
 sg13g2_dfrbp_1 _840_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(net130),
    .Q_N(_030_),
    .Q(\hopfield_inst.neuron_inst.u[6] ));
 sg13g2_dfrbp_1 _841_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net90),
    .D(net124),
    .Q_N(_416_),
    .Q(\hopfield_inst.neuron_inst.u[7] ));
 sg13g2_dfrbp_1 _842_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net92),
    .D(_019_),
    .Q_N(_376_),
    .Q(\hopfield_inst.neuron_inst.v[0] ));
 sg13g2_dfrbp_1 _843_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net92),
    .D(_046_),
    .Q_N(\hopfield_inst.neuron_inst.v[1] ),
    .Q(_040_));
 sg13g2_dfrbp_1 _844_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net92),
    .D(_047_),
    .Q_N(\hopfield_inst.neuron_inst.v[2] ),
    .Q(_041_));
 sg13g2_dfrbp_1 _845_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net93),
    .D(_020_),
    .Q_N(_375_),
    .Q(\hopfield_inst.neuron_inst.v[3] ));
 sg13g2_dfrbp_1 _846_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net92),
    .D(_048_),
    .Q_N(\hopfield_inst.neuron_inst.v[4] ),
    .Q(_042_));
 sg13g2_dfrbp_1 _847_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net93),
    .D(_021_),
    .Q_N(_374_),
    .Q(\hopfield_inst.neuron_inst.v[5] ));
 sg13g2_dfrbp_1 _848_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net93),
    .D(_049_),
    .Q_N(\hopfield_inst.neuron_inst.v[6] ),
    .Q(_043_));
 sg13g2_dfrbp_1 _849_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net93),
    .D(_050_),
    .Q_N(\hopfield_inst.neuron_inst.v[7] ),
    .Q(_044_));
 sg13g2_dfrbp_1 _850_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net92),
    .D(net46),
    .Q_N(_023_),
    .Q(\hopfield_inst.active_neuron[0] ));
 sg13g2_dfrbp_1 _851_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net92),
    .D(_009_),
    .Q_N(_417_),
    .Q(\hopfield_inst.active_neuron[1] ));
 sg13g2_dfrbp_1 _852_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net88),
    .D(net115),
    .Q_N(_418_),
    .Q(\hopfield_inst.active_neuron[2] ));
 sg13g2_dfrbp_1 _853_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net90),
    .D(net28),
    .Q_N(_419_),
    .Q(\hopfield_inst.currents[0] ));
 sg13g2_dfrbp_1 _854_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net90),
    .D(net30),
    .Q_N(_420_),
    .Q(\hopfield_inst.currents[1] ));
 sg13g2_dfrbp_1 _855_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net92),
    .D(net32),
    .Q_N(_421_),
    .Q(\hopfield_inst.currents[2] ));
 sg13g2_dfrbp_1 _856_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net89),
    .D(net34),
    .Q_N(_422_),
    .Q(\hopfield_inst.currents[3] ));
 sg13g2_dfrbp_1 _857_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(_015_),
    .Q_N(_423_),
    .Q(\hopfield_inst.currents[4] ));
 sg13g2_dfrbp_1 _858_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(_016_),
    .Q_N(_424_),
    .Q(\hopfield_inst.currents[5] ));
 sg13g2_dfrbp_1 _859_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(_017_),
    .Q_N(_425_),
    .Q(\hopfield_inst.currents[6] ));
 sg13g2_dfrbp_1 _860_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(net36),
    .Q_N(_426_),
    .Q(\hopfield_inst.currents[7] ));
 sg13g2_dfrbp_1 _861_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net86),
    .D(_001_),
    .Q_N(_427_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _862_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net86),
    .D(net104),
    .Q_N(_428_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _863_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net95),
    .D(net112),
    .Q_N(_429_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _864_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net86),
    .D(_004_),
    .Q_N(_430_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _865_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net92),
    .D(_005_),
    .Q_N(_431_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _866_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net88),
    .D(_006_),
    .Q_N(_432_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _867_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net88),
    .D(net121),
    .Q_N(_373_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _868_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net88),
    .D(_087_),
    .Q_N(_372_),
    .Q(\hopfield_inst.learning_inst.state[1] ));
 sg13g2_tiehi _799__17 (.L_HI(net17));
 sg13g2_tiehi _798__18 (.L_HI(net18));
 sg13g2_tiehi tt_um_cellular_alchemist_19 (.L_HI(net19));
 sg13g2_tiehi tt_um_cellular_alchemist_20 (.L_HI(net20));
 sg13g2_tiehi tt_um_cellular_alchemist_21 (.L_HI(net21));
 sg13g2_tiehi tt_um_cellular_alchemist_22 (.L_HI(net22));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_cellular_alchemist_7 (.L_LO(net7));
 sg13g2_tielo tt_um_cellular_alchemist_8 (.L_LO(net8));
 sg13g2_tielo tt_um_cellular_alchemist_9 (.L_LO(net9));
 sg13g2_tielo tt_um_cellular_alchemist_10 (.L_LO(net10));
 sg13g2_tielo tt_um_cellular_alchemist_11 (.L_LO(net11));
 sg13g2_tielo tt_um_cellular_alchemist_12 (.L_LO(net12));
 sg13g2_tielo tt_um_cellular_alchemist_13 (.L_LO(net13));
 sg13g2_tielo tt_um_cellular_alchemist_14 (.L_LO(net14));
 sg13g2_tielo tt_um_cellular_alchemist_15 (.L_LO(net15));
 sg13g2_tiehi _800__16 (.L_HI(net16));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(_347_));
 sg13g2_buf_2 fanout71 (.A(_347_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(net51));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_156_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(net41),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(\hopfield_inst.neuron_inst.v[4] ),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(\hopfield_inst.neuron_inst.v[3] ),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(net48),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_1 fanout80 (.A(net122),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(net1),
    .X(net81));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(net85));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(net85));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net85));
 sg13g2_buf_2 fanout85 (.A(net95),
    .X(net85));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(net87));
 sg13g2_buf_2 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(net95));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(net90));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(net94));
 sg13g2_buf_2 fanout91 (.A(net94),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(net94));
 sg13g2_buf_2 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(rst_n),
    .X(net95));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[3]),
    .X(net5));
 sg13g2_tielo tt_um_cellular_alchemist_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\temp_activity_count[2] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold2 (.A(\temp_activity_count[1] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold3 (.A(\temp_activity_count[0] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold4 (.A(_024_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold5 (.A(\hopfield_inst.learning_inst.temp_weight[0] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold6 (.A(_011_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold7 (.A(\hopfield_inst.learning_inst.temp_weight[1] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold8 (.A(_012_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold9 (.A(\hopfield_inst.learning_inst.temp_weight[2] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold10 (.A(_013_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold11 (.A(\hopfield_inst.learning_inst.temp_weight[3] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold12 (.A(_014_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hopfield_inst.learning_inst.temp_weight[5] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold14 (.A(_018_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hopfield_inst.learning_inst.temp_weight[4] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold16 (.A(\hopfield_inst.learning_inst.weights[25][3] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold17 (.A(\hopfield_inst.learning_inst.weights[33][3] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold18 (.A(uo_out[2]),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hopfield_inst.active_neuron[1] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold20 (.A(\hopfield_inst.learning_inst.weights[17][3] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold21 (.A(\hopfield_inst.learning_inst.weights[41][3] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hopfield_inst.learning_inst.weights[9][3] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold23 (.A(_023_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold24 (.A(_008_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold25 (.A(\hopfield_inst.learning_inst.state[2] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hopfield_inst.learning_inst.counter[2] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold27 (.A(_321_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold28 (.A(\hopfield_inst.learning_inst.weights[9][0] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold29 (.A(_339_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hopfield_inst.learning_inst.weights[41][1] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold31 (.A(\hopfield_inst.learning_inst.weights[1][1] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold32 (.A(_022_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold33 (.A(_062_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hopfield_inst.learning_inst.weights[1][2] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold35 (.A(\hopfield_inst.learning_inst.weights[9][1] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold36 (.A(\hopfield_inst.learning_inst.weights[1][3] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold37 (.A(uio_out[4]),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hopfield_inst.learning_inst.weights[9][2] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold39 (.A(\hopfield_inst.learning_inst.counter[1] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold40 (.A(\hopfield_inst.learning_inst.weights[17][0] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold41 (.A(\hopfield_inst.learning_inst.weights[17][1] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold42 (.A(\hopfield_inst.learning_inst.weights[1][0] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold43 (.A(\hopfield_inst.learning_inst.weights[33][2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold44 (.A(\hopfield_inst.learning_inst.weights[25][2] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold45 (.A(\hopfield_inst.learning_inst.weights[33][0] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold46 (.A(\hopfield_inst.learning_inst.state[1] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold47 (.A(\hopfield_inst.learning_inst.weights[25][1] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold48 (.A(\hopfield_inst.learning_inst.weights[17][2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold49 (.A(\hopfield_inst.learning_inst.weights[33][1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold50 (.A(\hopfield_inst.learning_inst.weights[41][0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold51 (.A(\hopfield_inst.learning_inst.state[0] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold52 (.A(\hopfield_inst.learning_inst.weights[41][2] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold53 (.A(\hopfield_inst.learning_inst.weights[25][0] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold54 (.A(uio_out[5]),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold55 (.A(_185_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold56 (.A(_002_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold57 (.A(\hopfield_inst.neuron_inst.v[7] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold58 (.A(_180_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold59 (.A(uo_out[1]),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold60 (.A(_192_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold61 (.A(uo_out[0]),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold62 (.A(uio_out[6]),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold63 (.A(_187_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold64 (.A(_003_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold65 (.A(uio_out[7]),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold66 (.A(\hopfield_inst.active_neuron[2] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold67 (.A(_010_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold68 (.A(\hopfield_inst.neuron_inst.u[0] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold69 (.A(_032_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold70 (.A(\hopfield_inst.neuron_inst.v[0] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold71 (.A(\hopfield_inst.active_neuron[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold72 (.A(_173_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold73 (.A(_007_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold74 (.A(\hopfield_inst.learning_inst.counter[0] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold75 (.A(\hopfield_inst.neuron_inst.u[6] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold76 (.A(_038_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold77 (.A(\hopfield_inst.neuron_inst.v[6] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold78 (.A(\hopfield_inst.neuron_inst.u[4] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold79 (.A(_036_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold80 (.A(\hopfield_inst.neuron_inst.v[1] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold81 (.A(_030_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold82 (.A(_037_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold83 (.A(\hopfield_inst.neuron_inst.u[2] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold84 (.A(\hopfield_inst.neuron_inst.v[2] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold85 (.A(\hopfield_inst.neuron_inst.u[3] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold86 (.A(_299_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold87 (.A(_035_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold88 (.A(_027_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold89 (.A(_294_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold90 (.A(\hopfield_inst.neuron_inst.v[5] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold91 (.A(\hopfield_inst.active_neuron[2] ),
    .X(net139));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_93 ();
 sg13g2_decap_8 FILLER_16_100 ();
 sg13g2_fill_2 FILLER_16_107 ();
 sg13g2_decap_8 FILLER_16_121 ();
 sg13g2_decap_8 FILLER_16_128 ();
 sg13g2_decap_8 FILLER_16_135 ();
 sg13g2_decap_8 FILLER_16_142 ();
 sg13g2_decap_8 FILLER_16_149 ();
 sg13g2_decap_8 FILLER_16_156 ();
 sg13g2_decap_8 FILLER_16_163 ();
 sg13g2_decap_8 FILLER_16_170 ();
 sg13g2_decap_8 FILLER_16_177 ();
 sg13g2_decap_8 FILLER_16_184 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_240 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_fill_2 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_108 ();
 sg13g2_decap_4 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_decap_8 FILLER_17_212 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_decap_8 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_111 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_decap_8 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_261 ();
 sg13g2_decap_8 FILLER_18_268 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_decap_8 FILLER_18_282 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_331 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_140 ();
 sg13g2_fill_1 FILLER_19_142 ();
 sg13g2_decap_4 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_171 ();
 sg13g2_decap_8 FILLER_19_191 ();
 sg13g2_decap_8 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_19_205 ();
 sg13g2_decap_8 FILLER_19_212 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_decap_8 FILLER_19_226 ();
 sg13g2_decap_8 FILLER_19_233 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_296 ();
 sg13g2_decap_8 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_fill_2 FILLER_20_74 ();
 sg13g2_fill_1 FILLER_20_76 ();
 sg13g2_fill_2 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_51 ();
 sg13g2_fill_2 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_fill_2 FILLER_21_66 ();
 sg13g2_decap_4 FILLER_21_92 ();
 sg13g2_fill_2 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_4 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_decap_8 FILLER_21_275 ();
 sg13g2_decap_8 FILLER_21_282 ();
 sg13g2_decap_8 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_296 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_72 ();
 sg13g2_fill_1 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_4 FILLER_22_204 ();
 sg13g2_decap_8 FILLER_22_213 ();
 sg13g2_decap_8 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_249 ();
 sg13g2_decap_4 FILLER_22_276 ();
 sg13g2_fill_1 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_4 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_68 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_decap_4 FILLER_23_139 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_decap_4 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_261 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_301 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_decap_4 FILLER_24_272 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_decap_8 FILLER_25_87 ();
 sg13g2_decap_4 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_decap_4 FILLER_25_140 ();
 sg13g2_fill_2 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_2 FILLER_25_208 ();
 sg13g2_decap_4 FILLER_25_216 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_fill_2 FILLER_25_339 ();
 sg13g2_decap_4 FILLER_25_362 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_118 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_2 FILLER_26_168 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_decap_4 FILLER_26_355 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_fill_1 FILLER_26_368 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_387 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_2 FILLER_27_138 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_157 ();
 sg13g2_decap_4 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_240 ();
 sg13g2_decap_4 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_83 ();
 sg13g2_decap_8 FILLER_28_90 ();
 sg13g2_decap_8 FILLER_28_97 ();
 sg13g2_decap_8 FILLER_28_104 ();
 sg13g2_fill_2 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_139 ();
 sg13g2_fill_2 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_387 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_86 ();
 sg13g2_fill_2 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_271 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_279 ();
 sg13g2_fill_1 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_decap_4 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_383 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_102 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_171 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_fill_2 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_decap_4 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_365 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_fill_2 FILLER_30_384 ();
 sg13g2_decap_4 FILLER_30_390 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_4 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_95 ();
 sg13g2_fill_2 FILLER_31_136 ();
 sg13g2_fill_2 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_decap_8 FILLER_31_232 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_248 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_decap_4 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_333 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_101 ();
 sg13g2_fill_1 FILLER_32_117 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_4 FILLER_32_245 ();
 sg13g2_fill_1 FILLER_32_249 ();
 sg13g2_fill_2 FILLER_32_267 ();
 sg13g2_fill_1 FILLER_32_269 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_282 ();
 sg13g2_decap_8 FILLER_32_309 ();
 sg13g2_decap_8 FILLER_32_316 ();
 sg13g2_decap_4 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_327 ();
 sg13g2_fill_2 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_decap_4 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_fill_2 FILLER_32_389 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_77 ();
 sg13g2_fill_2 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_118 ();
 sg13g2_fill_2 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_297 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_decap_4 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_decap_4 FILLER_34_242 ();
 sg13g2_fill_2 FILLER_34_246 ();
 sg13g2_decap_4 FILLER_34_262 ();
 sg13g2_fill_2 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_305 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_103 ();
 sg13g2_decap_4 FILLER_35_110 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_361 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_142 ();
 sg13g2_fill_1 FILLER_36_147 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_190 ();
 sg13g2_decap_8 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_229 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_279 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_fill_2 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_82 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_decap_4 FILLER_37_249 ();
 sg13g2_decap_8 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_decap_8 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_366 ();
 sg13g2_decap_8 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_2 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_255 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_fill_1 FILLER_38_264 ();
 sg13g2_decap_4 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net19;
 assign uio_oe[5] = net20;
 assign uio_oe[6] = net21;
 assign uio_oe[7] = net22;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uo_out[3] = net14;
 assign uo_out[4] = net15;
endmodule

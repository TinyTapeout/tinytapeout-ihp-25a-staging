module tt_um_udxs (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire \my_mlp.out[0] ;
 wire \my_mlp.out[10] ;
 wire \my_mlp.out[11] ;
 wire \my_mlp.out[12] ;
 wire \my_mlp.out[13] ;
 wire \my_mlp.out[14] ;
 wire net11;
 wire \my_mlp.out[1] ;
 wire \my_mlp.out[2] ;
 wire \my_mlp.out[3] ;
 wire \my_mlp.out[4] ;
 wire \my_mlp.out[5] ;
 wire \my_mlp.out[6] ;
 wire \my_mlp.out[7] ;
 wire \my_mlp.out[8] ;
 wire \my_mlp.out[9] ;
 wire \my_mlp.p0_bit_slice_47_comb[0] ;
 wire \my_mlp.p0_bit_slice_47_comb[10] ;
 wire \my_mlp.p0_bit_slice_47_comb[11] ;
 wire \my_mlp.p0_bit_slice_47_comb[12] ;
 wire \my_mlp.p0_bit_slice_47_comb[13] ;
 wire \my_mlp.p0_bit_slice_47_comb[14] ;
 wire \my_mlp.p0_bit_slice_47_comb[1] ;
 wire \my_mlp.p0_bit_slice_47_comb[2] ;
 wire \my_mlp.p0_bit_slice_47_comb[3] ;
 wire \my_mlp.p0_bit_slice_47_comb[4] ;
 wire \my_mlp.p0_bit_slice_47_comb[5] ;
 wire \my_mlp.p0_bit_slice_47_comb[6] ;
 wire \my_mlp.p0_bit_slice_47_comb[7] ;
 wire \my_mlp.p0_bit_slice_47_comb[8] ;
 wire \my_mlp.p0_bit_slice_47_comb[9] ;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net42;
 wire clknet_0_clk;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net43;
 wire net44;
 wire net45;

 sg13g2_inv_1 _196_ (.Y(_123_),
    .A(net9));
 sg13g2_inv_1 _197_ (.Y(_124_),
    .A(\my_mlp.p0_bit_slice_47_comb[3] ));
 sg13g2_inv_1 _198_ (.Y(_125_),
    .A(\my_mlp.p0_bit_slice_47_comb[5] ));
 sg13g2_inv_1 _199_ (.Y(_126_),
    .A(net1));
 sg13g2_nand3_1 _200_ (.B(net2),
    .C(net43),
    .A(net41),
    .Y(_127_));
 sg13g2_a21o_1 _201_ (.A2(net2),
    .A1(net41),
    .B1(net43),
    .X(_128_));
 sg13g2_and2_1 _202_ (.A(_127_),
    .B(_128_),
    .X(_129_));
 sg13g2_inv_1 _203_ (.Y(_130_),
    .A(_129_));
 sg13g2_nor2_1 _204_ (.A(net4),
    .B(_123_),
    .Y(_131_));
 sg13g2_nand3_1 _205_ (.B(net7),
    .C(net5),
    .A(net6),
    .Y(_132_));
 sg13g2_o21ai_1 _206_ (.B1(net5),
    .Y(_133_),
    .A1(net6),
    .A2(net7));
 sg13g2_nand2b_1 _207_ (.Y(_134_),
    .B(_132_),
    .A_N(_133_));
 sg13g2_nand2_1 _208_ (.Y(_135_),
    .A(net4),
    .B(net8));
 sg13g2_o21ai_1 _209_ (.B1(_132_),
    .Y(_136_),
    .A1(_133_),
    .A2(_135_));
 sg13g2_nand2_1 _210_ (.Y(_137_),
    .A(net8),
    .B(net5));
 sg13g2_xor2_1 _211_ (.B(_137_),
    .A(_134_),
    .X(_138_));
 sg13g2_xnor2_1 _212_ (.Y(_139_),
    .A(_136_),
    .B(_138_));
 sg13g2_nor3_1 _213_ (.A(net4),
    .B(_123_),
    .C(_139_),
    .Y(_140_));
 sg13g2_nand2b_1 _214_ (.Y(_141_),
    .B(net9),
    .A_N(net5));
 sg13g2_and3_1 _215_ (.X(_142_),
    .A(_133_),
    .B(_137_),
    .C(_141_));
 sg13g2_nor2_1 _216_ (.A(_140_),
    .B(_142_),
    .Y(_143_));
 sg13g2_nand3_1 _217_ (.B(net5),
    .C(net9),
    .A(net41),
    .Y(_144_));
 sg13g2_and2_1 _218_ (.A(net7),
    .B(net4),
    .X(_145_));
 sg13g2_a21o_1 _219_ (.A2(net5),
    .A1(net41),
    .B1(net9),
    .X(_146_));
 sg13g2_nand3_1 _220_ (.B(_145_),
    .C(_146_),
    .A(_144_),
    .Y(_147_));
 sg13g2_nand2_1 _221_ (.Y(_148_),
    .A(_144_),
    .B(_147_));
 sg13g2_xor2_1 _222_ (.B(_135_),
    .A(_134_),
    .X(_149_));
 sg13g2_and2_1 _223_ (.A(_148_),
    .B(_149_),
    .X(_150_));
 sg13g2_nand2b_1 _224_ (.Y(_151_),
    .B(net9),
    .A_N(net3));
 sg13g2_xnor2_1 _225_ (.Y(_152_),
    .A(_148_),
    .B(_149_));
 sg13g2_nor2_1 _226_ (.A(_151_),
    .B(_152_),
    .Y(_153_));
 sg13g2_xnor2_1 _227_ (.Y(_154_),
    .A(_131_),
    .B(_139_));
 sg13g2_o21ai_1 _228_ (.B1(_154_),
    .Y(_155_),
    .A1(_150_),
    .A2(_153_));
 sg13g2_or3_1 _229_ (.A(_150_),
    .B(_153_),
    .C(_154_),
    .X(_156_));
 sg13g2_nand2_1 _230_ (.Y(_157_),
    .A(_155_),
    .B(_156_));
 sg13g2_and4_1 _231_ (.A(net6),
    .B(net3),
    .C(net7),
    .D(net4),
    .X(_158_));
 sg13g2_nand4_1 _232_ (.B(net3),
    .C(net7),
    .A(net41),
    .Y(_159_),
    .D(net4));
 sg13g2_nand2_1 _233_ (.Y(_160_),
    .A(net2),
    .B(net8));
 sg13g2_a22oi_1 _234_ (.Y(_161_),
    .B1(net4),
    .B2(net41),
    .A2(net7),
    .A1(net3));
 sg13g2_nor3_1 _235_ (.A(_158_),
    .B(_160_),
    .C(_161_),
    .Y(_162_));
 sg13g2_o21ai_1 _236_ (.B1(_159_),
    .Y(_163_),
    .A1(_160_),
    .A2(_161_));
 sg13g2_a21o_1 _237_ (.A2(_146_),
    .A1(_144_),
    .B1(_145_),
    .X(_164_));
 sg13g2_and3_1 _238_ (.X(_165_),
    .A(_147_),
    .B(_163_),
    .C(_164_));
 sg13g2_nand2_1 _239_ (.Y(_015_),
    .A(net3),
    .B(net8));
 sg13g2_a21oi_1 _240_ (.A1(_147_),
    .A2(_164_),
    .Y(_016_),
    .B1(_163_));
 sg13g2_or3_1 _241_ (.A(_165_),
    .B(_015_),
    .C(_016_),
    .X(_017_));
 sg13g2_nand2b_1 _242_ (.Y(_018_),
    .B(_017_),
    .A_N(_165_));
 sg13g2_xor2_1 _243_ (.B(_152_),
    .A(_151_),
    .X(_019_));
 sg13g2_and2_1 _244_ (.A(_018_),
    .B(_019_),
    .X(_020_));
 sg13g2_nand4_1 _245_ (.B(net2),
    .C(net3),
    .A(net41),
    .Y(_021_),
    .D(net7));
 sg13g2_inv_1 _246_ (.Y(_022_),
    .A(_021_));
 sg13g2_o21ai_1 _247_ (.B1(_160_),
    .Y(_023_),
    .A1(_158_),
    .A2(_161_));
 sg13g2_nor2b_1 _248_ (.A(_162_),
    .B_N(_023_),
    .Y(_024_));
 sg13g2_and2_1 _249_ (.A(_022_),
    .B(_024_),
    .X(_025_));
 sg13g2_o21ai_1 _250_ (.B1(_015_),
    .Y(_026_),
    .A1(_165_),
    .A2(_016_));
 sg13g2_and3_1 _251_ (.X(_027_),
    .A(_017_),
    .B(_025_),
    .C(_026_));
 sg13g2_nand3_1 _252_ (.B(_025_),
    .C(_026_),
    .A(_017_),
    .Y(_028_));
 sg13g2_nor2_1 _253_ (.A(net2),
    .B(_123_),
    .Y(_029_));
 sg13g2_a21o_1 _254_ (.A2(_026_),
    .A1(_017_),
    .B1(_025_),
    .X(_030_));
 sg13g2_and3_1 _255_ (.X(_031_),
    .A(_028_),
    .B(_029_),
    .C(_030_));
 sg13g2_a21o_1 _256_ (.A2(_030_),
    .A1(_029_),
    .B1(_027_),
    .X(_032_));
 sg13g2_or2_1 _257_ (.X(_033_),
    .B(_019_),
    .A(_018_));
 sg13g2_xnor2_1 _258_ (.Y(_034_),
    .A(_018_),
    .B(_019_));
 sg13g2_a21oi_1 _259_ (.A1(_032_),
    .A2(_033_),
    .Y(_035_),
    .B1(_020_));
 sg13g2_o21ai_1 _260_ (.B1(_155_),
    .Y(_036_),
    .A1(_157_),
    .A2(_035_));
 sg13g2_nor3_1 _261_ (.A(_140_),
    .B(_142_),
    .C(_036_),
    .Y(_037_));
 sg13g2_nor2_1 _262_ (.A(\my_mlp.p0_bit_slice_47_comb[14] ),
    .B(net37),
    .Y(_038_));
 sg13g2_xnor2_1 _263_ (.Y(_039_),
    .A(\my_mlp.p0_bit_slice_47_comb[14] ),
    .B(net37));
 sg13g2_and2_1 _264_ (.A(\my_mlp.p0_bit_slice_47_comb[7] ),
    .B(net38),
    .X(_040_));
 sg13g2_xor2_1 _265_ (.B(_036_),
    .A(_143_),
    .X(_041_));
 sg13g2_nand2_1 _266_ (.Y(_042_),
    .A(\my_mlp.p0_bit_slice_47_comb[6] ),
    .B(_041_));
 sg13g2_xnor2_1 _267_ (.Y(_043_),
    .A(_157_),
    .B(_035_));
 sg13g2_nor2_1 _268_ (.A(_125_),
    .B(_043_),
    .Y(_044_));
 sg13g2_xnor2_1 _269_ (.Y(_045_),
    .A(_032_),
    .B(_034_));
 sg13g2_nand2_1 _270_ (.Y(_046_),
    .A(\my_mlp.p0_bit_slice_47_comb[4] ),
    .B(_045_));
 sg13g2_a21oi_1 _271_ (.A1(_028_),
    .A2(_030_),
    .Y(_047_),
    .B1(_029_));
 sg13g2_nor3_1 _272_ (.A(_124_),
    .B(_031_),
    .C(_047_),
    .Y(_048_));
 sg13g2_xnor2_1 _273_ (.Y(_049_),
    .A(_021_),
    .B(_024_));
 sg13g2_nand2_1 _274_ (.Y(_050_),
    .A(\my_mlp.p0_bit_slice_47_comb[2] ),
    .B(_049_));
 sg13g2_a22oi_1 _275_ (.Y(_051_),
    .B1(net7),
    .B2(net2),
    .A2(net3),
    .A1(net41));
 sg13g2_nor2_1 _276_ (.A(_022_),
    .B(_051_),
    .Y(_052_));
 sg13g2_xnor2_1 _277_ (.Y(_053_),
    .A(\my_mlp.p0_bit_slice_47_comb[1] ),
    .B(_052_));
 sg13g2_nor2_1 _278_ (.A(_127_),
    .B(_053_),
    .Y(_054_));
 sg13g2_a21oi_1 _279_ (.A1(\my_mlp.p0_bit_slice_47_comb[1] ),
    .A2(_052_),
    .Y(_055_),
    .B1(_054_));
 sg13g2_xnor2_1 _280_ (.Y(_056_),
    .A(net45),
    .B(_049_));
 sg13g2_o21ai_1 _281_ (.B1(_050_),
    .Y(_057_),
    .A1(_055_),
    .A2(_056_));
 sg13g2_o21ai_1 _282_ (.B1(_124_),
    .Y(_058_),
    .A1(_031_),
    .A2(_047_));
 sg13g2_nand2b_1 _283_ (.Y(_059_),
    .B(_058_),
    .A_N(_048_));
 sg13g2_a21oi_1 _284_ (.A1(_057_),
    .A2(_058_),
    .Y(_060_),
    .B1(_048_));
 sg13g2_xnor2_1 _285_ (.Y(_061_),
    .A(\my_mlp.p0_bit_slice_47_comb[4] ),
    .B(_045_));
 sg13g2_o21ai_1 _286_ (.B1(_046_),
    .Y(_062_),
    .A1(_060_),
    .A2(_061_));
 sg13g2_nand2_1 _287_ (.Y(_063_),
    .A(_125_),
    .B(_043_));
 sg13g2_nand2b_1 _288_ (.Y(_064_),
    .B(_063_),
    .A_N(_044_));
 sg13g2_a21oi_1 _289_ (.A1(_062_),
    .A2(_063_),
    .Y(_065_),
    .B1(_044_));
 sg13g2_xnor2_1 _290_ (.Y(_066_),
    .A(net44),
    .B(_041_));
 sg13g2_o21ai_1 _291_ (.B1(_042_),
    .Y(_067_),
    .A1(_065_),
    .A2(_066_));
 sg13g2_or2_1 _292_ (.X(_068_),
    .B(net38),
    .A(\my_mlp.p0_bit_slice_47_comb[7] ));
 sg13g2_nand2b_1 _293_ (.Y(_069_),
    .B(_068_),
    .A_N(_040_));
 sg13g2_a21oi_2 _294_ (.B1(_040_),
    .Y(_070_),
    .A2(_068_),
    .A1(_067_));
 sg13g2_xnor2_1 _295_ (.Y(_071_),
    .A(\my_mlp.p0_bit_slice_47_comb[11] ),
    .B(net38));
 sg13g2_and2_1 _296_ (.A(\my_mlp.p0_bit_slice_47_comb[10] ),
    .B(net38),
    .X(_072_));
 sg13g2_xnor2_1 _297_ (.Y(_073_),
    .A(\my_mlp.p0_bit_slice_47_comb[10] ),
    .B(net38));
 sg13g2_inv_1 _298_ (.Y(_074_),
    .A(_073_));
 sg13g2_xnor2_1 _299_ (.Y(_075_),
    .A(\my_mlp.p0_bit_slice_47_comb[9] ),
    .B(net37));
 sg13g2_nand2_1 _300_ (.Y(_076_),
    .A(\my_mlp.p0_bit_slice_47_comb[8] ),
    .B(_037_));
 sg13g2_xnor2_1 _301_ (.Y(_077_),
    .A(\my_mlp.p0_bit_slice_47_comb[8] ),
    .B(net38));
 sg13g2_or2_1 _302_ (.X(_078_),
    .B(_077_),
    .A(_075_));
 sg13g2_or3_1 _303_ (.A(_071_),
    .B(_073_),
    .C(_078_),
    .X(_079_));
 sg13g2_o21ai_1 _304_ (.B1(net37),
    .Y(_080_),
    .A1(\my_mlp.p0_bit_slice_47_comb[10] ),
    .A2(\my_mlp.p0_bit_slice_47_comb[11] ));
 sg13g2_o21ai_1 _305_ (.B1(net38),
    .Y(_081_),
    .A1(\my_mlp.p0_bit_slice_47_comb[8] ),
    .A2(\my_mlp.p0_bit_slice_47_comb[9] ));
 sg13g2_nor3_1 _306_ (.A(_071_),
    .B(_073_),
    .C(_081_),
    .Y(_082_));
 sg13g2_nor2b_1 _307_ (.A(_082_),
    .B_N(_080_),
    .Y(_083_));
 sg13g2_o21ai_1 _308_ (.B1(_083_),
    .Y(_084_),
    .A1(_070_),
    .A2(_079_));
 sg13g2_xnor2_1 _309_ (.Y(_085_),
    .A(\my_mlp.p0_bit_slice_47_comb[13] ),
    .B(net37));
 sg13g2_and2_1 _310_ (.A(\my_mlp.p0_bit_slice_47_comb[12] ),
    .B(net37),
    .X(_086_));
 sg13g2_xnor2_1 _311_ (.Y(_087_),
    .A(\my_mlp.p0_bit_slice_47_comb[12] ),
    .B(net37));
 sg13g2_inv_1 _312_ (.Y(_088_),
    .A(_087_));
 sg13g2_nor2_1 _313_ (.A(_085_),
    .B(_087_),
    .Y(_089_));
 sg13g2_a221oi_1 _314_ (.B2(_089_),
    .C1(_086_),
    .B1(_084_),
    .A1(\my_mlp.p0_bit_slice_47_comb[13] ),
    .Y(_090_),
    .A2(net37));
 sg13g2_nor2_1 _315_ (.A(_039_),
    .B(_090_),
    .Y(_091_));
 sg13g2_nor2_1 _316_ (.A(_038_),
    .B(_091_),
    .Y(_092_));
 sg13g2_xor2_1 _317_ (.B(_090_),
    .A(_039_),
    .X(_093_));
 sg13g2_inv_1 _318_ (.Y(_094_),
    .A(_093_));
 sg13g2_xnor2_1 _319_ (.Y(_095_),
    .A(_084_),
    .B(_088_));
 sg13g2_xor2_1 _320_ (.B(_077_),
    .A(_070_),
    .X(_096_));
 sg13g2_inv_1 _321_ (.Y(_097_),
    .A(_096_));
 sg13g2_xnor2_1 _322_ (.Y(_098_),
    .A(_065_),
    .B(_066_));
 sg13g2_xnor2_1 _323_ (.Y(_099_),
    .A(_062_),
    .B(_064_));
 sg13g2_inv_1 _324_ (.Y(_100_),
    .A(_099_));
 sg13g2_xor2_1 _325_ (.B(_061_),
    .A(_060_),
    .X(_101_));
 sg13g2_inv_1 _326_ (.Y(_102_),
    .A(_101_));
 sg13g2_xor2_1 _327_ (.B(_059_),
    .A(_057_),
    .X(_103_));
 sg13g2_xor2_1 _328_ (.B(_056_),
    .A(_055_),
    .X(_104_));
 sg13g2_inv_1 _329_ (.Y(_105_),
    .A(_104_));
 sg13g2_xor2_1 _330_ (.B(_053_),
    .A(_127_),
    .X(_106_));
 sg13g2_inv_1 _331_ (.Y(_107_),
    .A(_106_));
 sg13g2_nand2_1 _332_ (.Y(_108_),
    .A(_130_),
    .B(_103_));
 sg13g2_nor4_1 _333_ (.A(_101_),
    .B(_104_),
    .C(_106_),
    .D(_108_),
    .Y(_109_));
 sg13g2_xor2_1 _334_ (.B(_069_),
    .A(_067_),
    .X(_110_));
 sg13g2_nand4_1 _335_ (.B(_100_),
    .C(_109_),
    .A(_098_),
    .Y(_111_),
    .D(_110_));
 sg13g2_nor2_1 _336_ (.A(_096_),
    .B(_111_),
    .Y(_112_));
 sg13g2_o21ai_1 _337_ (.B1(_076_),
    .Y(_113_),
    .A1(_070_),
    .A2(_077_));
 sg13g2_xor2_1 _338_ (.B(_113_),
    .A(_075_),
    .X(_114_));
 sg13g2_o21ai_1 _339_ (.B1(_081_),
    .Y(_115_),
    .A1(_070_),
    .A2(_078_));
 sg13g2_xnor2_1 _340_ (.Y(_116_),
    .A(_074_),
    .B(_115_));
 sg13g2_nand4_1 _341_ (.B(_112_),
    .C(_114_),
    .A(_095_),
    .Y(_117_),
    .D(_116_));
 sg13g2_a21oi_1 _342_ (.A1(_074_),
    .A2(_115_),
    .Y(_118_),
    .B1(_072_));
 sg13g2_xor2_1 _343_ (.B(_118_),
    .A(_071_),
    .X(_119_));
 sg13g2_a21oi_1 _344_ (.A1(_084_),
    .A2(_088_),
    .Y(_120_),
    .B1(_086_));
 sg13g2_xor2_1 _345_ (.B(_120_),
    .A(_085_),
    .X(_121_));
 sg13g2_nor4_1 _346_ (.A(_093_),
    .B(_117_),
    .C(_119_),
    .D(_121_),
    .Y(_122_));
 sg13g2_nor3_1 _347_ (.A(_130_),
    .B(net36),
    .C(net34),
    .Y(\my_mlp.out[0] ));
 sg13g2_nor3_1 _348_ (.A(net36),
    .B(_107_),
    .C(net34),
    .Y(\my_mlp.out[1] ));
 sg13g2_nor3_1 _349_ (.A(net36),
    .B(_105_),
    .C(net34),
    .Y(\my_mlp.out[2] ));
 sg13g2_nor3_1 _350_ (.A(net36),
    .B(_103_),
    .C(net34),
    .Y(\my_mlp.out[3] ));
 sg13g2_nor3_1 _351_ (.A(net36),
    .B(_102_),
    .C(net34),
    .Y(\my_mlp.out[4] ));
 sg13g2_nor3_1 _352_ (.A(net36),
    .B(_100_),
    .C(net33),
    .Y(\my_mlp.out[5] ));
 sg13g2_nor3_1 _353_ (.A(net36),
    .B(_098_),
    .C(net33),
    .Y(\my_mlp.out[6] ));
 sg13g2_nor3_1 _354_ (.A(net35),
    .B(_110_),
    .C(net33),
    .Y(\my_mlp.out[7] ));
 sg13g2_nor3_1 _355_ (.A(net35),
    .B(_097_),
    .C(net33),
    .Y(\my_mlp.out[8] ));
 sg13g2_nor3_1 _356_ (.A(net35),
    .B(_114_),
    .C(net33),
    .Y(\my_mlp.out[9] ));
 sg13g2_nor3_1 _357_ (.A(net35),
    .B(_116_),
    .C(net33),
    .Y(\my_mlp.out[10] ));
 sg13g2_nor2b_1 _358_ (.A(net35),
    .B_N(_119_),
    .Y(\my_mlp.out[11] ));
 sg13g2_nor3_1 _359_ (.A(net35),
    .B(_095_),
    .C(net33),
    .Y(\my_mlp.out[12] ));
 sg13g2_nor2b_1 _360_ (.A(net35),
    .B_N(_121_),
    .Y(\my_mlp.out[13] ));
 sg13g2_nor3_1 _361_ (.A(net35),
    .B(_094_),
    .C(net33),
    .Y(\my_mlp.out[14] ));
 sg13g2_nor2_1 _362_ (.A(net40),
    .B(_130_),
    .Y(_000_));
 sg13g2_nor2_1 _363_ (.A(net40),
    .B(_107_),
    .Y(_001_));
 sg13g2_nor2_1 _364_ (.A(net40),
    .B(_105_),
    .Y(_002_));
 sg13g2_nor2_1 _365_ (.A(net40),
    .B(_103_),
    .Y(_003_));
 sg13g2_nor2_1 _366_ (.A(net39),
    .B(_102_),
    .Y(_004_));
 sg13g2_nor2_1 _367_ (.A(net39),
    .B(_100_),
    .Y(_005_));
 sg13g2_nor2_1 _368_ (.A(net39),
    .B(_098_),
    .Y(_006_));
 sg13g2_nor2_1 _369_ (.A(net40),
    .B(_110_),
    .Y(_007_));
 sg13g2_nor2_1 _370_ (.A(net39),
    .B(_097_),
    .Y(_008_));
 sg13g2_nor2_1 _371_ (.A(net39),
    .B(_114_),
    .Y(_009_));
 sg13g2_nor2_1 _372_ (.A(net39),
    .B(_116_),
    .Y(_010_));
 sg13g2_and2_1 _373_ (.A(net1),
    .B(_119_),
    .X(_011_));
 sg13g2_nor2_1 _374_ (.A(net39),
    .B(_095_),
    .Y(_012_));
 sg13g2_and2_1 _375_ (.A(net1),
    .B(_121_),
    .X(_013_));
 sg13g2_nor2_1 _376_ (.A(net39),
    .B(_094_),
    .Y(_014_));
 sg13g2_dfrbp_1 _377_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net19),
    .D(_000_),
    .Q_N(_180_),
    .Q(\my_mlp.p0_bit_slice_47_comb[0] ));
 sg13g2_dfrbp_1 _378_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net18),
    .D(_001_),
    .Q_N(_179_),
    .Q(\my_mlp.p0_bit_slice_47_comb[1] ));
 sg13g2_dfrbp_1 _379_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net17),
    .D(_002_),
    .Q_N(_178_),
    .Q(\my_mlp.p0_bit_slice_47_comb[2] ));
 sg13g2_dfrbp_1 _380_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net16),
    .D(_003_),
    .Q_N(_177_),
    .Q(\my_mlp.p0_bit_slice_47_comb[3] ));
 sg13g2_dfrbp_1 _381_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net15),
    .D(_004_),
    .Q_N(_176_),
    .Q(\my_mlp.p0_bit_slice_47_comb[4] ));
 sg13g2_dfrbp_1 _382_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net14),
    .D(_005_),
    .Q_N(_175_),
    .Q(\my_mlp.p0_bit_slice_47_comb[5] ));
 sg13g2_dfrbp_1 _383_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net13),
    .D(_006_),
    .Q_N(_174_),
    .Q(\my_mlp.p0_bit_slice_47_comb[6] ));
 sg13g2_dfrbp_1 _384_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net12),
    .D(_007_),
    .Q_N(_173_),
    .Q(\my_mlp.p0_bit_slice_47_comb[7] ));
 sg13g2_dfrbp_1 _385_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net11),
    .D(_008_),
    .Q_N(_172_),
    .Q(\my_mlp.p0_bit_slice_47_comb[8] ));
 sg13g2_dfrbp_1 _386_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net25),
    .D(_009_),
    .Q_N(_171_),
    .Q(\my_mlp.p0_bit_slice_47_comb[9] ));
 sg13g2_dfrbp_1 _387_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net24),
    .D(_010_),
    .Q_N(_170_),
    .Q(\my_mlp.p0_bit_slice_47_comb[10] ));
 sg13g2_dfrbp_1 _388_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net23),
    .D(_011_),
    .Q_N(_169_),
    .Q(\my_mlp.p0_bit_slice_47_comb[11] ));
 sg13g2_dfrbp_1 _389_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net22),
    .D(_012_),
    .Q_N(_168_),
    .Q(\my_mlp.p0_bit_slice_47_comb[12] ));
 sg13g2_dfrbp_1 _390_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net21),
    .D(_013_),
    .Q_N(_167_),
    .Q(\my_mlp.p0_bit_slice_47_comb[13] ));
 sg13g2_dfrbp_1 _391_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net20),
    .D(_014_),
    .Q_N(_166_),
    .Q(\my_mlp.p0_bit_slice_47_comb[14] ));
 sg13g2_tiehi _384__12 (.L_HI(net12));
 sg13g2_tiehi _383__13 (.L_HI(net13));
 sg13g2_tiehi _382__14 (.L_HI(net14));
 sg13g2_tiehi _381__15 (.L_HI(net15));
 sg13g2_tiehi _380__16 (.L_HI(net16));
 sg13g2_tiehi _379__17 (.L_HI(net17));
 sg13g2_tiehi _378__18 (.L_HI(net18));
 sg13g2_tiehi _377__19 (.L_HI(net19));
 sg13g2_tiehi _391__20 (.L_HI(net20));
 sg13g2_tiehi _390__21 (.L_HI(net21));
 sg13g2_tiehi _389__22 (.L_HI(net22));
 sg13g2_tiehi _388__23 (.L_HI(net23));
 sg13g2_tiehi _387__24 (.L_HI(net24));
 sg13g2_tiehi _386__25 (.L_HI(net25));
 sg13g2_tiehi tt_um_udxs_26 (.L_HI(net26));
 sg13g2_tiehi tt_um_udxs_27 (.L_HI(net27));
 sg13g2_tiehi tt_um_udxs_28 (.L_HI(net28));
 sg13g2_tiehi tt_um_udxs_29 (.L_HI(net29));
 sg13g2_tiehi tt_um_udxs_30 (.L_HI(net30));
 sg13g2_tiehi tt_um_udxs_31 (.L_HI(net31));
 sg13g2_tiehi tt_um_udxs_32 (.L_HI(net32));
 sg13g2_tiehi tt_um_udxs_33 (.L_HI(net42));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _385__11 (.L_HI(net11));
 sg13g2_buf_1 _416_ (.A(\my_mlp.out[8] ),
    .X(uio_out[0]));
 sg13g2_buf_1 _417_ (.A(\my_mlp.out[9] ),
    .X(uio_out[1]));
 sg13g2_buf_1 _418_ (.A(\my_mlp.out[10] ),
    .X(uio_out[2]));
 sg13g2_buf_1 _419_ (.A(\my_mlp.out[11] ),
    .X(uio_out[3]));
 sg13g2_buf_1 _420_ (.A(\my_mlp.out[12] ),
    .X(uio_out[4]));
 sg13g2_buf_1 _421_ (.A(\my_mlp.out[13] ),
    .X(uio_out[5]));
 sg13g2_buf_1 _422_ (.A(\my_mlp.out[14] ),
    .X(uio_out[6]));
 sg13g2_buf_1 _423_ (.A(net10),
    .X(uio_out[7]));
 sg13g2_buf_1 _424_ (.A(\my_mlp.out[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _425_ (.A(\my_mlp.out[1] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _426_ (.A(\my_mlp.out[2] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _427_ (.A(\my_mlp.out[3] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _428_ (.A(\my_mlp.out[4] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _429_ (.A(\my_mlp.out[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _430_ (.A(\my_mlp.out[6] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _431_ (.A(\my_mlp.out[7] ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout33 (.A(_122_),
    .X(net33));
 sg13g2_buf_1 fanout34 (.A(_122_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_092_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_092_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(net38),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_037_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_126_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_126_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(net6),
    .X(net41));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(uio_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(uio_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(uio_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[7]),
    .X(net9));
 sg13g2_tielo _423__10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\my_mlp.p0_bit_slice_47_comb[0] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold2 (.A(\my_mlp.p0_bit_slice_47_comb[6] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold3 (.A(\my_mlp.p0_bit_slice_47_comb[2] ),
    .X(net45));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_decap_8 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_decap_8 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_185 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_decap_8 FILLER_26_206 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_decap_8 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_227 ();
 sg13g2_decap_8 FILLER_26_234 ();
 sg13g2_decap_8 FILLER_26_241 ();
 sg13g2_decap_8 FILLER_26_248 ();
 sg13g2_decap_8 FILLER_26_255 ();
 sg13g2_decap_8 FILLER_26_262 ();
 sg13g2_decap_8 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_290 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_311 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_decap_8 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_decap_8 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_244 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_decap_8 FILLER_27_258 ();
 sg13g2_decap_8 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_decap_8 FILLER_27_293 ();
 sg13g2_decap_8 FILLER_27_300 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_decap_8 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_182 ();
 sg13g2_decap_4 FILLER_28_202 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_212 ();
 sg13g2_decap_8 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_240 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_261 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_decap_8 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_290 ();
 sg13g2_decap_4 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_120 ();
 sg13g2_decap_4 FILLER_30_127 ();
 sg13g2_decap_4 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_decap_8 FILLER_30_185 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_decap_8 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_324 ();
 sg13g2_decap_8 FILLER_30_331 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_decap_8 FILLER_31_152 ();
 sg13g2_decap_4 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_225 ();
 sg13g2_decap_4 FILLER_31_232 ();
 sg13g2_fill_2 FILLER_31_236 ();
 sg13g2_decap_4 FILLER_31_250 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_334 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_decap_8 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_116 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_4 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_decap_8 FILLER_32_267 ();
 sg13g2_decap_8 FILLER_32_274 ();
 sg13g2_decap_4 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_decap_8 FILLER_32_320 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_120 ();
 sg13g2_decap_4 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_decap_4 FILLER_33_149 ();
 sg13g2_fill_2 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_182 ();
 sg13g2_decap_4 FILLER_33_188 ();
 sg13g2_fill_1 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_204 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_219 ();
 sg13g2_decap_8 FILLER_33_225 ();
 sg13g2_decap_4 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_decap_8 FILLER_33_253 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_100 ();
 sg13g2_fill_2 FILLER_34_135 ();
 sg13g2_fill_1 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_197 ();
 sg13g2_fill_2 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_262 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_decap_8 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_8 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_4 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_fill_1 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_4 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_decap_4 FILLER_35_235 ();
 sg13g2_fill_2 FILLER_35_239 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_248 ();
 sg13g2_decap_4 FILLER_35_254 ();
 sg13g2_fill_2 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_274 ();
 sg13g2_fill_2 FILLER_35_281 ();
 sg13g2_decap_8 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_decap_8 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_4 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_decap_4 FILLER_36_144 ();
 sg13g2_decap_8 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_decap_4 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_fill_2 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_13 ();
 sg13g2_decap_8 FILLER_37_20 ();
 sg13g2_decap_8 FILLER_37_27 ();
 sg13g2_decap_8 FILLER_37_34 ();
 sg13g2_decap_8 FILLER_37_41 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_decap_8 FILLER_37_55 ();
 sg13g2_decap_8 FILLER_37_62 ();
 sg13g2_decap_8 FILLER_37_69 ();
 sg13g2_decap_8 FILLER_37_76 ();
 sg13g2_decap_8 FILLER_37_83 ();
 sg13g2_decap_8 FILLER_37_90 ();
 sg13g2_decap_8 FILLER_37_97 ();
 sg13g2_decap_8 FILLER_37_104 ();
 sg13g2_decap_8 FILLER_37_111 ();
 sg13g2_decap_8 FILLER_37_118 ();
 sg13g2_decap_4 FILLER_37_125 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_4 FILLER_37_196 ();
 sg13g2_fill_1 FILLER_37_204 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_251 ();
 sg13g2_fill_2 FILLER_37_258 ();
 sg13g2_decap_8 FILLER_37_269 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_decap_8 FILLER_37_283 ();
 sg13g2_decap_8 FILLER_37_290 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_decap_8 FILLER_38_130 ();
 sg13g2_decap_8 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_144 ();
 sg13g2_decap_8 FILLER_38_151 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_decap_4 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_decap_4 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_309 ();
 sg13g2_decap_8 FILLER_38_316 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_337 ();
 sg13g2_decap_8 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_4 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net26;
 assign uio_oe[1] = net27;
 assign uio_oe[2] = net28;
 assign uio_oe[3] = net29;
 assign uio_oe[4] = net30;
 assign uio_oe[5] = net31;
 assign uio_oe[6] = net32;
 assign uio_oe[7] = net42;
endmodule

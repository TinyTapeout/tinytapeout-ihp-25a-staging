module tt_um_uwasic_dinogame (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire \ai_controller_inst.button_down ;
 wire \ai_controller_inst.button_start ;
 wire \ai_controller_inst.button_up ;
 wire \ai_controller_inst.crash ;
 wire \ai_controller_inst.obstacle1_pos[2] ;
 wire \ai_controller_inst.obstacle1_pos[3] ;
 wire \ai_controller_inst.obstacle1_pos[4] ;
 wire \ai_controller_inst.obstacle1_pos[5] ;
 wire \ai_controller_inst.obstacle1_pos[6] ;
 wire \ai_controller_inst.obstacle1_pos[7] ;
 wire \ai_controller_inst.obstacle1_pos[8] ;
 wire \ai_controller_inst.obstacle1_pos[9] ;
 wire \ai_controller_inst.obstacle2_pos[2] ;
 wire \ai_controller_inst.obstacle2_pos[3] ;
 wire \ai_controller_inst.obstacle2_pos[4] ;
 wire \ai_controller_inst.obstacle2_pos[5] ;
 wire \ai_controller_inst.obstacle2_pos[6] ;
 wire \ai_controller_inst.obstacle2_pos[7] ;
 wire \ai_controller_inst.obstacle2_pos[8] ;
 wire \ai_controller_inst.obstacle2_pos[9] ;
 wire \ai_controller_inst.restart_counter[0] ;
 wire \ai_controller_inst.restart_counter[1] ;
 wire \ai_controller_inst.restart_counter[2] ;
 wire \ai_controller_inst.restart_counter[3] ;
 wire \ai_controller_inst.restart_counter[4] ;
 wire \ai_controller_inst.restart_counter[5] ;
 wire \ai_controller_inst.restart_counter[6] ;
 wire \ai_controller_inst.restart_counter[7] ;
 wire \audio_inst.game_over_sound ;
 wire \audio_inst.i_jump.active ;
 wire \audio_inst.i_jump.counter[0] ;
 wire \audio_inst.i_jump.counter[10] ;
 wire \audio_inst.i_jump.counter[11] ;
 wire \audio_inst.i_jump.counter[12] ;
 wire \audio_inst.i_jump.counter[13] ;
 wire \audio_inst.i_jump.counter[14] ;
 wire \audio_inst.i_jump.counter[15] ;
 wire \audio_inst.i_jump.counter[16] ;
 wire \audio_inst.i_jump.counter[17] ;
 wire \audio_inst.i_jump.counter[18] ;
 wire \audio_inst.i_jump.counter[1] ;
 wire \audio_inst.i_jump.counter[2] ;
 wire \audio_inst.i_jump.counter[3] ;
 wire \audio_inst.i_jump.counter[4] ;
 wire \audio_inst.i_jump.counter[5] ;
 wire \audio_inst.i_jump.counter[6] ;
 wire \audio_inst.i_jump.counter[7] ;
 wire \audio_inst.i_jump.counter[8] ;
 wire \audio_inst.i_jump.counter[9] ;
 wire \audio_inst.i_jump.decay_value[0] ;
 wire \audio_inst.i_jump.decay_value[10] ;
 wire \audio_inst.i_jump.decay_value[11] ;
 wire \audio_inst.i_jump.decay_value[12] ;
 wire \audio_inst.i_jump.decay_value[13] ;
 wire \audio_inst.i_jump.decay_value[14] ;
 wire \audio_inst.i_jump.decay_value[15] ;
 wire \audio_inst.i_jump.decay_value[16] ;
 wire \audio_inst.i_jump.decay_value[17] ;
 wire \audio_inst.i_jump.decay_value[1] ;
 wire \audio_inst.i_jump.decay_value[2] ;
 wire \audio_inst.i_jump.decay_value[3] ;
 wire \audio_inst.i_jump.decay_value[4] ;
 wire \audio_inst.i_jump.decay_value[5] ;
 wire \audio_inst.i_jump.decay_value[6] ;
 wire \audio_inst.i_jump.decay_value[7] ;
 wire \audio_inst.i_jump.decay_value[8] ;
 wire \audio_inst.i_jump.decay_value[9] ;
 wire \audio_inst.i_jump.stage_index[0] ;
 wire \audio_inst.i_jump.stage_index[1] ;
 wire \audio_inst.i_jump.stage_index[2] ;
 wire \audio_inst.i_jump.stage_index[3] ;
 wire \audio_inst.i_jump.stage_index[4] ;
 wire \audio_inst.i_jump.state[0] ;
 wire \audio_inst.i_jump.state[1] ;
 wire \audio_inst.i_jump.wave_out ;
 wire \audio_inst.i_over.active ;
 wire \audio_inst.i_over.counter[0] ;
 wire \audio_inst.i_over.counter[10] ;
 wire \audio_inst.i_over.counter[11] ;
 wire \audio_inst.i_over.counter[12] ;
 wire \audio_inst.i_over.counter[13] ;
 wire \audio_inst.i_over.counter[14] ;
 wire \audio_inst.i_over.counter[15] ;
 wire \audio_inst.i_over.counter[16] ;
 wire \audio_inst.i_over.counter[17] ;
 wire \audio_inst.i_over.counter[18] ;
 wire \audio_inst.i_over.counter[1] ;
 wire \audio_inst.i_over.counter[2] ;
 wire \audio_inst.i_over.counter[3] ;
 wire \audio_inst.i_over.counter[4] ;
 wire \audio_inst.i_over.counter[5] ;
 wire \audio_inst.i_over.counter[6] ;
 wire \audio_inst.i_over.counter[7] ;
 wire \audio_inst.i_over.counter[8] ;
 wire \audio_inst.i_over.counter[9] ;
 wire \audio_inst.i_over.decay_value[0] ;
 wire \audio_inst.i_over.decay_value[10] ;
 wire \audio_inst.i_over.decay_value[11] ;
 wire \audio_inst.i_over.decay_value[12] ;
 wire \audio_inst.i_over.decay_value[13] ;
 wire \audio_inst.i_over.decay_value[14] ;
 wire \audio_inst.i_over.decay_value[15] ;
 wire \audio_inst.i_over.decay_value[1] ;
 wire \audio_inst.i_over.decay_value[2] ;
 wire \audio_inst.i_over.decay_value[3] ;
 wire \audio_inst.i_over.decay_value[4] ;
 wire \audio_inst.i_over.decay_value[5] ;
 wire \audio_inst.i_over.decay_value[6] ;
 wire \audio_inst.i_over.decay_value[7] ;
 wire \audio_inst.i_over.decay_value[8] ;
 wire \audio_inst.i_over.decay_value[9] ;
 wire \audio_inst.i_over.stage_index[0] ;
 wire \audio_inst.i_over.stage_index[1] ;
 wire \audio_inst.i_over.stage_index[2] ;
 wire \audio_inst.i_over.stage_index[3] ;
 wire \audio_inst.i_over.stage_index[4] ;
 wire \audio_inst.i_over.state[0] ;
 wire \audio_inst.i_over.state[1] ;
 wire \audio_inst.sound ;
 wire \bg_line_inst.i_vpos[2] ;
 wire \bg_line_inst.i_vpos[3] ;
 wire \bg_line_inst.i_vpos[4] ;
 wire \bg_line_inst.i_vpos[5] ;
 wire \bg_line_inst.i_vpos[6] ;
 wire \bg_line_inst.i_vpos[7] ;
 wire \bg_line_inst.i_vpos[8] ;
 wire \bg_line_inst.i_vpos[9] ;
 wire \bg_object_inst.bg_object_pos[2] ;
 wire \bg_object_inst.bg_object_pos[3] ;
 wire \bg_object_inst.bg_object_pos[4] ;
 wire \bg_object_inst.bg_object_pos[5] ;
 wire \bg_object_inst.bg_object_pos[6] ;
 wire \bg_object_inst.bg_object_pos[7] ;
 wire \bg_object_inst.bg_object_pos[8] ;
 wire \bg_object_inst.bg_object_pos[9] ;
 wire \bg_object_rom_inst.i_rom_counter[0] ;
 wire \bg_object_rom_inst.i_rom_counter[1] ;
 wire \bg_object_rom_inst.i_rom_counter[2] ;
 wire \bg_object_rom_inst.i_rom_counter[3] ;
 wire \bg_object_rom_inst.i_rom_counter[4] ;
 wire \bg_object_rom_inst.i_rom_counter[5] ;
 wire \bg_render_inst.i_hpos[2] ;
 wire \bg_render_inst.i_hpos[3] ;
 wire \bg_render_inst.i_hpos[4] ;
 wire \bg_render_inst.i_hpos[5] ;
 wire \bg_render_inst.i_hpos[6] ;
 wire \bg_render_inst.i_hpos[7] ;
 wire \bg_render_inst.i_hpos[8] ;
 wire \bg_render_inst.i_hpos[9] ;
 wire \bg_render_inst.x_offset_r[5] ;
 wire \bg_render_inst.x_offset_r[6] ;
 wire \bg_render_inst.x_offset_r[7] ;
 wire \bg_render_inst.x_offset_r[8] ;
 wire \bg_render_inst.x_offset_r[9] ;
 wire \bg_render_inst.y_offset[2] ;
 wire \bg_render_inst.y_offset_r[5] ;
 wire \bg_render_inst.y_offset_r[6] ;
 wire \bg_render_inst.y_offset_r[7] ;
 wire \bg_render_inst.y_offset_r[8] ;
 wire \bg_render_inst.y_offset_r[9] ;
 wire \dino_inst.i_ypos[0] ;
 wire \dino_inst.i_ypos[1] ;
 wire \dino_inst.i_ypos[2] ;
 wire \dino_inst.i_ypos[3] ;
 wire \dino_inst.i_ypos[4] ;
 wire \dino_inst.i_ypos[5] ;
 wire \dino_inst.o_rom_counter[0] ;
 wire \dino_inst.o_rom_counter[1] ;
 wire \dino_inst.o_rom_counter[2] ;
 wire \dino_inst.o_rom_counter[3] ;
 wire \dino_inst.o_rom_counter[4] ;
 wire \dino_inst.o_rom_counter[5] ;
 wire \dino_inst.x_offset[3] ;
 wire \dino_inst.x_offset_r[5] ;
 wire \dino_inst.x_offset_r[6] ;
 wire \dino_inst.x_offset_r[7] ;
 wire \dino_inst.x_offset_r[8] ;
 wire \dino_inst.x_offset_r[9] ;
 wire \dino_inst.y_offset_r[5] ;
 wire \dino_inst.y_offset_r[6] ;
 wire \dino_inst.y_offset_r[7] ;
 wire \dino_inst.y_offset_r[8] ;
 wire \dino_inst.y_offset_r[9] ;
 wire \gamepad_pmod.decoder.data_reg[0] ;
 wire \gamepad_pmod.decoder.data_reg[10] ;
 wire \gamepad_pmod.decoder.data_reg[11] ;
 wire \gamepad_pmod.decoder.data_reg[1] ;
 wire \gamepad_pmod.decoder.data_reg[2] ;
 wire \gamepad_pmod.decoder.data_reg[3] ;
 wire \gamepad_pmod.decoder.data_reg[4] ;
 wire \gamepad_pmod.decoder.data_reg[5] ;
 wire \gamepad_pmod.decoder.data_reg[6] ;
 wire \gamepad_pmod.decoder.data_reg[7] ;
 wire \gamepad_pmod.decoder.data_reg[8] ;
 wire \gamepad_pmod.decoder.data_reg[9] ;
 wire \gamepad_pmod.driver.pmod_clk_prev ;
 wire \gamepad_pmod.driver.pmod_clk_sync[0] ;
 wire \gamepad_pmod.driver.pmod_clk_sync[1] ;
 wire \gamepad_pmod.driver.pmod_data_sync[0] ;
 wire \gamepad_pmod.driver.pmod_data_sync[1] ;
 wire \gamepad_pmod.driver.pmod_latch_prev ;
 wire \gamepad_pmod.driver.pmod_latch_sync[0] ;
 wire \gamepad_pmod.driver.pmod_latch_sync[1] ;
 wire \gamepad_pmod.driver.shift_reg[0] ;
 wire \gamepad_pmod.driver.shift_reg[10] ;
 wire \gamepad_pmod.driver.shift_reg[11] ;
 wire \gamepad_pmod.driver.shift_reg[1] ;
 wire \gamepad_pmod.driver.shift_reg[2] ;
 wire \gamepad_pmod.driver.shift_reg[3] ;
 wire \gamepad_pmod.driver.shift_reg[4] ;
 wire \gamepad_pmod.driver.shift_reg[5] ;
 wire \gamepad_pmod.driver.shift_reg[6] ;
 wire \gamepad_pmod.driver.shift_reg[7] ;
 wire \gamepad_pmod.driver.shift_reg[8] ;
 wire \gamepad_pmod.driver.shift_reg[9] ;
 wire \graphics_inst.B_r[0] ;
 wire \graphics_inst.B_r[1] ;
 wire \graphics_inst.G_r[0] ;
 wire \graphics_inst.G_r[1] ;
 wire \graphics_inst.R_r[1] ;
 wire \graphics_inst.color_decoder_inst.invert ;
 wire \graphics_inst.color_decoder_inst.rgb_scheme ;
 wire \graphics_inst.display_on_r ;
 wire \graphics_inst.display_on_r_r ;
 wire \graphics_inst.frame_counter[0] ;
 wire \graphics_inst.frame_counter[1] ;
 wire \graphics_inst.game_tick_r ;
 wire \graphics_inst.hpos[0] ;
 wire \graphics_inst.hpos[1] ;
 wire \graphics_inst.hsync_r ;
 wire \graphics_inst.hsync_r_r ;
 wire \graphics_inst.hvsync_gen.vpos[0] ;
 wire \graphics_inst.hvsync_gen.vpos[1] ;
 wire \graphics_inst.o_vsync ;
 wire \graphics_inst.vsync_r ;
 wire \lfsr_inst.r_lfsr[10] ;
 wire \lfsr_inst.r_lfsr[11] ;
 wire \lfsr_inst.r_lfsr[12] ;
 wire \lfsr_inst.r_lfsr[13] ;
 wire \lfsr_inst.r_lfsr[14] ;
 wire \lfsr_inst.r_lfsr[15] ;
 wire \lfsr_inst.r_lfsr[1] ;
 wire \lfsr_inst.r_lfsr[2] ;
 wire \lfsr_inst.r_lfsr[3] ;
 wire \lfsr_inst.r_lfsr[4] ;
 wire \lfsr_inst.r_lfsr[5] ;
 wire \lfsr_inst.r_lfsr[6] ;
 wire \lfsr_inst.r_lfsr[7] ;
 wire \lfsr_inst.r_lfsr[8] ;
 wire \lfsr_inst.r_lfsr[9] ;
 wire \obs_inst_1.o_rom_counter[0] ;
 wire \obs_inst_1.o_rom_counter[1] ;
 wire \obs_inst_1.o_rom_counter[2] ;
 wire \obs_inst_1.o_rom_counter[3] ;
 wire \obs_inst_1.o_rom_counter[4] ;
 wire \obs_inst_1.o_rom_counter[5] ;
 wire \obs_inst_1.o_rom_counter[6] ;
 wire \obs_inst_1.o_rom_counter[7] ;
 wire \obs_inst_1.x_offset_r[6] ;
 wire \obs_inst_1.x_offset_r[7] ;
 wire \obs_inst_1.x_offset_r[8] ;
 wire \obs_inst_1.x_offset_r[9] ;
 wire \obs_inst_1.y_offset[3] ;
 wire \obs_inst_1.y_offset_r[6] ;
 wire \obs_inst_1.y_offset_r[7] ;
 wire \obs_inst_1.y_offset_r[8] ;
 wire \obs_inst_1.y_offset_r[9] ;
 wire \obs_inst_2.o_rom_counter[0] ;
 wire \obs_inst_2.o_rom_counter[1] ;
 wire \obs_inst_2.o_rom_counter[2] ;
 wire \obs_inst_2.o_rom_counter[3] ;
 wire \obs_inst_2.x_offset_r[6] ;
 wire \obs_inst_2.x_offset_r[7] ;
 wire \obs_inst_2.x_offset_r[8] ;
 wire \obs_inst_2.x_offset_r[9] ;
 wire \obs_rom_inst_1.i_obs_type[0] ;
 wire \obs_rom_inst_1.i_obs_type[1] ;
 wire \obs_rom_inst_1.i_obs_type[2] ;
 wire \obs_rom_inst_2.i_obs_type[0] ;
 wire \obs_rom_inst_2.i_obs_type[1] ;
 wire \obs_rom_inst_2.i_obs_type[2] ;
 wire \obstacles_inst.obstacle1_cross_gen_line_reg ;
 wire \obstacles_inst.obstacle2_cross_gen_line_reg ;
 wire \player_constroller_inst.game_over ;
 wire \player_constroller_inst.game_state[0] ;
 wire \player_constroller_inst.game_state[1] ;
 wire \player_constroller_inst.game_state[2] ;
 wire \player_constroller_inst.game_state[3] ;
 wire \player_constroller_inst.game_state[5] ;
 wire \player_constroller_inst.u_player_physics.velocity[0] ;
 wire \player_constroller_inst.u_player_physics.velocity[1] ;
 wire \player_constroller_inst.u_player_physics.velocity[2] ;
 wire \player_constroller_inst.u_player_physics.velocity[3] ;
 wire \score[0] ;
 wire \score[11] ;
 wire \score[12] ;
 wire \score[13] ;
 wire \score[15] ;
 wire \score[16] ;
 wire \score[17] ;
 wire \score[18] ;
 wire \score[19] ;
 wire \score[1] ;
 wire \score[2] ;
 wire \score[3] ;
 wire \score[4] ;
 wire \score[5] ;
 wire \score[6] ;
 wire \score[7] ;
 wire \score[8] ;
 wire \score[9] ;
 wire \score_inst_1.num_r[0] ;
 wire \score_inst_1.num_r[1] ;
 wire \score_inst_1.num_r[2] ;
 wire \score_inst_1.num_r[3] ;
 wire \score_inst_1.x_offset[4] ;
 wire \score_inst_1.x_offset_r[3] ;
 wire \score_inst_1.x_offset_r[4] ;
 wire \score_inst_1.x_offset_r[5] ;
 wire \score_inst_1.x_offset_r[6] ;
 wire \score_inst_1.x_offset_r[7] ;
 wire \score_inst_1.x_offset_r[8] ;
 wire \score_inst_1.x_offset_r[9] ;
 wire \score_inst_1.y_offset_r[5] ;
 wire \score_inst_1.y_offset_r[6] ;
 wire \score_inst_1.y_offset_r[7] ;
 wire \score_inst_1.y_offset_r[8] ;
 wire \score_inst_1.y_offset_r[9] ;
 wire \score_inst_2.num_r[0] ;
 wire \score_inst_2.num_r[1] ;
 wire \score_inst_2.num_r[2] ;
 wire \score_inst_2.num_r[3] ;
 wire \score_inst_2.x_offset[2] ;
 wire \score_inst_2.x_offset_r[2] ;
 wire \score_inst_2.x_offset_r[3] ;
 wire \score_inst_2.x_offset_r[4] ;
 wire \score_inst_2.x_offset_r[5] ;
 wire \score_inst_2.x_offset_r[6] ;
 wire \score_inst_2.x_offset_r[7] ;
 wire \score_inst_2.x_offset_r[8] ;
 wire \score_inst_2.x_offset_r[9] ;
 wire \score_inst_3.num_r[0] ;
 wire \score_inst_3.num_r[1] ;
 wire \score_inst_3.num_r[2] ;
 wire \score_inst_3.num_r[3] ;
 wire \score_inst_3.x_offset_r[5] ;
 wire \score_inst_3.x_offset_r[6] ;
 wire \score_inst_3.x_offset_r[7] ;
 wire \score_inst_3.x_offset_r[8] ;
 wire \score_inst_3.x_offset_r[9] ;
 wire \score_inst_4.num_r[0] ;
 wire \score_inst_4.num_r[1] ;
 wire \score_inst_4.num_r[2] ;
 wire \score_inst_4.num_r[3] ;
 wire \score_inst_4.x_offset_r[3] ;
 wire \score_inst_4.x_offset_r[4] ;
 wire \score_inst_4.x_offset_r[5] ;
 wire \score_inst_4.x_offset_r[6] ;
 wire \score_inst_4.x_offset_r[7] ;
 wire \score_inst_4.x_offset_r[8] ;
 wire \score_inst_4.x_offset_r[9] ;
 wire \score_inst_5.num_r[0] ;
 wire \score_inst_5.num_r[1] ;
 wire \score_inst_5.num_r[2] ;
 wire \score_inst_5.num_r[3] ;
 wire \score_inst_5.x_offset[6] ;
 wire \score_inst_5.x_offset_r[4] ;
 wire \score_inst_5.x_offset_r[5] ;
 wire \score_inst_5.x_offset_r[6] ;
 wire \score_inst_5.x_offset_r[7] ;
 wire \score_inst_5.x_offset_r[8] ;
 wire \score_inst_5.x_offset_r[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_leaf_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;

 sg13g2_inv_1 _2902_ (.Y(_1993_),
    .A(net447));
 sg13g2_inv_1 _2903_ (.Y(_1994_),
    .A(net632));
 sg13g2_inv_1 _2904_ (.Y(_1995_),
    .A(net694));
 sg13g2_inv_1 _2905_ (.Y(_1996_),
    .A(net640));
 sg13g2_inv_1 _2906_ (.Y(_1997_),
    .A(net681));
 sg13g2_inv_1 _2907_ (.Y(_1998_),
    .A(net650));
 sg13g2_inv_1 _2908_ (.Y(_1999_),
    .A(net644));
 sg13g2_inv_1 _2909_ (.Y(_2000_),
    .A(net718));
 sg13g2_inv_1 _2910_ (.Y(_2001_),
    .A(net733));
 sg13g2_inv_1 _2911_ (.Y(_2002_),
    .A(net683));
 sg13g2_inv_1 _2912_ (.Y(_2003_),
    .A(net664));
 sg13g2_inv_1 _2913_ (.Y(_2004_),
    .A(net637));
 sg13g2_inv_1 _2914_ (.Y(_2005_),
    .A(\gamepad_pmod.driver.shift_reg[0] ));
 sg13g2_inv_2 _2915_ (.Y(_2006_),
    .A(net524));
 sg13g2_inv_1 _2916_ (.Y(_2007_),
    .A(net526));
 sg13g2_inv_1 _2917_ (.Y(_2008_),
    .A(net897));
 sg13g2_inv_1 _2918_ (.Y(_2009_),
    .A(\audio_inst.i_over.counter[14] ));
 sg13g2_inv_1 _2919_ (.Y(_2010_),
    .A(\audio_inst.i_over.counter[9] ));
 sg13g2_inv_1 _2920_ (.Y(_2011_),
    .A(\audio_inst.i_over.counter[8] ));
 sg13g2_inv_1 _2921_ (.Y(_2012_),
    .A(\audio_inst.i_over.counter[7] ));
 sg13g2_inv_1 _2922_ (.Y(_2013_),
    .A(\audio_inst.i_over.counter[5] ));
 sg13g2_inv_1 _2923_ (.Y(_2014_),
    .A(\audio_inst.i_over.counter[3] ));
 sg13g2_inv_1 _2924_ (.Y(_2015_),
    .A(\audio_inst.i_over.counter[2] ));
 sg13g2_inv_1 _2925_ (.Y(_2016_),
    .A(\audio_inst.i_over.counter[1] ));
 sg13g2_inv_1 _2926_ (.Y(_2017_),
    .A(\audio_inst.i_over.counter[0] ));
 sg13g2_inv_1 _2927_ (.Y(_2018_),
    .A(net536));
 sg13g2_inv_1 _2928_ (.Y(_2019_),
    .A(net466));
 sg13g2_inv_1 _2929_ (.Y(_2020_),
    .A(net673));
 sg13g2_inv_2 _2930_ (.Y(_2021_),
    .A(net463));
 sg13g2_inv_1 _2931_ (.Y(_2022_),
    .A(net668));
 sg13g2_inv_1 _2932_ (.Y(_2023_),
    .A(net771));
 sg13g2_inv_1 _2933_ (.Y(_2024_),
    .A(net461));
 sg13g2_inv_1 _2934_ (.Y(_2025_),
    .A(net457));
 sg13g2_inv_2 _2935_ (.Y(_2026_),
    .A(net462));
 sg13g2_inv_1 _2936_ (.Y(_2027_),
    .A(net392));
 sg13g2_inv_1 _2937_ (.Y(_2028_),
    .A(net869));
 sg13g2_inv_1 _2938_ (.Y(_2029_),
    .A(net824));
 sg13g2_inv_1 _2939_ (.Y(_2030_),
    .A(\ai_controller_inst.obstacle1_pos[6] ));
 sg13g2_inv_1 _2940_ (.Y(_2031_),
    .A(\ai_controller_inst.obstacle1_pos[5] ));
 sg13g2_inv_1 _2941_ (.Y(_2032_),
    .A(\obs_rom_inst_1.i_obs_type[1] ));
 sg13g2_inv_1 _2942_ (.Y(_2033_),
    .A(\obs_rom_inst_1.i_obs_type[0] ));
 sg13g2_inv_1 _2943_ (.Y(_2034_),
    .A(net574));
 sg13g2_inv_1 _2944_ (.Y(_2035_),
    .A(net711));
 sg13g2_inv_1 _2945_ (.Y(_2036_),
    .A(net766));
 sg13g2_inv_1 _2946_ (.Y(_2037_),
    .A(net699));
 sg13g2_inv_1 _2947_ (.Y(_2038_),
    .A(\dino_inst.i_ypos[1] ));
 sg13g2_inv_1 _2948_ (.Y(_2039_),
    .A(net420));
 sg13g2_inv_2 _2949_ (.Y(_2040_),
    .A(_0006_));
 sg13g2_inv_1 _2950_ (.Y(_2041_),
    .A(net556));
 sg13g2_inv_1 _2951_ (.Y(_2042_),
    .A(net554));
 sg13g2_inv_2 _2952_ (.Y(_2043_),
    .A(net873));
 sg13g2_inv_2 _2953_ (.Y(_2044_),
    .A(\bg_line_inst.i_vpos[8] ));
 sg13g2_inv_2 _2954_ (.Y(_2045_),
    .A(net859));
 sg13g2_inv_4 _2955_ (.A(net591),
    .Y(_2046_));
 sg13g2_inv_2 _2956_ (.Y(_2047_),
    .A(net583));
 sg13g2_inv_2 _2957_ (.Y(_2048_),
    .A(net579));
 sg13g2_inv_1 _2958_ (.Y(_2049_),
    .A(net547));
 sg13g2_inv_1 _2959_ (.Y(_2050_),
    .A(net798));
 sg13g2_inv_1 _2960_ (.Y(_2051_),
    .A(net620));
 sg13g2_inv_1 _2961_ (.Y(_2052_),
    .A(net449));
 sg13g2_inv_1 _2962_ (.Y(_2053_),
    .A(net430));
 sg13g2_inv_1 _2963_ (.Y(_2054_),
    .A(net418));
 sg13g2_inv_1 _2964_ (.Y(_2055_),
    .A(net468));
 sg13g2_inv_1 _2965_ (.Y(_2056_),
    .A(net411));
 sg13g2_inv_1 _2966_ (.Y(_2057_),
    .A(net439));
 sg13g2_inv_1 _2967_ (.Y(_2058_),
    .A(net654));
 sg13g2_inv_1 _2968_ (.Y(_2059_),
    .A(net671));
 sg13g2_inv_1 _2969_ (.Y(_2060_),
    .A(net655));
 sg13g2_inv_1 _2970_ (.Y(_2061_),
    .A(net428));
 sg13g2_inv_1 _2971_ (.Y(_2062_),
    .A(net436));
 sg13g2_inv_1 _2972_ (.Y(_2063_),
    .A(net642));
 sg13g2_inv_1 _2973_ (.Y(_2064_),
    .A(net465));
 sg13g2_inv_1 _2974_ (.Y(_2065_),
    .A(net634));
 sg13g2_inv_1 _2975_ (.Y(_2066_),
    .A(net685));
 sg13g2_inv_1 _2976_ (.Y(_2067_),
    .A(\audio_inst.i_jump.counter[4] ));
 sg13g2_inv_1 _2977_ (.Y(_2068_),
    .A(net639));
 sg13g2_inv_1 _2978_ (.Y(_2069_),
    .A(\audio_inst.i_jump.counter[16] ));
 sg13g2_inv_1 _2979_ (.Y(_2070_),
    .A(net774));
 sg13g2_inv_1 _2980_ (.Y(_2071_),
    .A(\audio_inst.i_jump.decay_value[2] ));
 sg13g2_inv_1 _2981_ (.Y(_2072_),
    .A(net666));
 sg13g2_inv_1 _2982_ (.Y(_2073_),
    .A(\audio_inst.i_jump.decay_value[6] ));
 sg13g2_inv_1 _2983_ (.Y(_2074_),
    .A(\audio_inst.i_jump.decay_value[7] ));
 sg13g2_inv_1 _2984_ (.Y(_2075_),
    .A(\audio_inst.i_jump.decay_value[4] ));
 sg13g2_inv_1 _2985_ (.Y(_2076_),
    .A(\audio_inst.i_jump.decay_value[5] ));
 sg13g2_inv_1 _2986_ (.Y(_2077_),
    .A(net661));
 sg13g2_inv_1 _2987_ (.Y(_2078_),
    .A(net464));
 sg13g2_inv_1 _2988_ (.Y(_2079_),
    .A(\audio_inst.i_jump.decay_value[10] ));
 sg13g2_inv_1 _2989_ (.Y(_2080_),
    .A(net680));
 sg13g2_inv_1 _2990_ (.Y(_2081_),
    .A(net772));
 sg13g2_inv_1 _2991_ (.Y(_2082_),
    .A(net763));
 sg13g2_inv_1 _2992_ (.Y(_2083_),
    .A(net749));
 sg13g2_inv_1 _2993_ (.Y(_2084_),
    .A(net709));
 sg13g2_inv_1 _2994_ (.Y(_2085_),
    .A(net696));
 sg13g2_inv_1 _2995_ (.Y(_2086_),
    .A(net407));
 sg13g2_inv_2 _2996_ (.Y(_2087_),
    .A(_0009_));
 sg13g2_inv_1 _2997_ (.Y(_2088_),
    .A(net576));
 sg13g2_inv_1 _2998_ (.Y(_2089_),
    .A(\obs_inst_1.o_rom_counter[2] ));
 sg13g2_inv_1 _2999_ (.Y(_2090_),
    .A(\obs_inst_1.o_rom_counter[3] ));
 sg13g2_inv_1 _3000_ (.Y(_2091_),
    .A(net559));
 sg13g2_inv_1 _3001_ (.Y(_2092_),
    .A(\obs_inst_1.o_rom_counter[1] ));
 sg13g2_inv_2 _3002_ (.Y(_2093_),
    .A(net561));
 sg13g2_inv_2 _3003_ (.Y(_2094_),
    .A(net564));
 sg13g2_inv_2 _3004_ (.Y(_2095_),
    .A(net565));
 sg13g2_inv_1 _3005_ (.Y(_2096_),
    .A(\obs_inst_2.o_rom_counter[3] ));
 sg13g2_inv_1 _3006_ (.Y(_2097_),
    .A(\obs_inst_2.o_rom_counter[2] ));
 sg13g2_inv_1 _3007_ (.Y(_2098_),
    .A(\obs_inst_2.o_rom_counter[1] ));
 sg13g2_inv_1 _3008_ (.Y(_2099_),
    .A(net571));
 sg13g2_inv_1 _3009_ (.Y(_2100_),
    .A(\dino_inst.o_rom_counter[1] ));
 sg13g2_inv_1 _3010_ (.Y(_2101_),
    .A(net569));
 sg13g2_inv_1 _3011_ (.Y(_2102_),
    .A(_0015_));
 sg13g2_inv_1 _3012_ (.Y(_2103_),
    .A(\bg_object_rom_inst.i_rom_counter[2] ));
 sg13g2_inv_1 _3013_ (.Y(_2104_),
    .A(\bg_object_rom_inst.i_rom_counter[0] ));
 sg13g2_inv_1 _3014_ (.Y(_2105_),
    .A(net558));
 sg13g2_inv_1 _3015_ (.Y(_2106_),
    .A(_0025_));
 sg13g2_inv_1 _3016_ (.Y(_2107_),
    .A(\score_inst_1.num_r[1] ));
 sg13g2_inv_1 _3017_ (.Y(_2108_),
    .A(\score_inst_2.num_r[3] ));
 sg13g2_inv_1 _3018_ (.Y(_2109_),
    .A(\score_inst_3.num_r[1] ));
 sg13g2_inv_1 _3019_ (.Y(_2110_),
    .A(\score_inst_3.num_r[0] ));
 sg13g2_inv_1 _3020_ (.Y(_2111_),
    .A(\score_inst_3.num_r[2] ));
 sg13g2_inv_1 _3021_ (.Y(_2112_),
    .A(\score_inst_3.num_r[3] ));
 sg13g2_inv_1 _3022_ (.Y(_2113_),
    .A(\score_inst_4.num_r[0] ));
 sg13g2_inv_1 _3023_ (.Y(_2114_),
    .A(\score_inst_4.num_r[2] ));
 sg13g2_inv_1 _3024_ (.Y(_2115_),
    .A(\score_inst_4.num_r[3] ));
 sg13g2_inv_1 _3025_ (.Y(_2116_),
    .A(\score_inst_5.num_r[1] ));
 sg13g2_inv_2 _3026_ (.Y(_2117_),
    .A(_0023_));
 sg13g2_inv_1 _3027_ (.Y(_2118_),
    .A(_0028_));
 sg13g2_inv_1 _3028_ (.Y(_2119_),
    .A(net845));
 sg13g2_inv_1 _3029_ (.Y(_2120_),
    .A(net830));
 sg13g2_inv_1 _3030_ (.Y(_2121_),
    .A(net855));
 sg13g2_inv_1 _3031_ (.Y(_2122_),
    .A(net901));
 sg13g2_nor2_2 _3032_ (.A(\player_constroller_inst.game_state[2] ),
    .B(\player_constroller_inst.game_state[5] ),
    .Y(_2123_));
 sg13g2_or2_1 _3033_ (.X(_2124_),
    .B(\player_constroller_inst.game_state[5] ),
    .A(\player_constroller_inst.game_state[2] ));
 sg13g2_or2_2 _3034_ (.X(_2125_),
    .B(net595),
    .A(net592));
 sg13g2_or2_2 _3035_ (.X(_2126_),
    .B(\bg_line_inst.i_vpos[9] ),
    .A(\bg_line_inst.i_vpos[8] ));
 sg13g2_nor4_1 _3036_ (.A(net581),
    .B(net578),
    .C(_2125_),
    .D(_2126_),
    .Y(_2127_));
 sg13g2_nor3_1 _3037_ (.A(net590),
    .B(net589),
    .C(net585),
    .Y(_2128_));
 sg13g2_or2_1 _3038_ (.X(_2129_),
    .B(net866),
    .A(net817));
 sg13g2_nor3_1 _3039_ (.A(\graphics_inst.hpos[0] ),
    .B(\graphics_inst.hpos[1] ),
    .C(net577),
    .Y(_2130_));
 sg13g2_nor2_1 _3040_ (.A(net549),
    .B(net551),
    .Y(_2131_));
 sg13g2_nor4_2 _3041_ (.A(net553),
    .B(net554),
    .C(net550),
    .Y(_2132_),
    .D(net551));
 sg13g2_nor4_2 _3042_ (.A(\graphics_inst.hvsync_gen.vpos[0] ),
    .B(\graphics_inst.hvsync_gen.vpos[1] ),
    .C(net555),
    .Y(_2133_),
    .D(net557));
 sg13g2_and4_1 _3043_ (.A(_2128_),
    .B(_2130_),
    .C(_2132_),
    .D(_2133_),
    .X(_2134_));
 sg13g2_and2_2 _3044_ (.A(_2127_),
    .B(_2134_),
    .X(_2135_));
 sg13g2_and4_1 _3045_ (.A(_2025_),
    .B(\graphics_inst.frame_counter[0] ),
    .C(_2127_),
    .D(_2134_),
    .X(_2136_));
 sg13g2_nand3_1 _3046_ (.B(\graphics_inst.frame_counter[0] ),
    .C(net501),
    .A(_2025_),
    .Y(_2137_));
 sg13g2_nor2_1 _3047_ (.A(_2123_),
    .B(net497),
    .Y(_2138_));
 sg13g2_nor2_1 _3048_ (.A(net795),
    .B(_2138_),
    .Y(_2139_));
 sg13g2_nor2_2 _3049_ (.A(net462),
    .B(net597),
    .Y(_2140_));
 sg13g2_nand2_2 _3050_ (.Y(_2141_),
    .A(_2026_),
    .B(net607));
 sg13g2_nor2_2 _3051_ (.A(net522),
    .B(net497),
    .Y(_2142_));
 sg13g2_nor3_1 _3052_ (.A(_2139_),
    .B(_2141_),
    .C(_2142_),
    .Y(_0001_));
 sg13g2_and2_1 _3053_ (.A(\ai_controller_inst.button_start ),
    .B(net499),
    .X(_2143_));
 sg13g2_nand2_1 _3054_ (.Y(_2144_),
    .A(net800),
    .B(net500));
 sg13g2_a21o_1 _3055_ (.A2(_2144_),
    .A1(net636),
    .B1(net597),
    .X(_0000_));
 sg13g2_o21ai_1 _3056_ (.B1(\player_constroller_inst.u_player_physics.velocity[3] ),
    .Y(_2145_),
    .A1(\dino_inst.i_ypos[4] ),
    .A2(_2049_));
 sg13g2_nand3_1 _3057_ (.B(\dino_inst.i_ypos[3] ),
    .C(net548),
    .A(\player_constroller_inst.u_player_physics.velocity[3] ),
    .Y(_2146_));
 sg13g2_nor2_1 _3058_ (.A(net521),
    .B(_2146_),
    .Y(_2147_));
 sg13g2_and2_1 _3059_ (.A(net521),
    .B(net547),
    .X(_2148_));
 sg13g2_nand2_1 _3060_ (.Y(_2149_),
    .A(net521),
    .B(net547));
 sg13g2_a22oi_1 _3061_ (.Y(_2150_),
    .B1(_2149_),
    .B2(\player_constroller_inst.u_player_physics.velocity[3] ),
    .A2(net548),
    .A1(\dino_inst.i_ypos[3] ));
 sg13g2_nor2_1 _3062_ (.A(_2147_),
    .B(_2150_),
    .Y(_2151_));
 sg13g2_and2_1 _3063_ (.A(\dino_inst.i_ypos[2] ),
    .B(net547),
    .X(_2152_));
 sg13g2_o21ai_1 _3064_ (.B1(_2152_),
    .Y(_2153_),
    .A1(net521),
    .A2(\player_constroller_inst.u_player_physics.velocity[2] ));
 sg13g2_nand2b_1 _3065_ (.Y(_2154_),
    .B(_2149_),
    .A_N(\player_constroller_inst.u_player_physics.velocity[2] ));
 sg13g2_o21ai_1 _3066_ (.B1(_2153_),
    .Y(_2155_),
    .A1(_2152_),
    .A2(_2154_));
 sg13g2_nor2_1 _3067_ (.A(net521),
    .B(\player_constroller_inst.u_player_physics.velocity[1] ),
    .Y(_2156_));
 sg13g2_nor3_1 _3068_ (.A(_2038_),
    .B(_2049_),
    .C(_2156_),
    .Y(_2157_));
 sg13g2_o21ai_1 _3069_ (.B1(net547),
    .Y(_2158_),
    .A1(net521),
    .A2(\dino_inst.i_ypos[1] ));
 sg13g2_nand2b_1 _3070_ (.Y(_2159_),
    .B(_2158_),
    .A_N(\player_constroller_inst.u_player_physics.velocity[1] ));
 sg13g2_nand2b_1 _3071_ (.Y(_2160_),
    .B(_2159_),
    .A_N(_2157_));
 sg13g2_nor2b_1 _3072_ (.A(\dino_inst.i_ypos[0] ),
    .B_N(net547),
    .Y(_2161_));
 sg13g2_nor3_2 _3073_ (.A(_2037_),
    .B(_2148_),
    .C(_2161_),
    .Y(_2162_));
 sg13g2_a21oi_1 _3074_ (.A1(_2159_),
    .A2(_2162_),
    .Y(_2163_),
    .B1(_2157_));
 sg13g2_o21ai_1 _3075_ (.B1(_2153_),
    .Y(_2164_),
    .A1(_2155_),
    .A2(_2163_));
 sg13g2_a21oi_1 _3076_ (.A1(_2151_),
    .A2(_2164_),
    .Y(_2165_),
    .B1(_2147_));
 sg13g2_and2_1 _3077_ (.A(\dino_inst.i_ypos[4] ),
    .B(net547),
    .X(_2166_));
 sg13g2_o21ai_1 _3078_ (.B1(_2145_),
    .Y(_2167_),
    .A1(\player_constroller_inst.u_player_physics.velocity[3] ),
    .A2(_2166_));
 sg13g2_o21ai_1 _3079_ (.B1(_2145_),
    .Y(_2168_),
    .A1(_2165_),
    .A2(_2167_));
 sg13g2_o21ai_1 _3080_ (.B1(net547),
    .Y(_2169_),
    .A1(\player_constroller_inst.u_player_physics.velocity[3] ),
    .A2(net575));
 sg13g2_a21oi_1 _3081_ (.A1(\player_constroller_inst.u_player_physics.velocity[3] ),
    .A2(net575),
    .Y(_2170_),
    .B1(_2169_));
 sg13g2_xnor2_1 _3082_ (.Y(_2171_),
    .A(_2168_),
    .B(_2170_));
 sg13g2_nand2_1 _3083_ (.Y(_2172_),
    .A(net838),
    .B(_2140_));
 sg13g2_nand4_1 _3084_ (.B(net838),
    .C(_2140_),
    .A(net548),
    .Y(_2173_),
    .D(_2171_));
 sg13g2_nand3_1 _3085_ (.B(net724),
    .C(_2143_),
    .A(net607),
    .Y(_2174_));
 sg13g2_nor4_1 _3086_ (.A(\ai_controller_inst.button_up ),
    .B(net521),
    .C(net497),
    .D(_2141_),
    .Y(_2175_));
 sg13g2_and3_1 _3087_ (.X(_2176_),
    .A(\player_constroller_inst.game_state[1] ),
    .B(_2140_),
    .C(_2142_));
 sg13g2_nor2_1 _3088_ (.A(net499),
    .B(_2141_),
    .Y(_2177_));
 sg13g2_a221oi_1 _3089_ (.B2(\player_constroller_inst.game_state[2] ),
    .C1(_2176_),
    .B1(_2177_),
    .A1(net757),
    .Y(_2178_),
    .A2(_2175_));
 sg13g2_nand3_1 _3090_ (.B(_2174_),
    .C(_2178_),
    .A(_2173_),
    .Y(_0002_));
 sg13g2_a22oi_1 _3091_ (.Y(_2179_),
    .B1(_2177_),
    .B2(net757),
    .A2(_2175_),
    .A1(\player_constroller_inst.game_state[2] ));
 sg13g2_inv_1 _3092_ (.Y(_0005_),
    .A(net758));
 sg13g2_a21oi_1 _3093_ (.A1(net548),
    .A2(_2171_),
    .Y(_2180_),
    .B1(_2172_));
 sg13g2_and2_2 _3094_ (.A(\ai_controller_inst.button_up ),
    .B(_2138_),
    .X(_2181_));
 sg13g2_nand2_2 _3095_ (.Y(_2182_),
    .A(\ai_controller_inst.button_up ),
    .B(_2138_));
 sg13g2_a21oi_1 _3096_ (.A1(net522),
    .A2(net499),
    .Y(_2183_),
    .B1(_2141_));
 sg13g2_a21oi_1 _3097_ (.A1(_2181_),
    .A2(_2183_),
    .Y(_2184_),
    .B1(net839));
 sg13g2_nand3_1 _3098_ (.B(net636),
    .C(_2143_),
    .A(net607),
    .Y(_2185_));
 sg13g2_nand2_1 _3099_ (.Y(_0003_),
    .A(_2184_),
    .B(_2185_));
 sg13g2_nor2_1 _3100_ (.A(\player_constroller_inst.game_state[1] ),
    .B(_2124_),
    .Y(_2186_));
 sg13g2_nand2b_2 _3101_ (.Y(_2187_),
    .B(_2123_),
    .A_N(\player_constroller_inst.game_state[1] ));
 sg13g2_nand2b_1 _3102_ (.Y(_2188_),
    .B(net513),
    .A_N(\player_constroller_inst.game_state[3] ));
 sg13g2_a22oi_1 _3103_ (.Y(_2189_),
    .B1(_2188_),
    .B2(net462),
    .A2(_2144_),
    .A1(net724));
 sg13g2_nor2_1 _3104_ (.A(net597),
    .B(net725),
    .Y(_0004_));
 sg13g2_and2_1 _3105_ (.A(\graphics_inst.display_on_r_r ),
    .B(\graphics_inst.B_r[1] ),
    .X(uo_out[4]));
 sg13g2_and2_1 _3106_ (.A(\graphics_inst.display_on_r_r ),
    .B(\graphics_inst.R_r[1] ),
    .X(uo_out[0]));
 sg13g2_and2_1 _3107_ (.A(\graphics_inst.display_on_r_r ),
    .B(\graphics_inst.G_r[0] ),
    .X(uo_out[5]));
 sg13g2_and2_1 _3108_ (.A(\graphics_inst.display_on_r_r ),
    .B(\graphics_inst.G_r[1] ),
    .X(uo_out[1]));
 sg13g2_and2_1 _3109_ (.A(\graphics_inst.display_on_r_r ),
    .B(\graphics_inst.B_r[0] ),
    .X(uo_out[6]));
 sg13g2_nor2b_2 _3110_ (.A(net535),
    .B_N(net532),
    .Y(_2190_));
 sg13g2_nand2b_1 _3111_ (.Y(_2191_),
    .B(net532),
    .A_N(net534));
 sg13g2_nand2_1 _3112_ (.Y(_2192_),
    .A(net527),
    .B(net530));
 sg13g2_inv_1 _3113_ (.Y(_2193_),
    .A(_2192_));
 sg13g2_nand3_1 _3114_ (.B(_2190_),
    .C(_2193_),
    .A(net525),
    .Y(_2194_));
 sg13g2_nor2_2 _3115_ (.A(_2050_),
    .B(net893),
    .Y(_2195_));
 sg13g2_nand2_1 _3116_ (.Y(_2196_),
    .A(net608),
    .B(_2195_));
 sg13g2_nor2_1 _3117_ (.A(_2194_),
    .B(_2196_),
    .Y(_0036_));
 sg13g2_nand2_1 _3118_ (.Y(_2197_),
    .A(_2194_),
    .B(_2195_));
 sg13g2_nand2b_1 _3119_ (.Y(_2198_),
    .B(net629),
    .A_N(\audio_inst.i_jump.state[1] ));
 sg13g2_o21ai_1 _3120_ (.B1(_2197_),
    .Y(_2199_),
    .A1(net798),
    .A2(_2198_));
 sg13g2_and2_1 _3121_ (.A(net608),
    .B(net799),
    .X(_0037_));
 sg13g2_nor2_2 _3122_ (.A(\audio_inst.i_over.state[1] ),
    .B(\audio_inst.i_over.state[0] ),
    .Y(_2200_));
 sg13g2_and2_2 _3123_ (.A(\audio_inst.i_over.state[1] ),
    .B(\audio_inst.i_over.state[0] ),
    .X(_2201_));
 sg13g2_nand2_2 _3124_ (.Y(_2202_),
    .A(\audio_inst.i_over.state[1] ),
    .B(\audio_inst.i_over.state[0] ));
 sg13g2_nor2_2 _3125_ (.A(_2200_),
    .B(_2201_),
    .Y(_2203_));
 sg13g2_nand2_1 _3126_ (.Y(_2204_),
    .A(net619),
    .B(_2203_));
 sg13g2_nand2_2 _3127_ (.Y(_2205_),
    .A(net541),
    .B(net545));
 sg13g2_nand4_1 _3128_ (.B(net543),
    .C(net544),
    .A(net538),
    .Y(_0394_),
    .D(net546));
 sg13g2_nor2_1 _3129_ (.A(\audio_inst.i_over.stage_index[4] ),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_nor2_1 _3130_ (.A(net867),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_nor2_1 _3131_ (.A(_2204_),
    .B(net868),
    .Y(_0038_));
 sg13g2_and2_1 _3132_ (.A(net422),
    .B(net611),
    .X(_0039_));
 sg13g2_and2_1 _3133_ (.A(net750),
    .B(net611),
    .X(_0040_));
 sg13g2_and2_1 _3134_ (.A(net715),
    .B(net611),
    .X(_0041_));
 sg13g2_nor2_1 _3135_ (.A(_2024_),
    .B(net596),
    .Y(_0042_));
 sg13g2_nand2_2 _3136_ (.Y(_0397_),
    .A(net817),
    .B(net866));
 sg13g2_nand2_2 _3137_ (.Y(_0398_),
    .A(net592),
    .B(net590));
 sg13g2_nand2_2 _3138_ (.Y(_0399_),
    .A(net592),
    .B(net595));
 sg13g2_nand3_1 _3139_ (.B(net595),
    .C(net590),
    .A(net592),
    .Y(_0400_));
 sg13g2_or2_2 _3140_ (.X(_0401_),
    .B(_0399_),
    .A(_0397_));
 sg13g2_nor2_1 _3141_ (.A(_0397_),
    .B(_0400_),
    .Y(_0402_));
 sg13g2_nor3_1 _3142_ (.A(net588),
    .B(net585),
    .C(net581),
    .Y(_0403_));
 sg13g2_nand2_1 _3143_ (.Y(_0404_),
    .A(net578),
    .B(net577));
 sg13g2_nand4_1 _3144_ (.B(net577),
    .C(_0402_),
    .A(net578),
    .Y(_0405_),
    .D(_0403_));
 sg13g2_and2_1 _3145_ (.A(net616),
    .B(_0405_),
    .X(_0406_));
 sg13g2_nand2_2 _3146_ (.Y(_0407_),
    .A(net612),
    .B(_0405_));
 sg13g2_and2_1 _3147_ (.A(net387),
    .B(_0406_),
    .X(_0043_));
 sg13g2_and3_1 _3148_ (.X(_0044_),
    .A(net612),
    .B(_2129_),
    .C(net818));
 sg13g2_xor2_1 _3149_ (.B(net818),
    .A(net595),
    .X(_0408_));
 sg13g2_nor2_1 _3150_ (.A(_0407_),
    .B(_0408_),
    .Y(_0045_));
 sg13g2_nor2_1 _3151_ (.A(net667),
    .B(_0397_),
    .Y(_0409_));
 sg13g2_xnor2_1 _3152_ (.Y(_0410_),
    .A(net592),
    .B(net819));
 sg13g2_nor2_1 _3153_ (.A(_0407_),
    .B(_0410_),
    .Y(_0046_));
 sg13g2_o21ai_1 _3154_ (.B1(net613),
    .Y(_0411_),
    .A1(net818),
    .A2(_0400_));
 sg13g2_a21oi_1 _3155_ (.A1(_2046_),
    .A2(_0401_),
    .Y(_0047_),
    .B1(_0411_));
 sg13g2_nor2_1 _3156_ (.A(net845),
    .B(_0399_),
    .Y(_0412_));
 sg13g2_nor2_1 _3157_ (.A(net845),
    .B(_0401_),
    .Y(_0413_));
 sg13g2_xnor2_1 _3158_ (.Y(_0414_),
    .A(net588),
    .B(_0413_));
 sg13g2_nor2_1 _3159_ (.A(_0407_),
    .B(_0414_),
    .Y(_0048_));
 sg13g2_and2_2 _3160_ (.A(net590),
    .B(net588),
    .X(_0415_));
 sg13g2_nand2_2 _3161_ (.Y(_0416_),
    .A(net590),
    .B(net589));
 sg13g2_nand2_1 _3162_ (.Y(_0417_),
    .A(net594),
    .B(_0415_));
 sg13g2_nor2_2 _3163_ (.A(_0401_),
    .B(_0416_),
    .Y(_0418_));
 sg13g2_xnor2_1 _3164_ (.Y(_0419_),
    .A(net585),
    .B(_0418_));
 sg13g2_nor2_1 _3165_ (.A(_0407_),
    .B(_0419_),
    .Y(_0049_));
 sg13g2_nor3_1 _3166_ (.A(net830),
    .B(_0401_),
    .C(_0416_),
    .Y(_0420_));
 sg13g2_o21ai_1 _3167_ (.B1(_0406_),
    .Y(_0421_),
    .A1(net581),
    .A2(_0420_));
 sg13g2_a21oi_1 _3168_ (.A1(net581),
    .A2(_0420_),
    .Y(_0050_),
    .B1(_0421_));
 sg13g2_nor2_1 _3169_ (.A(_2048_),
    .B(_0418_),
    .Y(_0422_));
 sg13g2_nand2_2 _3170_ (.Y(_0423_),
    .A(net584),
    .B(net582));
 sg13g2_xnor2_1 _3171_ (.Y(_0424_),
    .A(net579),
    .B(_0423_));
 sg13g2_a21oi_1 _3172_ (.A1(_0418_),
    .A2(_0424_),
    .Y(_0425_),
    .B1(_0422_));
 sg13g2_nor2_1 _3173_ (.A(_0407_),
    .B(_0425_),
    .Y(_0051_));
 sg13g2_nor2_2 _3174_ (.A(net884),
    .B(_0423_),
    .Y(_0426_));
 sg13g2_nand2_1 _3175_ (.Y(_0427_),
    .A(_0418_),
    .B(_0426_));
 sg13g2_xor2_1 _3176_ (.B(_0427_),
    .A(net577),
    .X(_0428_));
 sg13g2_nor2_1 _3177_ (.A(_0407_),
    .B(_0428_),
    .Y(_0052_));
 sg13g2_nand2_2 _3178_ (.Y(_0429_),
    .A(net608),
    .B(_2182_));
 sg13g2_nand2b_1 _3179_ (.Y(_0430_),
    .B(_2182_),
    .A_N(_2196_));
 sg13g2_nor2_2 _3180_ (.A(net524),
    .B(net528),
    .Y(_0431_));
 sg13g2_nand2_1 _3181_ (.Y(_0432_),
    .A(_2006_),
    .B(net520));
 sg13g2_nor2_1 _3182_ (.A(net529),
    .B(_2040_),
    .Y(_0433_));
 sg13g2_nor4_1 _3183_ (.A(net531),
    .B(_2040_),
    .C(net480),
    .D(_0432_),
    .Y(_0434_));
 sg13g2_a21o_1 _3184_ (.A2(net481),
    .A1(net657),
    .B1(_0434_),
    .X(_0053_));
 sg13g2_nor2b_1 _3185_ (.A(\gamepad_pmod.driver.pmod_clk_prev ),
    .B_N(\gamepad_pmod.driver.pmod_clk_sync[1] ),
    .Y(_0435_));
 sg13g2_nor2_1 _3186_ (.A(net598),
    .B(net517),
    .Y(_0436_));
 sg13g2_a22oi_1 _3187_ (.Y(_0054_),
    .B1(net512),
    .B2(_2005_),
    .A2(net518),
    .A1(_2039_));
 sg13g2_a22oi_1 _3188_ (.Y(_0055_),
    .B1(net511),
    .B2(_2004_),
    .A2(net518),
    .A1(_2005_));
 sg13g2_a22oi_1 _3189_ (.Y(_0056_),
    .B1(net512),
    .B2(_2003_),
    .A2(net518),
    .A1(_2004_));
 sg13g2_a22oi_1 _3190_ (.Y(_0057_),
    .B1(net511),
    .B2(_2002_),
    .A2(net517),
    .A1(_2003_));
 sg13g2_a22oi_1 _3191_ (.Y(_0058_),
    .B1(net512),
    .B2(_2001_),
    .A2(net518),
    .A1(_2002_));
 sg13g2_a22oi_1 _3192_ (.Y(_0059_),
    .B1(net512),
    .B2(_2000_),
    .A2(net518),
    .A1(_2001_));
 sg13g2_a22oi_1 _3193_ (.Y(_0060_),
    .B1(net511),
    .B2(_1999_),
    .A2(net517),
    .A1(_2000_));
 sg13g2_a22oi_1 _3194_ (.Y(_0061_),
    .B1(net511),
    .B2(_1998_),
    .A2(net517),
    .A1(_1999_));
 sg13g2_a22oi_1 _3195_ (.Y(_0062_),
    .B1(net511),
    .B2(_1997_),
    .A2(net517),
    .A1(_1998_));
 sg13g2_a22oi_1 _3196_ (.Y(_0063_),
    .B1(net511),
    .B2(_1996_),
    .A2(net517),
    .A1(_1997_));
 sg13g2_a22oi_1 _3197_ (.Y(_0064_),
    .B1(net511),
    .B2(_1995_),
    .A2(net517),
    .A1(_1996_));
 sg13g2_a22oi_1 _3198_ (.Y(_0065_),
    .B1(net511),
    .B2(_1994_),
    .A2(net517),
    .A1(_1995_));
 sg13g2_and2_1 _3199_ (.A(net623),
    .B(net3),
    .X(_0066_));
 sg13g2_and2_1 _3200_ (.A(net623),
    .B(net394),
    .X(_0067_));
 sg13g2_and2_1 _3201_ (.A(net622),
    .B(net2),
    .X(_0068_));
 sg13g2_and2_1 _3202_ (.A(net623),
    .B(net402),
    .X(_0069_));
 sg13g2_a21o_1 _3203_ (.A2(_2143_),
    .A1(\player_constroller_inst.game_over ),
    .B1(net597),
    .X(_0437_));
 sg13g2_o21ai_1 _3204_ (.B1(_2161_),
    .Y(_0438_),
    .A1(_2037_),
    .A2(_2148_));
 sg13g2_nor2b_1 _3205_ (.A(_2162_),
    .B_N(_0438_),
    .Y(_0439_));
 sg13g2_or3_2 _3206_ (.A(_2049_),
    .B(\player_constroller_inst.game_over ),
    .C(net499),
    .X(_0440_));
 sg13g2_nor2_2 _3207_ (.A(_2171_),
    .B(_0440_),
    .Y(_0441_));
 sg13g2_a22oi_1 _3208_ (.Y(_0442_),
    .B1(_0441_),
    .B2(_0439_),
    .A2(_0440_),
    .A1(net794));
 sg13g2_nor2_1 _3209_ (.A(net492),
    .B(_0442_),
    .Y(_0070_));
 sg13g2_xnor2_1 _3210_ (.Y(_0443_),
    .A(_2160_),
    .B(_2162_));
 sg13g2_a22oi_1 _3211_ (.Y(_0444_),
    .B1(_0441_),
    .B2(_0443_),
    .A2(_0440_),
    .A1(net860));
 sg13g2_nor2_1 _3212_ (.A(net493),
    .B(_0444_),
    .Y(_0071_));
 sg13g2_xor2_1 _3213_ (.B(_2163_),
    .A(_2155_),
    .X(_0445_));
 sg13g2_a22oi_1 _3214_ (.Y(_0446_),
    .B1(_0441_),
    .B2(_0445_),
    .A2(_0440_),
    .A1(net756));
 sg13g2_nor2_1 _3215_ (.A(net493),
    .B(_0446_),
    .Y(_0072_));
 sg13g2_xor2_1 _3216_ (.B(_2164_),
    .A(_2151_),
    .X(_0447_));
 sg13g2_a22oi_1 _3217_ (.Y(_0448_),
    .B1(_0441_),
    .B2(_0447_),
    .A2(_0440_),
    .A1(net826));
 sg13g2_nor2_1 _3218_ (.A(net492),
    .B(_0448_),
    .Y(_0073_));
 sg13g2_xor2_1 _3219_ (.B(_2167_),
    .A(_2165_),
    .X(_0449_));
 sg13g2_a22oi_1 _3220_ (.Y(_0450_),
    .B1(_0441_),
    .B2(_0449_),
    .A2(_0440_),
    .A1(net848));
 sg13g2_nor2_1 _3221_ (.A(net492),
    .B(_0450_),
    .Y(_0074_));
 sg13g2_a21oi_1 _3222_ (.A1(net575),
    .A2(_0440_),
    .Y(_0451_),
    .B1(_0441_));
 sg13g2_nor2_1 _3223_ (.A(net492),
    .B(_0451_),
    .Y(_0075_));
 sg13g2_a21oi_1 _3224_ (.A1(net548),
    .A2(_2171_),
    .Y(_0452_),
    .B1(net499));
 sg13g2_nor4_2 _3225_ (.A(net521),
    .B(net575),
    .C(net497),
    .Y(_0453_),
    .D(_2181_));
 sg13g2_nor3_2 _3226_ (.A(\player_constroller_inst.game_over ),
    .B(_0452_),
    .C(_0453_),
    .Y(_0454_));
 sg13g2_or3_1 _3227_ (.A(\player_constroller_inst.game_over ),
    .B(_0452_),
    .C(_0453_),
    .X(_0455_));
 sg13g2_o21ai_1 _3228_ (.B1(_2142_),
    .Y(_0456_),
    .A1(_2181_),
    .A2(_0439_));
 sg13g2_a21o_1 _3229_ (.A2(_0456_),
    .A1(_0454_),
    .B1(net492),
    .X(_0457_));
 sg13g2_a21oi_1 _3230_ (.A1(_2037_),
    .A2(_0455_),
    .Y(_0076_),
    .B1(_0457_));
 sg13g2_nand4_1 _3231_ (.B(_2182_),
    .C(_0443_),
    .A(_2142_),
    .Y(_0458_),
    .D(_0454_));
 sg13g2_nand2_1 _3232_ (.Y(_0459_),
    .A(net669),
    .B(_0455_));
 sg13g2_a21oi_1 _3233_ (.A1(_0458_),
    .A2(_0459_),
    .Y(_0077_),
    .B1(net492));
 sg13g2_nand4_1 _3234_ (.B(_2182_),
    .C(_0445_),
    .A(_2142_),
    .Y(_0460_),
    .D(_0454_));
 sg13g2_nand2_1 _3235_ (.Y(_0461_),
    .A(net652),
    .B(_0455_));
 sg13g2_a21oi_1 _3236_ (.A1(_0460_),
    .A2(_0461_),
    .Y(_0078_),
    .B1(net492));
 sg13g2_nor2_1 _3237_ (.A(net841),
    .B(_0454_),
    .Y(_0462_));
 sg13g2_o21ai_1 _3238_ (.B1(_2142_),
    .Y(_0463_),
    .A1(_2181_),
    .A2(_0447_));
 sg13g2_a21oi_1 _3239_ (.A1(_0454_),
    .A2(_0463_),
    .Y(_0464_),
    .B1(net492));
 sg13g2_nor2b_1 _3240_ (.A(net842),
    .B_N(_0464_),
    .Y(_0079_));
 sg13g2_nor2_2 _3241_ (.A(\player_constroller_inst.game_state[0] ),
    .B(\player_constroller_inst.game_over ),
    .Y(_0465_));
 sg13g2_a21oi_2 _3242_ (.B1(net493),
    .Y(_0466_),
    .A2(_2143_),
    .A1(\player_constroller_inst.game_state[0] ));
 sg13g2_o21ai_1 _3243_ (.B1(net607),
    .Y(_0467_),
    .A1(_2144_),
    .A2(_0465_));
 sg13g2_nor2_1 _3244_ (.A(\ai_controller_inst.obstacle1_pos[9] ),
    .B(\ai_controller_inst.obstacle1_pos[8] ),
    .Y(_0468_));
 sg13g2_nor3_2 _3245_ (.A(\ai_controller_inst.obstacle1_pos[7] ),
    .B(net908),
    .C(net792),
    .Y(_0469_));
 sg13g2_nor2_1 _3246_ (.A(\ai_controller_inst.obstacle1_pos[3] ),
    .B(\ai_controller_inst.obstacle1_pos[2] ),
    .Y(_0470_));
 sg13g2_nor3_2 _3247_ (.A(\ai_controller_inst.obstacle1_pos[4] ),
    .B(\ai_controller_inst.obstacle1_pos[3] ),
    .C(\ai_controller_inst.obstacle1_pos[2] ),
    .Y(_0471_));
 sg13g2_and3_1 _3248_ (.X(_0472_),
    .A(_0468_),
    .B(_0469_),
    .C(_0471_));
 sg13g2_nand2_1 _3249_ (.Y(_0473_),
    .A(\obstacles_inst.obstacle2_cross_gen_line_reg ),
    .B(_0472_));
 sg13g2_nand2_2 _3250_ (.Y(_0474_),
    .A(net501),
    .B(_0465_));
 sg13g2_nor2_2 _3251_ (.A(net498),
    .B(net495),
    .Y(_0475_));
 sg13g2_nand2_1 _3252_ (.Y(_0476_),
    .A(net865),
    .B(net822));
 sg13g2_nand3_1 _3253_ (.B(\ai_controller_inst.obstacle2_pos[3] ),
    .C(net913),
    .A(\ai_controller_inst.obstacle2_pos[4] ),
    .Y(_0477_));
 sg13g2_or3_1 _3254_ (.A(\ai_controller_inst.obstacle2_pos[7] ),
    .B(\ai_controller_inst.obstacle2_pos[6] ),
    .C(\ai_controller_inst.obstacle2_pos[5] ),
    .X(_0478_));
 sg13g2_nand2b_1 _3255_ (.Y(_0479_),
    .B(\ai_controller_inst.obstacle2_pos[8] ),
    .A_N(\ai_controller_inst.obstacle2_pos[9] ));
 sg13g2_nor4_1 _3256_ (.A(net495),
    .B(_0477_),
    .C(_0478_),
    .D(_0479_),
    .Y(_0480_));
 sg13g2_nor2_1 _3257_ (.A(net766),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_o21ai_1 _3258_ (.B1(_0466_),
    .Y(_0080_),
    .A1(_0475_),
    .A2(_0481_));
 sg13g2_nand2_1 _3259_ (.Y(_0482_),
    .A(net861),
    .B(\ai_controller_inst.obstacle1_pos[2] ));
 sg13g2_nand3_1 _3260_ (.B(\ai_controller_inst.obstacle1_pos[3] ),
    .C(\ai_controller_inst.obstacle1_pos[2] ),
    .A(\ai_controller_inst.obstacle1_pos[4] ),
    .Y(_0483_));
 sg13g2_nand2_1 _3261_ (.Y(_0484_),
    .A(\ai_controller_inst.obstacle1_pos[8] ),
    .B(_0469_));
 sg13g2_nor4_1 _3262_ (.A(\ai_controller_inst.obstacle1_pos[9] ),
    .B(net496),
    .C(_0483_),
    .D(_0484_),
    .Y(_0485_));
 sg13g2_nor2_1 _3263_ (.A(net711),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_nor2_1 _3264_ (.A(\ai_controller_inst.obstacle2_pos[3] ),
    .B(\ai_controller_inst.obstacle2_pos[2] ),
    .Y(_0487_));
 sg13g2_nor3_1 _3265_ (.A(\ai_controller_inst.obstacle2_pos[4] ),
    .B(\ai_controller_inst.obstacle2_pos[3] ),
    .C(net918),
    .Y(_0488_));
 sg13g2_inv_1 _3266_ (.Y(_0489_),
    .A(_0488_));
 sg13g2_nor2_1 _3267_ (.A(\ai_controller_inst.obstacle2_pos[9] ),
    .B(\ai_controller_inst.obstacle2_pos[8] ),
    .Y(_0490_));
 sg13g2_nor4_2 _3268_ (.A(\ai_controller_inst.obstacle2_pos[9] ),
    .B(\ai_controller_inst.obstacle2_pos[8] ),
    .C(_0478_),
    .Y(_0491_),
    .D(_0489_));
 sg13g2_nand2_1 _3269_ (.Y(_0492_),
    .A(net711),
    .B(_0491_));
 sg13g2_nor2_2 _3270_ (.A(net495),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_nor3_1 _3271_ (.A(net489),
    .B(net712),
    .C(_0493_),
    .Y(_0081_));
 sg13g2_o21ai_1 _3272_ (.B1(net453),
    .Y(_0494_),
    .A1(net495),
    .A2(net494));
 sg13g2_nand2_1 _3273_ (.Y(_0495_),
    .A(\lfsr_inst.r_lfsr[6] ),
    .B(_0493_));
 sg13g2_a21oi_1 _3274_ (.A1(_0494_),
    .A2(_0495_),
    .Y(_0082_),
    .B1(net489));
 sg13g2_o21ai_1 _3275_ (.B1(net789),
    .Y(_0496_),
    .A1(net495),
    .A2(net494));
 sg13g2_nand2_1 _3276_ (.Y(_0497_),
    .A(net736),
    .B(_0493_));
 sg13g2_a21oi_1 _3277_ (.A1(_0496_),
    .A2(_0497_),
    .Y(_0083_),
    .B1(net491));
 sg13g2_o21ai_1 _3278_ (.B1(net720),
    .Y(_0498_),
    .A1(net495),
    .A2(net494));
 sg13g2_nand2_1 _3279_ (.Y(_0499_),
    .A(\lfsr_inst.r_lfsr[8] ),
    .B(_0493_));
 sg13g2_a21oi_1 _3280_ (.A1(_0498_),
    .A2(_0499_),
    .Y(_0084_),
    .B1(net491));
 sg13g2_o21ai_1 _3281_ (.B1(\obs_rom_inst_1.i_obs_type[0] ),
    .Y(_0500_),
    .A1(_0473_),
    .A2(net496));
 sg13g2_nand2_1 _3282_ (.Y(_0501_),
    .A(net713),
    .B(_0475_));
 sg13g2_a21oi_1 _3283_ (.A1(_0500_),
    .A2(_0501_),
    .Y(_0085_),
    .B1(net491));
 sg13g2_o21ai_1 _3284_ (.B1(net572),
    .Y(_0502_),
    .A1(net498),
    .A2(net496));
 sg13g2_nand2_1 _3285_ (.Y(_0503_),
    .A(net736),
    .B(_0475_));
 sg13g2_a21oi_1 _3286_ (.A1(_0502_),
    .A2(_0503_),
    .Y(_0086_),
    .B1(net490));
 sg13g2_o21ai_1 _3287_ (.B1(\obs_rom_inst_1.i_obs_type[2] ),
    .Y(_0504_),
    .A1(net498),
    .A2(net495));
 sg13g2_nand2_1 _3288_ (.Y(_0505_),
    .A(net747),
    .B(_0475_));
 sg13g2_a21oi_1 _3289_ (.A1(_0504_),
    .A2(_0505_),
    .Y(_0087_),
    .B1(net490));
 sg13g2_a21oi_2 _3290_ (.B1(net495),
    .Y(_0506_),
    .A2(_0491_),
    .A1(_2035_));
 sg13g2_nand2b_1 _3291_ (.Y(_0507_),
    .B(net822),
    .A_N(_0506_));
 sg13g2_mux2_1 _3292_ (.A0(net423),
    .A1(_0017_),
    .S(net494),
    .X(_0508_));
 sg13g2_nand2_1 _3293_ (.Y(_0509_),
    .A(_0506_),
    .B(_0508_));
 sg13g2_a21oi_1 _3294_ (.A1(_0507_),
    .A2(_0509_),
    .Y(_0088_),
    .B1(net491));
 sg13g2_nand2_1 _3295_ (.Y(_0510_),
    .A(_0487_),
    .B(_0506_));
 sg13g2_nand2_1 _3296_ (.Y(_0511_),
    .A(_0476_),
    .B(_0510_));
 sg13g2_o21ai_1 _3297_ (.B1(_0511_),
    .Y(_0512_),
    .A1(net857),
    .A2(net494));
 sg13g2_nand2b_1 _3298_ (.Y(_0513_),
    .B(net865),
    .A_N(_0506_));
 sg13g2_a21oi_1 _3299_ (.A1(_0512_),
    .A2(_0513_),
    .Y(_0089_),
    .B1(net489));
 sg13g2_nor2_1 _3300_ (.A(net760),
    .B(net494),
    .Y(_0514_));
 sg13g2_nand2_1 _3301_ (.Y(_0515_),
    .A(_0488_),
    .B(_0506_));
 sg13g2_nor2_1 _3302_ (.A(_0514_),
    .B(_0515_),
    .Y(_0516_));
 sg13g2_a21oi_1 _3303_ (.A1(net827),
    .A2(_0510_),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_nor2_1 _3304_ (.A(net489),
    .B(_0517_),
    .Y(_0090_));
 sg13g2_nand2_1 _3305_ (.Y(_0518_),
    .A(\ai_controller_inst.obstacle2_pos[5] ),
    .B(_0489_));
 sg13g2_o21ai_1 _3306_ (.B1(_0518_),
    .Y(_0519_),
    .A1(\ai_controller_inst.obstacle2_pos[5] ),
    .A2(_0515_));
 sg13g2_o21ai_1 _3307_ (.B1(_0519_),
    .Y(_0520_),
    .A1(net813),
    .A2(net494));
 sg13g2_nand2b_1 _3308_ (.Y(_0521_),
    .B(net876),
    .A_N(_0506_));
 sg13g2_a21oi_1 _3309_ (.A1(_0520_),
    .A2(_0521_),
    .Y(_0091_),
    .B1(net489));
 sg13g2_o21ai_1 _3310_ (.B1(net834),
    .Y(_0522_),
    .A1(\ai_controller_inst.obstacle2_pos[5] ),
    .A2(_0515_));
 sg13g2_or4_2 _3311_ (.A(\ai_controller_inst.obstacle2_pos[6] ),
    .B(\ai_controller_inst.obstacle2_pos[5] ),
    .C(\ai_controller_inst.obstacle2_pos[4] ),
    .D(_0510_),
    .X(_0523_));
 sg13g2_inv_1 _3312_ (.Y(_0524_),
    .A(_0523_));
 sg13g2_o21ai_1 _3313_ (.B1(_0524_),
    .Y(_0525_),
    .A1(net784),
    .A2(net494));
 sg13g2_a21oi_1 _3314_ (.A1(net835),
    .A2(_0525_),
    .Y(_0092_),
    .B1(net489));
 sg13g2_nor2_1 _3315_ (.A(\ai_controller_inst.obstacle2_pos[7] ),
    .B(_0523_),
    .Y(_0526_));
 sg13g2_xor2_1 _3316_ (.B(_0523_),
    .A(net889),
    .X(_0527_));
 sg13g2_nor2_1 _3317_ (.A(net489),
    .B(_0527_),
    .Y(_0093_));
 sg13g2_nor3_1 _3318_ (.A(\ai_controller_inst.obstacle2_pos[8] ),
    .B(net906),
    .C(_0523_),
    .Y(_0528_));
 sg13g2_xnor2_1 _3319_ (.Y(_0529_),
    .A(net887),
    .B(_0526_));
 sg13g2_nor3_1 _3320_ (.A(net489),
    .B(_0493_),
    .C(net888),
    .Y(_0094_));
 sg13g2_o21ai_1 _3321_ (.B1(_0466_),
    .Y(_0530_),
    .A1(net803),
    .A2(net907));
 sg13g2_a21oi_1 _3322_ (.A1(net803),
    .A2(net907),
    .Y(_0095_),
    .B1(_0530_));
 sg13g2_a21oi_2 _3323_ (.B1(net496),
    .Y(_0531_),
    .A2(_0472_),
    .A1(_2036_));
 sg13g2_nand2b_1 _3324_ (.Y(_0532_),
    .B(\ai_controller_inst.obstacle1_pos[2] ),
    .A_N(_0531_));
 sg13g2_mux2_1 _3325_ (.A0(net423),
    .A1(net849),
    .S(net498),
    .X(_0533_));
 sg13g2_nand2_1 _3326_ (.Y(_0534_),
    .A(_0531_),
    .B(_0533_));
 sg13g2_a21oi_1 _3327_ (.A1(_0532_),
    .A2(_0534_),
    .Y(_0096_),
    .B1(net490));
 sg13g2_nand2_1 _3328_ (.Y(_0535_),
    .A(_0470_),
    .B(_0531_));
 sg13g2_nand2_1 _3329_ (.Y(_0536_),
    .A(_0482_),
    .B(_0535_));
 sg13g2_o21ai_1 _3330_ (.B1(_0536_),
    .Y(_0537_),
    .A1(net857),
    .A2(net498));
 sg13g2_nand2b_1 _3331_ (.Y(_0538_),
    .B(net861),
    .A_N(_0531_));
 sg13g2_a21oi_1 _3332_ (.A1(_0537_),
    .A2(_0538_),
    .Y(_0097_),
    .B1(net490));
 sg13g2_nand2_1 _3333_ (.Y(_0539_),
    .A(net815),
    .B(_0535_));
 sg13g2_nor2_1 _3334_ (.A(net815),
    .B(_0535_),
    .Y(_0540_));
 sg13g2_o21ai_1 _3335_ (.B1(_0540_),
    .Y(_0541_),
    .A1(net760),
    .A2(net498));
 sg13g2_a21oi_1 _3336_ (.A1(_0539_),
    .A2(_0541_),
    .Y(_0098_),
    .B1(net491));
 sg13g2_nand3_1 _3337_ (.B(_0471_),
    .C(_0531_),
    .A(_2031_),
    .Y(_0542_));
 sg13g2_o21ai_1 _3338_ (.B1(_0542_),
    .Y(_0543_),
    .A1(_2031_),
    .A2(_0471_));
 sg13g2_o21ai_1 _3339_ (.B1(_0543_),
    .Y(_0544_),
    .A1(\lfsr_inst.r_lfsr[4] ),
    .A2(net498));
 sg13g2_nand2b_1 _3340_ (.Y(_0545_),
    .B(net792),
    .A_N(_0531_));
 sg13g2_a21oi_1 _3341_ (.A1(_0544_),
    .A2(_0545_),
    .Y(_0099_),
    .B1(net490));
 sg13g2_nor2_1 _3342_ (.A(net784),
    .B(net498),
    .Y(_0546_));
 sg13g2_nor3_1 _3343_ (.A(net871),
    .B(_0542_),
    .C(_0546_),
    .Y(_0547_));
 sg13g2_a21oi_1 _3344_ (.A1(net871),
    .A2(_0542_),
    .Y(_0548_),
    .B1(_0547_));
 sg13g2_nor2_1 _3345_ (.A(net490),
    .B(_0548_),
    .Y(_0100_));
 sg13g2_o21ai_1 _3346_ (.B1(net820),
    .Y(_0549_),
    .A1(\ai_controller_inst.obstacle1_pos[6] ),
    .A2(_0542_));
 sg13g2_nand2_1 _3347_ (.Y(_0550_),
    .A(_0469_),
    .B(_0540_));
 sg13g2_a21oi_1 _3348_ (.A1(net821),
    .A2(_0550_),
    .Y(_0101_),
    .B1(net490));
 sg13g2_nor2_1 _3349_ (.A(\ai_controller_inst.obstacle1_pos[8] ),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_xor2_1 _3350_ (.B(_0550_),
    .A(net885),
    .X(_0552_));
 sg13g2_nor3_1 _3351_ (.A(net490),
    .B(_0475_),
    .C(_0552_),
    .Y(_0102_));
 sg13g2_o21ai_1 _3352_ (.B1(_0466_),
    .Y(_0553_),
    .A1(net726),
    .A2(_0551_));
 sg13g2_a21oi_1 _3353_ (.A1(net726),
    .A2(_0551_),
    .Y(_0103_),
    .B1(_0553_));
 sg13g2_nor3_1 _3354_ (.A(\bg_object_inst.bg_object_pos[4] ),
    .B(\bg_object_inst.bg_object_pos[3] ),
    .C(\bg_object_inst.bg_object_pos[2] ),
    .Y(_0554_));
 sg13g2_nor4_1 _3355_ (.A(\bg_object_inst.bg_object_pos[9] ),
    .B(\bg_object_inst.bg_object_pos[8] ),
    .C(\bg_object_inst.bg_object_pos[7] ),
    .D(\bg_object_inst.bg_object_pos[5] ),
    .Y(_0555_));
 sg13g2_nand3b_1 _3356_ (.B(_0554_),
    .C(_0555_),
    .Y(_0556_),
    .A_N(\bg_object_inst.bg_object_pos[6] ));
 sg13g2_mux2_1 _3357_ (.A0(net760),
    .A1(_0018_),
    .S(_0556_),
    .X(_0557_));
 sg13g2_o21ai_1 _3358_ (.B1(net622),
    .Y(_0558_),
    .A1(_2137_),
    .A2(_0557_));
 sg13g2_a21oi_1 _3359_ (.A1(_2029_),
    .A2(net497),
    .Y(_0104_),
    .B1(_0558_));
 sg13g2_a21oi_1 _3360_ (.A1(_2029_),
    .A2(net500),
    .Y(_0559_),
    .B1(_2028_));
 sg13g2_nor3_2 _3361_ (.A(net869),
    .B(net824),
    .C(_2137_),
    .Y(_0560_));
 sg13g2_nor2_1 _3362_ (.A(_0559_),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_nor3_1 _3363_ (.A(net813),
    .B(net497),
    .C(_0556_),
    .Y(_0562_));
 sg13g2_nor3_1 _3364_ (.A(net604),
    .B(_0561_),
    .C(_0562_),
    .Y(_0105_));
 sg13g2_nand2b_1 _3365_ (.Y(_0563_),
    .B(net761),
    .A_N(_0560_));
 sg13g2_nor2b_1 _3366_ (.A(net761),
    .B_N(_0560_),
    .Y(_0564_));
 sg13g2_o21ai_1 _3367_ (.B1(_0564_),
    .Y(_0565_),
    .A1(\lfsr_inst.r_lfsr[5] ),
    .A2(_0556_));
 sg13g2_nand2_1 _3368_ (.Y(_0566_),
    .A(net500),
    .B(_0554_));
 sg13g2_a21oi_1 _3369_ (.A1(_0563_),
    .A2(_0565_),
    .Y(_0106_),
    .B1(net604));
 sg13g2_nor2_1 _3370_ (.A(net713),
    .B(_0556_),
    .Y(_0567_));
 sg13g2_nand2b_1 _3371_ (.Y(_0568_),
    .B(_0564_),
    .A_N(\bg_object_inst.bg_object_pos[5] ));
 sg13g2_nor2_1 _3372_ (.A(_0567_),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_a21oi_1 _3373_ (.A1(net828),
    .A2(_0566_),
    .Y(_0570_),
    .B1(_0569_));
 sg13g2_nor2_1 _3374_ (.A(net603),
    .B(net829),
    .Y(_0107_));
 sg13g2_nor4_1 _3375_ (.A(\bg_object_inst.bg_object_pos[9] ),
    .B(\bg_object_inst.bg_object_pos[8] ),
    .C(\bg_object_inst.bg_object_pos[7] ),
    .D(\lfsr_inst.r_lfsr[7] ),
    .Y(_0571_));
 sg13g2_nor3_1 _3376_ (.A(net836),
    .B(_0568_),
    .C(_0571_),
    .Y(_0572_));
 sg13g2_a21oi_1 _3377_ (.A1(net836),
    .A2(_0568_),
    .Y(_0573_),
    .B1(_0572_));
 sg13g2_nor2_1 _3378_ (.A(net604),
    .B(net837),
    .Y(_0108_));
 sg13g2_o21ai_1 _3379_ (.B1(net853),
    .Y(_0574_),
    .A1(net836),
    .A2(_0568_));
 sg13g2_or4_2 _3380_ (.A(net853),
    .B(\bg_object_inst.bg_object_pos[6] ),
    .C(net828),
    .D(_0566_),
    .X(_0575_));
 sg13g2_a21oi_1 _3381_ (.A1(_0574_),
    .A2(_0575_),
    .Y(_0109_),
    .B1(net604));
 sg13g2_nor2_1 _3382_ (.A(\bg_object_inst.bg_object_pos[8] ),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_xor2_1 _3383_ (.B(_0575_),
    .A(net879),
    .X(_0577_));
 sg13g2_nor2_1 _3384_ (.A(net603),
    .B(_0577_),
    .Y(_0110_));
 sg13g2_o21ai_1 _3385_ (.B1(net624),
    .Y(_0578_),
    .A1(net737),
    .A2(_0576_));
 sg13g2_a21oi_1 _3386_ (.A1(net737),
    .A2(_0576_),
    .Y(_0111_),
    .B1(_0578_));
 sg13g2_nor2_1 _3387_ (.A(net587),
    .B(_0398_),
    .Y(_0579_));
 sg13g2_xor2_1 _3388_ (.B(_0398_),
    .A(net587),
    .X(_0580_));
 sg13g2_nor2_1 _3389_ (.A(net599),
    .B(_0580_),
    .Y(_0112_));
 sg13g2_a21oi_1 _3390_ (.A1(net587),
    .A2(_0398_),
    .Y(_0581_),
    .B1(net585));
 sg13g2_and3_1 _3391_ (.X(_0582_),
    .A(net585),
    .B(net587),
    .C(_0398_));
 sg13g2_nor3_1 _3392_ (.A(net599),
    .B(_0581_),
    .C(_0582_),
    .Y(_0113_));
 sg13g2_nand2b_1 _3393_ (.Y(_0583_),
    .B(_0398_),
    .A_N(net588));
 sg13g2_nand2_1 _3394_ (.Y(_0584_),
    .A(_0398_),
    .B(_0403_));
 sg13g2_o21ai_1 _3395_ (.B1(net581),
    .Y(_0585_),
    .A1(net585),
    .A2(_0583_));
 sg13g2_a21oi_1 _3396_ (.A1(_0584_),
    .A2(_0585_),
    .Y(_0114_),
    .B1(net599));
 sg13g2_nor2_1 _3397_ (.A(net578),
    .B(_0584_),
    .Y(_0586_));
 sg13g2_xnor2_1 _3398_ (.Y(_0587_),
    .A(_2048_),
    .B(_0584_));
 sg13g2_nor2_1 _3399_ (.A(net599),
    .B(_0587_),
    .Y(_0115_));
 sg13g2_nor2b_1 _3400_ (.A(net578),
    .B_N(net577),
    .Y(_0588_));
 sg13g2_o21ai_1 _3401_ (.B1(net607),
    .Y(_0589_),
    .A1(net577),
    .A2(_0586_));
 sg13g2_a21oi_1 _3402_ (.A1(net577),
    .A2(_0586_),
    .Y(_0116_),
    .B1(_0589_));
 sg13g2_nor2_2 _3403_ (.A(net530),
    .B(net532),
    .Y(_0590_));
 sg13g2_or2_2 _3404_ (.X(_0591_),
    .B(net533),
    .A(net531));
 sg13g2_nand2_2 _3405_ (.Y(_0592_),
    .A(net530),
    .B(net533));
 sg13g2_nand3_1 _3406_ (.B(_0591_),
    .C(_0592_),
    .A(_0431_),
    .Y(_0593_));
 sg13g2_nand2_1 _3407_ (.Y(_0594_),
    .A(net438),
    .B(net480));
 sg13g2_o21ai_1 _3408_ (.B1(_0594_),
    .Y(_0117_),
    .A1(net480),
    .A2(_0593_));
 sg13g2_nand2b_1 _3409_ (.Y(_0595_),
    .B(net822),
    .A_N(\bg_render_inst.i_hpos[2] ));
 sg13g2_nand2b_1 _3410_ (.Y(_0596_),
    .B(net595),
    .A_N(net822));
 sg13g2_a21oi_1 _3411_ (.A1(_0595_),
    .A2(_0596_),
    .Y(_0118_),
    .B1(net602));
 sg13g2_nor2b_1 _3412_ (.A(\ai_controller_inst.obstacle2_pos[3] ),
    .B_N(net593),
    .Y(_0597_));
 sg13g2_nand2b_1 _3413_ (.Y(_0598_),
    .B(net593),
    .A_N(\ai_controller_inst.obstacle2_pos[3] ));
 sg13g2_nand2b_1 _3414_ (.Y(_0599_),
    .B(\ai_controller_inst.obstacle2_pos[3] ),
    .A_N(net593));
 sg13g2_and2_1 _3415_ (.A(_0598_),
    .B(_0599_),
    .X(_0600_));
 sg13g2_nor2_1 _3416_ (.A(_0595_),
    .B(_0600_),
    .Y(_0601_));
 sg13g2_nand2_1 _3417_ (.Y(_0602_),
    .A(_0595_),
    .B(_0600_));
 sg13g2_nand2_1 _3418_ (.Y(_0603_),
    .A(net621),
    .B(_0602_));
 sg13g2_nor2_1 _3419_ (.A(_0601_),
    .B(_0603_),
    .Y(_0119_));
 sg13g2_nor2_1 _3420_ (.A(\ai_controller_inst.obstacle2_pos[4] ),
    .B(_2046_),
    .Y(_0604_));
 sg13g2_xnor2_1 _3421_ (.Y(_0605_),
    .A(\ai_controller_inst.obstacle2_pos[4] ),
    .B(net591));
 sg13g2_nand2_1 _3422_ (.Y(_0606_),
    .A(_0597_),
    .B(_0605_));
 sg13g2_xnor2_1 _3423_ (.Y(_0607_),
    .A(_0597_),
    .B(_0605_));
 sg13g2_nand4_1 _3424_ (.B(_0598_),
    .C(_0599_),
    .A(_0595_),
    .Y(_0608_),
    .D(_0605_));
 sg13g2_nand2_1 _3425_ (.Y(_0609_),
    .A(net621),
    .B(_0608_));
 sg13g2_a21oi_1 _3426_ (.A1(_0602_),
    .A2(_0607_),
    .Y(_0120_),
    .B1(_0609_));
 sg13g2_nand2b_1 _3427_ (.Y(_0610_),
    .B(net589),
    .A_N(\ai_controller_inst.obstacle2_pos[5] ));
 sg13g2_xnor2_1 _3428_ (.Y(_0611_),
    .A(\ai_controller_inst.obstacle2_pos[5] ),
    .B(net589));
 sg13g2_and2_1 _3429_ (.A(_0604_),
    .B(_0611_),
    .X(_0612_));
 sg13g2_xnor2_1 _3430_ (.Y(_0613_),
    .A(_0604_),
    .B(_0611_));
 sg13g2_and3_1 _3431_ (.X(_0614_),
    .A(_0606_),
    .B(_0608_),
    .C(_0613_));
 sg13g2_a21oi_1 _3432_ (.A1(_0606_),
    .A2(_0608_),
    .Y(_0615_),
    .B1(_0613_));
 sg13g2_nor3_1 _3433_ (.A(net602),
    .B(_0614_),
    .C(_0615_),
    .Y(_0121_));
 sg13g2_nand2b_1 _3434_ (.Y(_0616_),
    .B(\ai_controller_inst.obstacle2_pos[6] ),
    .A_N(net586));
 sg13g2_xnor2_1 _3435_ (.Y(_0617_),
    .A(\ai_controller_inst.obstacle2_pos[6] ),
    .B(net586));
 sg13g2_nor2_1 _3436_ (.A(_0610_),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_xor2_1 _3437_ (.B(_0617_),
    .A(_0610_),
    .X(_0619_));
 sg13g2_nor3_1 _3438_ (.A(_0612_),
    .B(_0615_),
    .C(_0619_),
    .Y(_0620_));
 sg13g2_o21ai_1 _3439_ (.B1(_0619_),
    .Y(_0621_),
    .A1(_0612_),
    .A2(_0615_));
 sg13g2_nand2_1 _3440_ (.Y(_0622_),
    .A(net621),
    .B(_0621_));
 sg13g2_nor2_1 _3441_ (.A(_0620_),
    .B(_0622_),
    .Y(_0122_));
 sg13g2_nor2b_1 _3442_ (.A(_0618_),
    .B_N(_0621_),
    .Y(_0623_));
 sg13g2_nor2_1 _3443_ (.A(\ai_controller_inst.obstacle2_pos[7] ),
    .B(_2047_),
    .Y(_0624_));
 sg13g2_xnor2_1 _3444_ (.Y(_0625_),
    .A(\ai_controller_inst.obstacle2_pos[7] ),
    .B(net583));
 sg13g2_nand2_1 _3445_ (.Y(_0626_),
    .A(_0616_),
    .B(_0625_));
 sg13g2_xnor2_1 _3446_ (.Y(_0627_),
    .A(_0616_),
    .B(_0625_));
 sg13g2_or2_1 _3447_ (.X(_0628_),
    .B(_0627_),
    .A(_0623_));
 sg13g2_nand2_1 _3448_ (.Y(_0629_),
    .A(net621),
    .B(_0628_));
 sg13g2_a21oi_1 _3449_ (.A1(_0623_),
    .A2(_0627_),
    .Y(_0123_),
    .B1(_0629_));
 sg13g2_and2_1 _3450_ (.A(_0626_),
    .B(_0628_),
    .X(_0630_));
 sg13g2_nand2b_1 _3451_ (.Y(_0631_),
    .B(net580),
    .A_N(\ai_controller_inst.obstacle2_pos[8] ));
 sg13g2_xnor2_1 _3452_ (.Y(_0632_),
    .A(\ai_controller_inst.obstacle2_pos[8] ),
    .B(net580));
 sg13g2_nand2_1 _3453_ (.Y(_0633_),
    .A(_0624_),
    .B(_0632_));
 sg13g2_xnor2_1 _3454_ (.Y(_0634_),
    .A(_0624_),
    .B(_0632_));
 sg13g2_or2_1 _3455_ (.X(_0635_),
    .B(_0634_),
    .A(_0630_));
 sg13g2_nand2_1 _3456_ (.Y(_0636_),
    .A(net623),
    .B(_0635_));
 sg13g2_a21oi_1 _3457_ (.A1(_0630_),
    .A2(_0634_),
    .Y(_0124_),
    .B1(_0636_));
 sg13g2_xor2_1 _3458_ (.B(\bg_render_inst.i_hpos[9] ),
    .A(\ai_controller_inst.obstacle2_pos[9] ),
    .X(_0637_));
 sg13g2_xnor2_1 _3459_ (.Y(_0638_),
    .A(_0631_),
    .B(_0637_));
 sg13g2_a21oi_1 _3460_ (.A1(_0633_),
    .A2(_0635_),
    .Y(_0639_),
    .B1(_0638_));
 sg13g2_and3_1 _3461_ (.X(_0640_),
    .A(_0633_),
    .B(_0635_),
    .C(_0638_));
 sg13g2_nor3_1 _3462_ (.A(net602),
    .B(_0639_),
    .C(_0640_),
    .Y(_0125_));
 sg13g2_nand2_2 _3463_ (.Y(_0641_),
    .A(_2050_),
    .B(\audio_inst.i_jump.state[1] ));
 sg13g2_o21ai_1 _3464_ (.B1(net608),
    .Y(_0642_),
    .A1(_2181_),
    .A2(_0641_));
 sg13g2_inv_1 _3465_ (.Y(_0643_),
    .A(net476));
 sg13g2_o21ai_1 _3466_ (.B1(\audio_inst.i_jump.counter[2] ),
    .Y(_0644_),
    .A1(\audio_inst.i_jump.counter[1] ),
    .A2(\audio_inst.i_jump.counter[0] ));
 sg13g2_a21o_1 _3467_ (.A2(_0644_),
    .A1(_2064_),
    .B1(_2067_),
    .X(_0645_));
 sg13g2_nor4_1 _3468_ (.A(\audio_inst.i_jump.counter[7] ),
    .B(\audio_inst.i_jump.counter[6] ),
    .C(\audio_inst.i_jump.counter[5] ),
    .D(\audio_inst.i_jump.counter[8] ),
    .Y(_0646_));
 sg13g2_nand2_1 _3469_ (.Y(_0647_),
    .A(\audio_inst.i_jump.counter[10] ),
    .B(\audio_inst.i_jump.counter[9] ));
 sg13g2_a21oi_1 _3470_ (.A1(_0645_),
    .A2(_0646_),
    .Y(_0648_),
    .B1(_0647_));
 sg13g2_o21ai_1 _3471_ (.B1(\audio_inst.i_jump.counter[12] ),
    .Y(_0649_),
    .A1(\audio_inst.i_jump.counter[11] ),
    .A2(_0648_));
 sg13g2_nor3_1 _3472_ (.A(\audio_inst.i_jump.counter[15] ),
    .B(\audio_inst.i_jump.counter[14] ),
    .C(\audio_inst.i_jump.counter[13] ),
    .Y(_0650_));
 sg13g2_a21oi_1 _3473_ (.A1(_0649_),
    .A2(_0650_),
    .Y(_0651_),
    .B1(_2069_));
 sg13g2_o21ai_1 _3474_ (.B1(\audio_inst.i_jump.counter[18] ),
    .Y(_0652_),
    .A1(\audio_inst.i_jump.counter[17] ),
    .A2(_0651_));
 sg13g2_nand2_2 _3475_ (.Y(_0653_),
    .A(_2195_),
    .B(_0652_));
 sg13g2_nor2_1 _3476_ (.A(_2181_),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_nor3_2 _3477_ (.A(_2181_),
    .B(net476),
    .C(_0653_),
    .Y(_0655_));
 sg13g2_nand4_1 _3478_ (.B(_2195_),
    .C(_0643_),
    .A(_2182_),
    .Y(_0656_),
    .D(_0652_));
 sg13g2_a22oi_1 _3479_ (.Y(_0657_),
    .B1(_0655_),
    .B2(net389),
    .A2(net474),
    .A1(\audio_inst.i_jump.counter[0] ));
 sg13g2_inv_1 _3480_ (.Y(_0126_),
    .A(net390));
 sg13g2_nand2_1 _3481_ (.Y(_0658_),
    .A(net831),
    .B(net474));
 sg13g2_xnor2_1 _3482_ (.Y(_0659_),
    .A(net831),
    .B(\audio_inst.i_jump.counter[0] ));
 sg13g2_o21ai_1 _3483_ (.B1(_0658_),
    .Y(_0127_),
    .A1(net469),
    .A2(_0659_));
 sg13g2_nand2_1 _3484_ (.Y(_0660_),
    .A(net780),
    .B(net474));
 sg13g2_nand3_1 _3485_ (.B(\audio_inst.i_jump.counter[0] ),
    .C(net904),
    .A(net903),
    .Y(_0661_));
 sg13g2_a21o_1 _3486_ (.A2(\audio_inst.i_jump.counter[0] ),
    .A1(net903),
    .B1(net780),
    .X(_0662_));
 sg13g2_nand2_1 _3487_ (.Y(_0663_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_o21ai_1 _3488_ (.B1(_0660_),
    .Y(_0128_),
    .A1(net469),
    .A2(_0663_));
 sg13g2_nand2_1 _3489_ (.Y(_0664_),
    .A(net465),
    .B(net474));
 sg13g2_and4_2 _3490_ (.A(\audio_inst.i_jump.counter[1] ),
    .B(\audio_inst.i_jump.counter[0] ),
    .C(\audio_inst.i_jump.counter[2] ),
    .D(\audio_inst.i_jump.counter[3] ),
    .X(_0665_));
 sg13g2_xnor2_1 _3491_ (.Y(_0666_),
    .A(_2064_),
    .B(net905));
 sg13g2_o21ai_1 _3492_ (.B1(_0664_),
    .Y(_0129_),
    .A1(net469),
    .A2(_0666_));
 sg13g2_nand2_1 _3493_ (.Y(_0667_),
    .A(net805),
    .B(net474));
 sg13g2_xnor2_1 _3494_ (.Y(_0668_),
    .A(net805),
    .B(_0665_));
 sg13g2_o21ai_1 _3495_ (.B1(_0667_),
    .Y(_0130_),
    .A1(net469),
    .A2(_0668_));
 sg13g2_nand2_1 _3496_ (.Y(_0669_),
    .A(net787),
    .B(net474));
 sg13g2_nand3_1 _3497_ (.B(\audio_inst.i_jump.counter[4] ),
    .C(_0665_),
    .A(\audio_inst.i_jump.counter[5] ),
    .Y(_0670_));
 sg13g2_a21o_1 _3498_ (.A2(_0665_),
    .A1(\audio_inst.i_jump.counter[4] ),
    .B1(net787),
    .X(_0671_));
 sg13g2_nand2_1 _3499_ (.Y(_0672_),
    .A(_0670_),
    .B(_0671_));
 sg13g2_o21ai_1 _3500_ (.B1(_0669_),
    .Y(_0131_),
    .A1(net469),
    .A2(_0672_));
 sg13g2_nand2_1 _3501_ (.Y(_0673_),
    .A(net685),
    .B(net474));
 sg13g2_nand4_1 _3502_ (.B(\audio_inst.i_jump.counter[5] ),
    .C(\audio_inst.i_jump.counter[4] ),
    .A(\audio_inst.i_jump.counter[6] ),
    .Y(_0674_),
    .D(_0665_));
 sg13g2_xnor2_1 _3503_ (.Y(_0675_),
    .A(_2066_),
    .B(_0670_));
 sg13g2_o21ai_1 _3504_ (.B1(_0673_),
    .Y(_0132_),
    .A1(net469),
    .A2(_0675_));
 sg13g2_nand2_1 _3505_ (.Y(_0676_),
    .A(net634),
    .B(net474));
 sg13g2_nor2_1 _3506_ (.A(_2065_),
    .B(_0674_),
    .Y(_0677_));
 sg13g2_xnor2_1 _3507_ (.Y(_0678_),
    .A(_2065_),
    .B(_0674_));
 sg13g2_o21ai_1 _3508_ (.B1(_0676_),
    .Y(_0133_),
    .A1(net469),
    .A2(_0678_));
 sg13g2_nand2_1 _3509_ (.Y(_0679_),
    .A(net812),
    .B(net475));
 sg13g2_xnor2_1 _3510_ (.Y(_0680_),
    .A(net812),
    .B(_0677_));
 sg13g2_o21ai_1 _3511_ (.B1(_0679_),
    .Y(_0134_),
    .A1(net469),
    .A2(_0680_));
 sg13g2_and3_1 _3512_ (.X(_0681_),
    .A(net769),
    .B(\audio_inst.i_jump.counter[8] ),
    .C(_0677_));
 sg13g2_a21oi_1 _3513_ (.A1(\audio_inst.i_jump.counter[8] ),
    .A2(_0677_),
    .Y(_0682_),
    .B1(net769));
 sg13g2_nor3_1 _3514_ (.A(net470),
    .B(_0681_),
    .C(_0682_),
    .Y(_0683_));
 sg13g2_a21o_1 _3515_ (.A2(net475),
    .A1(net769),
    .B1(_0683_),
    .X(_0135_));
 sg13g2_nand2_1 _3516_ (.Y(_0684_),
    .A(net810),
    .B(net475));
 sg13g2_xnor2_1 _3517_ (.Y(_0685_),
    .A(net810),
    .B(_0681_));
 sg13g2_o21ai_1 _3518_ (.B1(_0684_),
    .Y(_0136_),
    .A1(net470),
    .A2(_0685_));
 sg13g2_nand2_1 _3519_ (.Y(_0686_),
    .A(net710),
    .B(net475));
 sg13g2_a21oi_1 _3520_ (.A1(net902),
    .A2(_0681_),
    .Y(_0687_),
    .B1(net710));
 sg13g2_and3_2 _3521_ (.X(_0688_),
    .A(net915),
    .B(net710),
    .C(_0681_));
 sg13g2_or2_1 _3522_ (.X(_0689_),
    .B(_0688_),
    .A(_0687_));
 sg13g2_o21ai_1 _3523_ (.B1(_0686_),
    .Y(_0137_),
    .A1(net470),
    .A2(_0689_));
 sg13g2_nand2_1 _3524_ (.Y(_0690_),
    .A(net814),
    .B(_0642_));
 sg13g2_xnor2_1 _3525_ (.Y(_0691_),
    .A(net814),
    .B(_0688_));
 sg13g2_o21ai_1 _3526_ (.B1(_0690_),
    .Y(_0138_),
    .A1(net470),
    .A2(_0691_));
 sg13g2_nand2_1 _3527_ (.Y(_0692_),
    .A(net742),
    .B(net476));
 sg13g2_a21oi_1 _3528_ (.A1(\audio_inst.i_jump.counter[12] ),
    .A2(_0688_),
    .Y(_0693_),
    .B1(net742));
 sg13g2_nand3_1 _3529_ (.B(\audio_inst.i_jump.counter[12] ),
    .C(_0688_),
    .A(net911),
    .Y(_0694_));
 sg13g2_nand2b_1 _3530_ (.Y(_0695_),
    .B(_0694_),
    .A_N(_0693_));
 sg13g2_o21ai_1 _3531_ (.B1(_0692_),
    .Y(_0139_),
    .A1(net470),
    .A2(_0695_));
 sg13g2_nand2_1 _3532_ (.Y(_0696_),
    .A(net639),
    .B(net476));
 sg13g2_nor2_1 _3533_ (.A(_2068_),
    .B(_0694_),
    .Y(_0697_));
 sg13g2_xnor2_1 _3534_ (.Y(_0698_),
    .A(_2068_),
    .B(_0694_));
 sg13g2_o21ai_1 _3535_ (.B1(_0696_),
    .Y(_0140_),
    .A1(net470),
    .A2(_0698_));
 sg13g2_nand2_1 _3536_ (.Y(_0699_),
    .A(net775),
    .B(net476));
 sg13g2_and2_1 _3537_ (.A(\audio_inst.i_jump.counter[15] ),
    .B(_0697_),
    .X(_0700_));
 sg13g2_o21ai_1 _3538_ (.B1(_0655_),
    .Y(_0701_),
    .A1(net775),
    .A2(_0697_));
 sg13g2_o21ai_1 _3539_ (.B1(_0699_),
    .Y(_0141_),
    .A1(_0700_),
    .A2(_0701_));
 sg13g2_nand2_1 _3540_ (.Y(_0702_),
    .A(net678),
    .B(net476));
 sg13g2_and2_1 _3541_ (.A(net678),
    .B(_0700_),
    .X(_0703_));
 sg13g2_o21ai_1 _3542_ (.B1(_0655_),
    .Y(_0704_),
    .A1(net678),
    .A2(_0700_));
 sg13g2_o21ai_1 _3543_ (.B1(_0702_),
    .Y(_0142_),
    .A1(_0703_),
    .A2(_0704_));
 sg13g2_nand3_1 _3544_ (.B(\audio_inst.i_jump.counter[17] ),
    .C(_0700_),
    .A(net678),
    .Y(_0705_));
 sg13g2_a21oi_1 _3545_ (.A1(_0654_),
    .A2(_0705_),
    .Y(_0706_),
    .B1(net476));
 sg13g2_a21oi_1 _3546_ (.A1(_0643_),
    .A2(_0703_),
    .Y(_0707_),
    .B1(net754));
 sg13g2_nor2_1 _3547_ (.A(_0706_),
    .B(_0707_),
    .Y(_0143_));
 sg13g2_nand4_1 _3548_ (.B(_2070_),
    .C(_0655_),
    .A(net754),
    .Y(_0708_),
    .D(_0703_));
 sg13g2_o21ai_1 _3549_ (.B1(_0708_),
    .Y(_0144_),
    .A1(_2070_),
    .A2(_0706_));
 sg13g2_nor2b_2 _3550_ (.A(\audio_inst.i_over.state[0] ),
    .B_N(\audio_inst.i_over.state[1] ),
    .Y(_0709_));
 sg13g2_nand2b_2 _3551_ (.Y(_0710_),
    .B(\audio_inst.i_over.state[1] ),
    .A_N(\audio_inst.i_over.state[0] ));
 sg13g2_xor2_1 _3552_ (.B(_0394_),
    .A(\audio_inst.i_over.stage_index[4] ),
    .X(_0711_));
 sg13g2_nor2_2 _3553_ (.A(_2087_),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_nand2_2 _3554_ (.Y(_0713_),
    .A(net544),
    .B(net546));
 sg13g2_nor2_1 _3555_ (.A(net539),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_xor2_1 _3556_ (.B(_0713_),
    .A(net539),
    .X(_0715_));
 sg13g2_and2_2 _3557_ (.A(_0712_),
    .B(_0715_),
    .X(_0716_));
 sg13g2_nand2_2 _3558_ (.Y(_0717_),
    .A(_0712_),
    .B(_0715_));
 sg13g2_and2_2 _3559_ (.A(_0712_),
    .B(_0714_),
    .X(_0718_));
 sg13g2_nor2_1 _3560_ (.A(_0009_),
    .B(_0711_),
    .Y(_0719_));
 sg13g2_nand2_2 _3561_ (.Y(_0720_),
    .A(_0715_),
    .B(_0719_));
 sg13g2_nor2_1 _3562_ (.A(_0713_),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_nor2_1 _3563_ (.A(_0718_),
    .B(_0721_),
    .Y(_0722_));
 sg13g2_o21ai_1 _3564_ (.B1(_0722_),
    .Y(_0723_),
    .A1(net544),
    .A2(_0717_));
 sg13g2_o21ai_1 _3565_ (.B1(net462),
    .Y(_0724_),
    .A1(\player_constroller_inst.game_state[0] ),
    .A2(_2188_));
 sg13g2_nor2_2 _3566_ (.A(_2137_),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_nor2b_1 _3567_ (.A(\audio_inst.i_over.state[0] ),
    .B_N(_0711_),
    .Y(_0726_));
 sg13g2_or3_1 _3568_ (.A(_2204_),
    .B(_0725_),
    .C(_0726_),
    .X(_0727_));
 sg13g2_inv_1 _3569_ (.Y(_0728_),
    .A(net484));
 sg13g2_nor2b_2 _3570_ (.A(net546),
    .B_N(net544),
    .Y(_0729_));
 sg13g2_nor2b_2 _3571_ (.A(net544),
    .B_N(net546),
    .Y(_0730_));
 sg13g2_or2_2 _3572_ (.X(_0731_),
    .B(_0730_),
    .A(_0729_));
 sg13g2_inv_1 _3573_ (.Y(_0732_),
    .A(_0731_));
 sg13g2_and2_1 _3574_ (.A(net917),
    .B(_0710_),
    .X(_0733_));
 sg13g2_nand2_1 _3575_ (.Y(_0734_),
    .A(_0026_),
    .B(_0710_));
 sg13g2_nor2_2 _3576_ (.A(net544),
    .B(net546),
    .Y(_0735_));
 sg13g2_inv_1 _3577_ (.Y(_0736_),
    .A(_0735_));
 sg13g2_nor2_1 _3578_ (.A(net538),
    .B(net539),
    .Y(_0737_));
 sg13g2_a22oi_1 _3579_ (.Y(_0738_),
    .B1(_0737_),
    .B2(_0731_),
    .A2(_0735_),
    .A1(net538));
 sg13g2_nor2_1 _3580_ (.A(_0734_),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_a21oi_2 _3581_ (.B1(_0739_),
    .Y(_0740_),
    .A2(_0723_),
    .A1(_0709_));
 sg13g2_nor2_1 _3582_ (.A(net459),
    .B(net473),
    .Y(_0741_));
 sg13g2_a21oi_1 _3583_ (.A1(net473),
    .A2(_0740_),
    .Y(_0145_),
    .B1(_0741_));
 sg13g2_nand3_1 _3584_ (.B(net539),
    .C(_0729_),
    .A(\audio_inst.i_over.stage_index[4] ),
    .Y(_0742_));
 sg13g2_nor2_2 _3585_ (.A(_2087_),
    .B(_0742_),
    .Y(_0743_));
 sg13g2_nand3_1 _3586_ (.B(_0712_),
    .C(_0730_),
    .A(net539),
    .Y(_0744_));
 sg13g2_nand2b_1 _3587_ (.Y(_0745_),
    .B(_0744_),
    .A_N(_0743_));
 sg13g2_nor2_1 _3588_ (.A(_0716_),
    .B(_0745_),
    .Y(_0746_));
 sg13g2_and3_1 _3589_ (.X(_0747_),
    .A(net539),
    .B(_0719_),
    .C(_0730_));
 sg13g2_nor2_1 _3590_ (.A(_0009_),
    .B(_0742_),
    .Y(_0748_));
 sg13g2_nor3_2 _3591_ (.A(_0718_),
    .B(_0747_),
    .C(_0748_),
    .Y(_0749_));
 sg13g2_nand2_1 _3592_ (.Y(_0750_),
    .A(\audio_inst.i_over.stage_index[4] ),
    .B(_0735_));
 sg13g2_nand3_1 _3593_ (.B(net539),
    .C(_0735_),
    .A(\audio_inst.i_over.stage_index[4] ),
    .Y(_0751_));
 sg13g2_nand4_1 _3594_ (.B(_0746_),
    .C(_0749_),
    .A(_0720_),
    .Y(_0752_),
    .D(_0751_));
 sg13g2_and2_2 _3595_ (.A(_0709_),
    .B(_0752_),
    .X(_0753_));
 sg13g2_or2_1 _3596_ (.X(_0754_),
    .B(_0751_),
    .A(_2087_));
 sg13g2_nor2_2 _3597_ (.A(_0009_),
    .B(_0751_),
    .Y(_0755_));
 sg13g2_inv_1 _3598_ (.Y(_0756_),
    .A(_0755_));
 sg13g2_nand3_1 _3599_ (.B(_0751_),
    .C(_0753_),
    .A(_0722_),
    .Y(_0757_));
 sg13g2_nand2_1 _3600_ (.Y(_0758_),
    .A(_0713_),
    .B(_0716_));
 sg13g2_nor2b_1 _3601_ (.A(_0757_),
    .B_N(_0758_),
    .Y(_0759_));
 sg13g2_nor2_1 _3602_ (.A(\audio_inst.i_over.stage_index[4] ),
    .B(_0709_),
    .Y(_0760_));
 sg13g2_nand2b_2 _3603_ (.Y(_0761_),
    .B(_0710_),
    .A_N(\audio_inst.i_over.stage_index[4] ));
 sg13g2_o21ai_1 _3604_ (.B1(_0760_),
    .Y(_0762_),
    .A1(_2018_),
    .A2(net546));
 sg13g2_nor2b_1 _3605_ (.A(net545),
    .B_N(net541),
    .Y(_0763_));
 sg13g2_o21ai_1 _3606_ (.B1(_0762_),
    .Y(_0764_),
    .A1(_0761_),
    .A2(_0763_));
 sg13g2_nand2_1 _3607_ (.Y(_0765_),
    .A(net542),
    .B(_0736_));
 sg13g2_nor2_1 _3608_ (.A(net536),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_nand2b_1 _3609_ (.Y(_0767_),
    .B(_0027_),
    .A_N(net541));
 sg13g2_nand2_1 _3610_ (.Y(_0768_),
    .A(_0764_),
    .B(_0767_));
 sg13g2_o21ai_1 _3611_ (.B1(net473),
    .Y(_0769_),
    .A1(_0766_),
    .A2(_0768_));
 sg13g2_nand2_1 _3612_ (.Y(_0770_),
    .A(net455),
    .B(net483));
 sg13g2_o21ai_1 _3613_ (.B1(_0770_),
    .Y(_0146_),
    .A1(_0759_),
    .A2(_0769_));
 sg13g2_nand2_1 _3614_ (.Y(_0771_),
    .A(_0720_),
    .B(_0753_));
 sg13g2_nor2_1 _3615_ (.A(net539),
    .B(_0750_),
    .Y(_0772_));
 sg13g2_a221oi_1 _3616_ (.B2(_0009_),
    .C1(_0743_),
    .B1(_0772_),
    .A1(_0716_),
    .Y(_0773_),
    .A2(_0729_));
 sg13g2_nand4_1 _3617_ (.B(_0749_),
    .C(_0753_),
    .A(_0720_),
    .Y(_0774_),
    .D(_0773_));
 sg13g2_nand3_1 _3618_ (.B(net540),
    .C(_0730_),
    .A(net538),
    .Y(_0775_));
 sg13g2_a21oi_1 _3619_ (.A1(net542),
    .A2(\audio_inst.i_over.stage_index[0] ),
    .Y(_0776_),
    .B1(net537));
 sg13g2_o21ai_1 _3620_ (.B1(_0776_),
    .Y(_0777_),
    .A1(net542),
    .A2(_0731_));
 sg13g2_a21oi_1 _3621_ (.A1(_0775_),
    .A2(_0777_),
    .Y(_0778_),
    .B1(_0761_));
 sg13g2_nor2_1 _3622_ (.A(net482),
    .B(_0778_),
    .Y(_0779_));
 sg13g2_a22oi_1 _3623_ (.Y(_0780_),
    .B1(_0774_),
    .B2(_0779_),
    .A2(net483),
    .A1(net732));
 sg13g2_inv_1 _3624_ (.Y(_0147_),
    .A(_0780_));
 sg13g2_nor2b_1 _3625_ (.A(_0720_),
    .B_N(_0730_),
    .Y(_0781_));
 sg13g2_nor2_1 _3626_ (.A(_0718_),
    .B(_0781_),
    .Y(_0782_));
 sg13g2_nand2b_1 _3627_ (.Y(_0783_),
    .B(_0716_),
    .A_N(_0713_));
 sg13g2_nand4_1 _3628_ (.B(_0756_),
    .C(_0782_),
    .A(_0742_),
    .Y(_0784_),
    .D(_0783_));
 sg13g2_nand2_1 _3629_ (.Y(_0785_),
    .A(net542),
    .B(_0729_));
 sg13g2_xor2_1 _3630_ (.B(_0729_),
    .A(net543),
    .X(_0786_));
 sg13g2_nor2_2 _3631_ (.A(net542),
    .B(net544),
    .Y(_0787_));
 sg13g2_nor2_1 _3632_ (.A(net541),
    .B(net546),
    .Y(_0788_));
 sg13g2_nor2_1 _3633_ (.A(_0787_),
    .B(_0788_),
    .Y(_0789_));
 sg13g2_a21oi_1 _3634_ (.A1(_0765_),
    .A2(_0789_),
    .Y(_0790_),
    .B1(net537));
 sg13g2_a21oi_1 _3635_ (.A1(net537),
    .A2(_0786_),
    .Y(_0791_),
    .B1(_0790_));
 sg13g2_a221oi_1 _3636_ (.B2(_0733_),
    .C1(net482),
    .B1(_0791_),
    .A1(_0709_),
    .Y(_0792_),
    .A2(_0784_));
 sg13g2_a21oi_1 _3637_ (.A1(_2085_),
    .A2(net483),
    .Y(_0148_),
    .B1(_0792_));
 sg13g2_nor2b_2 _3638_ (.A(_0729_),
    .B_N(net540),
    .Y(_0793_));
 sg13g2_nand2_1 _3639_ (.Y(_0794_),
    .A(net537),
    .B(_0767_));
 sg13g2_o21ai_1 _3640_ (.B1(_0794_),
    .Y(_0795_),
    .A1(net537),
    .A2(_0793_));
 sg13g2_a21oi_1 _3641_ (.A1(_0764_),
    .A2(_0795_),
    .Y(_0796_),
    .B1(net482));
 sg13g2_o21ai_1 _3642_ (.B1(_0796_),
    .Y(_0797_),
    .A1(_0743_),
    .A2(_0757_));
 sg13g2_o21ai_1 _3643_ (.B1(_0797_),
    .Y(_0149_),
    .A1(_2084_),
    .A2(net473));
 sg13g2_nor3_1 _3644_ (.A(net540),
    .B(_0009_),
    .C(_0750_),
    .Y(_0798_));
 sg13g2_or3_1 _3645_ (.A(_0710_),
    .B(_0747_),
    .C(_0798_),
    .X(_0799_));
 sg13g2_a21oi_1 _3646_ (.A1(_0716_),
    .A2(_0730_),
    .Y(_0800_),
    .B1(_0799_));
 sg13g2_nand4_1 _3647_ (.B(_0752_),
    .C(_0754_),
    .A(_0742_),
    .Y(_0801_),
    .D(_0800_));
 sg13g2_nand2_1 _3648_ (.Y(_0802_),
    .A(net536),
    .B(_2205_));
 sg13g2_nor2_1 _3649_ (.A(_0787_),
    .B(_0802_),
    .Y(_0803_));
 sg13g2_o21ai_1 _3650_ (.B1(_0760_),
    .Y(_0804_),
    .A1(net537),
    .A2(_0786_));
 sg13g2_a21oi_1 _3651_ (.A1(_0736_),
    .A2(_0803_),
    .Y(_0805_),
    .B1(_0804_));
 sg13g2_nor2_1 _3652_ (.A(net482),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_a22oi_1 _3653_ (.Y(_0807_),
    .B1(_0801_),
    .B2(_0806_),
    .A2(net483),
    .A1(net688));
 sg13g2_inv_1 _3654_ (.Y(_0150_),
    .A(_0807_));
 sg13g2_o21ai_1 _3655_ (.B1(_0756_),
    .Y(_0808_),
    .A1(_0717_),
    .A2(_0735_));
 sg13g2_nor2_1 _3656_ (.A(_0799_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_o21ai_1 _3657_ (.B1(_2205_),
    .Y(_0810_),
    .A1(net545),
    .A2(_2118_));
 sg13g2_nand2b_1 _3658_ (.Y(_0811_),
    .B(_0731_),
    .A_N(_0802_));
 sg13g2_a21oi_1 _3659_ (.A1(_2018_),
    .A2(_0810_),
    .Y(_0812_),
    .B1(_0761_));
 sg13g2_a221oi_1 _3660_ (.B2(_0812_),
    .C1(net482),
    .B1(_0811_),
    .A1(_0752_),
    .Y(_0813_),
    .A2(_0809_));
 sg13g2_a21o_1 _3661_ (.A2(net485),
    .A1(net716),
    .B1(_0813_),
    .X(_0151_));
 sg13g2_nor2_1 _3662_ (.A(_0717_),
    .B(_0731_),
    .Y(_0814_));
 sg13g2_nor4_2 _3663_ (.A(_0748_),
    .B(_0755_),
    .C(_0771_),
    .Y(_0815_),
    .D(_0814_));
 sg13g2_a21oi_1 _3664_ (.A1(net541),
    .A2(_0027_),
    .Y(_0816_),
    .B1(net536));
 sg13g2_nand2b_1 _3665_ (.Y(_0817_),
    .B(_0735_),
    .A_N(net542));
 sg13g2_a22oi_1 _3666_ (.Y(_0818_),
    .B1(_0816_),
    .B2(_0817_),
    .A2(_0788_),
    .A1(net536));
 sg13g2_o21ai_1 _3667_ (.B1(net473),
    .Y(_0819_),
    .A1(_0761_),
    .A2(_0818_));
 sg13g2_nand2_1 _3668_ (.Y(_0820_),
    .A(net446),
    .B(net484));
 sg13g2_o21ai_1 _3669_ (.B1(_0820_),
    .Y(_0152_),
    .A1(_0815_),
    .A2(_0819_));
 sg13g2_nor4_1 _3670_ (.A(_0710_),
    .B(_0743_),
    .C(_0747_),
    .D(_0814_),
    .Y(_0821_));
 sg13g2_and3_1 _3671_ (.X(_0822_),
    .A(_0752_),
    .B(_0782_),
    .C(_0821_));
 sg13g2_o21ai_1 _3672_ (.B1(_0816_),
    .Y(_0823_),
    .A1(net541),
    .A2(_0731_));
 sg13g2_nand2b_1 _3673_ (.Y(_0824_),
    .B(_0028_),
    .A_N(net541));
 sg13g2_nand3_1 _3674_ (.B(_0785_),
    .C(_0824_),
    .A(net536),
    .Y(_0825_));
 sg13g2_a21oi_1 _3675_ (.A1(_0823_),
    .A2(_0825_),
    .Y(_0826_),
    .B1(_0761_));
 sg13g2_nor3_1 _3676_ (.A(net482),
    .B(_0822_),
    .C(_0826_),
    .Y(_0827_));
 sg13g2_a21o_1 _3677_ (.A2(net484),
    .A1(net687),
    .B1(_0827_),
    .X(_0153_));
 sg13g2_nor2_1 _3678_ (.A(_0721_),
    .B(_0798_),
    .Y(_0828_));
 sg13g2_nand2_1 _3679_ (.Y(_0829_),
    .A(_0749_),
    .B(_0828_));
 sg13g2_or2_1 _3680_ (.X(_0830_),
    .B(_0829_),
    .A(_0781_));
 sg13g2_nand3_1 _3681_ (.B(_0753_),
    .C(_0758_),
    .A(_0744_),
    .Y(_0831_));
 sg13g2_nor2_1 _3682_ (.A(net537),
    .B(_0824_),
    .Y(_0832_));
 sg13g2_nor4_1 _3683_ (.A(_0762_),
    .B(_0766_),
    .C(_0803_),
    .D(_0832_),
    .Y(_0833_));
 sg13g2_nor2_1 _3684_ (.A(net482),
    .B(_0833_),
    .Y(_0834_));
 sg13g2_o21ai_1 _3685_ (.B1(_0834_),
    .Y(_0835_),
    .A1(_0830_),
    .A2(_0831_));
 sg13g2_o21ai_1 _3686_ (.B1(_0835_),
    .Y(_0154_),
    .A1(_2083_),
    .A2(_0728_));
 sg13g2_nor2_2 _3687_ (.A(_0720_),
    .B(_0732_),
    .Y(_0836_));
 sg13g2_o21ai_1 _3688_ (.B1(_0709_),
    .Y(_0837_),
    .A1(_0793_),
    .A2(_0836_));
 sg13g2_o21ai_1 _3689_ (.B1(_0765_),
    .Y(_0838_),
    .A1(net543),
    .A2(_0731_));
 sg13g2_o21ai_1 _3690_ (.B1(_0838_),
    .Y(_0839_),
    .A1(_2018_),
    .A2(_2205_));
 sg13g2_a21oi_1 _3691_ (.A1(_0733_),
    .A2(_0839_),
    .Y(_0840_),
    .B1(net484));
 sg13g2_a22oi_1 _3692_ (.Y(_0155_),
    .B1(_0837_),
    .B2(_0840_),
    .A2(net484),
    .A1(_2082_));
 sg13g2_a21oi_1 _3693_ (.A1(net546),
    .A2(_0716_),
    .Y(_0841_),
    .B1(_0743_));
 sg13g2_nand3b_1 _3694_ (.B(_0841_),
    .C(_0749_),
    .Y(_0842_),
    .A_N(_0836_));
 sg13g2_nand2_1 _3695_ (.Y(_0843_),
    .A(_0709_),
    .B(_0842_));
 sg13g2_nand2b_1 _3696_ (.Y(_0844_),
    .B(_0730_),
    .A_N(net542));
 sg13g2_a21oi_1 _3697_ (.A1(net541),
    .A2(_0027_),
    .Y(_0845_),
    .B1(_2018_));
 sg13g2_a22oi_1 _3698_ (.Y(_0846_),
    .B1(_0844_),
    .B2(_0845_),
    .A2(_0789_),
    .A1(_0776_));
 sg13g2_nor2_1 _3699_ (.A(_0734_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_nor2_1 _3700_ (.A(net484),
    .B(_0847_),
    .Y(_0848_));
 sg13g2_a22oi_1 _3701_ (.Y(_0156_),
    .B1(_0843_),
    .B2(_0848_),
    .A2(net484),
    .A1(_2081_));
 sg13g2_nor4_1 _3702_ (.A(_0718_),
    .B(_0755_),
    .C(_0814_),
    .D(_0836_),
    .Y(_0849_));
 sg13g2_nand3_1 _3703_ (.B(_0753_),
    .C(_0849_),
    .A(_0744_),
    .Y(_0850_));
 sg13g2_nor3_1 _3704_ (.A(net536),
    .B(_0763_),
    .C(_0788_),
    .Y(_0851_));
 sg13g2_o21ai_1 _3705_ (.B1(_0733_),
    .Y(_0852_),
    .A1(_0803_),
    .A2(_0851_));
 sg13g2_nand3_1 _3706_ (.B(_0850_),
    .C(_0852_),
    .A(net473),
    .Y(_0853_));
 sg13g2_o21ai_1 _3707_ (.B1(_0853_),
    .Y(_0157_),
    .A1(_2080_),
    .A2(_0728_));
 sg13g2_nor3_1 _3708_ (.A(_0745_),
    .B(_0755_),
    .C(_0829_),
    .Y(_0854_));
 sg13g2_nand2b_1 _3709_ (.Y(_0855_),
    .B(_0009_),
    .A_N(net545));
 sg13g2_nand3_1 _3710_ (.B(_0733_),
    .C(_0855_),
    .A(_2205_),
    .Y(_0856_));
 sg13g2_o21ai_1 _3711_ (.B1(_0856_),
    .Y(_0857_),
    .A1(_0710_),
    .A2(_0854_));
 sg13g2_mux2_1 _3712_ (.A0(net679),
    .A1(_0857_),
    .S(net473),
    .X(_0158_));
 sg13g2_or3_1 _3713_ (.A(net536),
    .B(_0734_),
    .C(_0787_),
    .X(_0858_));
 sg13g2_o21ai_1 _3714_ (.B1(_0858_),
    .Y(_0859_),
    .A1(_0710_),
    .A2(_0746_));
 sg13g2_mux2_1 _3715_ (.A0(net693),
    .A1(_0859_),
    .S(net473),
    .X(_0159_));
 sg13g2_nand2_1 _3716_ (.Y(_0860_),
    .A(_0009_),
    .B(_0787_));
 sg13g2_a221oi_1 _3717_ (.B2(_0860_),
    .C1(net482),
    .B1(_0760_),
    .A1(_0753_),
    .Y(_0861_),
    .A2(_0754_));
 sg13g2_a21o_1 _3718_ (.A2(net484),
    .A1(net746),
    .B1(_0861_),
    .X(_0160_));
 sg13g2_nand2b_1 _3719_ (.Y(_0862_),
    .B(net534),
    .A_N(net529));
 sg13g2_nor2b_2 _3720_ (.A(net534),
    .B_N(net529),
    .Y(_0863_));
 sg13g2_nand2b_2 _3721_ (.Y(_0864_),
    .B(net535),
    .A_N(net533));
 sg13g2_o21ai_1 _3722_ (.B1(_0864_),
    .Y(_0865_),
    .A1(net531),
    .A2(_2190_));
 sg13g2_nand2b_1 _3723_ (.Y(_0866_),
    .B(net520),
    .A_N(_0865_));
 sg13g2_nand3_1 _3724_ (.B(_0591_),
    .C(_0592_),
    .A(net528),
    .Y(_0867_));
 sg13g2_a21oi_1 _3725_ (.A1(_0866_),
    .A2(_0867_),
    .Y(_0868_),
    .B1(net525));
 sg13g2_mux2_1 _3726_ (.A0(_0868_),
    .A1(net752),
    .S(net480),
    .X(_0161_));
 sg13g2_nand2_2 _3727_ (.Y(_0869_),
    .A(net520),
    .B(net532));
 sg13g2_a21oi_1 _3728_ (.A1(_0591_),
    .A2(_0869_),
    .Y(_0870_),
    .B1(net525));
 sg13g2_o21ai_1 _3729_ (.B1(_0870_),
    .Y(_0871_),
    .A1(net528),
    .A2(_0864_));
 sg13g2_nand2_1 _3730_ (.Y(_0872_),
    .A(net444),
    .B(net481));
 sg13g2_o21ai_1 _3731_ (.B1(_0872_),
    .Y(_0162_),
    .A1(net480),
    .A2(_0871_));
 sg13g2_nor2_1 _3732_ (.A(net532),
    .B(net534),
    .Y(_0873_));
 sg13g2_or2_1 _3733_ (.X(_0874_),
    .B(net535),
    .A(net533));
 sg13g2_nand2_1 _3734_ (.Y(_0875_),
    .A(net529),
    .B(_0874_));
 sg13g2_nand2_1 _3735_ (.Y(_0876_),
    .A(net520),
    .B(_0875_));
 sg13g2_nor2b_2 _3736_ (.A(net529),
    .B_N(_0864_),
    .Y(_0877_));
 sg13g2_nand2_2 _3737_ (.Y(_0878_),
    .A(net533),
    .B(net535));
 sg13g2_nand3b_1 _3738_ (.B(_0878_),
    .C(net527),
    .Y(_0879_),
    .A_N(net529));
 sg13g2_nand2_1 _3739_ (.Y(_0880_),
    .A(net523),
    .B(_0879_));
 sg13g2_inv_1 _3740_ (.Y(_0881_),
    .A(_0880_));
 sg13g2_o21ai_1 _3741_ (.B1(_0881_),
    .Y(_0882_),
    .A1(_0876_),
    .A2(_0877_));
 sg13g2_nand2_1 _3742_ (.Y(_0883_),
    .A(net530),
    .B(_0006_));
 sg13g2_nor2_1 _3743_ (.A(net526),
    .B(_0862_),
    .Y(_0884_));
 sg13g2_a21oi_1 _3744_ (.A1(_0862_),
    .A2(_0883_),
    .Y(_0885_),
    .B1(net526));
 sg13g2_or2_2 _3745_ (.X(_0886_),
    .B(_0878_),
    .A(_2192_));
 sg13g2_nand2_1 _3746_ (.Y(_0887_),
    .A(_0879_),
    .B(_0886_));
 sg13g2_a21oi_1 _3747_ (.A1(_0591_),
    .A2(_0885_),
    .Y(_0888_),
    .B1(_0887_));
 sg13g2_o21ai_1 _3748_ (.B1(_0882_),
    .Y(_0889_),
    .A1(net523),
    .A2(_0888_));
 sg13g2_mux2_1 _3749_ (.A0(_0889_),
    .A1(net675),
    .S(net477),
    .X(_0163_));
 sg13g2_nor2_1 _3750_ (.A(net526),
    .B(_0592_),
    .Y(_0890_));
 sg13g2_nor2_1 _3751_ (.A(net523),
    .B(_0890_),
    .Y(_0891_));
 sg13g2_nor3_1 _3752_ (.A(net523),
    .B(_0884_),
    .C(_0890_),
    .Y(_0892_));
 sg13g2_nor2_1 _3753_ (.A(_2007_),
    .B(_2190_),
    .Y(_0893_));
 sg13g2_o21ai_1 _3754_ (.B1(_0893_),
    .Y(_0894_),
    .A1(net532),
    .A2(_0021_));
 sg13g2_nand2_1 _3755_ (.Y(_0895_),
    .A(_2007_),
    .B(_0590_));
 sg13g2_nand3_1 _3756_ (.B(_0894_),
    .C(_0895_),
    .A(_0892_),
    .Y(_0896_));
 sg13g2_nand2_1 _3757_ (.Y(_0897_),
    .A(net527),
    .B(_0592_));
 sg13g2_nand2_2 _3758_ (.Y(_0898_),
    .A(_2191_),
    .B(_0864_));
 sg13g2_nand3_1 _3759_ (.B(_0592_),
    .C(_0864_),
    .A(net527),
    .Y(_0899_));
 sg13g2_nor2_1 _3760_ (.A(net526),
    .B(_0863_),
    .Y(_0900_));
 sg13g2_nor3_2 _3761_ (.A(net526),
    .B(_0863_),
    .C(_0873_),
    .Y(_0901_));
 sg13g2_o21ai_1 _3762_ (.B1(net523),
    .Y(_0902_),
    .A1(_0897_),
    .A2(_0898_));
 sg13g2_o21ai_1 _3763_ (.B1(_0896_),
    .Y(_0903_),
    .A1(_0901_),
    .A2(_0902_));
 sg13g2_nand2_1 _3764_ (.Y(_0904_),
    .A(net425),
    .B(net477));
 sg13g2_o21ai_1 _3765_ (.B1(_0904_),
    .Y(_0164_),
    .A1(net477),
    .A2(_0903_));
 sg13g2_nor2_1 _3766_ (.A(net535),
    .B(_0591_),
    .Y(_0905_));
 sg13g2_a21oi_1 _3767_ (.A1(net526),
    .A2(_0905_),
    .Y(_0906_),
    .B1(_2006_));
 sg13g2_nand2b_1 _3768_ (.Y(_0907_),
    .B(_0906_),
    .A_N(_0885_));
 sg13g2_a21oi_1 _3769_ (.A1(_2192_),
    .A2(_0869_),
    .Y(_0908_),
    .B1(_0863_));
 sg13g2_o21ai_1 _3770_ (.B1(_0907_),
    .Y(_0909_),
    .A1(net523),
    .A2(_0908_));
 sg13g2_nand2_1 _3771_ (.Y(_0910_),
    .A(net424),
    .B(net477));
 sg13g2_o21ai_1 _3772_ (.B1(_0910_),
    .Y(_0165_),
    .A1(net478),
    .A2(_0909_));
 sg13g2_nand2_1 _3773_ (.Y(_0911_),
    .A(net520),
    .B(_2040_));
 sg13g2_a221oi_1 _3774_ (.B2(_0911_),
    .C1(net478),
    .B1(_0906_),
    .A1(_0891_),
    .Y(_0912_),
    .A2(_0899_));
 sg13g2_a21oi_1 _3775_ (.A1(_2072_),
    .A2(net477),
    .Y(_0166_),
    .B1(_0912_));
 sg13g2_o21ai_1 _3776_ (.B1(net523),
    .Y(_0913_),
    .A1(_0873_),
    .A2(_0879_));
 sg13g2_and2_1 _3777_ (.A(net529),
    .B(_0898_),
    .X(_0914_));
 sg13g2_nor3_1 _3778_ (.A(net526),
    .B(_0433_),
    .C(_0914_),
    .Y(_0915_));
 sg13g2_nor2_1 _3779_ (.A(_0877_),
    .B(_0914_),
    .Y(_0916_));
 sg13g2_o21ai_1 _3780_ (.B1(net520),
    .Y(_0917_),
    .A1(net529),
    .A2(_0873_));
 sg13g2_a21oi_1 _3781_ (.A1(_0916_),
    .A2(_0917_),
    .Y(_0918_),
    .B1(net523));
 sg13g2_o21ai_1 _3782_ (.B1(_0918_),
    .Y(_0919_),
    .A1(_0916_),
    .A2(_0917_));
 sg13g2_o21ai_1 _3783_ (.B1(_0919_),
    .Y(_0920_),
    .A1(_0913_),
    .A2(_0915_));
 sg13g2_mux2_1 _3784_ (.A0(_0920_),
    .A1(net706),
    .S(net477),
    .X(_0167_));
 sg13g2_a21oi_1 _3785_ (.A1(_2191_),
    .A2(_0877_),
    .Y(_0921_),
    .B1(_0876_));
 sg13g2_nand2_1 _3786_ (.Y(_0922_),
    .A(_2006_),
    .B(net528));
 sg13g2_nor3_1 _3787_ (.A(_0590_),
    .B(_0898_),
    .C(_0922_),
    .Y(_0923_));
 sg13g2_a22oi_1 _3788_ (.Y(_0924_),
    .B1(_0863_),
    .B2(net532),
    .A2(_0590_),
    .A1(net534));
 sg13g2_nand2_1 _3789_ (.Y(_0925_),
    .A(_0431_),
    .B(_0924_));
 sg13g2_o21ai_1 _3790_ (.B1(_0925_),
    .Y(_0926_),
    .A1(_0880_),
    .A2(_0921_));
 sg13g2_nor3_1 _3791_ (.A(net479),
    .B(_0923_),
    .C(_0926_),
    .Y(_0927_));
 sg13g2_a21o_1 _3792_ (.A2(net478),
    .A1(net458),
    .B1(_0927_),
    .X(_0168_));
 sg13g2_a21oi_1 _3793_ (.A1(net534),
    .A2(_0006_),
    .Y(_0928_),
    .B1(_0863_));
 sg13g2_o21ai_1 _3794_ (.B1(_0879_),
    .Y(_0929_),
    .A1(_2007_),
    .A2(_0883_));
 sg13g2_nand2_1 _3795_ (.Y(_0930_),
    .A(_0021_),
    .B(_0874_));
 sg13g2_and2_1 _3796_ (.A(net525),
    .B(_0020_),
    .X(_0931_));
 sg13g2_a22oi_1 _3797_ (.Y(_0932_),
    .B1(_0930_),
    .B2(_0931_),
    .A2(_0929_),
    .A1(_2006_));
 sg13g2_o21ai_1 _3798_ (.B1(_0932_),
    .Y(_0933_),
    .A1(_0432_),
    .A2(_0928_));
 sg13g2_mux2_1 _3799_ (.A0(_0933_),
    .A1(net702),
    .S(net477),
    .X(_0169_));
 sg13g2_a22oi_1 _3800_ (.Y(_0934_),
    .B1(_0877_),
    .B2(_2191_),
    .A2(_0863_),
    .A1(net532));
 sg13g2_o21ai_1 _3801_ (.B1(_0892_),
    .Y(_0935_),
    .A1(net520),
    .A2(_0934_));
 sg13g2_o21ai_1 _3802_ (.B1(_0935_),
    .Y(_0936_),
    .A1(_0900_),
    .A2(_0913_));
 sg13g2_nand2_1 _3803_ (.Y(_0937_),
    .A(net451),
    .B(net477));
 sg13g2_o21ai_1 _3804_ (.B1(_0937_),
    .Y(_0170_),
    .A1(net478),
    .A2(_0936_));
 sg13g2_nand2_1 _3805_ (.Y(_0938_),
    .A(net527),
    .B(_0875_));
 sg13g2_nor2_1 _3806_ (.A(_0905_),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_nor2_1 _3807_ (.A(_2006_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_a21oi_1 _3808_ (.A1(net520),
    .A2(_0914_),
    .Y(_0941_),
    .B1(_0884_));
 sg13g2_nand3_1 _3809_ (.B(_0864_),
    .C(_0869_),
    .A(_2192_),
    .Y(_0942_));
 sg13g2_a21oi_1 _3810_ (.A1(net534),
    .A2(_2193_),
    .Y(_0943_),
    .B1(net524));
 sg13g2_a221oi_1 _3811_ (.B2(_0943_),
    .C1(net478),
    .B1(_0942_),
    .A1(_0940_),
    .Y(_0944_),
    .A2(_0941_));
 sg13g2_a21o_1 _3812_ (.A2(net479),
    .A1(net677),
    .B1(_0944_),
    .X(_0171_));
 sg13g2_nand4_1 _3813_ (.B(net527),
    .C(_0875_),
    .A(_2006_),
    .Y(_0945_),
    .D(_0878_));
 sg13g2_a21oi_1 _3814_ (.A1(net534),
    .A2(_0590_),
    .Y(_0946_),
    .B1(_2190_));
 sg13g2_nor2_1 _3815_ (.A(net527),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_o21ai_1 _3816_ (.B1(_0945_),
    .Y(_0948_),
    .A1(_0880_),
    .A2(_0947_));
 sg13g2_a21oi_1 _3817_ (.A1(_0431_),
    .A2(_0916_),
    .Y(_0949_),
    .B1(_0948_));
 sg13g2_mux2_1 _3818_ (.A0(_0949_),
    .A1(net689),
    .S(net479),
    .X(_0172_));
 sg13g2_nor3_1 _3819_ (.A(net524),
    .B(_0901_),
    .C(_0929_),
    .Y(_0950_));
 sg13g2_a21oi_1 _3820_ (.A1(_0866_),
    .A2(_0940_),
    .Y(_0951_),
    .B1(_0950_));
 sg13g2_mux2_1 _3821_ (.A0(_0951_),
    .A1(net707),
    .S(net479),
    .X(_0173_));
 sg13g2_a21oi_1 _3822_ (.A1(_0591_),
    .A2(_0869_),
    .Y(_0952_),
    .B1(_2006_));
 sg13g2_a22oi_1 _3823_ (.Y(_0953_),
    .B1(_0864_),
    .B2(_0952_),
    .A2(_0431_),
    .A1(_0022_));
 sg13g2_o21ai_1 _3824_ (.B1(_0953_),
    .Y(_0954_),
    .A1(_0922_),
    .A2(_0924_));
 sg13g2_mux2_1 _3825_ (.A0(_0954_),
    .A1(net697),
    .S(net478),
    .X(_0174_));
 sg13g2_nor2_1 _3826_ (.A(_0865_),
    .B(_0922_),
    .Y(_0955_));
 sg13g2_and3_1 _3827_ (.X(_0956_),
    .A(_0591_),
    .B(_0592_),
    .C(_0931_));
 sg13g2_nor3_1 _3828_ (.A(_0021_),
    .B(_0432_),
    .C(_0864_),
    .Y(_0957_));
 sg13g2_nor4_1 _3829_ (.A(net480),
    .B(_0955_),
    .C(_0956_),
    .D(_0957_),
    .Y(_0958_));
 sg13g2_a21oi_1 _3830_ (.A1(_2078_),
    .A2(net480),
    .Y(_0175_),
    .B1(_0958_));
 sg13g2_nor2_1 _3831_ (.A(_0877_),
    .B(_0897_),
    .Y(_0959_));
 sg13g2_a21oi_1 _3832_ (.A1(net524),
    .A2(_0895_),
    .Y(_0960_),
    .B1(_0959_));
 sg13g2_a21oi_1 _3833_ (.A1(_0925_),
    .A2(_0960_),
    .Y(_0961_),
    .B1(net478));
 sg13g2_a21oi_1 _3834_ (.A1(_2077_),
    .A2(net480),
    .Y(_0176_),
    .B1(_0961_));
 sg13g2_nand3_1 _3835_ (.B(net619),
    .C(_2200_),
    .A(net433),
    .Y(_0962_));
 sg13g2_nand2b_1 _3836_ (.Y(_0963_),
    .B(_0394_),
    .A_N(\audio_inst.i_over.state[0] ));
 sg13g2_nand3_1 _3837_ (.B(_2203_),
    .C(_0963_),
    .A(net619),
    .Y(_0964_));
 sg13g2_o21ai_1 _3838_ (.B1(_0962_),
    .Y(_0177_),
    .A1(_0395_),
    .A2(_0964_));
 sg13g2_nor2_1 _3839_ (.A(net598),
    .B(_2119_),
    .Y(_0178_));
 sg13g2_o21ai_1 _3840_ (.B1(net613),
    .Y(_0965_),
    .A1(net590),
    .A2(net588));
 sg13g2_nor2_1 _3841_ (.A(_0415_),
    .B(_0965_),
    .Y(_0179_));
 sg13g2_xnor2_1 _3842_ (.Y(_0966_),
    .A(net830),
    .B(_0415_));
 sg13g2_nor2_1 _3843_ (.A(net602),
    .B(_0966_),
    .Y(_0180_));
 sg13g2_a21oi_1 _3844_ (.A1(net830),
    .A2(_0416_),
    .Y(_0967_),
    .B1(net581));
 sg13g2_nor3_1 _3845_ (.A(_2047_),
    .B(_2120_),
    .C(_0415_),
    .Y(_0968_));
 sg13g2_nor3_1 _3846_ (.A(net602),
    .B(_0967_),
    .C(_0968_),
    .Y(_0181_));
 sg13g2_nor3_1 _3847_ (.A(net584),
    .B(net582),
    .C(_0415_),
    .Y(_0969_));
 sg13g2_and2_1 _3848_ (.A(_2048_),
    .B(_0969_),
    .X(_0970_));
 sg13g2_xnor2_1 _3849_ (.Y(_0971_),
    .A(net579),
    .B(_0969_));
 sg13g2_nor2_1 _3850_ (.A(net598),
    .B(_0971_),
    .Y(_0182_));
 sg13g2_o21ai_1 _3851_ (.B1(net614),
    .Y(_0972_),
    .A1(net576),
    .A2(_0970_));
 sg13g2_a21oi_1 _3852_ (.A1(net576),
    .A2(_0970_),
    .Y(_0183_),
    .B1(_0972_));
 sg13g2_and2_1 _3853_ (.A(net556),
    .B(net557),
    .X(_0973_));
 sg13g2_nand2_1 _3854_ (.Y(_0974_),
    .A(net555),
    .B(net557));
 sg13g2_nor2_2 _3855_ (.A(_2042_),
    .B(_0974_),
    .Y(_0975_));
 sg13g2_nand2_1 _3856_ (.Y(_0976_),
    .A(net554),
    .B(_0973_));
 sg13g2_xnor2_1 _3857_ (.Y(_0977_),
    .A(net759),
    .B(_0975_));
 sg13g2_nor2_1 _3858_ (.A(net600),
    .B(_0977_),
    .Y(_0184_));
 sg13g2_o21ai_1 _3859_ (.B1(net875),
    .Y(_0978_),
    .A1(net552),
    .A2(_0976_));
 sg13g2_xnor2_1 _3860_ (.Y(_0979_),
    .A(_2043_),
    .B(_0978_));
 sg13g2_nor2_1 _3861_ (.A(net600),
    .B(_0979_),
    .Y(_0185_));
 sg13g2_nor3_2 _3862_ (.A(net550),
    .B(net872),
    .C(_0978_),
    .Y(_0980_));
 sg13g2_o21ai_1 _3863_ (.B1(net550),
    .Y(_0981_),
    .A1(net872),
    .A2(_0978_));
 sg13g2_nor2b_1 _3864_ (.A(_0980_),
    .B_N(_0981_),
    .Y(_0982_));
 sg13g2_nor2_1 _3865_ (.A(net600),
    .B(_0982_),
    .Y(_0186_));
 sg13g2_and2_1 _3866_ (.A(_2044_),
    .B(_0980_),
    .X(_0983_));
 sg13g2_xnor2_1 _3867_ (.Y(_0984_),
    .A(net882),
    .B(_0980_));
 sg13g2_nor2_1 _3868_ (.A(net600),
    .B(_0984_),
    .Y(_0187_));
 sg13g2_o21ai_1 _3869_ (.B1(net617),
    .Y(_0985_),
    .A1(net859),
    .A2(_0983_));
 sg13g2_a21oi_1 _3870_ (.A1(net859),
    .A2(_0983_),
    .Y(_0188_),
    .B1(_0985_));
 sg13g2_a21oi_1 _3871_ (.A1(_2125_),
    .A2(_0399_),
    .Y(_0189_),
    .B1(net606));
 sg13g2_o21ai_1 _3872_ (.B1(net613),
    .Y(_0986_),
    .A1(_2119_),
    .A2(_2125_));
 sg13g2_a21oi_1 _3873_ (.A1(_2119_),
    .A2(_2125_),
    .Y(_0190_),
    .B1(_0986_));
 sg13g2_nand2_1 _3874_ (.Y(_0987_),
    .A(net590),
    .B(_2125_));
 sg13g2_xor2_1 _3875_ (.B(_0987_),
    .A(net587),
    .X(_0988_));
 sg13g2_nor2_1 _3876_ (.A(net598),
    .B(_0988_),
    .Y(_0191_));
 sg13g2_o21ai_1 _3877_ (.B1(net587),
    .Y(_0989_),
    .A1(net588),
    .A2(_0987_));
 sg13g2_xor2_1 _3878_ (.B(_0989_),
    .A(net584),
    .X(_0990_));
 sg13g2_nor2_1 _3879_ (.A(net599),
    .B(_0990_),
    .Y(_0192_));
 sg13g2_or3_1 _3880_ (.A(net584),
    .B(net582),
    .C(_0989_),
    .X(_0991_));
 sg13g2_o21ai_1 _3881_ (.B1(net582),
    .Y(_0992_),
    .A1(net584),
    .A2(_0989_));
 sg13g2_a21oi_1 _3882_ (.A1(_0991_),
    .A2(_0992_),
    .Y(_0193_),
    .B1(net599));
 sg13g2_nor2_1 _3883_ (.A(net578),
    .B(_0991_),
    .Y(_0993_));
 sg13g2_xnor2_1 _3884_ (.Y(_0994_),
    .A(_2048_),
    .B(_0991_));
 sg13g2_nor2_1 _3885_ (.A(net598),
    .B(_0994_),
    .Y(_0194_));
 sg13g2_o21ai_1 _3886_ (.B1(net615),
    .Y(_0995_),
    .A1(net691),
    .A2(_0993_));
 sg13g2_a21oi_1 _3887_ (.A1(net691),
    .A2(_0993_),
    .Y(_0195_),
    .B1(_0995_));
 sg13g2_and2_1 _3888_ (.A(net406),
    .B(net609),
    .X(_0196_));
 sg13g2_and2_1 _3889_ (.A(net426),
    .B(net609),
    .X(_0197_));
 sg13g2_and2_1 _3890_ (.A(net403),
    .B(net609),
    .X(_0198_));
 sg13g2_and2_1 _3891_ (.A(net405),
    .B(net609),
    .X(_0199_));
 sg13g2_and2_1 _3892_ (.A(net613),
    .B(net388),
    .X(_0200_));
 sg13g2_and2_1 _3893_ (.A(net592),
    .B(net613),
    .X(_0224_));
 sg13g2_nor2_1 _3894_ (.A(_2046_),
    .B(net598),
    .Y(_0225_));
 sg13g2_nor2_1 _3895_ (.A(_0224_),
    .B(_0225_),
    .Y(_0996_));
 sg13g2_a21oi_1 _3896_ (.A1(net592),
    .A2(net590),
    .Y(_0201_),
    .B1(_0996_));
 sg13g2_and3_1 _3897_ (.X(_0202_),
    .A(net612),
    .B(_0417_),
    .C(_0583_));
 sg13g2_o21ai_1 _3898_ (.B1(net612),
    .Y(_0997_),
    .A1(net584),
    .A2(_0579_));
 sg13g2_a21oi_1 _3899_ (.A1(net584),
    .A2(_0579_),
    .Y(_0203_),
    .B1(_0997_));
 sg13g2_a21oi_1 _3900_ (.A1(net592),
    .A2(_0415_),
    .Y(_0998_),
    .B1(net582));
 sg13g2_nor2_1 _3901_ (.A(_0417_),
    .B(_0423_),
    .Y(_0999_));
 sg13g2_o21ai_1 _3902_ (.B1(net612),
    .Y(_1000_),
    .A1(net584),
    .A2(net582));
 sg13g2_nor3_1 _3903_ (.A(_0998_),
    .B(_0999_),
    .C(_1000_),
    .Y(_0204_));
 sg13g2_nor3_1 _3904_ (.A(_2048_),
    .B(_0417_),
    .C(_0423_),
    .Y(_1001_));
 sg13g2_o21ai_1 _3905_ (.B1(net614),
    .Y(_1002_),
    .A1(net578),
    .A2(_0999_));
 sg13g2_nor2_1 _3906_ (.A(_1001_),
    .B(_1002_),
    .Y(_0205_));
 sg13g2_o21ai_1 _3907_ (.B1(net612),
    .Y(_1003_),
    .A1(net576),
    .A2(_1001_));
 sg13g2_a21oi_1 _3908_ (.A1(net576),
    .A2(_1001_),
    .Y(_0206_),
    .B1(_1003_));
 sg13g2_nor2_1 _3909_ (.A(_2021_),
    .B(net596),
    .Y(_0207_));
 sg13g2_nor2_1 _3910_ (.A(_2020_),
    .B(net596),
    .Y(_0208_));
 sg13g2_and2_1 _3911_ (.A(net452),
    .B(net609),
    .X(_0209_));
 sg13g2_and2_1 _3912_ (.A(net649),
    .B(net609),
    .X(_0210_));
 sg13g2_and2_1 _3913_ (.A(net613),
    .B(net667),
    .X(_0211_));
 sg13g2_and3_1 _3914_ (.X(_0212_),
    .A(net610),
    .B(_2125_),
    .C(_0399_));
 sg13g2_nand2_1 _3915_ (.Y(_1004_),
    .A(net613),
    .B(_0400_));
 sg13g2_a21oi_1 _3916_ (.A1(_2046_),
    .A2(_0399_),
    .Y(_0213_),
    .B1(_1004_));
 sg13g2_o21ai_1 _3917_ (.B1(net613),
    .Y(_1005_),
    .A1(net587),
    .A2(_0412_));
 sg13g2_a21oi_1 _3918_ (.A1(net587),
    .A2(_0412_),
    .Y(_0214_),
    .B1(_1005_));
 sg13g2_o21ai_1 _3919_ (.B1(net811),
    .Y(_1006_),
    .A1(net588),
    .A2(_0400_));
 sg13g2_o21ai_1 _3920_ (.B1(net612),
    .Y(_1007_),
    .A1(_2120_),
    .A2(_1006_));
 sg13g2_a21oi_1 _3921_ (.A1(_2120_),
    .A2(_1006_),
    .Y(_0215_),
    .B1(_1007_));
 sg13g2_nand2b_1 _3922_ (.Y(_1008_),
    .B(_1006_),
    .A_N(_0423_));
 sg13g2_o21ai_1 _3923_ (.B1(_1008_),
    .Y(_1009_),
    .A1(net582),
    .A2(_1006_));
 sg13g2_nor2_1 _3924_ (.A(_1000_),
    .B(_1009_),
    .Y(_0216_));
 sg13g2_o21ai_1 _3925_ (.B1(net612),
    .Y(_1010_),
    .A1(_2048_),
    .A2(_1008_));
 sg13g2_a21oi_1 _3926_ (.A1(_2048_),
    .A2(_1008_),
    .Y(_0217_),
    .B1(_1010_));
 sg13g2_o21ai_1 _3927_ (.B1(net614),
    .Y(_1011_),
    .A1(net576),
    .A2(_0426_));
 sg13g2_nand3_1 _3928_ (.B(_0426_),
    .C(_1006_),
    .A(net576),
    .Y(_1012_));
 sg13g2_o21ai_1 _3929_ (.B1(_1012_),
    .Y(_1013_),
    .A1(net576),
    .A2(_1006_));
 sg13g2_nor2_1 _3930_ (.A(_1011_),
    .B(_1013_),
    .Y(_0218_));
 sg13g2_and2_1 _3931_ (.A(net684),
    .B(net609),
    .X(_0219_));
 sg13g2_and2_1 _3932_ (.A(net628),
    .B(net609),
    .X(_0220_));
 sg13g2_and2_1 _3933_ (.A(net427),
    .B(net610),
    .X(_0221_));
 sg13g2_nor2_1 _3934_ (.A(_2022_),
    .B(net596),
    .Y(_0222_));
 sg13g2_and2_1 _3935_ (.A(net595),
    .B(net614),
    .X(_0223_));
 sg13g2_and2_1 _3936_ (.A(net588),
    .B(net614),
    .X(_0226_));
 sg13g2_nor2_1 _3937_ (.A(net606),
    .B(_2120_),
    .Y(_0227_));
 sg13g2_nor2b_1 _3938_ (.A(_1000_),
    .B_N(_0423_),
    .Y(_0228_));
 sg13g2_and2_1 _3939_ (.A(net621),
    .B(_0424_),
    .X(_0229_));
 sg13g2_a21oi_1 _3940_ (.A1(net691),
    .A2(_0426_),
    .Y(_0230_),
    .B1(_1011_));
 sg13g2_and2_1 _3941_ (.A(net410),
    .B(net610),
    .X(_0231_));
 sg13g2_and2_1 _3942_ (.A(net413),
    .B(net610),
    .X(_0232_));
 sg13g2_nor2_1 _3943_ (.A(_2023_),
    .B(net596),
    .Y(_0233_));
 sg13g2_and2_1 _3944_ (.A(net435),
    .B(net610),
    .X(_0234_));
 sg13g2_nor2b_1 _3945_ (.A(net557),
    .B_N(net833),
    .Y(_1014_));
 sg13g2_xnor2_1 _3946_ (.Y(_1015_),
    .A(net794),
    .B(net557));
 sg13g2_nor2_1 _3947_ (.A(net596),
    .B(_1015_),
    .Y(_0235_));
 sg13g2_nand2b_1 _3948_ (.Y(_1016_),
    .B(\dino_inst.i_ypos[1] ),
    .A_N(net556));
 sg13g2_xnor2_1 _3949_ (.Y(_1017_),
    .A(\dino_inst.i_ypos[1] ),
    .B(net556));
 sg13g2_and2_1 _3950_ (.A(_1014_),
    .B(_1017_),
    .X(_1018_));
 sg13g2_nor2_1 _3951_ (.A(_1014_),
    .B(_1017_),
    .Y(_1019_));
 sg13g2_nor3_1 _3952_ (.A(net597),
    .B(_1018_),
    .C(_1019_),
    .Y(_0236_));
 sg13g2_nor2b_1 _3953_ (.A(net554),
    .B_N(net756),
    .Y(_1020_));
 sg13g2_xnor2_1 _3954_ (.Y(_1021_),
    .A(\dino_inst.i_ypos[2] ),
    .B(net554));
 sg13g2_a21oi_1 _3955_ (.A1(\dino_inst.i_ypos[1] ),
    .A2(_2041_),
    .Y(_1022_),
    .B1(_1021_));
 sg13g2_xnor2_1 _3956_ (.Y(_1023_),
    .A(_1016_),
    .B(_1021_));
 sg13g2_o21ai_1 _3957_ (.B1(net607),
    .Y(_1024_),
    .A1(_1019_),
    .A2(_1023_));
 sg13g2_a21oi_1 _3958_ (.A1(_1019_),
    .A2(_1023_),
    .Y(_0237_),
    .B1(_1024_));
 sg13g2_a21oi_1 _3959_ (.A1(_1019_),
    .A2(_1023_),
    .Y(_1025_),
    .B1(_1022_));
 sg13g2_nand2b_1 _3960_ (.Y(_1026_),
    .B(\dino_inst.i_ypos[3] ),
    .A_N(net553));
 sg13g2_xnor2_1 _3961_ (.Y(_1027_),
    .A(\dino_inst.i_ypos[3] ),
    .B(net553));
 sg13g2_or2_1 _3962_ (.X(_1028_),
    .B(_1027_),
    .A(_1020_));
 sg13g2_xnor2_1 _3963_ (.Y(_1029_),
    .A(_1020_),
    .B(_1027_));
 sg13g2_or2_1 _3964_ (.X(_1030_),
    .B(_1029_),
    .A(_1025_));
 sg13g2_nand2_1 _3965_ (.Y(_1031_),
    .A(net608),
    .B(_1030_));
 sg13g2_a21oi_1 _3966_ (.A1(_1025_),
    .A2(_1029_),
    .Y(_0238_),
    .B1(_1031_));
 sg13g2_nor2_1 _3967_ (.A(\dino_inst.i_ypos[4] ),
    .B(_2043_),
    .Y(_1032_));
 sg13g2_xnor2_1 _3968_ (.Y(_1033_),
    .A(\dino_inst.i_ypos[4] ),
    .B(net551));
 sg13g2_nand2_1 _3969_ (.Y(_1034_),
    .A(_1026_),
    .B(_1033_));
 sg13g2_xnor2_1 _3970_ (.Y(_1035_),
    .A(_1026_),
    .B(_1033_));
 sg13g2_nand3_1 _3971_ (.B(_1030_),
    .C(_1035_),
    .A(_1028_),
    .Y(_1036_));
 sg13g2_a21o_1 _3972_ (.A2(_1030_),
    .A1(_1028_),
    .B1(_1035_),
    .X(_1037_));
 sg13g2_and3_1 _3973_ (.X(_0239_),
    .A(net608),
    .B(_1036_),
    .C(_1037_));
 sg13g2_and2_1 _3974_ (.A(_1034_),
    .B(_1037_),
    .X(_1038_));
 sg13g2_nor2b_1 _3975_ (.A(net575),
    .B_N(net550),
    .Y(_1039_));
 sg13g2_xnor2_1 _3976_ (.Y(_1040_),
    .A(net912),
    .B(net550));
 sg13g2_nand2_1 _3977_ (.Y(_1041_),
    .A(_1032_),
    .B(_1040_));
 sg13g2_xnor2_1 _3978_ (.Y(_1042_),
    .A(_1032_),
    .B(_1040_));
 sg13g2_or2_1 _3979_ (.X(_1043_),
    .B(_1042_),
    .A(_1038_));
 sg13g2_nand2_1 _3980_ (.Y(_1044_),
    .A(net607),
    .B(_1043_));
 sg13g2_a21oi_1 _3981_ (.A1(_1038_),
    .A2(_1042_),
    .Y(_0240_),
    .B1(_1044_));
 sg13g2_nor2_1 _3982_ (.A(net575),
    .B(net550),
    .Y(_1045_));
 sg13g2_xnor2_1 _3983_ (.Y(_1046_),
    .A(_2044_),
    .B(_1045_));
 sg13g2_and3_1 _3984_ (.X(_1047_),
    .A(_1041_),
    .B(_1043_),
    .C(_1046_));
 sg13g2_a21oi_1 _3985_ (.A1(_1041_),
    .A2(_1043_),
    .Y(_1048_),
    .B1(_1046_));
 sg13g2_nor3_1 _3986_ (.A(net597),
    .B(_1047_),
    .C(_1048_),
    .Y(_0241_));
 sg13g2_a21oi_1 _3987_ (.A1(net882),
    .A2(_1039_),
    .Y(_1049_),
    .B1(_1048_));
 sg13g2_xnor2_1 _3988_ (.Y(_1050_),
    .A(\bg_line_inst.i_vpos[8] ),
    .B(net900));
 sg13g2_nor2_1 _3989_ (.A(net575),
    .B(net859),
    .Y(_1051_));
 sg13g2_a21oi_1 _3990_ (.A1(net575),
    .A2(_1050_),
    .Y(_1052_),
    .B1(_1051_));
 sg13g2_o21ai_1 _3991_ (.B1(net608),
    .Y(_1053_),
    .A1(_1049_),
    .A2(_1052_));
 sg13g2_a21oi_1 _3992_ (.A1(_1049_),
    .A2(_1052_),
    .Y(_0242_),
    .B1(_1053_));
 sg13g2_nand2b_1 _3993_ (.Y(_1054_),
    .B(net824),
    .A_N(\bg_render_inst.i_hpos[2] ));
 sg13g2_nand2_1 _3994_ (.Y(_1055_),
    .A(_2029_),
    .B(net881));
 sg13g2_a21oi_1 _3995_ (.A1(_1054_),
    .A2(_1055_),
    .Y(_0243_),
    .B1(net604));
 sg13g2_nor2b_1 _3996_ (.A(net869),
    .B_N(net594),
    .Y(_1056_));
 sg13g2_nand2b_1 _3997_ (.Y(_1057_),
    .B(net593),
    .A_N(\bg_object_inst.bg_object_pos[3] ));
 sg13g2_nand2b_1 _3998_ (.Y(_1058_),
    .B(net899),
    .A_N(net593));
 sg13g2_and2_1 _3999_ (.A(_1057_),
    .B(_1058_),
    .X(_1059_));
 sg13g2_nor2_1 _4000_ (.A(_1054_),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_nand2_1 _4001_ (.Y(_1061_),
    .A(_1054_),
    .B(_1059_));
 sg13g2_nand2_1 _4002_ (.Y(_1062_),
    .A(net618),
    .B(_1061_));
 sg13g2_nor2_1 _4003_ (.A(_1060_),
    .B(_1062_),
    .Y(_0244_));
 sg13g2_nand2b_1 _4004_ (.Y(_1063_),
    .B(net591),
    .A_N(\bg_object_inst.bg_object_pos[4] ));
 sg13g2_xnor2_1 _4005_ (.Y(_1064_),
    .A(\bg_object_inst.bg_object_pos[4] ),
    .B(net591));
 sg13g2_nand2_1 _4006_ (.Y(_1065_),
    .A(_1056_),
    .B(_1064_));
 sg13g2_xnor2_1 _4007_ (.Y(_1066_),
    .A(_1056_),
    .B(_1064_));
 sg13g2_nand4_1 _4008_ (.B(_1057_),
    .C(_1058_),
    .A(_1054_),
    .Y(_1067_),
    .D(_1064_));
 sg13g2_nand2_1 _4009_ (.Y(_1068_),
    .A(net618),
    .B(_1067_));
 sg13g2_a21oi_1 _4010_ (.A1(_1061_),
    .A2(_1066_),
    .Y(_0245_),
    .B1(_1068_));
 sg13g2_nand2b_1 _4011_ (.Y(_1069_),
    .B(\bg_object_inst.bg_object_pos[5] ),
    .A_N(\bg_render_inst.i_hpos[5] ));
 sg13g2_xnor2_1 _4012_ (.Y(_1070_),
    .A(\bg_object_inst.bg_object_pos[5] ),
    .B(net589));
 sg13g2_nor2_1 _4013_ (.A(_1063_),
    .B(_1070_),
    .Y(_1071_));
 sg13g2_xnor2_1 _4014_ (.Y(_1072_),
    .A(_1063_),
    .B(_1070_));
 sg13g2_and3_1 _4015_ (.X(_1073_),
    .A(_1065_),
    .B(_1067_),
    .C(_1072_));
 sg13g2_a21oi_1 _4016_ (.A1(_1065_),
    .A2(_1067_),
    .Y(_1074_),
    .B1(_1072_));
 sg13g2_nor3_1 _4017_ (.A(net604),
    .B(_1073_),
    .C(_1074_),
    .Y(_0246_));
 sg13g2_nor2b_1 _4018_ (.A(\bg_object_inst.bg_object_pos[6] ),
    .B_N(net586),
    .Y(_1075_));
 sg13g2_xnor2_1 _4019_ (.Y(_1076_),
    .A(\bg_object_inst.bg_object_pos[6] ),
    .B(net586));
 sg13g2_nand2_1 _4020_ (.Y(_1077_),
    .A(_1069_),
    .B(_1076_));
 sg13g2_xor2_1 _4021_ (.B(_1076_),
    .A(_1069_),
    .X(_1078_));
 sg13g2_nor3_1 _4022_ (.A(_1071_),
    .B(_1074_),
    .C(_1078_),
    .Y(_1079_));
 sg13g2_o21ai_1 _4023_ (.B1(_1078_),
    .Y(_1080_),
    .A1(_1071_),
    .A2(_1074_));
 sg13g2_nand2_1 _4024_ (.Y(_1081_),
    .A(net620),
    .B(_1080_));
 sg13g2_nor2_1 _4025_ (.A(_1079_),
    .B(_1081_),
    .Y(_0247_));
 sg13g2_and2_1 _4026_ (.A(_1077_),
    .B(_1080_),
    .X(_1082_));
 sg13g2_nor2_1 _4027_ (.A(\bg_object_inst.bg_object_pos[7] ),
    .B(_2047_),
    .Y(_1083_));
 sg13g2_xnor2_1 _4028_ (.Y(_1084_),
    .A(\bg_object_inst.bg_object_pos[7] ),
    .B(net583));
 sg13g2_nand2_1 _4029_ (.Y(_1085_),
    .A(_1075_),
    .B(_1084_));
 sg13g2_xnor2_1 _4030_ (.Y(_1086_),
    .A(_1075_),
    .B(_1084_));
 sg13g2_or2_1 _4031_ (.X(_1087_),
    .B(_1086_),
    .A(_1082_));
 sg13g2_nand2_1 _4032_ (.Y(_1088_),
    .A(net620),
    .B(_1087_));
 sg13g2_a21oi_1 _4033_ (.A1(_1082_),
    .A2(_1086_),
    .Y(_0248_),
    .B1(_1088_));
 sg13g2_and2_1 _4034_ (.A(_1085_),
    .B(_1087_),
    .X(_1089_));
 sg13g2_nand2b_1 _4035_ (.Y(_1090_),
    .B(net580),
    .A_N(\bg_object_inst.bg_object_pos[8] ));
 sg13g2_xnor2_1 _4036_ (.Y(_1091_),
    .A(\bg_object_inst.bg_object_pos[8] ),
    .B(net580));
 sg13g2_nand2_1 _4037_ (.Y(_1092_),
    .A(_1083_),
    .B(_1091_));
 sg13g2_xnor2_1 _4038_ (.Y(_1093_),
    .A(_1083_),
    .B(_1091_));
 sg13g2_or2_1 _4039_ (.X(_1094_),
    .B(_1093_),
    .A(_1089_));
 sg13g2_nand2_1 _4040_ (.Y(_1095_),
    .A(net620),
    .B(_1094_));
 sg13g2_a21oi_1 _4041_ (.A1(_1089_),
    .A2(_1093_),
    .Y(_0249_),
    .B1(_1095_));
 sg13g2_xor2_1 _4042_ (.B(\bg_render_inst.i_hpos[9] ),
    .A(\bg_object_inst.bg_object_pos[9] ),
    .X(_1096_));
 sg13g2_xnor2_1 _4043_ (.Y(_1097_),
    .A(_1090_),
    .B(_1096_));
 sg13g2_a21oi_1 _4044_ (.A1(_1092_),
    .A2(_1094_),
    .Y(_1098_),
    .B1(_1097_));
 sg13g2_and3_1 _4045_ (.X(_1099_),
    .A(_1092_),
    .B(_1094_),
    .C(_1097_));
 sg13g2_nor3_1 _4046_ (.A(net603),
    .B(_1098_),
    .C(_1099_),
    .Y(_0250_));
 sg13g2_and2_1 _4047_ (.A(net432),
    .B(net621),
    .X(_0251_));
 sg13g2_and2_1 _4048_ (.A(net621),
    .B(net397),
    .X(_0252_));
 sg13g2_nor2_1 _4049_ (.A(net555),
    .B(net554),
    .Y(_1100_));
 sg13g2_xor2_1 _4050_ (.B(net816),
    .A(net555),
    .X(_1101_));
 sg13g2_nor2_1 _4051_ (.A(net602),
    .B(_1101_),
    .Y(_0253_));
 sg13g2_o21ai_1 _4052_ (.B1(net618),
    .Y(_1102_),
    .A1(net759),
    .A2(_1100_));
 sg13g2_a21oi_1 _4053_ (.A1(net759),
    .A2(_1100_),
    .Y(_0254_),
    .B1(_1102_));
 sg13g2_o21ai_1 _4054_ (.B1(net553),
    .Y(_1103_),
    .A1(net555),
    .A2(net554));
 sg13g2_o21ai_1 _4055_ (.B1(net618),
    .Y(_1104_),
    .A1(_2121_),
    .A2(_1103_));
 sg13g2_a21oi_1 _4056_ (.A1(_2121_),
    .A2(_1103_),
    .Y(_0255_),
    .B1(_1104_));
 sg13g2_o21ai_1 _4057_ (.B1(net855),
    .Y(_1105_),
    .A1(net551),
    .A2(_1103_));
 sg13g2_nor2_1 _4058_ (.A(net549),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_and2_1 _4059_ (.A(net549),
    .B(_1105_),
    .X(_1107_));
 sg13g2_nor3_1 _4060_ (.A(net601),
    .B(_1106_),
    .C(_1107_),
    .Y(_0256_));
 sg13g2_o21ai_1 _4061_ (.B1(net619),
    .Y(_1108_),
    .A1(net717),
    .A2(_1107_));
 sg13g2_a21oi_1 _4062_ (.A1(net717),
    .A2(_1107_),
    .Y(_0257_),
    .B1(_1108_));
 sg13g2_a21oi_1 _4063_ (.A1(_2044_),
    .A2(_1107_),
    .Y(_1109_),
    .B1(_2122_));
 sg13g2_xnor2_1 _4064_ (.Y(_1110_),
    .A(_2045_),
    .B(_1109_));
 sg13g2_and2_1 _4065_ (.A(net619),
    .B(_1110_),
    .X(_0258_));
 sg13g2_xor2_1 _4066_ (.B(net735),
    .A(net404),
    .X(_1111_));
 sg13g2_nand2_1 _4067_ (.Y(_0259_),
    .A(net626),
    .B(_1111_));
 sg13g2_and2_1 _4068_ (.A(net423),
    .B(net625),
    .X(_0260_));
 sg13g2_nand2b_1 _4069_ (.Y(_0261_),
    .B(net625),
    .A_N(net857));
 sg13g2_and2_1 _4070_ (.A(net760),
    .B(net625),
    .X(_0262_));
 sg13g2_nand2b_1 _4071_ (.Y(_0263_),
    .B(net625),
    .A_N(net813));
 sg13g2_and2_1 _4072_ (.A(net784),
    .B(net625),
    .X(_0264_));
 sg13g2_nand2b_1 _4073_ (.Y(_0265_),
    .B(net625),
    .A_N(net713));
 sg13g2_and2_1 _4074_ (.A(net736),
    .B(net625),
    .X(_0266_));
 sg13g2_nand2b_1 _4075_ (.Y(_0267_),
    .B(net626),
    .A_N(net747));
 sg13g2_and2_1 _4076_ (.A(net626),
    .B(net401),
    .X(_0268_));
 sg13g2_nand2b_1 _4077_ (.Y(_0269_),
    .B(net626),
    .A_N(net414));
 sg13g2_and2_1 _4078_ (.A(net626),
    .B(net391),
    .X(_0270_));
 sg13g2_nand2b_1 _4079_ (.Y(_0271_),
    .B(net626),
    .A_N(net417));
 sg13g2_and2_1 _4080_ (.A(net626),
    .B(net400),
    .X(_0272_));
 sg13g2_nand2b_1 _4081_ (.Y(_0273_),
    .B(net625),
    .A_N(net404));
 sg13g2_nand2b_1 _4082_ (.Y(_1112_),
    .B(net896),
    .A_N(net595));
 sg13g2_nand2b_1 _4083_ (.Y(_1113_),
    .B(net595),
    .A_N(net896));
 sg13g2_a21oi_1 _4084_ (.A1(_1112_),
    .A2(_1113_),
    .Y(_0274_),
    .B1(net605));
 sg13g2_nor2b_1 _4085_ (.A(\ai_controller_inst.obstacle1_pos[3] ),
    .B_N(net593),
    .Y(_1114_));
 sg13g2_nand2b_1 _4086_ (.Y(_1115_),
    .B(net593),
    .A_N(\ai_controller_inst.obstacle1_pos[3] ));
 sg13g2_nand2b_1 _4087_ (.Y(_1116_),
    .B(\ai_controller_inst.obstacle1_pos[3] ),
    .A_N(net593));
 sg13g2_and2_1 _4088_ (.A(_1115_),
    .B(_1116_),
    .X(_1117_));
 sg13g2_nor2_1 _4089_ (.A(_1112_),
    .B(_1117_),
    .Y(_1118_));
 sg13g2_nand2_1 _4090_ (.Y(_1119_),
    .A(_1112_),
    .B(_1117_));
 sg13g2_nand2_1 _4091_ (.Y(_1120_),
    .A(net622),
    .B(_1119_));
 sg13g2_nor2_1 _4092_ (.A(_1118_),
    .B(_1120_),
    .Y(_0275_));
 sg13g2_nor2_1 _4093_ (.A(\ai_controller_inst.obstacle1_pos[4] ),
    .B(_2046_),
    .Y(_1121_));
 sg13g2_xnor2_1 _4094_ (.Y(_1122_),
    .A(\ai_controller_inst.obstacle1_pos[4] ),
    .B(net591));
 sg13g2_nand2_1 _4095_ (.Y(_1123_),
    .A(_1114_),
    .B(_1122_));
 sg13g2_xnor2_1 _4096_ (.Y(_1124_),
    .A(_1114_),
    .B(_1122_));
 sg13g2_nand4_1 _4097_ (.B(_1115_),
    .C(_1116_),
    .A(_1112_),
    .Y(_1125_),
    .D(_1122_));
 sg13g2_nand2_1 _4098_ (.Y(_1126_),
    .A(net622),
    .B(_1125_));
 sg13g2_a21oi_1 _4099_ (.A1(_1119_),
    .A2(_1124_),
    .Y(_0276_),
    .B1(_1126_));
 sg13g2_nand2_1 _4100_ (.Y(_1127_),
    .A(_2031_),
    .B(net589));
 sg13g2_xnor2_1 _4101_ (.Y(_1128_),
    .A(\ai_controller_inst.obstacle1_pos[5] ),
    .B(net589));
 sg13g2_and2_1 _4102_ (.A(_1121_),
    .B(_1128_),
    .X(_1129_));
 sg13g2_xnor2_1 _4103_ (.Y(_1130_),
    .A(_1121_),
    .B(_1128_));
 sg13g2_and3_1 _4104_ (.X(_1131_),
    .A(_1123_),
    .B(_1125_),
    .C(_1130_));
 sg13g2_a21oi_1 _4105_ (.A1(_1123_),
    .A2(_1125_),
    .Y(_1132_),
    .B1(_1130_));
 sg13g2_nor3_1 _4106_ (.A(net605),
    .B(_1131_),
    .C(_1132_),
    .Y(_0277_));
 sg13g2_nand2b_1 _4107_ (.Y(_1133_),
    .B(\ai_controller_inst.obstacle1_pos[6] ),
    .A_N(net586));
 sg13g2_xnor2_1 _4108_ (.Y(_1134_),
    .A(\ai_controller_inst.obstacle1_pos[6] ),
    .B(net586));
 sg13g2_nor2_1 _4109_ (.A(_1127_),
    .B(_1134_),
    .Y(_1135_));
 sg13g2_xor2_1 _4110_ (.B(_1134_),
    .A(_1127_),
    .X(_1136_));
 sg13g2_nor3_1 _4111_ (.A(_1129_),
    .B(_1132_),
    .C(_1136_),
    .Y(_1137_));
 sg13g2_o21ai_1 _4112_ (.B1(_1136_),
    .Y(_1138_),
    .A1(_1129_),
    .A2(_1132_));
 sg13g2_nand2_1 _4113_ (.Y(_1139_),
    .A(net622),
    .B(_1138_));
 sg13g2_nor2_1 _4114_ (.A(_1137_),
    .B(_1139_),
    .Y(_0278_));
 sg13g2_nor2b_1 _4115_ (.A(_1135_),
    .B_N(_1138_),
    .Y(_1140_));
 sg13g2_nor2_1 _4116_ (.A(\ai_controller_inst.obstacle1_pos[7] ),
    .B(_2047_),
    .Y(_1141_));
 sg13g2_xnor2_1 _4117_ (.Y(_1142_),
    .A(\ai_controller_inst.obstacle1_pos[7] ),
    .B(net583));
 sg13g2_nand2_1 _4118_ (.Y(_1143_),
    .A(_1133_),
    .B(_1142_));
 sg13g2_xnor2_1 _4119_ (.Y(_1144_),
    .A(_1133_),
    .B(_1142_));
 sg13g2_or2_1 _4120_ (.X(_1145_),
    .B(_1144_),
    .A(_1140_));
 sg13g2_nand2_1 _4121_ (.Y(_1146_),
    .A(net622),
    .B(_1145_));
 sg13g2_a21oi_1 _4122_ (.A1(_1140_),
    .A2(_1144_),
    .Y(_0279_),
    .B1(_1146_));
 sg13g2_and2_1 _4123_ (.A(_1143_),
    .B(_1145_),
    .X(_1147_));
 sg13g2_nand2b_1 _4124_ (.Y(_1148_),
    .B(net580),
    .A_N(\ai_controller_inst.obstacle1_pos[8] ));
 sg13g2_xnor2_1 _4125_ (.Y(_1149_),
    .A(\ai_controller_inst.obstacle1_pos[8] ),
    .B(net580));
 sg13g2_nand2_1 _4126_ (.Y(_1150_),
    .A(_1141_),
    .B(_1149_));
 sg13g2_xnor2_1 _4127_ (.Y(_1151_),
    .A(_1141_),
    .B(_1149_));
 sg13g2_or2_1 _4128_ (.X(_1152_),
    .B(_1151_),
    .A(_1147_));
 sg13g2_nand2_1 _4129_ (.Y(_1153_),
    .A(net622),
    .B(_1152_));
 sg13g2_a21oi_1 _4130_ (.A1(_1147_),
    .A2(_1151_),
    .Y(_0280_),
    .B1(_1153_));
 sg13g2_xor2_1 _4131_ (.B(\bg_render_inst.i_hpos[9] ),
    .A(\ai_controller_inst.obstacle1_pos[9] ),
    .X(_1154_));
 sg13g2_xnor2_1 _4132_ (.Y(_1155_),
    .A(_1148_),
    .B(_1154_));
 sg13g2_a21oi_1 _4133_ (.A1(_1150_),
    .A2(_1152_),
    .Y(_1156_),
    .B1(_1155_));
 sg13g2_and3_1 _4134_ (.X(_1157_),
    .A(_1150_),
    .B(_1152_),
    .C(_1155_));
 sg13g2_nor3_1 _4135_ (.A(net605),
    .B(_1156_),
    .C(_1157_),
    .Y(_0281_));
 sg13g2_and2_1 _4136_ (.A(net617),
    .B(net396),
    .X(_0282_));
 sg13g2_o21ai_1 _4137_ (.B1(net617),
    .Y(_1158_),
    .A1(net555),
    .A2(net557));
 sg13g2_nor2_1 _4138_ (.A(_0973_),
    .B(_1158_),
    .Y(_0283_));
 sg13g2_nor2_1 _4139_ (.A(net557),
    .B(net816),
    .Y(_1159_));
 sg13g2_nor4_1 _4140_ (.A(net600),
    .B(_0975_),
    .C(_1100_),
    .D(_1159_),
    .Y(_0284_));
 sg13g2_nand2_2 _4141_ (.Y(_1160_),
    .A(net553),
    .B(_0975_));
 sg13g2_o21ai_1 _4142_ (.B1(net617),
    .Y(_1161_),
    .A1(net552),
    .A2(_0975_));
 sg13g2_nor2b_1 _4143_ (.A(_1161_),
    .B_N(_1160_),
    .Y(_0285_));
 sg13g2_xnor2_1 _4144_ (.Y(_1162_),
    .A(_2121_),
    .B(_1160_));
 sg13g2_nor2_1 _4145_ (.A(net601),
    .B(_1162_),
    .Y(_0286_));
 sg13g2_a21oi_1 _4146_ (.A1(net855),
    .A2(_1160_),
    .Y(_1163_),
    .B1(net549));
 sg13g2_and3_1 _4147_ (.X(_1164_),
    .A(net549),
    .B(net855),
    .C(_1160_));
 sg13g2_nor3_1 _4148_ (.A(net601),
    .B(_1163_),
    .C(_1164_),
    .Y(_0287_));
 sg13g2_nand3_1 _4149_ (.B(_2131_),
    .C(_1160_),
    .A(_2044_),
    .Y(_1165_));
 sg13g2_a21o_1 _4150_ (.A2(_1160_),
    .A1(_2131_),
    .B1(_2044_),
    .X(_1166_));
 sg13g2_a21oi_1 _4151_ (.A1(_1165_),
    .A2(_1166_),
    .Y(_0288_),
    .B1(net601));
 sg13g2_o21ai_1 _4152_ (.B1(net618),
    .Y(_1167_),
    .A1(_2045_),
    .A2(_1165_));
 sg13g2_a21oi_1 _4153_ (.A1(_2045_),
    .A2(_1165_),
    .Y(_0289_),
    .B1(_1167_));
 sg13g2_nand2_1 _4154_ (.Y(_1168_),
    .A(\graphics_inst.hvsync_gen.vpos[0] ),
    .B(_0406_));
 sg13g2_nor4_1 _4155_ (.A(\graphics_inst.hvsync_gen.vpos[0] ),
    .B(\graphics_inst.hvsync_gen.vpos[1] ),
    .C(\bg_line_inst.i_vpos[8] ),
    .D(_2045_),
    .Y(_1169_));
 sg13g2_nand3_1 _4156_ (.B(_0973_),
    .C(_1169_),
    .A(_2132_),
    .Y(_1170_));
 sg13g2_nand2_1 _4157_ (.Y(_1171_),
    .A(net617),
    .B(_1170_));
 sg13g2_or2_1 _4158_ (.X(_1172_),
    .B(_1171_),
    .A(_0405_));
 sg13g2_o21ai_1 _4159_ (.B1(_1168_),
    .Y(_0290_),
    .A1(_2027_),
    .A2(_1172_));
 sg13g2_nand2_1 _4160_ (.Y(_1173_),
    .A(net781),
    .B(_0406_));
 sg13g2_xnor2_1 _4161_ (.Y(_1174_),
    .A(net672),
    .B(net781));
 sg13g2_o21ai_1 _4162_ (.B1(_1173_),
    .Y(_0291_),
    .A1(_1172_),
    .A2(_1174_));
 sg13g2_o21ai_1 _4163_ (.B1(net617),
    .Y(_1175_),
    .A1(_0405_),
    .A2(_1170_));
 sg13g2_nand3_1 _4164_ (.B(\graphics_inst.hvsync_gen.vpos[1] ),
    .C(_0407_),
    .A(\graphics_inst.hvsync_gen.vpos[0] ),
    .Y(_1176_));
 sg13g2_inv_1 _4165_ (.Y(_1177_),
    .A(_1176_));
 sg13g2_xor2_1 _4166_ (.B(_1176_),
    .A(net557),
    .X(_1178_));
 sg13g2_nor2_1 _4167_ (.A(_1175_),
    .B(_1178_),
    .Y(_0292_));
 sg13g2_nor2_1 _4168_ (.A(net396),
    .B(_1176_),
    .Y(_1179_));
 sg13g2_xnor2_1 _4169_ (.Y(_1180_),
    .A(net555),
    .B(_1179_));
 sg13g2_nor2_1 _4170_ (.A(_1175_),
    .B(_1180_),
    .Y(_0293_));
 sg13g2_a21oi_1 _4171_ (.A1(_0973_),
    .A2(_1177_),
    .Y(_1181_),
    .B1(net554));
 sg13g2_nor2_2 _4172_ (.A(_0976_),
    .B(_1176_),
    .Y(_1182_));
 sg13g2_nor3_1 _4173_ (.A(_1175_),
    .B(_1181_),
    .C(_1182_),
    .Y(_0294_));
 sg13g2_nand2_1 _4174_ (.Y(_1183_),
    .A(net552),
    .B(_1182_));
 sg13g2_nand2b_1 _4175_ (.Y(_1184_),
    .B(_1183_),
    .A_N(_1175_));
 sg13g2_nor2_1 _4176_ (.A(net552),
    .B(_1182_),
    .Y(_1185_));
 sg13g2_nor2_1 _4177_ (.A(_1184_),
    .B(_1185_),
    .Y(_0295_));
 sg13g2_nand3_1 _4178_ (.B(net617),
    .C(_1170_),
    .A(_2043_),
    .Y(_1186_));
 sg13g2_a22oi_1 _4179_ (.Y(_0296_),
    .B1(_1184_),
    .B2(_1186_),
    .A2(_1183_),
    .A1(_2043_));
 sg13g2_nor2_1 _4180_ (.A(net855),
    .B(_1183_),
    .Y(_1187_));
 sg13g2_xnor2_1 _4181_ (.Y(_1188_),
    .A(net549),
    .B(_1187_));
 sg13g2_nor2_1 _4182_ (.A(_1175_),
    .B(_1188_),
    .Y(_0297_));
 sg13g2_nand4_1 _4183_ (.B(net549),
    .C(net551),
    .A(net552),
    .Y(_1189_),
    .D(_1182_));
 sg13g2_nand3_1 _4184_ (.B(net551),
    .C(\bg_line_inst.i_vpos[8] ),
    .A(net549),
    .Y(_1190_));
 sg13g2_xnor2_1 _4185_ (.Y(_1191_),
    .A(_2044_),
    .B(_1189_));
 sg13g2_nor2_1 _4186_ (.A(_1175_),
    .B(_1191_),
    .Y(_0298_));
 sg13g2_nor2_1 _4187_ (.A(net717),
    .B(_1189_),
    .Y(_1192_));
 sg13g2_xnor2_1 _4188_ (.Y(_1193_),
    .A(net859),
    .B(_1192_));
 sg13g2_nor2_1 _4189_ (.A(_1175_),
    .B(_1193_),
    .Y(_0299_));
 sg13g2_and2_1 _4190_ (.A(net620),
    .B(net409),
    .X(_0300_));
 sg13g2_nand4_1 _4191_ (.B(_2042_),
    .C(net550),
    .A(net552),
    .Y(_1194_),
    .D(net551));
 sg13g2_nand3_1 _4192_ (.B(_2045_),
    .C(_2133_),
    .A(\bg_line_inst.i_vpos[8] ),
    .Y(_1195_));
 sg13g2_nor2_1 _4193_ (.A(net759),
    .B(_1190_),
    .Y(_1196_));
 sg13g2_nand2_1 _4194_ (.Y(_1197_),
    .A(_2045_),
    .B(net617));
 sg13g2_o21ai_1 _4195_ (.B1(_2088_),
    .Y(_1198_),
    .A1(net581),
    .A2(net578));
 sg13g2_o21ai_1 _4196_ (.B1(_1198_),
    .Y(_1199_),
    .A1(_1194_),
    .A2(_1195_));
 sg13g2_nor3_2 _4197_ (.A(_1196_),
    .B(_1197_),
    .C(_1199_),
    .Y(_0301_));
 sg13g2_and2_1 _4198_ (.A(net620),
    .B(net395),
    .X(_0302_));
 sg13g2_and2_1 _4199_ (.A(net620),
    .B(net398),
    .X(_0303_));
 sg13g2_nand3_1 _4200_ (.B(net555),
    .C(_1159_),
    .A(net781),
    .Y(_1200_));
 sg13g2_or2_1 _4201_ (.X(_1201_),
    .B(_1197_),
    .A(_1190_));
 sg13g2_nand2b_1 _4202_ (.Y(_1202_),
    .B(net552),
    .A_N(net895));
 sg13g2_a221oi_1 _4203_ (.B2(net759),
    .C1(_1201_),
    .B1(_1202_),
    .A1(net552),
    .Y(_0304_),
    .A2(_1200_));
 sg13g2_o21ai_1 _4204_ (.B1(_0588_),
    .Y(_1203_),
    .A1(_0416_),
    .A2(_0423_));
 sg13g2_nand3b_1 _4205_ (.B(net577),
    .C(net581),
    .Y(_1204_),
    .A_N(_2128_));
 sg13g2_a221oi_1 _4206_ (.B2(_0404_),
    .C1(net600),
    .B1(_1204_),
    .A1(_2088_),
    .Y(_0305_),
    .A2(_1203_));
 sg13g2_nor2_1 _4207_ (.A(\score_inst_1.y_offset_r[5] ),
    .B(\score_inst_1.y_offset_r[7] ),
    .Y(_1205_));
 sg13g2_nor3_2 _4208_ (.A(\score_inst_1.y_offset_r[6] ),
    .B(\score_inst_1.y_offset_r[9] ),
    .C(\score_inst_1.y_offset_r[8] ),
    .Y(_1206_));
 sg13g2_nand2_2 _4209_ (.Y(_1207_),
    .A(\bg_object_rom_inst.i_rom_counter[4] ),
    .B(\bg_object_rom_inst.i_rom_counter[3] ));
 sg13g2_nand3_1 _4210_ (.B(\bg_object_rom_inst.i_rom_counter[4] ),
    .C(\bg_object_rom_inst.i_rom_counter[3] ),
    .A(net558),
    .Y(_1208_));
 sg13g2_and3_2 _4211_ (.X(_1209_),
    .A(_1205_),
    .B(_1206_),
    .C(_1208_));
 sg13g2_or4_1 _4212_ (.A(\score_inst_2.x_offset_r[7] ),
    .B(\score_inst_2.x_offset_r[6] ),
    .C(\score_inst_2.x_offset_r[9] ),
    .D(\score_inst_2.x_offset_r[8] ),
    .X(_1210_));
 sg13g2_nor3_2 _4213_ (.A(\score_inst_2.x_offset_r[5] ),
    .B(\score_inst_2.x_offset_r[4] ),
    .C(_1210_),
    .Y(_1211_));
 sg13g2_nand3_1 _4214_ (.B(_1205_),
    .C(_1206_),
    .A(_2105_),
    .Y(_1212_));
 sg13g2_nand4_1 _4215_ (.B(_1205_),
    .C(_1206_),
    .A(_2105_),
    .Y(_1213_),
    .D(_1207_));
 sg13g2_nor2_1 _4216_ (.A(\score_inst_2.x_offset_r[3] ),
    .B(\score_inst_2.x_offset_r[2] ),
    .Y(_1214_));
 sg13g2_nand2_1 _4217_ (.Y(_1215_),
    .A(_1211_),
    .B(_1214_));
 sg13g2_or2_1 _4218_ (.X(_1216_),
    .B(\score_inst_2.num_r[2] ),
    .A(\score_inst_2.num_r[1] ));
 sg13g2_nor2_1 _4219_ (.A(\score_inst_2.num_r[0] ),
    .B(\score_inst_2.num_r[2] ),
    .Y(_1217_));
 sg13g2_nor4_1 _4220_ (.A(\score_inst_2.num_r[0] ),
    .B(net508),
    .C(_1215_),
    .D(_1216_),
    .Y(_1218_));
 sg13g2_and2_1 _4221_ (.A(\score_inst_2.x_offset_r[3] ),
    .B(\score_inst_2.x_offset_r[2] ),
    .X(_1219_));
 sg13g2_nand2_1 _4222_ (.Y(_1220_),
    .A(_1211_),
    .B(_1219_));
 sg13g2_nor2_1 _4223_ (.A(\score_inst_2.num_r[1] ),
    .B(\score_inst_2.num_r[0] ),
    .Y(_1221_));
 sg13g2_nor2b_1 _4224_ (.A(_1221_),
    .B_N(\score_inst_2.num_r[2] ),
    .Y(_1222_));
 sg13g2_nand3_1 _4225_ (.B(\score_inst_2.x_offset_r[2] ),
    .C(_1211_),
    .A(\score_inst_2.x_offset_r[3] ),
    .Y(_1223_));
 sg13g2_nor3_1 _4226_ (.A(net508),
    .B(_1222_),
    .C(_1223_),
    .Y(_1224_));
 sg13g2_o21ai_1 _4227_ (.B1(_2108_),
    .Y(_1225_),
    .A1(_1218_),
    .A2(_1224_));
 sg13g2_or2_1 _4228_ (.X(_1226_),
    .B(_1216_),
    .A(_2108_));
 sg13g2_nand2_1 _4229_ (.Y(_1227_),
    .A(\score_inst_2.num_r[2] ),
    .B(_2108_));
 sg13g2_nand2_1 _4230_ (.Y(_1228_),
    .A(\score_inst_2.num_r[1] ),
    .B(\score_inst_2.num_r[0] ));
 sg13g2_o21ai_1 _4231_ (.B1(_1226_),
    .Y(_1229_),
    .A1(_1227_),
    .A2(_1228_));
 sg13g2_nor2_2 _4232_ (.A(\bg_object_rom_inst.i_rom_counter[4] ),
    .B(\bg_object_rom_inst.i_rom_counter[3] ),
    .Y(_1230_));
 sg13g2_nor2b_1 _4233_ (.A(net509),
    .B_N(_1230_),
    .Y(_1231_));
 sg13g2_nand2b_2 _4234_ (.Y(_1232_),
    .B(_1230_),
    .A_N(net509));
 sg13g2_o21ai_1 _4235_ (.B1(_1232_),
    .Y(_1233_),
    .A1(net508),
    .A2(_1220_));
 sg13g2_nand2b_1 _4236_ (.Y(_1234_),
    .B(_1228_),
    .A_N(_1227_));
 sg13g2_nor2_2 _4237_ (.A(_1207_),
    .B(net510),
    .Y(_1235_));
 sg13g2_a221oi_1 _4238_ (.B2(_1234_),
    .C1(net510),
    .B1(_1226_),
    .A1(_1207_),
    .Y(_1236_),
    .A2(_1215_));
 sg13g2_a21oi_1 _4239_ (.A1(_1229_),
    .A2(_1233_),
    .Y(_1237_),
    .B1(_1236_));
 sg13g2_nand2b_1 _4240_ (.Y(_1238_),
    .B(\score_inst_2.num_r[1] ),
    .A_N(\score_inst_2.num_r[3] ));
 sg13g2_a21o_1 _4241_ (.A2(_1238_),
    .A1(_1216_),
    .B1(\score_inst_2.num_r[0] ),
    .X(_1239_));
 sg13g2_o21ai_1 _4242_ (.B1(_1216_),
    .Y(_1240_),
    .A1(\score_inst_2.num_r[3] ),
    .A2(_1217_));
 sg13g2_nand3_1 _4243_ (.B(_1219_),
    .C(_1240_),
    .A(_1211_),
    .Y(_1241_));
 sg13g2_o21ai_1 _4244_ (.B1(_1241_),
    .Y(_1242_),
    .A1(_1215_),
    .A2(_1239_));
 sg13g2_nor2_1 _4245_ (.A(\score_inst_2.num_r[2] ),
    .B(_1238_),
    .Y(_1243_));
 sg13g2_nor2b_1 _4246_ (.A(\bg_object_rom_inst.i_rom_counter[3] ),
    .B_N(\bg_object_rom_inst.i_rom_counter[4] ),
    .Y(_1244_));
 sg13g2_nand2_1 _4247_ (.Y(_1245_),
    .A(\bg_object_rom_inst.i_rom_counter[5] ),
    .B(_1244_));
 sg13g2_nand4_1 _4248_ (.B(_1205_),
    .C(_1206_),
    .A(net558),
    .Y(_1246_),
    .D(_1244_));
 sg13g2_nor3_1 _4249_ (.A(\score_inst_2.num_r[0] ),
    .B(_1226_),
    .C(_1246_),
    .Y(_1247_));
 sg13g2_a21oi_1 _4250_ (.A1(_1235_),
    .A2(_1243_),
    .Y(_1248_),
    .B1(_1247_));
 sg13g2_nand2_2 _4251_ (.Y(_1249_),
    .A(_1232_),
    .B(_1246_));
 sg13g2_a21oi_1 _4252_ (.A1(_2108_),
    .A2(_1217_),
    .Y(_1250_),
    .B1(_1243_));
 sg13g2_o21ai_1 _4253_ (.B1(_1250_),
    .Y(_1251_),
    .A1(_1221_),
    .A2(_1234_));
 sg13g2_a22oi_1 _4254_ (.Y(_1252_),
    .B1(_1249_),
    .B2(_1251_),
    .A2(_1242_),
    .A1(net510));
 sg13g2_nand4_1 _4255_ (.B(_1237_),
    .C(_1248_),
    .A(_1225_),
    .Y(_1253_),
    .D(_1252_));
 sg13g2_nor2_1 _4256_ (.A(\score_inst_1.x_offset_r[5] ),
    .B(\score_inst_1.x_offset_r[4] ),
    .Y(_1254_));
 sg13g2_nor4_2 _4257_ (.A(\score_inst_1.x_offset_r[7] ),
    .B(\score_inst_1.x_offset_r[6] ),
    .C(\score_inst_1.x_offset_r[9] ),
    .Y(_1255_),
    .D(\score_inst_1.x_offset_r[8] ));
 sg13g2_nand2_1 _4258_ (.Y(_1256_),
    .A(_1254_),
    .B(_1255_));
 sg13g2_nor2_1 _4259_ (.A(\score_inst_1.num_r[1] ),
    .B(\score_inst_1.num_r[0] ),
    .Y(_1257_));
 sg13g2_nor2b_1 _4260_ (.A(\score_inst_1.num_r[3] ),
    .B_N(\score_inst_1.num_r[2] ),
    .Y(_1258_));
 sg13g2_nand2b_1 _4261_ (.Y(_1259_),
    .B(\score_inst_1.num_r[2] ),
    .A_N(\score_inst_1.num_r[3] ));
 sg13g2_nand2_1 _4262_ (.Y(_1260_),
    .A(\score_inst_1.num_r[1] ),
    .B(\score_inst_1.num_r[0] ));
 sg13g2_nand2_1 _4263_ (.Y(_1261_),
    .A(_1258_),
    .B(_1260_));
 sg13g2_nor2_1 _4264_ (.A(\score_inst_1.num_r[2] ),
    .B(\score_inst_1.num_r[3] ),
    .Y(_1262_));
 sg13g2_nand2_1 _4265_ (.Y(_1263_),
    .A(\score_inst_1.num_r[1] ),
    .B(_1262_));
 sg13g2_nor3_1 _4266_ (.A(\score_inst_1.num_r[0] ),
    .B(\score_inst_1.num_r[2] ),
    .C(\score_inst_1.num_r[3] ),
    .Y(_1264_));
 sg13g2_o21ai_1 _4267_ (.B1(_1263_),
    .Y(_1265_),
    .A1(_1257_),
    .A2(_1261_));
 sg13g2_o21ai_1 _4268_ (.B1(_1249_),
    .Y(_1266_),
    .A1(_1264_),
    .A2(_1265_));
 sg13g2_nor2_1 _4269_ (.A(_2107_),
    .B(\score_inst_1.num_r[0] ),
    .Y(_1267_));
 sg13g2_nand2b_1 _4270_ (.Y(_1268_),
    .B(\score_inst_1.num_r[1] ),
    .A_N(\score_inst_1.num_r[0] ));
 sg13g2_nor2b_1 _4271_ (.A(\score_inst_1.num_r[2] ),
    .B_N(\score_inst_1.num_r[3] ),
    .Y(_1269_));
 sg13g2_nand2_1 _4272_ (.Y(_1270_),
    .A(_2107_),
    .B(_1269_));
 sg13g2_a221oi_1 _4273_ (.B2(_1257_),
    .C1(_1264_),
    .B1(_1269_),
    .A1(_1258_),
    .Y(_1271_),
    .A2(_1267_));
 sg13g2_nor4_1 _4274_ (.A(net569),
    .B(\score_inst_1.x_offset_r[3] ),
    .C(_1256_),
    .D(_1271_),
    .Y(_1272_));
 sg13g2_nand2_1 _4275_ (.Y(_1273_),
    .A(net569),
    .B(\score_inst_1.x_offset_r[3] ));
 sg13g2_o21ai_1 _4276_ (.B1(_1270_),
    .Y(_1274_),
    .A1(_1259_),
    .A2(_1260_));
 sg13g2_a221oi_1 _4277_ (.B2(_2107_),
    .C1(_1258_),
    .B1(_1269_),
    .A1(_1262_),
    .Y(_1275_),
    .A2(_1268_));
 sg13g2_nor3_1 _4278_ (.A(_1256_),
    .B(_1273_),
    .C(_1275_),
    .Y(_1276_));
 sg13g2_o21ai_1 _4279_ (.B1(net510),
    .Y(_1277_),
    .A1(_1272_),
    .A2(_1276_));
 sg13g2_nor3_1 _4280_ (.A(net508),
    .B(_1256_),
    .C(_1273_),
    .Y(_1278_));
 sg13g2_nor3_1 _4281_ (.A(\score_inst_1.num_r[1] ),
    .B(\score_inst_1.num_r[0] ),
    .C(\score_inst_1.num_r[3] ),
    .Y(_1279_));
 sg13g2_o21ai_1 _4282_ (.B1(_1278_),
    .Y(_1280_),
    .A1(_1262_),
    .A2(_1279_));
 sg13g2_o21ai_1 _4283_ (.B1(_1274_),
    .Y(_1281_),
    .A1(_1231_),
    .A2(_1278_));
 sg13g2_o21ai_1 _4284_ (.B1(_1270_),
    .Y(_1282_),
    .A1(_1259_),
    .A2(_1268_));
 sg13g2_o21ai_1 _4285_ (.B1(_2107_),
    .Y(_1283_),
    .A1(_1258_),
    .A2(_1264_));
 sg13g2_o21ai_1 _4286_ (.B1(_1263_),
    .Y(_1284_),
    .A1(\score_inst_1.num_r[1] ),
    .A2(_1259_));
 sg13g2_nor3_1 _4287_ (.A(\score_inst_1.num_r[0] ),
    .B(_1246_),
    .C(_1270_),
    .Y(_1285_));
 sg13g2_a21oi_1 _4288_ (.A1(_1235_),
    .A2(_1284_),
    .Y(_1286_),
    .B1(_1285_));
 sg13g2_nor4_1 _4289_ (.A(net569),
    .B(\score_inst_1.x_offset_r[3] ),
    .C(net508),
    .D(_1256_),
    .Y(_1287_));
 sg13g2_o21ai_1 _4290_ (.B1(_1282_),
    .Y(_1288_),
    .A1(_1235_),
    .A2(_1287_));
 sg13g2_nand2b_1 _4291_ (.Y(_1289_),
    .B(_1287_),
    .A_N(_1283_));
 sg13g2_and4_1 _4292_ (.A(_1281_),
    .B(_1286_),
    .C(_1288_),
    .D(_1289_),
    .X(_1290_));
 sg13g2_nand4_1 _4293_ (.B(_1277_),
    .C(_1280_),
    .A(_1266_),
    .Y(_1291_),
    .D(_1290_));
 sg13g2_nor2_1 _4294_ (.A(\score_inst_5.x_offset_r[5] ),
    .B(\score_inst_5.x_offset_r[4] ),
    .Y(_1292_));
 sg13g2_nor4_2 _4295_ (.A(\score_inst_5.x_offset_r[7] ),
    .B(\score_inst_5.x_offset_r[6] ),
    .C(\score_inst_5.x_offset_r[9] ),
    .Y(_1293_),
    .D(\score_inst_5.x_offset_r[8] ));
 sg13g2_nand2_1 _4296_ (.Y(_1294_),
    .A(_1292_),
    .B(_1293_));
 sg13g2_nor2_1 _4297_ (.A(\score_inst_5.num_r[1] ),
    .B(\score_inst_5.num_r[0] ),
    .Y(_1295_));
 sg13g2_nor2b_2 _4298_ (.A(\score_inst_5.num_r[3] ),
    .B_N(\score_inst_5.num_r[2] ),
    .Y(_1296_));
 sg13g2_xor2_1 _4299_ (.B(\score_inst_5.num_r[0] ),
    .A(\score_inst_5.num_r[1] ),
    .X(_1297_));
 sg13g2_nor2_1 _4300_ (.A(\score_inst_5.num_r[2] ),
    .B(\score_inst_5.num_r[3] ),
    .Y(_1298_));
 sg13g2_nor3_1 _4301_ (.A(\score_inst_5.num_r[0] ),
    .B(\score_inst_5.num_r[2] ),
    .C(\score_inst_5.num_r[3] ),
    .Y(_1299_));
 sg13g2_a221oi_1 _4302_ (.B2(\score_inst_5.num_r[1] ),
    .C1(_1299_),
    .B1(_1298_),
    .A1(_1296_),
    .Y(_1300_),
    .A2(_1297_));
 sg13g2_a21oi_1 _4303_ (.A1(_1232_),
    .A2(_1246_),
    .Y(_1301_),
    .B1(_1300_));
 sg13g2_nand4_1 _4304_ (.B(\score_inst_1.x_offset_r[3] ),
    .C(_1292_),
    .A(net570),
    .Y(_1302_),
    .D(_1293_));
 sg13g2_nor2b_1 _4305_ (.A(_1295_),
    .B_N(\score_inst_5.num_r[2] ),
    .Y(_1303_));
 sg13g2_or3_1 _4306_ (.A(net570),
    .B(\score_inst_1.x_offset_r[3] ),
    .C(_1294_),
    .X(_1304_));
 sg13g2_o21ai_1 _4307_ (.B1(_2116_),
    .Y(_1305_),
    .A1(_1296_),
    .A2(_1299_));
 sg13g2_nor3_1 _4308_ (.A(net507),
    .B(_1304_),
    .C(_1305_),
    .Y(_1306_));
 sg13g2_nor2b_1 _4309_ (.A(\score_inst_5.num_r[0] ),
    .B_N(\score_inst_5.num_r[1] ),
    .Y(_1307_));
 sg13g2_nand2b_1 _4310_ (.Y(_1308_),
    .B(\score_inst_5.num_r[1] ),
    .A_N(\score_inst_5.num_r[0] ));
 sg13g2_nand2_1 _4311_ (.Y(_1309_),
    .A(_1296_),
    .B(_1307_));
 sg13g2_nor2b_1 _4312_ (.A(\score_inst_5.num_r[2] ),
    .B_N(\score_inst_5.num_r[3] ),
    .Y(_1310_));
 sg13g2_nand2_1 _4313_ (.Y(_1311_),
    .A(_2116_),
    .B(_1310_));
 sg13g2_a221oi_1 _4314_ (.B2(_1311_),
    .C1(net510),
    .B1(_1309_),
    .A1(_1207_),
    .Y(_1312_),
    .A2(_1304_));
 sg13g2_nand3_1 _4315_ (.B(\score_inst_5.num_r[0] ),
    .C(_1296_),
    .A(\score_inst_5.num_r[1] ),
    .Y(_1313_));
 sg13g2_nand2_1 _4316_ (.Y(_1314_),
    .A(_1311_),
    .B(_1313_));
 sg13g2_o21ai_1 _4317_ (.B1(_1232_),
    .Y(_1315_),
    .A1(net507),
    .A2(_1302_));
 sg13g2_a221oi_1 _4318_ (.B2(_1295_),
    .C1(_1299_),
    .B1(_1310_),
    .A1(_1296_),
    .Y(_1316_),
    .A2(_1307_));
 sg13g2_nor4_1 _4319_ (.A(net570),
    .B(\score_inst_1.x_offset_r[3] ),
    .C(_1294_),
    .D(_1316_),
    .Y(_1317_));
 sg13g2_a221oi_1 _4320_ (.B2(_2116_),
    .C1(_1296_),
    .B1(_1310_),
    .A1(_1298_),
    .Y(_1318_),
    .A2(_1308_));
 sg13g2_nor2_1 _4321_ (.A(_1302_),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_o21ai_1 _4322_ (.B1(net509),
    .Y(_1320_),
    .A1(_1317_),
    .A2(_1319_));
 sg13g2_nor3_1 _4323_ (.A(\score_inst_5.num_r[0] ),
    .B(_1246_),
    .C(_1311_),
    .Y(_1321_));
 sg13g2_mux2_1 _4324_ (.A0(_1296_),
    .A1(_1298_),
    .S(\score_inst_5.num_r[1] ),
    .X(_1322_));
 sg13g2_nor4_1 _4325_ (.A(\score_inst_5.num_r[3] ),
    .B(net508),
    .C(_1302_),
    .D(_1303_),
    .Y(_1323_));
 sg13g2_nor4_1 _4326_ (.A(_1301_),
    .B(_1312_),
    .C(_1321_),
    .D(_1323_),
    .Y(_1324_));
 sg13g2_nor2b_1 _4327_ (.A(_1306_),
    .B_N(_1320_),
    .Y(_1325_));
 sg13g2_a22oi_1 _4328_ (.Y(_1326_),
    .B1(_1322_),
    .B2(_1235_),
    .A2(_1315_),
    .A1(_1314_));
 sg13g2_nand3_1 _4329_ (.B(_1325_),
    .C(_1326_),
    .A(_1324_),
    .Y(_1327_));
 sg13g2_or4_1 _4330_ (.A(\score_inst_4.x_offset_r[7] ),
    .B(\score_inst_4.x_offset_r[6] ),
    .C(\score_inst_4.x_offset_r[9] ),
    .D(\score_inst_4.x_offset_r[8] ),
    .X(_1328_));
 sg13g2_nor3_2 _4331_ (.A(\score_inst_4.x_offset_r[5] ),
    .B(\score_inst_4.x_offset_r[4] ),
    .C(_1328_),
    .Y(_1329_));
 sg13g2_nand3_1 _4332_ (.B(\score_inst_4.x_offset_r[3] ),
    .C(_1329_),
    .A(\score_inst_2.x_offset_r[2] ),
    .Y(_1330_));
 sg13g2_o21ai_1 _4333_ (.B1(\score_inst_4.num_r[2] ),
    .Y(_1331_),
    .A1(\score_inst_4.num_r[1] ),
    .A2(\score_inst_4.num_r[0] ));
 sg13g2_inv_1 _4334_ (.Y(_1332_),
    .A(_1331_));
 sg13g2_o21ai_1 _4335_ (.B1(_2113_),
    .Y(_1333_),
    .A1(\score_inst_4.num_r[1] ),
    .A2(_2114_));
 sg13g2_nor2_1 _4336_ (.A(\score_inst_4.num_r[1] ),
    .B(\score_inst_4.num_r[2] ),
    .Y(_1334_));
 sg13g2_xor2_1 _4337_ (.B(\score_inst_4.num_r[2] ),
    .A(\score_inst_4.num_r[1] ),
    .X(_1335_));
 sg13g2_nand2_1 _4338_ (.Y(_1336_),
    .A(\score_inst_4.num_r[0] ),
    .B(_1335_));
 sg13g2_a221oi_1 _4339_ (.B2(_1336_),
    .C1(\score_inst_4.num_r[3] ),
    .B1(_1333_),
    .A1(_1232_),
    .Y(_1337_),
    .A2(_1246_));
 sg13g2_nor4_1 _4340_ (.A(\score_inst_4.num_r[3] ),
    .B(net507),
    .C(_1330_),
    .D(_1332_),
    .Y(_1338_));
 sg13g2_nand2_1 _4341_ (.Y(_1339_),
    .A(\score_inst_4.num_r[3] ),
    .B(_1334_));
 sg13g2_nand3_1 _4342_ (.B(\score_inst_4.num_r[0] ),
    .C(\score_inst_4.num_r[2] ),
    .A(\score_inst_4.num_r[1] ),
    .Y(_1340_));
 sg13g2_o21ai_1 _4343_ (.B1(_1339_),
    .Y(_1341_),
    .A1(\score_inst_4.num_r[3] ),
    .A2(_1340_));
 sg13g2_or2_1 _4344_ (.X(_1342_),
    .B(\score_inst_4.num_r[2] ),
    .A(\score_inst_4.num_r[0] ));
 sg13g2_a21oi_1 _4345_ (.A1(_2115_),
    .A2(_1342_),
    .Y(_1343_),
    .B1(_1334_));
 sg13g2_nor2_1 _4346_ (.A(_1330_),
    .B(_1343_),
    .Y(_1344_));
 sg13g2_nor2_1 _4347_ (.A(\score_inst_2.x_offset_r[2] ),
    .B(\score_inst_4.x_offset_r[3] ),
    .Y(_1345_));
 sg13g2_nand2_1 _4348_ (.Y(_1346_),
    .A(_1329_),
    .B(_1345_));
 sg13g2_and2_1 _4349_ (.A(\score_inst_4.num_r[1] ),
    .B(\score_inst_4.num_r[3] ),
    .X(_1347_));
 sg13g2_nor3_1 _4350_ (.A(_1333_),
    .B(_1346_),
    .C(_1347_),
    .Y(_1348_));
 sg13g2_o21ai_1 _4351_ (.B1(net509),
    .Y(_1349_),
    .A1(_1344_),
    .A2(_1348_));
 sg13g2_nand4_1 _4352_ (.B(_2113_),
    .C(\score_inst_4.num_r[2] ),
    .A(\score_inst_4.num_r[1] ),
    .Y(_1350_),
    .D(_2115_));
 sg13g2_nor2_1 _4353_ (.A(\score_inst_4.num_r[1] ),
    .B(\score_inst_4.num_r[3] ),
    .Y(_1351_));
 sg13g2_o21ai_1 _4354_ (.B1(_1351_),
    .Y(_1352_),
    .A1(_2113_),
    .A2(\score_inst_4.num_r[2] ));
 sg13g2_o21ai_1 _4355_ (.B1(_1232_),
    .Y(_1353_),
    .A1(net507),
    .A2(_1330_));
 sg13g2_nor3_1 _4356_ (.A(\score_inst_4.num_r[3] ),
    .B(_1207_),
    .C(net509),
    .Y(_1354_));
 sg13g2_nor3_1 _4357_ (.A(\score_inst_4.num_r[0] ),
    .B(_1246_),
    .C(_1339_),
    .Y(_1355_));
 sg13g2_a221oi_1 _4358_ (.B2(_1335_),
    .C1(_1355_),
    .B1(_1354_),
    .A1(_1341_),
    .Y(_1356_),
    .A2(_1353_));
 sg13g2_nor3_1 _4359_ (.A(net507),
    .B(_1346_),
    .C(_1352_),
    .Y(_1357_));
 sg13g2_a221oi_1 _4360_ (.B2(_1339_),
    .C1(net509),
    .B1(_1350_),
    .A1(_1207_),
    .Y(_1358_),
    .A2(_1346_));
 sg13g2_nor4_1 _4361_ (.A(_1337_),
    .B(_1338_),
    .C(_1357_),
    .D(_1358_),
    .Y(_1359_));
 sg13g2_nand3_1 _4362_ (.B(_1356_),
    .C(_1359_),
    .A(_1349_),
    .Y(_1360_));
 sg13g2_nor2_1 _4363_ (.A(\dino_inst.o_rom_counter[2] ),
    .B(\score_inst_3.x_offset_r[5] ),
    .Y(_1361_));
 sg13g2_nor4_2 _4364_ (.A(\score_inst_3.x_offset_r[7] ),
    .B(\score_inst_3.x_offset_r[6] ),
    .C(\score_inst_3.x_offset_r[9] ),
    .Y(_1362_),
    .D(\score_inst_3.x_offset_r[8] ));
 sg13g2_nor2_1 _4365_ (.A(\score_inst_3.num_r[2] ),
    .B(\score_inst_3.num_r[3] ),
    .Y(_1363_));
 sg13g2_nor2_2 _4366_ (.A(\dino_inst.o_rom_counter[1] ),
    .B(net569),
    .Y(_1364_));
 sg13g2_nand3_1 _4367_ (.B(_1362_),
    .C(_1364_),
    .A(_1361_),
    .Y(_1365_));
 sg13g2_nor2_1 _4368_ (.A(net507),
    .B(_1365_),
    .Y(_1366_));
 sg13g2_nor2_2 _4369_ (.A(\score_inst_3.num_r[1] ),
    .B(\score_inst_3.num_r[0] ),
    .Y(_1367_));
 sg13g2_a22oi_1 _4370_ (.Y(_1368_),
    .B1(_1366_),
    .B2(_1367_),
    .A2(_1235_),
    .A1(\score_inst_3.num_r[1] ));
 sg13g2_nor2b_1 _4371_ (.A(_1368_),
    .B_N(_1363_),
    .Y(_1369_));
 sg13g2_nand4_1 _4372_ (.B(net570),
    .C(_1361_),
    .A(\dino_inst.o_rom_counter[1] ),
    .Y(_1370_),
    .D(_1362_));
 sg13g2_nor2_1 _4373_ (.A(_2111_),
    .B(_1367_),
    .Y(_1371_));
 sg13g2_nor4_1 _4374_ (.A(\score_inst_3.num_r[3] ),
    .B(net507),
    .C(_1370_),
    .D(_1371_),
    .Y(_1372_));
 sg13g2_nor2_1 _4375_ (.A(_2111_),
    .B(\score_inst_3.num_r[3] ),
    .Y(_1373_));
 sg13g2_o21ai_1 _4376_ (.B1(_1373_),
    .Y(_1374_),
    .A1(_2109_),
    .A2(_2110_));
 sg13g2_o21ai_1 _4377_ (.B1(_1363_),
    .Y(_1375_),
    .A1(\score_inst_3.num_r[1] ),
    .A2(_2110_));
 sg13g2_o21ai_1 _4378_ (.B1(_1375_),
    .Y(_1376_),
    .A1(_1367_),
    .A2(_1374_));
 sg13g2_a21oi_1 _4379_ (.A1(_1249_),
    .A2(_1376_),
    .Y(_1377_),
    .B1(_1372_));
 sg13g2_nor2_1 _4380_ (.A(_2109_),
    .B(\score_inst_3.num_r[0] ),
    .Y(_1378_));
 sg13g2_nand2_1 _4381_ (.Y(_1379_),
    .A(\score_inst_3.num_r[1] ),
    .B(_2110_));
 sg13g2_a22oi_1 _4382_ (.Y(_1380_),
    .B1(_1378_),
    .B2(_2112_),
    .A2(_1367_),
    .A1(_2111_));
 sg13g2_nor2_1 _4383_ (.A(_1365_),
    .B(_1380_),
    .Y(_1381_));
 sg13g2_nor2_1 _4384_ (.A(\score_inst_3.num_r[2] ),
    .B(_2112_),
    .Y(_1382_));
 sg13g2_nand2_1 _4385_ (.Y(_1383_),
    .A(_2109_),
    .B(_1382_));
 sg13g2_nand3_1 _4386_ (.B(\score_inst_3.num_r[0] ),
    .C(_1373_),
    .A(\score_inst_3.num_r[1] ),
    .Y(_1384_));
 sg13g2_nand2_1 _4387_ (.Y(_1385_),
    .A(_1383_),
    .B(_1384_));
 sg13g2_a221oi_1 _4388_ (.B2(_2109_),
    .C1(_1373_),
    .B1(_1382_),
    .A1(_1363_),
    .Y(_1386_),
    .A2(_1379_));
 sg13g2_nor2_1 _4389_ (.A(_1370_),
    .B(_1386_),
    .Y(_1387_));
 sg13g2_o21ai_1 _4390_ (.B1(net509),
    .Y(_1388_),
    .A1(_1381_),
    .A2(_1387_));
 sg13g2_nand3b_1 _4391_ (.B(_1367_),
    .C(_1382_),
    .Y(_1389_),
    .A_N(_1246_));
 sg13g2_o21ai_1 _4392_ (.B1(_1232_),
    .Y(_1390_),
    .A1(net507),
    .A2(_1370_));
 sg13g2_a221oi_1 _4393_ (.B2(_1383_),
    .C1(net509),
    .B1(_1374_),
    .A1(_1207_),
    .Y(_1391_),
    .A2(_1365_));
 sg13g2_a21oi_1 _4394_ (.A1(_1385_),
    .A2(_1390_),
    .Y(_1392_),
    .B1(_1391_));
 sg13g2_nand4_1 _4395_ (.B(_1388_),
    .C(_1389_),
    .A(_1377_),
    .Y(_1393_),
    .D(_1392_));
 sg13g2_nand3_1 _4396_ (.B(_1329_),
    .C(_1360_),
    .A(_1209_),
    .Y(_1394_));
 sg13g2_and3_1 _4397_ (.X(_1395_),
    .A(_1209_),
    .B(_1254_),
    .C(_1255_));
 sg13g2_and2_1 _4398_ (.A(_1209_),
    .B(_1211_),
    .X(_1396_));
 sg13g2_a22oi_1 _4399_ (.Y(_1397_),
    .B1(_1396_),
    .B2(_1253_),
    .A2(_1395_),
    .A1(_1291_));
 sg13g2_and3_1 _4400_ (.X(_1398_),
    .A(_1209_),
    .B(_1361_),
    .C(_1362_));
 sg13g2_o21ai_1 _4401_ (.B1(_1398_),
    .Y(_1399_),
    .A1(_1369_),
    .A2(_1393_));
 sg13g2_nand4_1 _4402_ (.B(_1292_),
    .C(_1293_),
    .A(_1209_),
    .Y(_1400_),
    .D(_1327_));
 sg13g2_and4_2 _4403_ (.A(_1394_),
    .B(_1397_),
    .C(_1399_),
    .D(_1400_),
    .X(_1401_));
 sg13g2_nor2b_1 _4404_ (.A(\obs_rom_inst_2.i_obs_type[2] ),
    .B_N(\obs_rom_inst_2.i_obs_type[1] ),
    .Y(_1402_));
 sg13g2_nand2b_2 _4405_ (.Y(_1403_),
    .B(\obs_rom_inst_2.i_obs_type[1] ),
    .A_N(\obs_rom_inst_2.i_obs_type[2] ));
 sg13g2_and2_1 _4406_ (.A(_0013_),
    .B(_1403_),
    .X(_1404_));
 sg13g2_nand2_1 _4407_ (.Y(_1405_),
    .A(_0013_),
    .B(_1403_));
 sg13g2_nor2b_1 _4408_ (.A(net563),
    .B_N(net561),
    .Y(_1406_));
 sg13g2_nand2b_2 _4409_ (.Y(_1407_),
    .B(net560),
    .A_N(net563));
 sg13g2_nor2_1 _4410_ (.A(_2094_),
    .B(_1407_),
    .Y(_1408_));
 sg13g2_nand3b_1 _4411_ (.B(net564),
    .C(net560),
    .Y(_1409_),
    .A_N(net563));
 sg13g2_and2_1 _4412_ (.A(net564),
    .B(net566),
    .X(_1410_));
 sg13g2_nor2_1 _4413_ (.A(_2095_),
    .B(_1409_),
    .Y(_1411_));
 sg13g2_nand2_2 _4414_ (.Y(_1412_),
    .A(_1406_),
    .B(_1410_));
 sg13g2_a21oi_1 _4415_ (.A1(net506),
    .A2(_1412_),
    .Y(_1413_),
    .B1(net519));
 sg13g2_nand2b_2 _4416_ (.Y(_1414_),
    .B(\obs_rom_inst_2.i_obs_type[1] ),
    .A_N(_0013_));
 sg13g2_nor2_1 _4417_ (.A(net574),
    .B(_1414_),
    .Y(_1415_));
 sg13g2_nand2b_1 _4418_ (.Y(_1416_),
    .B(net563),
    .A_N(net560));
 sg13g2_nand2b_2 _4419_ (.Y(_1417_),
    .B(net565),
    .A_N(net564));
 sg13g2_nor4_2 _4420_ (.A(net573),
    .B(_1414_),
    .C(_1416_),
    .Y(_1418_),
    .D(_1417_));
 sg13g2_nor2_2 _4421_ (.A(net505),
    .B(_1418_),
    .Y(_1419_));
 sg13g2_nand2_1 _4422_ (.Y(_1420_),
    .A(net560),
    .B(\obs_inst_1.o_rom_counter[6] ));
 sg13g2_nor2_2 _4423_ (.A(net564),
    .B(_1420_),
    .Y(_1421_));
 sg13g2_nand3b_1 _4424_ (.B(net563),
    .C(net560),
    .Y(_1422_),
    .A_N(net564));
 sg13g2_nor2_2 _4425_ (.A(net573),
    .B(_1403_),
    .Y(_1423_));
 sg13g2_nor3_2 _4426_ (.A(net574),
    .B(_1403_),
    .C(_1422_),
    .Y(_1424_));
 sg13g2_nand3b_1 _4427_ (.B(net573),
    .C(\obs_rom_inst_2.i_obs_type[1] ),
    .Y(_1425_),
    .A_N(_0013_));
 sg13g2_or2_2 _4428_ (.X(_1426_),
    .B(net563),
    .A(net560));
 sg13g2_nor3_1 _4429_ (.A(_2094_),
    .B(_1425_),
    .C(_1426_),
    .Y(_1427_));
 sg13g2_nor4_1 _4430_ (.A(_2094_),
    .B(_2095_),
    .C(_1425_),
    .D(_1426_),
    .Y(_1428_));
 sg13g2_a21oi_2 _4431_ (.B1(_1428_),
    .Y(_1429_),
    .A2(_1424_),
    .A1(_2095_));
 sg13g2_nand2_1 _4432_ (.Y(_1430_),
    .A(_1419_),
    .B(_1429_));
 sg13g2_nor2_2 _4433_ (.A(net564),
    .B(net566),
    .Y(_1431_));
 sg13g2_nor2_2 _4434_ (.A(net565),
    .B(_1422_),
    .Y(_1432_));
 sg13g2_o21ai_1 _4435_ (.B1(_1423_),
    .Y(_1433_),
    .A1(net504),
    .A2(_1432_));
 sg13g2_nand2_1 _4436_ (.Y(_1434_),
    .A(_1419_),
    .B(_1433_));
 sg13g2_a21oi_1 _4437_ (.A1(_2093_),
    .A2(net506),
    .Y(_1435_),
    .B1(net571));
 sg13g2_a221oi_1 _4438_ (.B2(_1435_),
    .C1(_2098_),
    .B1(_1434_),
    .A1(_1413_),
    .Y(_1436_),
    .A2(_1430_));
 sg13g2_a21oi_1 _4439_ (.A1(net519),
    .A2(net504),
    .Y(_1437_),
    .B1(_1405_));
 sg13g2_nand2b_1 _4440_ (.Y(_1438_),
    .B(_1437_),
    .A_N(_1432_));
 sg13g2_nand3b_1 _4441_ (.B(net563),
    .C(net564),
    .Y(_1439_),
    .A_N(net560));
 sg13g2_nor3_1 _4442_ (.A(net573),
    .B(_1414_),
    .C(_1439_),
    .Y(_1440_));
 sg13g2_nor4_2 _4443_ (.A(net573),
    .B(net566),
    .C(_1414_),
    .Y(_1441_),
    .D(_1439_));
 sg13g2_nor2_1 _4444_ (.A(net519),
    .B(_1441_),
    .Y(_1442_));
 sg13g2_a21oi_1 _4445_ (.A1(net566),
    .A2(_1440_),
    .Y(_1443_),
    .B1(net505));
 sg13g2_nor2_1 _4446_ (.A(net505),
    .B(_1441_),
    .Y(_1444_));
 sg13g2_o21ai_1 _4447_ (.B1(net571),
    .Y(_1445_),
    .A1(net505),
    .A2(_1441_));
 sg13g2_o21ai_1 _4448_ (.B1(_1445_),
    .Y(_1446_),
    .A1(net571),
    .A2(_1443_));
 sg13g2_a21oi_1 _4449_ (.A1(_1438_),
    .A2(_1446_),
    .Y(_1447_),
    .B1(\obs_inst_2.o_rom_counter[1] ));
 sg13g2_nor3_1 _4450_ (.A(\obs_inst_2.o_rom_counter[2] ),
    .B(_1436_),
    .C(_1447_),
    .Y(_1448_));
 sg13g2_nor3_2 _4451_ (.A(_1417_),
    .B(_1425_),
    .C(_1426_),
    .Y(_1449_));
 sg13g2_o21ai_1 _4452_ (.B1(net566),
    .Y(_1450_),
    .A1(_1424_),
    .A2(_1449_));
 sg13g2_nor2_2 _4453_ (.A(_1407_),
    .B(_1431_),
    .Y(_1451_));
 sg13g2_o21ai_1 _4454_ (.B1(_1420_),
    .Y(_1452_),
    .A1(_1407_),
    .A2(_1431_));
 sg13g2_nand2_1 _4455_ (.Y(_1453_),
    .A(_1423_),
    .B(_1452_));
 sg13g2_nor4_2 _4456_ (.A(_2094_),
    .B(net566),
    .C(_1425_),
    .Y(_1454_),
    .D(_1426_));
 sg13g2_nor3_1 _4457_ (.A(\obs_inst_2.o_rom_counter[0] ),
    .B(_1440_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_a22oi_1 _4458_ (.Y(_1456_),
    .B1(_1453_),
    .B2(_1455_),
    .A2(_1450_),
    .A1(_1442_));
 sg13g2_nor3_2 _4459_ (.A(\obs_rom_inst_2.i_obs_type[1] ),
    .B(net573),
    .C(_0013_),
    .Y(_1457_));
 sg13g2_o21ai_1 _4460_ (.B1(_1409_),
    .Y(_1458_),
    .A1(net565),
    .A2(_1422_));
 sg13g2_nor2_2 _4461_ (.A(_2034_),
    .B(_1403_),
    .Y(_1459_));
 sg13g2_a22oi_1 _4462_ (.Y(_1460_),
    .B1(_1459_),
    .B2(_1451_),
    .A2(_1458_),
    .A1(_1457_));
 sg13g2_nand2_1 _4463_ (.Y(_1461_),
    .A(_1405_),
    .B(_1460_));
 sg13g2_nand3_1 _4464_ (.B(net505),
    .C(_1409_),
    .A(net519),
    .Y(_1462_));
 sg13g2_nand3_1 _4465_ (.B(net506),
    .C(_1422_),
    .A(net571),
    .Y(_1463_));
 sg13g2_and2_1 _4466_ (.A(_1462_),
    .B(_1463_),
    .X(_1464_));
 sg13g2_o21ai_1 _4467_ (.B1(_1464_),
    .Y(_1465_),
    .A1(_1456_),
    .A2(_1461_));
 sg13g2_a21oi_2 _4468_ (.B1(net560),
    .Y(_1466_),
    .A2(_1410_),
    .A1(net563));
 sg13g2_a22oi_1 _4469_ (.Y(_1467_),
    .B1(_1457_),
    .B2(net561),
    .A2(_1402_),
    .A1(net573));
 sg13g2_or2_1 _4470_ (.X(_1468_),
    .B(_1467_),
    .A(_1466_));
 sg13g2_nor3_2 _4471_ (.A(\obs_rom_inst_2.i_obs_type[1] ),
    .B(_2034_),
    .C(_0013_),
    .Y(_1469_));
 sg13g2_nor2_2 _4472_ (.A(_2095_),
    .B(_1422_),
    .Y(_1470_));
 sg13g2_a21oi_1 _4473_ (.A1(_1469_),
    .A2(_1470_),
    .Y(_1471_),
    .B1(_1427_));
 sg13g2_nand3_1 _4474_ (.B(_1468_),
    .C(_1471_),
    .A(_1419_),
    .Y(_1472_));
 sg13g2_a21oi_1 _4475_ (.A1(net505),
    .A2(_1466_),
    .Y(_1473_),
    .B1(net519));
 sg13g2_a22oi_1 _4476_ (.Y(_1474_),
    .B1(_1469_),
    .B2(_1421_),
    .A2(_1457_),
    .A1(_1432_));
 sg13g2_a221oi_1 _4477_ (.B2(net504),
    .C1(_1449_),
    .B1(_1459_),
    .A1(_1421_),
    .Y(_1475_),
    .A2(_1423_));
 sg13g2_nand3_1 _4478_ (.B(_1474_),
    .C(_1475_),
    .A(_1419_),
    .Y(_1476_));
 sg13g2_nand2b_1 _4479_ (.Y(_1477_),
    .B(net506),
    .A_N(_1470_));
 sg13g2_nand3_1 _4480_ (.B(_1476_),
    .C(_1477_),
    .A(net519),
    .Y(_1478_));
 sg13g2_a21oi_1 _4481_ (.A1(_1472_),
    .A2(_1473_),
    .Y(_1479_),
    .B1(_2098_));
 sg13g2_a221oi_1 _4482_ (.B2(_1479_),
    .C1(_2097_),
    .B1(_1478_),
    .A1(_2098_),
    .Y(_1480_),
    .A2(_1465_));
 sg13g2_nor3_1 _4483_ (.A(\obs_inst_2.o_rom_counter[3] ),
    .B(_1448_),
    .C(_1480_),
    .Y(_1481_));
 sg13g2_nor2_2 _4484_ (.A(net565),
    .B(_1409_),
    .Y(_1482_));
 sg13g2_nand2_1 _4485_ (.Y(_1483_),
    .A(_1457_),
    .B(_1482_));
 sg13g2_a22oi_1 _4486_ (.Y(_1484_),
    .B1(_1469_),
    .B2(net504),
    .A2(_1459_),
    .A1(net561));
 sg13g2_nand4_1 _4487_ (.B(_1450_),
    .C(_1483_),
    .A(_1443_),
    .Y(_1485_),
    .D(_1484_));
 sg13g2_a221oi_1 _4488_ (.B2(net561),
    .C1(_1424_),
    .B1(_1469_),
    .A1(_2095_),
    .Y(_1486_),
    .A2(_1427_));
 sg13g2_nand3_1 _4489_ (.B(_1468_),
    .C(_1486_),
    .A(_1444_),
    .Y(_1487_));
 sg13g2_a21oi_1 _4490_ (.A1(net505),
    .A2(_1466_),
    .Y(_1488_),
    .B1(net571));
 sg13g2_a22oi_1 _4491_ (.Y(_1489_),
    .B1(_1487_),
    .B2(_1488_),
    .A2(_1485_),
    .A1(_1413_));
 sg13g2_o21ai_1 _4492_ (.B1(_1459_),
    .Y(_1490_),
    .A1(net504),
    .A2(_1421_));
 sg13g2_nor3_1 _4493_ (.A(_2099_),
    .B(_1418_),
    .C(_1454_),
    .Y(_1491_));
 sg13g2_a22oi_1 _4494_ (.Y(_1492_),
    .B1(_1470_),
    .B2(_1459_),
    .A2(_1469_),
    .A1(_1408_));
 sg13g2_nor3_1 _4495_ (.A(net571),
    .B(net505),
    .C(_1449_),
    .Y(_1493_));
 sg13g2_a22oi_1 _4496_ (.Y(_1494_),
    .B1(_1492_),
    .B2(_1493_),
    .A2(_1491_),
    .A1(_1490_));
 sg13g2_nor3_2 _4497_ (.A(_1407_),
    .B(_1410_),
    .C(_1431_),
    .Y(_1495_));
 sg13g2_a22oi_1 _4498_ (.Y(_1496_),
    .B1(_1457_),
    .B2(_1495_),
    .A2(_1423_),
    .A1(net561));
 sg13g2_inv_1 _4499_ (.Y(_1497_),
    .A(_1496_));
 sg13g2_and2_1 _4500_ (.A(\obs_inst_2.o_rom_counter[1] ),
    .B(_1462_),
    .X(_1498_));
 sg13g2_o21ai_1 _4501_ (.B1(_1498_),
    .Y(_1499_),
    .A1(_1494_),
    .A2(_1497_));
 sg13g2_o21ai_1 _4502_ (.B1(_1499_),
    .Y(_1500_),
    .A1(\obs_inst_2.o_rom_counter[1] ),
    .A2(_1489_));
 sg13g2_nand3_1 _4503_ (.B(_1444_),
    .C(_1490_),
    .A(_1429_),
    .Y(_1501_));
 sg13g2_nand3_1 _4504_ (.B(_1415_),
    .C(_1431_),
    .A(_1406_),
    .Y(_1502_));
 sg13g2_nand3_1 _4505_ (.B(_1433_),
    .C(_1502_),
    .A(_1419_),
    .Y(_1503_));
 sg13g2_and2_1 _4506_ (.A(net571),
    .B(_1477_),
    .X(_1504_));
 sg13g2_a22oi_1 _4507_ (.Y(_1505_),
    .B1(_1503_),
    .B2(_1504_),
    .A2(_1501_),
    .A1(_1435_));
 sg13g2_nor4_1 _4508_ (.A(net573),
    .B(_1407_),
    .C(_1414_),
    .D(_1417_),
    .Y(_1506_));
 sg13g2_mux2_1 _4509_ (.A0(_1458_),
    .A1(_1506_),
    .S(_1405_),
    .X(_1507_));
 sg13g2_a21oi_1 _4510_ (.A1(net519),
    .A2(_1507_),
    .Y(_1508_),
    .B1(_2098_));
 sg13g2_o21ai_1 _4511_ (.B1(_1508_),
    .Y(_1509_),
    .A1(net519),
    .A2(_1502_));
 sg13g2_a21oi_1 _4512_ (.A1(_2098_),
    .A2(_1505_),
    .Y(_1510_),
    .B1(_2097_));
 sg13g2_a221oi_1 _4513_ (.B2(_1510_),
    .C1(_2096_),
    .B1(_1509_),
    .A1(_2097_),
    .Y(_1511_),
    .A2(_1500_));
 sg13g2_o21ai_1 _4514_ (.B1(_1404_),
    .Y(_1512_),
    .A1(\obs_rom_inst_2.i_obs_type[2] ),
    .A2(_2034_));
 sg13g2_nor4_1 _4515_ (.A(\obs_inst_2.x_offset_r[9] ),
    .B(\obs_inst_2.x_offset_r[8] ),
    .C(\obs_inst_2.x_offset_r[7] ),
    .D(\obs_inst_2.x_offset_r[6] ),
    .Y(_1513_));
 sg13g2_nor4_2 _4516_ (.A(\obs_inst_1.y_offset_r[9] ),
    .B(\obs_inst_1.y_offset_r[8] ),
    .C(\obs_inst_1.y_offset_r[7] ),
    .Y(_1514_),
    .D(\obs_inst_1.y_offset_r[6] ));
 sg13g2_nand3_1 _4517_ (.B(_1513_),
    .C(_1514_),
    .A(_1512_),
    .Y(_1515_));
 sg13g2_or3_2 _4518_ (.A(_1481_),
    .B(_1511_),
    .C(_1515_),
    .X(_1516_));
 sg13g2_nand2_2 _4519_ (.Y(_1517_),
    .A(net572),
    .B(_0012_));
 sg13g2_a21oi_2 _4520_ (.B1(\obs_rom_inst_1.i_obs_type[2] ),
    .Y(_1518_),
    .A2(_0012_),
    .A1(net572));
 sg13g2_a21o_2 _4521_ (.A2(_0012_),
    .A1(net572),
    .B1(\obs_rom_inst_1.i_obs_type[2] ),
    .X(_1519_));
 sg13g2_nand3b_1 _4522_ (.B(net572),
    .C(\obs_rom_inst_1.i_obs_type[2] ),
    .Y(_1520_),
    .A_N(\obs_rom_inst_1.i_obs_type[0] ));
 sg13g2_nor3_1 _4523_ (.A(net566),
    .B(_1439_),
    .C(_1520_),
    .Y(_1521_));
 sg13g2_nor2_1 _4524_ (.A(_1518_),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_nor2_2 _4525_ (.A(_2033_),
    .B(_1517_),
    .Y(_1523_));
 sg13g2_nand2b_1 _4526_ (.Y(_1524_),
    .B(_1523_),
    .A_N(_1466_));
 sg13g2_nand3_1 _4527_ (.B(net572),
    .C(\obs_rom_inst_1.i_obs_type[0] ),
    .A(\obs_rom_inst_1.i_obs_type[2] ),
    .Y(_1525_));
 sg13g2_nor3_2 _4528_ (.A(_2094_),
    .B(_1426_),
    .C(_1525_),
    .Y(_1526_));
 sg13g2_inv_1 _4529_ (.Y(_1527_),
    .A(_1526_));
 sg13g2_nand2_1 _4530_ (.Y(_1528_),
    .A(_2095_),
    .B(_1526_));
 sg13g2_nor2_2 _4531_ (.A(\obs_rom_inst_1.i_obs_type[0] ),
    .B(_1517_),
    .Y(_1529_));
 sg13g2_nor3_1 _4532_ (.A(\obs_rom_inst_1.i_obs_type[0] ),
    .B(_1422_),
    .C(_1517_),
    .Y(_1530_));
 sg13g2_nor2b_1 _4533_ (.A(net572),
    .B_N(\obs_rom_inst_1.i_obs_type[2] ),
    .Y(_1531_));
 sg13g2_a21oi_1 _4534_ (.A1(net562),
    .A2(_1531_),
    .Y(_1532_),
    .B1(_1530_));
 sg13g2_nand4_1 _4535_ (.B(_1524_),
    .C(_1528_),
    .A(_1522_),
    .Y(_1533_),
    .D(_1532_));
 sg13g2_a21oi_1 _4536_ (.A1(_1466_),
    .A2(net516),
    .Y(_1534_),
    .B1(net559));
 sg13g2_a21oi_1 _4537_ (.A1(_1412_),
    .A2(net516),
    .Y(_1535_),
    .B1(_2091_));
 sg13g2_and2_1 _4538_ (.A(_2033_),
    .B(_1531_),
    .X(_1536_));
 sg13g2_nand3b_1 _4539_ (.B(\obs_rom_inst_1.i_obs_type[0] ),
    .C(\obs_rom_inst_1.i_obs_type[2] ),
    .Y(_1537_),
    .A_N(net572));
 sg13g2_or2_1 _4540_ (.X(_1538_),
    .B(_1537_),
    .A(_1412_));
 sg13g2_o21ai_1 _4541_ (.B1(_1519_),
    .Y(_1539_),
    .A1(_1439_),
    .A2(_1520_));
 sg13g2_o21ai_1 _4542_ (.B1(_1539_),
    .Y(_1540_),
    .A1(net565),
    .A2(net516));
 sg13g2_nor3_2 _4543_ (.A(_1417_),
    .B(_1426_),
    .C(_1525_),
    .Y(_1541_));
 sg13g2_o21ai_1 _4544_ (.B1(\obs_inst_1.o_rom_counter[4] ),
    .Y(_1542_),
    .A1(_1530_),
    .A2(_1541_));
 sg13g2_a22oi_1 _4545_ (.Y(_1543_),
    .B1(_1536_),
    .B2(_1482_),
    .A2(_1523_),
    .A1(net562));
 sg13g2_nand4_1 _4546_ (.B(_1540_),
    .C(_1542_),
    .A(_1538_),
    .Y(_1544_),
    .D(_1543_));
 sg13g2_a221oi_1 _4547_ (.B2(_1544_),
    .C1(\obs_inst_1.o_rom_counter[1] ),
    .B1(_1535_),
    .A1(_1533_),
    .Y(_1545_),
    .A2(_1534_));
 sg13g2_nand3_1 _4548_ (.B(_1409_),
    .C(net516),
    .A(_2091_),
    .Y(_1546_));
 sg13g2_nor2_1 _4549_ (.A(_1409_),
    .B(_1537_),
    .Y(_1547_));
 sg13g2_nor4_1 _4550_ (.A(_2033_),
    .B(_2095_),
    .C(_1422_),
    .D(_1517_),
    .Y(_1548_));
 sg13g2_nor4_1 _4551_ (.A(net516),
    .B(_1541_),
    .C(_1547_),
    .D(_1548_),
    .Y(_1549_));
 sg13g2_a22oi_1 _4552_ (.Y(_1550_),
    .B1(_1536_),
    .B2(_1495_),
    .A2(_1529_),
    .A1(net562));
 sg13g2_o21ai_1 _4553_ (.B1(_1550_),
    .Y(_1551_),
    .A1(net559),
    .A2(_1549_));
 sg13g2_o21ai_1 _4554_ (.B1(_1523_),
    .Y(_1552_),
    .A1(net504),
    .A2(_1421_));
 sg13g2_or3_1 _4555_ (.A(_1416_),
    .B(_1417_),
    .C(_1520_),
    .X(_1553_));
 sg13g2_nand3_1 _4556_ (.B(_1552_),
    .C(_1553_),
    .A(_1528_),
    .Y(_1554_));
 sg13g2_a221oi_1 _4557_ (.B2(\obs_inst_1.o_rom_counter[0] ),
    .C1(_2092_),
    .B1(_1554_),
    .A1(_1546_),
    .Y(_1555_),
    .A2(_1551_));
 sg13g2_nor3_1 _4558_ (.A(\obs_inst_1.o_rom_counter[2] ),
    .B(_1545_),
    .C(_1555_),
    .Y(_1556_));
 sg13g2_nor4_2 _4559_ (.A(\obs_inst_1.o_rom_counter[5] ),
    .B(\obs_inst_1.o_rom_counter[4] ),
    .C(_1407_),
    .Y(_1557_),
    .D(_1520_));
 sg13g2_and2_1 _4560_ (.A(_1519_),
    .B(_1553_),
    .X(_1558_));
 sg13g2_o21ai_1 _4561_ (.B1(_1529_),
    .Y(_1559_),
    .A1(net504),
    .A2(_1432_));
 sg13g2_nand2_1 _4562_ (.Y(_1560_),
    .A(_1558_),
    .B(_1559_));
 sg13g2_a21oi_1 _4563_ (.A1(_1558_),
    .A2(_1559_),
    .Y(_1561_),
    .B1(\obs_inst_1.o_rom_counter[1] ));
 sg13g2_nor2_1 _4564_ (.A(_1470_),
    .B(_1519_),
    .Y(_1562_));
 sg13g2_nand2_1 _4565_ (.Y(_1563_),
    .A(_2092_),
    .B(_1562_));
 sg13g2_o21ai_1 _4566_ (.B1(_1563_),
    .Y(_1564_),
    .A1(_1557_),
    .A2(_1561_));
 sg13g2_a22oi_1 _4567_ (.Y(_1565_),
    .B1(_1529_),
    .B2(_1432_),
    .A2(_1526_),
    .A1(net565));
 sg13g2_nand3_1 _4568_ (.B(_1552_),
    .C(_1565_),
    .A(_1522_),
    .Y(_1566_));
 sg13g2_a21oi_1 _4569_ (.A1(_2093_),
    .A2(net516),
    .Y(_1567_),
    .B1(\obs_inst_1.o_rom_counter[1] ));
 sg13g2_nand2_1 _4570_ (.Y(_1568_),
    .A(_1566_),
    .B(_1567_));
 sg13g2_nand2b_1 _4571_ (.Y(_1569_),
    .B(net516),
    .A_N(_1458_));
 sg13g2_or3_1 _4572_ (.A(_1407_),
    .B(_1417_),
    .C(_1520_),
    .X(_1570_));
 sg13g2_a21oi_1 _4573_ (.A1(_1519_),
    .A2(_1570_),
    .Y(_1571_),
    .B1(_2092_));
 sg13g2_a21oi_1 _4574_ (.A1(_1569_),
    .A2(_1571_),
    .Y(_1572_),
    .B1(net559));
 sg13g2_a221oi_1 _4575_ (.B2(_1572_),
    .C1(_2089_),
    .B1(_1568_),
    .A1(\obs_inst_1.o_rom_counter[0] ),
    .Y(_1573_),
    .A2(_1564_));
 sg13g2_nor3_1 _4576_ (.A(_2090_),
    .B(_1556_),
    .C(_1573_),
    .Y(_1574_));
 sg13g2_a22oi_1 _4577_ (.Y(_1575_),
    .B1(_1536_),
    .B2(_1458_),
    .A2(_1523_),
    .A1(_1451_));
 sg13g2_a21oi_1 _4578_ (.A1(_1421_),
    .A2(net516),
    .Y(_1576_),
    .B1(_2091_));
 sg13g2_a221oi_1 _4579_ (.B2(_1452_),
    .C1(_1539_),
    .B1(_1529_),
    .A1(_2095_),
    .Y(_1577_),
    .A2(_1526_));
 sg13g2_o21ai_1 _4580_ (.B1(_1575_),
    .Y(_1578_),
    .A1(_1576_),
    .A2(_1577_));
 sg13g2_nand2b_1 _4581_ (.Y(_1579_),
    .B(_1542_),
    .A_N(_1521_));
 sg13g2_a221oi_1 _4582_ (.B2(\obs_inst_1.o_rom_counter[0] ),
    .C1(\obs_inst_1.o_rom_counter[1] ),
    .B1(_1579_),
    .A1(_1546_),
    .Y(_1580_),
    .A2(_1578_));
 sg13g2_nor2_1 _4583_ (.A(_1422_),
    .B(_1537_),
    .Y(_1581_));
 sg13g2_a21oi_1 _4584_ (.A1(_1432_),
    .A2(_1536_),
    .Y(_1582_),
    .B1(_1581_));
 sg13g2_a221oi_1 _4585_ (.B2(_1421_),
    .C1(_1541_),
    .B1(_1529_),
    .A1(_1411_),
    .Y(_1583_),
    .A2(_1523_));
 sg13g2_nand3_1 _4586_ (.B(_1582_),
    .C(_1583_),
    .A(_1558_),
    .Y(_1584_));
 sg13g2_nor2_1 _4587_ (.A(net559),
    .B(_1562_),
    .Y(_1585_));
 sg13g2_a22oi_1 _4588_ (.Y(_1586_),
    .B1(_1581_),
    .B2(net565),
    .A2(_1536_),
    .A1(net562));
 sg13g2_nand4_1 _4589_ (.B(_1527_),
    .C(_1558_),
    .A(_1524_),
    .Y(_1587_),
    .D(_1586_));
 sg13g2_a21oi_1 _4590_ (.A1(_1466_),
    .A2(_1518_),
    .Y(_1588_),
    .B1(_2091_));
 sg13g2_a221oi_1 _4591_ (.B2(_1588_),
    .C1(_2092_),
    .B1(_1587_),
    .A1(_1584_),
    .Y(_1589_),
    .A2(_1585_));
 sg13g2_nor3_1 _4592_ (.A(_2089_),
    .B(_1580_),
    .C(_1589_),
    .Y(_1590_));
 sg13g2_nand2_1 _4593_ (.Y(_1591_),
    .A(_1558_),
    .B(_1565_));
 sg13g2_a21oi_1 _4594_ (.A1(_2093_),
    .A2(_1518_),
    .Y(_1592_),
    .B1(net559));
 sg13g2_a221oi_1 _4595_ (.B2(_1560_),
    .C1(_2092_),
    .B1(_1592_),
    .A1(_1535_),
    .Y(_1593_),
    .A2(_1591_));
 sg13g2_o21ai_1 _4596_ (.B1(net559),
    .Y(_1594_),
    .A1(_1432_),
    .A2(_1519_));
 sg13g2_nor2_1 _4597_ (.A(_1522_),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_nor3_1 _4598_ (.A(net504),
    .B(_1432_),
    .C(_1519_),
    .Y(_1596_));
 sg13g2_nor3_1 _4599_ (.A(net559),
    .B(_1540_),
    .C(_1596_),
    .Y(_1597_));
 sg13g2_nor3_1 _4600_ (.A(\obs_inst_1.o_rom_counter[1] ),
    .B(_1595_),
    .C(_1597_),
    .Y(_1598_));
 sg13g2_nor3_1 _4601_ (.A(\obs_inst_1.o_rom_counter[2] ),
    .B(_1593_),
    .C(_1598_),
    .Y(_1599_));
 sg13g2_nor3_1 _4602_ (.A(\obs_inst_1.o_rom_counter[3] ),
    .B(_1590_),
    .C(_1599_),
    .Y(_1600_));
 sg13g2_a21oi_1 _4603_ (.A1(_2032_),
    .A2(\obs_rom_inst_1.i_obs_type[0] ),
    .Y(_1601_),
    .B1(_1519_));
 sg13g2_nor4_1 _4604_ (.A(\obs_inst_1.x_offset_r[9] ),
    .B(\obs_inst_1.x_offset_r[8] ),
    .C(\obs_inst_1.x_offset_r[7] ),
    .D(\obs_inst_1.x_offset_r[6] ),
    .Y(_1602_));
 sg13g2_nand2_1 _4605_ (.Y(_1603_),
    .A(_1514_),
    .B(_1602_));
 sg13g2_or4_2 _4606_ (.A(_1574_),
    .B(_1600_),
    .C(_1601_),
    .D(_1603_),
    .X(_1604_));
 sg13g2_and2_1 _4607_ (.A(_1516_),
    .B(_1604_),
    .X(_1605_));
 sg13g2_nand2_1 _4608_ (.Y(_1606_),
    .A(_1516_),
    .B(_1604_));
 sg13g2_or3_2 _4609_ (.A(net567),
    .B(net568),
    .C(_0014_),
    .X(_1607_));
 sg13g2_inv_1 _4610_ (.Y(_1608_),
    .A(_1607_));
 sg13g2_o21ai_1 _4611_ (.B1(\dino_inst.o_rom_counter[5] ),
    .Y(_1609_),
    .A1(net567),
    .A2(net568));
 sg13g2_and2_1 _4612_ (.A(\dino_inst.o_rom_counter[4] ),
    .B(\dino_inst.o_rom_counter[3] ),
    .X(_1610_));
 sg13g2_nand2_2 _4613_ (.Y(_1611_),
    .A(net567),
    .B(net568));
 sg13g2_nor2_1 _4614_ (.A(_1609_),
    .B(_1610_),
    .Y(_1612_));
 sg13g2_and3_1 _4615_ (.X(_1613_),
    .A(net567),
    .B(net568),
    .C(_0014_));
 sg13g2_nand3_1 _4616_ (.B(net568),
    .C(_0014_),
    .A(net567),
    .Y(_1614_));
 sg13g2_a21oi_1 _4617_ (.A1(_1609_),
    .A2(_1611_),
    .Y(_1615_),
    .B1(_1613_));
 sg13g2_nand3_1 _4618_ (.B(_1609_),
    .C(_1611_),
    .A(_1607_),
    .Y(_1616_));
 sg13g2_o21ai_1 _4619_ (.B1(_1609_),
    .Y(_1617_),
    .A1(\dino_inst.o_rom_counter[5] ),
    .A2(_1610_));
 sg13g2_o21ai_1 _4620_ (.B1(_0014_),
    .Y(_1618_),
    .A1(net567),
    .A2(net568));
 sg13g2_nand2b_1 _4621_ (.Y(_1619_),
    .B(_1611_),
    .A_N(_1618_));
 sg13g2_nand3b_1 _4622_ (.B(_1617_),
    .C(_1619_),
    .Y(_1620_),
    .A_N(_1615_));
 sg13g2_nand4_1 _4623_ (.B(_1614_),
    .C(_1616_),
    .A(_2186_),
    .Y(_1621_),
    .D(_1620_));
 sg13g2_o21ai_1 _4624_ (.B1(\player_constroller_inst.game_state[5] ),
    .Y(_1622_),
    .A1(_1608_),
    .A2(_1612_));
 sg13g2_a22oi_1 _4625_ (.Y(_1623_),
    .B1(_2102_),
    .B2(_1615_),
    .A2(\dino_inst.o_rom_counter[5] ),
    .A1(\player_constroller_inst.game_state[2] ));
 sg13g2_a21o_1 _4626_ (.A2(_1623_),
    .A1(_1622_),
    .B1(net513),
    .X(_1624_));
 sg13g2_a21oi_1 _4627_ (.A1(_1621_),
    .A2(_1624_),
    .Y(_1625_),
    .B1(net569));
 sg13g2_nor2b_1 _4628_ (.A(net567),
    .B_N(net568),
    .Y(_1626_));
 sg13g2_nand3b_1 _4629_ (.B(net568),
    .C(\dino_inst.o_rom_counter[5] ),
    .Y(_1627_),
    .A_N(net567));
 sg13g2_nand2_1 _4630_ (.Y(_1628_),
    .A(_1607_),
    .B(_1627_));
 sg13g2_nand3_1 _4631_ (.B(_1614_),
    .C(_1627_),
    .A(_1607_),
    .Y(_1629_));
 sg13g2_o21ai_1 _4632_ (.B1(_2187_),
    .Y(_1630_),
    .A1(_0015_),
    .A2(_1607_));
 sg13g2_nor3_1 _4633_ (.A(_0015_),
    .B(_1609_),
    .C(_1610_),
    .Y(_1631_));
 sg13g2_a221oi_1 _4634_ (.B2(_2124_),
    .C1(_1630_),
    .B1(_1629_),
    .A1(_2102_),
    .Y(_1632_),
    .A2(_1612_));
 sg13g2_nand3_1 _4635_ (.B(_1617_),
    .C(_1627_),
    .A(net513),
    .Y(_1633_));
 sg13g2_nand2_1 _4636_ (.Y(_1634_),
    .A(net569),
    .B(_1633_));
 sg13g2_o21ai_1 _4637_ (.B1(\dino_inst.o_rom_counter[1] ),
    .Y(_1635_),
    .A1(_1632_),
    .A2(_1634_));
 sg13g2_or2_1 _4638_ (.X(_1636_),
    .B(_1635_),
    .A(_1625_));
 sg13g2_nand4_1 _4639_ (.B(_1609_),
    .C(_1611_),
    .A(_1607_),
    .Y(_1637_),
    .D(_1618_));
 sg13g2_nor2_1 _4640_ (.A(_2123_),
    .B(_1617_),
    .Y(_1638_));
 sg13g2_a221oi_1 _4641_ (.B2(_1638_),
    .C1(net513),
    .B1(_1637_),
    .A1(_2102_),
    .Y(_1639_),
    .A2(_1628_));
 sg13g2_a21o_1 _4642_ (.A2(_1617_),
    .A1(net513),
    .B1(_1639_),
    .X(_1640_));
 sg13g2_a21oi_1 _4643_ (.A1(net513),
    .A2(_1620_),
    .Y(_1641_),
    .B1(_2124_));
 sg13g2_a21o_1 _4644_ (.A2(_1627_),
    .A1(_1607_),
    .B1(_1641_),
    .X(_1642_));
 sg13g2_nand2_1 _4645_ (.Y(_1643_),
    .A(_2100_),
    .B(net569));
 sg13g2_a21oi_1 _4646_ (.A1(_2187_),
    .A2(_1631_),
    .Y(_1644_),
    .B1(_1643_));
 sg13g2_a22oi_1 _4647_ (.Y(_1645_),
    .B1(_1642_),
    .B2(_1644_),
    .A2(_1640_),
    .A1(_1364_));
 sg13g2_a21o_1 _4648_ (.A2(_1645_),
    .A1(_1636_),
    .B1(\dino_inst.o_rom_counter[2] ),
    .X(_1646_));
 sg13g2_nor4_1 _4649_ (.A(\dino_inst.y_offset_r[6] ),
    .B(\dino_inst.y_offset_r[9] ),
    .C(\dino_inst.y_offset_r[8] ),
    .D(\dino_inst.y_offset_r[5] ),
    .Y(_1647_));
 sg13g2_nor4_1 _4650_ (.A(\dino_inst.x_offset_r[9] ),
    .B(\dino_inst.x_offset_r[8] ),
    .C(\dino_inst.x_offset_r[7] ),
    .D(\dino_inst.y_offset_r[7] ),
    .Y(_1648_));
 sg13g2_nand2_1 _4651_ (.Y(_1649_),
    .A(_1647_),
    .B(_1648_));
 sg13g2_nor3_1 _4652_ (.A(\dino_inst.x_offset_r[6] ),
    .B(\dino_inst.x_offset_r[5] ),
    .C(_1649_),
    .Y(_1650_));
 sg13g2_nor2_1 _4653_ (.A(_2123_),
    .B(_1637_),
    .Y(_1651_));
 sg13g2_nand2_1 _4654_ (.Y(_1652_),
    .A(_0014_),
    .B(_1626_));
 sg13g2_nor2_1 _4655_ (.A(_2123_),
    .B(_1652_),
    .Y(_1653_));
 sg13g2_o21ai_1 _4656_ (.B1(_2187_),
    .Y(_1654_),
    .A1(_0015_),
    .A2(_1617_));
 sg13g2_or3_1 _4657_ (.A(_1651_),
    .B(_1653_),
    .C(_1654_),
    .X(_1655_));
 sg13g2_nand3_1 _4658_ (.B(_1620_),
    .C(_1652_),
    .A(net513),
    .Y(_1656_));
 sg13g2_nand3_1 _4659_ (.B(_1655_),
    .C(_1656_),
    .A(_2101_),
    .Y(_1657_));
 sg13g2_or2_1 _4660_ (.X(_1658_),
    .B(_1653_),
    .A(_1630_));
 sg13g2_nand2b_1 _4661_ (.Y(_1659_),
    .B(_1626_),
    .A_N(\dino_inst.o_rom_counter[5] ));
 sg13g2_a21oi_1 _4662_ (.A1(net513),
    .A2(_1659_),
    .Y(_1660_),
    .B1(_2101_));
 sg13g2_a21oi_1 _4663_ (.A1(_1658_),
    .A2(_1660_),
    .Y(_1661_),
    .B1(_2100_));
 sg13g2_a21o_1 _4664_ (.A2(_1611_),
    .A1(_1609_),
    .B1(_0014_),
    .X(_1662_));
 sg13g2_nor3_1 _4665_ (.A(_0014_),
    .B(_2187_),
    .C(_1609_),
    .Y(_1663_));
 sg13g2_a22oi_1 _4666_ (.Y(_1664_),
    .B1(_1662_),
    .B2(_2124_),
    .A2(_1629_),
    .A1(_2102_));
 sg13g2_a21oi_1 _4667_ (.A1(_2187_),
    .A2(_1664_),
    .Y(_1665_),
    .B1(_1663_));
 sg13g2_nor2_1 _4668_ (.A(_1643_),
    .B(_1665_),
    .Y(_1666_));
 sg13g2_o21ai_1 _4669_ (.B1(\player_constroller_inst.game_state[2] ),
    .Y(_1667_),
    .A1(_0014_),
    .A2(_1611_));
 sg13g2_nand3b_1 _4670_ (.B(_1364_),
    .C(_1667_),
    .Y(_1668_),
    .A_N(\player_constroller_inst.game_state[5] ));
 sg13g2_a21oi_1 _4671_ (.A1(\player_constroller_inst.game_state[1] ),
    .A2(_1616_),
    .Y(_1669_),
    .B1(_1668_));
 sg13g2_a221oi_1 _4672_ (.B2(_2187_),
    .C1(_1666_),
    .B1(_1669_),
    .A1(_1657_),
    .Y(_1670_),
    .A2(_1661_));
 sg13g2_nand2b_1 _4673_ (.Y(_1671_),
    .B(\dino_inst.o_rom_counter[2] ),
    .A_N(_1670_));
 sg13g2_nand3_1 _4674_ (.B(_1650_),
    .C(_1671_),
    .A(_1646_),
    .Y(_1672_));
 sg13g2_inv_1 _4675_ (.Y(_1673_),
    .A(_1672_));
 sg13g2_nor3_2 _4676_ (.A(_2126_),
    .B(_0974_),
    .C(_1194_),
    .Y(_1674_));
 sg13g2_nor4_1 _4677_ (.A(\bg_render_inst.y_offset_r[8] ),
    .B(\bg_render_inst.y_offset_r[7] ),
    .C(\bg_render_inst.y_offset_r[6] ),
    .D(\bg_render_inst.y_offset_r[5] ),
    .Y(_1675_));
 sg13g2_nor2_1 _4678_ (.A(\bg_render_inst.x_offset_r[9] ),
    .B(\bg_render_inst.x_offset_r[8] ),
    .Y(_1676_));
 sg13g2_nor4_1 _4679_ (.A(\bg_render_inst.x_offset_r[7] ),
    .B(\bg_render_inst.x_offset_r[6] ),
    .C(\bg_render_inst.x_offset_r[5] ),
    .D(\bg_render_inst.y_offset_r[9] ),
    .Y(_1677_));
 sg13g2_nand3_1 _4680_ (.B(_1676_),
    .C(_1677_),
    .A(_1675_),
    .Y(_1678_));
 sg13g2_nor2_1 _4681_ (.A(\bg_object_rom_inst.i_rom_counter[3] ),
    .B(_0024_),
    .Y(_1679_));
 sg13g2_nand2_1 _4682_ (.Y(_1680_),
    .A(\bg_object_rom_inst.i_rom_counter[4] ),
    .B(_1679_));
 sg13g2_a22oi_1 _4683_ (.Y(_1681_),
    .B1(_1679_),
    .B2(\bg_object_rom_inst.i_rom_counter[4] ),
    .A2(_1230_),
    .A1(net558));
 sg13g2_and2_1 _4684_ (.A(_1208_),
    .B(_1681_),
    .X(_1682_));
 sg13g2_or2_1 _4685_ (.X(_1683_),
    .B(_1682_),
    .A(\bg_object_rom_inst.i_rom_counter[0] ));
 sg13g2_nand3b_1 _4686_ (.B(\bg_object_rom_inst.i_rom_counter[3] ),
    .C(net558),
    .Y(_1684_),
    .A_N(\bg_object_rom_inst.i_rom_counter[4] ));
 sg13g2_nand4_1 _4687_ (.B(_1680_),
    .C(_1683_),
    .A(\bg_object_rom_inst.i_rom_counter[1] ),
    .Y(_1685_),
    .D(_1684_));
 sg13g2_o21ai_1 _4688_ (.B1(_1245_),
    .Y(_1686_),
    .A1(net558),
    .A2(_1207_));
 sg13g2_a21oi_1 _4689_ (.A1(_2104_),
    .A2(_1686_),
    .Y(_1687_),
    .B1(\bg_object_rom_inst.i_rom_counter[1] ));
 sg13g2_o21ai_1 _4690_ (.B1(_1687_),
    .Y(_1688_),
    .A1(_2104_),
    .A2(_1682_));
 sg13g2_nand3_1 _4691_ (.B(_1685_),
    .C(_1688_),
    .A(\bg_object_rom_inst.i_rom_counter[2] ),
    .Y(_1689_));
 sg13g2_and2_1 _4692_ (.A(_1681_),
    .B(_1684_),
    .X(_1690_));
 sg13g2_a21oi_1 _4693_ (.A1(\bg_object_rom_inst.i_rom_counter[1] ),
    .A2(\bg_object_rom_inst.i_rom_counter[4] ),
    .Y(_1691_),
    .B1(\bg_object_rom_inst.i_rom_counter[0] ));
 sg13g2_o21ai_1 _4694_ (.B1(_1691_),
    .Y(_1692_),
    .A1(\bg_object_rom_inst.i_rom_counter[1] ),
    .A2(_1690_));
 sg13g2_a21oi_1 _4695_ (.A1(\bg_object_rom_inst.i_rom_counter[3] ),
    .A2(_2106_),
    .Y(_1693_),
    .B1(_1679_));
 sg13g2_o21ai_1 _4696_ (.B1(\bg_object_rom_inst.i_rom_counter[1] ),
    .Y(_1694_),
    .A1(net558),
    .A2(_2106_));
 sg13g2_a21oi_1 _4697_ (.A1(net558),
    .A2(\bg_object_rom_inst.i_rom_counter[3] ),
    .Y(_1695_),
    .B1(_1694_));
 sg13g2_nor2_1 _4698_ (.A(_2104_),
    .B(_1695_),
    .Y(_1696_));
 sg13g2_o21ai_1 _4699_ (.B1(_1696_),
    .Y(_1697_),
    .A1(\bg_object_rom_inst.i_rom_counter[1] ),
    .A2(_1693_));
 sg13g2_nand3_1 _4700_ (.B(_1692_),
    .C(_1697_),
    .A(_2103_),
    .Y(_1698_));
 sg13g2_a21oi_1 _4701_ (.A1(_1689_),
    .A2(_1698_),
    .Y(_1699_),
    .B1(_1678_));
 sg13g2_nor2_1 _4702_ (.A(_1674_),
    .B(_1699_),
    .Y(_1700_));
 sg13g2_and4_1 _4703_ (.A(_1516_),
    .B(_1604_),
    .C(_1672_),
    .D(_1700_),
    .X(_1701_));
 sg13g2_a21oi_1 _4704_ (.A1(_1685_),
    .A2(_1688_),
    .Y(_1702_),
    .B1(_2103_));
 sg13g2_a21oi_1 _4705_ (.A1(_1692_),
    .A2(_1697_),
    .Y(_1703_),
    .B1(\bg_object_rom_inst.i_rom_counter[2] ));
 sg13g2_nor3_1 _4706_ (.A(_1678_),
    .B(_1702_),
    .C(_1703_),
    .Y(_1704_));
 sg13g2_nand3_1 _4707_ (.B(_1650_),
    .C(_1671_),
    .A(_1646_),
    .Y(_1705_));
 sg13g2_nor2_1 _4708_ (.A(_1674_),
    .B(_1704_),
    .Y(_1706_));
 sg13g2_and3_2 _4709_ (.X(_1707_),
    .A(_1401_),
    .B(_1705_),
    .C(_1706_));
 sg13g2_a21oi_1 _4710_ (.A1(_1605_),
    .A2(_1707_),
    .Y(_1708_),
    .B1(_2117_));
 sg13g2_and3_1 _4711_ (.X(_1709_),
    .A(_2117_),
    .B(_1605_),
    .C(_1707_));
 sg13g2_nor3_1 _4712_ (.A(net603),
    .B(_1708_),
    .C(_1709_),
    .Y(_0306_));
 sg13g2_and2_1 _4713_ (.A(\graphics_inst.color_decoder_inst.rgb_scheme ),
    .B(_1401_),
    .X(_1710_));
 sg13g2_and3_1 _4714_ (.X(_1711_),
    .A(\graphics_inst.color_decoder_inst.rgb_scheme ),
    .B(_1401_),
    .C(_1672_));
 sg13g2_nand3_1 _4715_ (.B(_1401_),
    .C(_1672_),
    .A(\graphics_inst.color_decoder_inst.rgb_scheme ),
    .Y(_1712_));
 sg13g2_a221oi_1 _4716_ (.B2(_1605_),
    .C1(_2117_),
    .B1(_1711_),
    .A1(_1401_),
    .Y(_1713_),
    .A2(_1701_));
 sg13g2_nor3_1 _4717_ (.A(_0023_),
    .B(_1606_),
    .C(_1712_),
    .Y(_1714_));
 sg13g2_nor4_1 _4718_ (.A(net603),
    .B(_1709_),
    .C(_1713_),
    .D(_1714_),
    .Y(_0307_));
 sg13g2_a221oi_1 _4719_ (.B2(_1606_),
    .C1(_2117_),
    .B1(_1711_),
    .A1(_1401_),
    .Y(_1715_),
    .A2(_1701_));
 sg13g2_nor3_1 _4720_ (.A(_0023_),
    .B(_1605_),
    .C(_1712_),
    .Y(_1716_));
 sg13g2_nor4_1 _4721_ (.A(net603),
    .B(_1709_),
    .C(_1715_),
    .D(_1716_),
    .Y(_0308_));
 sg13g2_a221oi_1 _4722_ (.B2(_1707_),
    .C1(_2117_),
    .B1(_1605_),
    .A1(\graphics_inst.color_decoder_inst.rgb_scheme ),
    .Y(_1717_),
    .A2(_1401_));
 sg13g2_and2_1 _4723_ (.A(_2117_),
    .B(_1710_),
    .X(_1718_));
 sg13g2_nor4_1 _4724_ (.A(net603),
    .B(_1709_),
    .C(_1717_),
    .D(_1718_),
    .Y(_0309_));
 sg13g2_a221oi_1 _4725_ (.B2(_1673_),
    .C1(_2117_),
    .B1(_1710_),
    .A1(_1605_),
    .Y(_1719_),
    .A2(_1707_));
 sg13g2_and3_1 _4726_ (.X(_1720_),
    .A(_2117_),
    .B(_1673_),
    .C(_1710_));
 sg13g2_nor4_1 _4727_ (.A(net603),
    .B(_1709_),
    .C(_1719_),
    .D(_1720_),
    .Y(_0310_));
 sg13g2_nor2_1 _4728_ (.A(net596),
    .B(net497),
    .Y(_0311_));
 sg13g2_nand3_1 _4729_ (.B(_1606_),
    .C(_1673_),
    .A(net409),
    .Y(_1721_));
 sg13g2_a21oi_1 _4730_ (.A1(_2026_),
    .A2(_1721_),
    .Y(_0312_),
    .B1(_0467_));
 sg13g2_and2_1 _4731_ (.A(net622),
    .B(net1),
    .X(_0313_));
 sg13g2_and2_1 _4732_ (.A(net621),
    .B(net399),
    .X(_0314_));
 sg13g2_a21oi_1 _4733_ (.A1(_2025_),
    .A2(net501),
    .Y(_1722_),
    .B1(net808));
 sg13g2_a21oi_1 _4734_ (.A1(net808),
    .A2(net501),
    .Y(_1723_),
    .B1(_1722_));
 sg13g2_and2_1 _4735_ (.A(net607),
    .B(_1723_),
    .X(_0315_));
 sg13g2_nand2b_1 _4736_ (.Y(_1724_),
    .B(net457),
    .A_N(net501));
 sg13g2_a21oi_1 _4737_ (.A1(net497),
    .A2(_1724_),
    .Y(_0316_),
    .B1(net597));
 sg13g2_nand2_1 _4738_ (.Y(_1725_),
    .A(net435),
    .B(_2023_));
 sg13g2_nand2b_1 _4739_ (.Y(_1726_),
    .B(net668),
    .A_N(net427));
 sg13g2_nand2b_1 _4740_ (.Y(_1727_),
    .B(net684),
    .A_N(net628));
 sg13g2_nor2_1 _4741_ (.A(_1726_),
    .B(_1727_),
    .Y(_1728_));
 sg13g2_nand2b_1 _4742_ (.Y(_1729_),
    .B(net703),
    .A_N(\score[6] ));
 sg13g2_and3_1 _4743_ (.X(_1730_),
    .A(net406),
    .B(net499),
    .C(_0465_));
 sg13g2_nand2b_1 _4744_ (.Y(_1731_),
    .B(net405),
    .A_N(net403));
 sg13g2_nor2_1 _4745_ (.A(net426),
    .B(_1731_),
    .Y(_1732_));
 sg13g2_and2_1 _4746_ (.A(_1730_),
    .B(_1732_),
    .X(_1733_));
 sg13g2_nand4_1 _4747_ (.B(net499),
    .C(_0465_),
    .A(net722),
    .Y(_1734_),
    .D(_1732_));
 sg13g2_nor2_2 _4748_ (.A(_2021_),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_nor4_2 _4749_ (.A(net673),
    .B(_2021_),
    .C(_1729_),
    .Y(_1736_),
    .D(_1734_));
 sg13g2_nand3_1 _4750_ (.B(_1728_),
    .C(_1736_),
    .A(net410),
    .Y(_1737_));
 sg13g2_nor3_2 _4751_ (.A(net413),
    .B(_1725_),
    .C(_1737_),
    .Y(_1738_));
 sg13g2_and2_1 _4752_ (.A(net422),
    .B(_1738_),
    .X(_1739_));
 sg13g2_nor4_2 _4753_ (.A(net673),
    .B(_2021_),
    .C(_1729_),
    .Y(_1740_),
    .D(_1734_));
 sg13g2_and2_1 _4754_ (.A(_1728_),
    .B(_1740_),
    .X(_1741_));
 sg13g2_and2_1 _4755_ (.A(net410),
    .B(_1741_),
    .X(_1742_));
 sg13g2_nor2_1 _4756_ (.A(net422),
    .B(_1738_),
    .Y(_1743_));
 sg13g2_nor3_1 _4757_ (.A(net488),
    .B(_1739_),
    .C(_1743_),
    .Y(_0317_));
 sg13g2_and2_1 _4758_ (.A(net750),
    .B(_1739_),
    .X(_1744_));
 sg13g2_nor3_1 _4759_ (.A(_2024_),
    .B(net715),
    .C(net750),
    .Y(_1745_));
 sg13g2_nor2_1 _4760_ (.A(net750),
    .B(_1739_),
    .Y(_1746_));
 sg13g2_nor4_1 _4761_ (.A(net488),
    .B(_1744_),
    .C(_1745_),
    .D(_1746_),
    .Y(_0318_));
 sg13g2_or2_1 _4762_ (.X(_1747_),
    .B(_1744_),
    .A(net715));
 sg13g2_nand2_1 _4763_ (.Y(_1748_),
    .A(net715),
    .B(_1744_));
 sg13g2_and3_1 _4764_ (.X(_0319_),
    .A(_0466_),
    .B(_1747_),
    .C(_1748_));
 sg13g2_xor2_1 _4765_ (.B(net750),
    .A(net715),
    .X(_1749_));
 sg13g2_nor2_1 _4766_ (.A(_2024_),
    .B(_1749_),
    .Y(_1750_));
 sg13g2_a221oi_1 _4767_ (.B2(_1739_),
    .C1(net488),
    .B1(_1750_),
    .A1(_2024_),
    .Y(_0320_),
    .A2(_1748_));
 sg13g2_nor2_1 _4768_ (.A(net410),
    .B(_1741_),
    .Y(_1751_));
 sg13g2_nor3_1 _4769_ (.A(net487),
    .B(_1742_),
    .C(_1751_),
    .Y(_0321_));
 sg13g2_a21oi_1 _4770_ (.A1(_1725_),
    .A2(_1742_),
    .Y(_1752_),
    .B1(net413));
 sg13g2_and2_1 _4771_ (.A(net413),
    .B(_1742_),
    .X(_1753_));
 sg13g2_nor3_1 _4772_ (.A(net487),
    .B(_1752_),
    .C(_1753_),
    .Y(_0322_));
 sg13g2_o21ai_1 _4773_ (.B1(_0466_),
    .Y(_1754_),
    .A1(\graphics_inst.color_decoder_inst.rgb_scheme ),
    .A2(_1753_));
 sg13g2_nand2_1 _4774_ (.Y(_1755_),
    .A(\graphics_inst.color_decoder_inst.rgb_scheme ),
    .B(_1753_));
 sg13g2_nor2b_1 _4775_ (.A(_1754_),
    .B_N(_1755_),
    .Y(_0323_));
 sg13g2_xor2_1 _4776_ (.B(_1755_),
    .A(net435),
    .X(_1756_));
 sg13g2_nor3_1 _4777_ (.A(net488),
    .B(_1738_),
    .C(_1756_),
    .Y(_0324_));
 sg13g2_or2_1 _4778_ (.X(_1757_),
    .B(_1736_),
    .A(net684));
 sg13g2_nand2_1 _4779_ (.Y(_1758_),
    .A(net684),
    .B(_1736_));
 sg13g2_and3_1 _4780_ (.X(_0325_),
    .A(_0466_),
    .B(_1757_),
    .C(_1758_));
 sg13g2_nand2_1 _4781_ (.Y(_1759_),
    .A(net628),
    .B(_1758_));
 sg13g2_nand3b_1 _4782_ (.B(net723),
    .C(_1726_),
    .Y(_1760_),
    .A_N(_1727_));
 sg13g2_a21oi_1 _4783_ (.A1(_1759_),
    .A2(_1760_),
    .Y(_0326_),
    .B1(net486));
 sg13g2_nand2_1 _4784_ (.Y(_1761_),
    .A(\score[9] ),
    .B(net790));
 sg13g2_xnor2_1 _4785_ (.Y(_1762_),
    .A(_0023_),
    .B(net791));
 sg13g2_o21ai_1 _4786_ (.B1(_1740_),
    .Y(_1763_),
    .A1(_1728_),
    .A2(_1762_));
 sg13g2_o21ai_1 _4787_ (.B1(_1763_),
    .Y(_1764_),
    .A1(net427),
    .A2(net705));
 sg13g2_nor2_1 _4788_ (.A(net487),
    .B(_1764_),
    .Y(_0327_));
 sg13g2_nand4_1 _4789_ (.B(net628),
    .C(net684),
    .A(net427),
    .Y(_1765_),
    .D(_1740_));
 sg13g2_nor2_1 _4790_ (.A(net487),
    .B(_1741_),
    .Y(_1766_));
 sg13g2_o21ai_1 _4791_ (.B1(_1766_),
    .Y(_1767_),
    .A1(_2022_),
    .A2(_1765_));
 sg13g2_a21oi_1 _4792_ (.A1(_2022_),
    .A2(_1765_),
    .Y(_0328_),
    .B1(_1767_));
 sg13g2_nor2_1 _4793_ (.A(net463),
    .B(_1733_),
    .Y(_1768_));
 sg13g2_nor3_1 _4794_ (.A(net486),
    .B(_1735_),
    .C(_1768_),
    .Y(_0329_));
 sg13g2_nor3_1 _4795_ (.A(_2020_),
    .B(net486),
    .C(_1735_),
    .Y(_1769_));
 sg13g2_nand4_1 _4796_ (.B(_0466_),
    .C(net704),
    .A(_2020_),
    .Y(_1770_),
    .D(_1735_));
 sg13g2_nand2b_1 _4797_ (.Y(_0330_),
    .B(_1770_),
    .A_N(_1769_));
 sg13g2_a21oi_1 _4798_ (.A1(net673),
    .A2(_1735_),
    .Y(_1771_),
    .B1(net452));
 sg13g2_and3_1 _4799_ (.X(_1772_),
    .A(net452),
    .B(net673),
    .C(_1735_));
 sg13g2_nor3_1 _4800_ (.A(net486),
    .B(net674),
    .C(_1772_),
    .Y(_0331_));
 sg13g2_nor2_1 _4801_ (.A(net649),
    .B(_1772_),
    .Y(_1773_));
 sg13g2_and2_1 _4802_ (.A(net649),
    .B(_1772_),
    .X(_1774_));
 sg13g2_nor4_1 _4803_ (.A(net486),
    .B(_1736_),
    .C(_1773_),
    .D(_1774_),
    .Y(_0332_));
 sg13g2_a21oi_1 _4804_ (.A1(net499),
    .A2(_0465_),
    .Y(_1775_),
    .B1(net406));
 sg13g2_nor3_1 _4805_ (.A(net487),
    .B(_1730_),
    .C(_1775_),
    .Y(_0333_));
 sg13g2_and2_1 _4806_ (.A(net426),
    .B(_1730_),
    .X(_1776_));
 sg13g2_a21oi_1 _4807_ (.A1(_1730_),
    .A2(_1731_),
    .Y(_1777_),
    .B1(net426));
 sg13g2_nor3_1 _4808_ (.A(net486),
    .B(_1776_),
    .C(_1777_),
    .Y(_0334_));
 sg13g2_nor2_1 _4809_ (.A(net403),
    .B(_1776_),
    .Y(_1778_));
 sg13g2_and2_1 _4810_ (.A(net403),
    .B(_1776_),
    .X(_1779_));
 sg13g2_nor3_1 _4811_ (.A(net486),
    .B(_1778_),
    .C(_1779_),
    .Y(_0335_));
 sg13g2_nor2_1 _4812_ (.A(net405),
    .B(_1779_),
    .Y(_1780_));
 sg13g2_and2_1 _4813_ (.A(net405),
    .B(_1779_),
    .X(_1781_));
 sg13g2_nor4_1 _4814_ (.A(net486),
    .B(_1733_),
    .C(_1780_),
    .D(_1781_),
    .Y(_0336_));
 sg13g2_a22oi_1 _4815_ (.Y(_1782_),
    .B1(_2082_),
    .B2(\audio_inst.i_over.counter[10] ),
    .A2(_2081_),
    .A1(\audio_inst.i_over.counter[11] ));
 sg13g2_nand2b_1 _4816_ (.Y(_1783_),
    .B(\audio_inst.i_over.decay_value[6] ),
    .A_N(\audio_inst.i_over.counter[6] ));
 sg13g2_nand2b_1 _4817_ (.Y(_1784_),
    .B(\audio_inst.i_over.counter[1] ),
    .A_N(\audio_inst.i_over.decay_value[1] ));
 sg13g2_a22oi_1 _4818_ (.Y(_1785_),
    .B1(\audio_inst.i_over.decay_value[0] ),
    .B2(_2017_),
    .A2(\audio_inst.i_over.decay_value[1] ),
    .A1(_2016_));
 sg13g2_o21ai_1 _4819_ (.B1(_1784_),
    .Y(_1786_),
    .A1(_2015_),
    .A2(\audio_inst.i_over.decay_value[2] ));
 sg13g2_a22oi_1 _4820_ (.Y(_1787_),
    .B1(\audio_inst.i_over.decay_value[2] ),
    .B2(_2015_),
    .A2(\audio_inst.i_over.decay_value[3] ),
    .A1(_2014_));
 sg13g2_o21ai_1 _4821_ (.B1(_1787_),
    .Y(_1788_),
    .A1(_1785_),
    .A2(_1786_));
 sg13g2_a22oi_1 _4822_ (.Y(_1789_),
    .B1(_2085_),
    .B2(\audio_inst.i_over.counter[3] ),
    .A2(_2084_),
    .A1(\audio_inst.i_over.counter[4] ));
 sg13g2_nor2_1 _4823_ (.A(\audio_inst.i_over.counter[4] ),
    .B(_2084_),
    .Y(_1790_));
 sg13g2_a221oi_1 _4824_ (.B2(_1789_),
    .C1(_1790_),
    .B1(_1788_),
    .A1(_2013_),
    .Y(_1791_),
    .A2(\audio_inst.i_over.decay_value[5] ));
 sg13g2_nor2_1 _4825_ (.A(_2013_),
    .B(\audio_inst.i_over.decay_value[5] ),
    .Y(_1792_));
 sg13g2_o21ai_1 _4826_ (.B1(_1783_),
    .Y(_1793_),
    .A1(_1791_),
    .A2(_1792_));
 sg13g2_nand2b_1 _4827_ (.Y(_1794_),
    .B(\audio_inst.i_over.counter[7] ),
    .A_N(\audio_inst.i_over.decay_value[7] ));
 sg13g2_nand2b_1 _4828_ (.Y(_1795_),
    .B(\audio_inst.i_over.counter[6] ),
    .A_N(\audio_inst.i_over.decay_value[6] ));
 sg13g2_nand3_1 _4829_ (.B(_1794_),
    .C(_1795_),
    .A(_1793_),
    .Y(_1796_));
 sg13g2_nand2b_1 _4830_ (.Y(_1797_),
    .B(\audio_inst.i_over.counter[8] ),
    .A_N(\audio_inst.i_over.decay_value[8] ));
 sg13g2_o21ai_1 _4831_ (.B1(_1797_),
    .Y(_1798_),
    .A1(\audio_inst.i_over.counter[9] ),
    .A2(_2083_));
 sg13g2_a221oi_1 _4832_ (.B2(_2012_),
    .C1(_1798_),
    .B1(\audio_inst.i_over.decay_value[7] ),
    .A1(_2011_),
    .Y(_1799_),
    .A2(\audio_inst.i_over.decay_value[8] ));
 sg13g2_a21oi_1 _4833_ (.A1(_2010_),
    .A2(\audio_inst.i_over.decay_value[9] ),
    .Y(_1800_),
    .B1(_1797_));
 sg13g2_a221oi_1 _4834_ (.B2(_1799_),
    .C1(_1800_),
    .B1(_1796_),
    .A1(\audio_inst.i_over.counter[9] ),
    .Y(_1801_),
    .A2(_2083_));
 sg13g2_nor2_1 _4835_ (.A(\audio_inst.i_over.counter[10] ),
    .B(_2082_),
    .Y(_1802_));
 sg13g2_o21ai_1 _4836_ (.B1(_1782_),
    .Y(_1803_),
    .A1(_1801_),
    .A2(_1802_));
 sg13g2_nor2_1 _4837_ (.A(_2008_),
    .B(\audio_inst.i_over.decay_value[15] ),
    .Y(_1804_));
 sg13g2_xnor2_1 _4838_ (.Y(_1805_),
    .A(\audio_inst.i_over.counter[15] ),
    .B(\audio_inst.i_over.decay_value[15] ));
 sg13g2_xnor2_1 _4839_ (.Y(_1806_),
    .A(\audio_inst.i_over.counter[14] ),
    .B(\audio_inst.i_over.decay_value[14] ));
 sg13g2_nor2b_1 _4840_ (.A(\audio_inst.i_over.decay_value[13] ),
    .B_N(\audio_inst.i_over.counter[13] ),
    .Y(_1807_));
 sg13g2_nand2b_1 _4841_ (.Y(_1808_),
    .B(\audio_inst.i_over.counter[13] ),
    .A_N(\audio_inst.i_over.decay_value[13] ));
 sg13g2_nand2b_1 _4842_ (.Y(_1809_),
    .B(\audio_inst.i_over.decay_value[12] ),
    .A_N(\audio_inst.i_over.counter[12] ));
 sg13g2_nand2b_1 _4843_ (.Y(_1810_),
    .B(\audio_inst.i_over.counter[12] ),
    .A_N(\audio_inst.i_over.decay_value[12] ));
 sg13g2_nor2b_1 _4844_ (.A(\audio_inst.i_over.counter[13] ),
    .B_N(\audio_inst.i_over.decay_value[13] ),
    .Y(_1811_));
 sg13g2_nor2_1 _4845_ (.A(\audio_inst.i_over.counter[11] ),
    .B(_2081_),
    .Y(_1812_));
 sg13g2_nand4_1 _4846_ (.B(_1806_),
    .C(_1809_),
    .A(_1805_),
    .Y(_1813_),
    .D(_1810_));
 sg13g2_nor4_1 _4847_ (.A(_1807_),
    .B(_1811_),
    .C(_1812_),
    .D(_1813_),
    .Y(_1814_));
 sg13g2_o21ai_1 _4848_ (.B1(_1808_),
    .Y(_1815_),
    .A1(_1810_),
    .A2(_1811_));
 sg13g2_nand3_1 _4849_ (.B(_1806_),
    .C(_1815_),
    .A(_1805_),
    .Y(_1816_));
 sg13g2_nand3b_1 _4850_ (.B(_1805_),
    .C(\audio_inst.i_over.counter[14] ),
    .Y(_1817_),
    .A_N(\audio_inst.i_over.decay_value[14] ));
 sg13g2_nor4_1 _4851_ (.A(\audio_inst.i_over.counter[18] ),
    .B(\audio_inst.i_over.counter[17] ),
    .C(\audio_inst.i_over.counter[16] ),
    .D(_1804_),
    .Y(_1818_));
 sg13g2_nand4_1 _4852_ (.B(_1816_),
    .C(_1817_),
    .A(_2203_),
    .Y(_1819_),
    .D(_1818_));
 sg13g2_a21oi_1 _4853_ (.A1(_1803_),
    .A2(_1814_),
    .Y(_1820_),
    .B1(_1819_));
 sg13g2_nand2_1 _4854_ (.Y(_1821_),
    .A(\audio_inst.i_over.counter[11] ),
    .B(\audio_inst.i_over.counter[10] ));
 sg13g2_nor4_1 _4855_ (.A(\audio_inst.i_over.counter[5] ),
    .B(\audio_inst.i_over.counter[4] ),
    .C(\audio_inst.i_over.counter[1] ),
    .D(\audio_inst.i_over.counter[0] ),
    .Y(_1822_));
 sg13g2_nand4_1 _4856_ (.B(_2015_),
    .C(_2086_),
    .A(_2014_),
    .Y(_1823_),
    .D(_1822_));
 sg13g2_a21o_1 _4857_ (.A2(_1823_),
    .A1(\audio_inst.i_over.counter[6] ),
    .B1(\audio_inst.i_over.counter[7] ),
    .X(_1824_));
 sg13g2_a21oi_1 _4858_ (.A1(\audio_inst.i_over.counter[8] ),
    .A2(_1824_),
    .Y(_1825_),
    .B1(\audio_inst.i_over.counter[9] ));
 sg13g2_nor4_1 _4859_ (.A(\audio_inst.i_over.counter[15] ),
    .B(\audio_inst.i_over.counter[14] ),
    .C(\audio_inst.i_over.counter[13] ),
    .D(\audio_inst.i_over.counter[12] ),
    .Y(_1826_));
 sg13g2_o21ai_1 _4860_ (.B1(_1826_),
    .Y(_1827_),
    .A1(_1821_),
    .A2(_1825_));
 sg13g2_nand3_1 _4861_ (.B(\audio_inst.i_over.counter[16] ),
    .C(_1827_),
    .A(\audio_inst.i_over.counter[17] ),
    .Y(_1828_));
 sg13g2_nand2b_2 _4862_ (.Y(_1829_),
    .B(_1828_),
    .A_N(\audio_inst.i_over.counter[18] ));
 sg13g2_nand2_2 _4863_ (.Y(_1830_),
    .A(_2202_),
    .B(_1829_));
 sg13g2_nor2_2 _4864_ (.A(net600),
    .B(_0725_),
    .Y(_1831_));
 sg13g2_nand2b_2 _4865_ (.Y(_1832_),
    .B(_1831_),
    .A_N(_2200_));
 sg13g2_nor2_2 _4866_ (.A(_1830_),
    .B(_1832_),
    .Y(_1833_));
 sg13g2_or2_2 _4867_ (.X(_1834_),
    .B(_1832_),
    .A(_1830_));
 sg13g2_nand2_1 _4868_ (.Y(_1835_),
    .A(_1820_),
    .B(_1831_));
 sg13g2_a22oi_1 _4869_ (.Y(_0337_),
    .B1(_1834_),
    .B2(_1835_),
    .A2(_1820_),
    .A1(_2019_));
 sg13g2_a21oi_1 _4870_ (.A1(_2202_),
    .A2(_1829_),
    .Y(_1836_),
    .B1(_1832_));
 sg13g2_nand2b_2 _4871_ (.Y(_1837_),
    .B(_1830_),
    .A_N(_1832_));
 sg13g2_a22oi_1 _4872_ (.Y(_1838_),
    .B1(net471),
    .B2(\audio_inst.i_over.stage_index[0] ),
    .A2(_1833_),
    .A1(net415));
 sg13g2_inv_1 _4873_ (.Y(_0338_),
    .A(net416));
 sg13g2_nand2_1 _4874_ (.Y(_1839_),
    .A(net544),
    .B(net471));
 sg13g2_o21ai_1 _4875_ (.B1(_1839_),
    .Y(_0339_),
    .A1(_0732_),
    .A2(_1834_));
 sg13g2_a22oi_1 _4876_ (.Y(_1840_),
    .B1(net471),
    .B2(net543),
    .A2(_1833_),
    .A1(_0715_));
 sg13g2_inv_1 _4877_ (.Y(_0340_),
    .A(_1840_));
 sg13g2_nand2_1 _4878_ (.Y(_1841_),
    .A(net538),
    .B(net471));
 sg13g2_xnor2_1 _4879_ (.Y(_1842_),
    .A(_2087_),
    .B(_0714_));
 sg13g2_o21ai_1 _4880_ (.B1(_1841_),
    .Y(_0341_),
    .A1(_1834_),
    .A2(_1842_));
 sg13g2_nand2_1 _4881_ (.Y(_1843_),
    .A(\audio_inst.i_over.stage_index[4] ),
    .B(net471));
 sg13g2_xnor2_1 _4882_ (.Y(_1844_),
    .A(net782),
    .B(_0394_));
 sg13g2_o21ai_1 _4883_ (.B1(_1843_),
    .Y(_0342_),
    .A1(_1834_),
    .A2(_1844_));
 sg13g2_nor3_2 _4884_ (.A(_2200_),
    .B(_2201_),
    .C(_1829_),
    .Y(_1845_));
 sg13g2_o21ai_1 _4885_ (.B1(_1831_),
    .Y(_1846_),
    .A1(net785),
    .A2(_1845_));
 sg13g2_a21oi_1 _4886_ (.A1(net785),
    .A2(_2202_),
    .Y(_0343_),
    .B1(_1846_));
 sg13g2_and3_1 _4887_ (.X(_1847_),
    .A(net740),
    .B(net914),
    .C(_2202_));
 sg13g2_a21oi_1 _4888_ (.A1(\audio_inst.i_over.counter[0] ),
    .A2(_2202_),
    .Y(_1848_),
    .B1(net740));
 sg13g2_nor3_1 _4889_ (.A(_1837_),
    .B(_1847_),
    .C(net741),
    .Y(_0344_));
 sg13g2_o21ai_1 _4890_ (.B1(net471),
    .Y(_1849_),
    .A1(net676),
    .A2(_1847_));
 sg13g2_a21oi_1 _4891_ (.A1(net676),
    .A2(_1847_),
    .Y(_0345_),
    .B1(_1849_));
 sg13g2_a21oi_1 _4892_ (.A1(net676),
    .A2(_1847_),
    .Y(_1850_),
    .B1(net739));
 sg13g2_and4_1 _4893_ (.A(\audio_inst.i_over.counter[3] ),
    .B(\audio_inst.i_over.counter[2] ),
    .C(\audio_inst.i_over.counter[1] ),
    .D(\audio_inst.i_over.counter[0] ),
    .X(_1851_));
 sg13g2_and2_2 _4894_ (.A(_2202_),
    .B(_1851_),
    .X(_1852_));
 sg13g2_nor3_1 _4895_ (.A(_1837_),
    .B(_1850_),
    .C(_1852_),
    .Y(_0346_));
 sg13g2_o21ai_1 _4896_ (.B1(net472),
    .Y(_1853_),
    .A1(net851),
    .A2(_1852_));
 sg13g2_a21oi_1 _4897_ (.A1(net851),
    .A2(_1852_),
    .Y(_0347_),
    .B1(_1853_));
 sg13g2_and3_1 _4898_ (.X(_1854_),
    .A(net730),
    .B(\audio_inst.i_over.counter[4] ),
    .C(_1852_));
 sg13g2_a21oi_1 _4899_ (.A1(\audio_inst.i_over.counter[4] ),
    .A2(_1852_),
    .Y(_1855_),
    .B1(net730));
 sg13g2_nor3_1 _4900_ (.A(_1837_),
    .B(_1854_),
    .C(net731),
    .Y(_0348_));
 sg13g2_o21ai_1 _4901_ (.B1(net472),
    .Y(_1856_),
    .A1(net809),
    .A2(_1854_));
 sg13g2_a21oi_1 _4902_ (.A1(net809),
    .A2(_1854_),
    .Y(_0349_),
    .B1(_1856_));
 sg13g2_and4_1 _4903_ (.A(\audio_inst.i_over.counter[7] ),
    .B(\audio_inst.i_over.counter[6] ),
    .C(\audio_inst.i_over.counter[5] ),
    .D(\audio_inst.i_over.counter[4] ),
    .X(_1857_));
 sg13g2_and2_1 _4904_ (.A(_1852_),
    .B(_1857_),
    .X(_1858_));
 sg13g2_a21oi_1 _4905_ (.A1(\audio_inst.i_over.counter[6] ),
    .A2(_1854_),
    .Y(_1859_),
    .B1(net728));
 sg13g2_nor3_1 _4906_ (.A(_1837_),
    .B(_1858_),
    .C(net729),
    .Y(_0350_));
 sg13g2_o21ai_1 _4907_ (.B1(net472),
    .Y(_1860_),
    .A1(net804),
    .A2(_1858_));
 sg13g2_a21oi_1 _4908_ (.A1(net804),
    .A2(_1858_),
    .Y(_0351_),
    .B1(_1860_));
 sg13g2_a21oi_1 _4909_ (.A1(net804),
    .A2(_1858_),
    .Y(_1861_),
    .B1(net807));
 sg13g2_nand4_1 _4910_ (.B(\audio_inst.i_over.counter[8] ),
    .C(_1851_),
    .A(\audio_inst.i_over.counter[9] ),
    .Y(_1862_),
    .D(_1857_));
 sg13g2_nor2_2 _4911_ (.A(_2201_),
    .B(_1862_),
    .Y(_1863_));
 sg13g2_nor3_1 _4912_ (.A(_1837_),
    .B(_1861_),
    .C(_1863_),
    .Y(_0352_));
 sg13g2_and2_1 _4913_ (.A(net870),
    .B(_1863_),
    .X(_1864_));
 sg13g2_o21ai_1 _4914_ (.B1(net472),
    .Y(_1865_),
    .A1(net870),
    .A2(_1863_));
 sg13g2_nor2_1 _4915_ (.A(_1864_),
    .B(_1865_),
    .Y(_0353_));
 sg13g2_and2_1 _4916_ (.A(net863),
    .B(_1864_),
    .X(_1866_));
 sg13g2_o21ai_1 _4917_ (.B1(net472),
    .Y(_1867_),
    .A1(net863),
    .A2(_1864_));
 sg13g2_nor2_1 _4918_ (.A(_1866_),
    .B(net864),
    .Y(_0354_));
 sg13g2_and2_1 _4919_ (.A(net846),
    .B(_1866_),
    .X(_1868_));
 sg13g2_o21ai_1 _4920_ (.B1(net472),
    .Y(_1869_),
    .A1(net846),
    .A2(_1866_));
 sg13g2_nor2_1 _4921_ (.A(_1868_),
    .B(net847),
    .Y(_0355_));
 sg13g2_nand4_1 _4922_ (.B(net846),
    .C(net909),
    .A(net858),
    .Y(_1870_),
    .D(\audio_inst.i_over.counter[10] ));
 sg13g2_nor3_2 _4923_ (.A(_2201_),
    .B(_1862_),
    .C(net910),
    .Y(_1871_));
 sg13g2_o21ai_1 _4924_ (.B1(net471),
    .Y(_1872_),
    .A1(net858),
    .A2(_1868_));
 sg13g2_nor2_1 _4925_ (.A(_1871_),
    .B(_1872_),
    .Y(_0356_));
 sg13g2_nand2_1 _4926_ (.Y(_1873_),
    .A(net880),
    .B(_1871_));
 sg13g2_o21ai_1 _4927_ (.B1(net471),
    .Y(_1874_),
    .A1(net880),
    .A2(_1871_));
 sg13g2_nor2b_1 _4928_ (.A(_1874_),
    .B_N(_1873_),
    .Y(_0357_));
 sg13g2_xnor2_1 _4929_ (.Y(_1875_),
    .A(_2008_),
    .B(_1873_));
 sg13g2_nor2_1 _4930_ (.A(_1837_),
    .B(_1875_),
    .Y(_0358_));
 sg13g2_nor3_1 _4931_ (.A(_2008_),
    .B(_2009_),
    .C(_1870_),
    .Y(_1876_));
 sg13g2_nor2b_1 _4932_ (.A(_1862_),
    .B_N(_1876_),
    .Y(_1877_));
 sg13g2_a21oi_1 _4933_ (.A1(_1845_),
    .A2(_1877_),
    .Y(_1878_),
    .B1(net708));
 sg13g2_and3_1 _4934_ (.X(_1879_),
    .A(net708),
    .B(_1863_),
    .C(_1876_));
 sg13g2_nor3_1 _4935_ (.A(_1837_),
    .B(_1878_),
    .C(_1879_),
    .Y(_0359_));
 sg13g2_xnor2_1 _4936_ (.Y(_1880_),
    .A(net765),
    .B(_1879_));
 sg13g2_nor2_1 _4937_ (.A(_1837_),
    .B(_1880_),
    .Y(_0360_));
 sg13g2_a22oi_1 _4938_ (.Y(_1881_),
    .B1(_1845_),
    .B2(_2086_),
    .A2(_2201_),
    .A1(\audio_inst.i_over.counter[18] ));
 sg13g2_nor2b_1 _4939_ (.A(net408),
    .B_N(_1831_),
    .Y(_0361_));
 sg13g2_a21oi_1 _4940_ (.A1(net433),
    .A2(_2202_),
    .Y(_1882_),
    .B1(_0725_));
 sg13g2_nor2_1 _4941_ (.A(net600),
    .B(_1882_),
    .Y(_0362_));
 sg13g2_nor2b_1 _4942_ (.A(\audio_inst.i_jump.decay_value[10] ),
    .B_N(\audio_inst.i_jump.counter[10] ),
    .Y(_1883_));
 sg13g2_nor2b_1 _4943_ (.A(\audio_inst.i_jump.decay_value[11] ),
    .B_N(\audio_inst.i_jump.counter[11] ),
    .Y(_1884_));
 sg13g2_nand2b_1 _4944_ (.Y(_1885_),
    .B(\audio_inst.i_jump.decay_value[11] ),
    .A_N(\audio_inst.i_jump.counter[11] ));
 sg13g2_o21ai_1 _4945_ (.B1(_1885_),
    .Y(_1886_),
    .A1(_1883_),
    .A2(_1884_));
 sg13g2_o21ai_1 _4946_ (.B1(_1885_),
    .Y(_1887_),
    .A1(\audio_inst.i_jump.counter[10] ),
    .A2(_2079_));
 sg13g2_nor3_1 _4947_ (.A(_1883_),
    .B(_1884_),
    .C(_1887_),
    .Y(_1888_));
 sg13g2_nand2b_1 _4948_ (.Y(_1889_),
    .B(\audio_inst.i_jump.counter[9] ),
    .A_N(\audio_inst.i_jump.decay_value[9] ));
 sg13g2_nand2b_1 _4949_ (.Y(_1890_),
    .B(\audio_inst.i_jump.decay_value[9] ),
    .A_N(\audio_inst.i_jump.counter[9] ));
 sg13g2_nand3b_1 _4950_ (.B(_1890_),
    .C(\audio_inst.i_jump.counter[8] ),
    .Y(_1891_),
    .A_N(\audio_inst.i_jump.decay_value[8] ));
 sg13g2_nand2_1 _4951_ (.Y(_1892_),
    .A(_1889_),
    .B(_1891_));
 sg13g2_nor2_1 _4952_ (.A(\audio_inst.i_jump.counter[5] ),
    .B(_2076_),
    .Y(_1893_));
 sg13g2_nor2_1 _4953_ (.A(\audio_inst.i_jump.counter[2] ),
    .B(_2071_),
    .Y(_1894_));
 sg13g2_nand2b_1 _4954_ (.Y(_1895_),
    .B(\audio_inst.i_jump.decay_value[1] ),
    .A_N(\audio_inst.i_jump.counter[1] ));
 sg13g2_nand2b_1 _4955_ (.Y(_1896_),
    .B(\audio_inst.i_jump.decay_value[0] ),
    .A_N(\audio_inst.i_jump.counter[0] ));
 sg13g2_nor2b_1 _4956_ (.A(\audio_inst.i_jump.decay_value[1] ),
    .B_N(\audio_inst.i_jump.counter[1] ),
    .Y(_1897_));
 sg13g2_a221oi_1 _4957_ (.B2(_1896_),
    .C1(_1897_),
    .B1(_1895_),
    .A1(\audio_inst.i_jump.counter[2] ),
    .Y(_1898_),
    .A2(_2071_));
 sg13g2_nand2_1 _4958_ (.Y(_1899_),
    .A(\audio_inst.i_jump.counter[3] ),
    .B(_2072_));
 sg13g2_o21ai_1 _4959_ (.B1(_1899_),
    .Y(_1900_),
    .A1(_1894_),
    .A2(_1898_));
 sg13g2_a22oi_1 _4960_ (.Y(_1901_),
    .B1(\audio_inst.i_jump.decay_value[4] ),
    .B2(_2067_),
    .A2(\audio_inst.i_jump.decay_value[3] ),
    .A1(_2064_));
 sg13g2_a22oi_1 _4961_ (.Y(_1902_),
    .B1(_1900_),
    .B2(_1901_),
    .A2(_2075_),
    .A1(\audio_inst.i_jump.counter[4] ));
 sg13g2_a22oi_1 _4962_ (.Y(_1903_),
    .B1(_2076_),
    .B2(\audio_inst.i_jump.counter[5] ),
    .A2(_2073_),
    .A1(\audio_inst.i_jump.counter[6] ));
 sg13g2_o21ai_1 _4963_ (.B1(_1903_),
    .Y(_1904_),
    .A1(_1893_),
    .A2(_1902_));
 sg13g2_a22oi_1 _4964_ (.Y(_1905_),
    .B1(\audio_inst.i_jump.decay_value[7] ),
    .B2(_2065_),
    .A2(\audio_inst.i_jump.decay_value[6] ),
    .A1(_2066_));
 sg13g2_a22oi_1 _4965_ (.Y(_1906_),
    .B1(_1904_),
    .B2(_1905_),
    .A2(_2074_),
    .A1(\audio_inst.i_jump.counter[7] ));
 sg13g2_xnor2_1 _4966_ (.Y(_1907_),
    .A(\audio_inst.i_jump.counter[8] ),
    .B(\audio_inst.i_jump.decay_value[8] ));
 sg13g2_nand4_1 _4967_ (.B(_1889_),
    .C(_1890_),
    .A(_1888_),
    .Y(_1908_),
    .D(_1907_));
 sg13g2_nand2_1 _4968_ (.Y(_1909_),
    .A(_1888_),
    .B(_1892_));
 sg13g2_and2_1 _4969_ (.A(_1886_),
    .B(_1909_),
    .X(_1910_));
 sg13g2_o21ai_1 _4970_ (.B1(_1910_),
    .Y(_1911_),
    .A1(_1906_),
    .A2(_1908_));
 sg13g2_nand2_1 _4971_ (.Y(_1912_),
    .A(_2068_),
    .B(\audio_inst.i_jump.decay_value[14] ));
 sg13g2_o21ai_1 _4972_ (.B1(_1912_),
    .Y(_1913_),
    .A1(\audio_inst.i_jump.counter[13] ),
    .A2(_2077_));
 sg13g2_nor2b_1 _4973_ (.A(\audio_inst.i_jump.counter[12] ),
    .B_N(\audio_inst.i_jump.decay_value[12] ),
    .Y(_1914_));
 sg13g2_nand2b_1 _4974_ (.Y(_1915_),
    .B(\audio_inst.i_jump.decay_value[15] ),
    .A_N(\audio_inst.i_jump.counter[15] ));
 sg13g2_nor2b_1 _4975_ (.A(\audio_inst.i_jump.decay_value[12] ),
    .B_N(\audio_inst.i_jump.counter[12] ),
    .Y(_1916_));
 sg13g2_a21o_1 _4976_ (.A2(_2077_),
    .A1(\audio_inst.i_jump.counter[13] ),
    .B1(_1916_),
    .X(_1917_));
 sg13g2_nand2b_1 _4977_ (.Y(_1918_),
    .B(\audio_inst.i_jump.counter[15] ),
    .A_N(\audio_inst.i_jump.decay_value[15] ));
 sg13g2_nand2b_1 _4978_ (.Y(_1919_),
    .B(\audio_inst.i_jump.counter[14] ),
    .A_N(\audio_inst.i_jump.decay_value[14] ));
 sg13g2_nand3_1 _4979_ (.B(_1918_),
    .C(_1919_),
    .A(_1915_),
    .Y(_1920_));
 sg13g2_nor4_1 _4980_ (.A(_1913_),
    .B(_1914_),
    .C(_1917_),
    .D(_1920_),
    .Y(_1921_));
 sg13g2_nand2b_1 _4981_ (.Y(_1922_),
    .B(_1917_),
    .A_N(_1913_));
 sg13g2_nand3_1 _4982_ (.B(_1919_),
    .C(_1922_),
    .A(_1918_),
    .Y(_1923_));
 sg13g2_a22oi_1 _4983_ (.Y(_1924_),
    .B1(_1923_),
    .B2(_1915_),
    .A2(_1921_),
    .A1(_1911_));
 sg13g2_nand2b_1 _4984_ (.Y(_1925_),
    .B(\audio_inst.i_jump.counter[17] ),
    .A_N(\audio_inst.i_jump.decay_value[17] ));
 sg13g2_o21ai_1 _4985_ (.B1(_1925_),
    .Y(_1926_),
    .A1(_2069_),
    .A2(\audio_inst.i_jump.decay_value[16] ));
 sg13g2_nand2_1 _4986_ (.Y(_1927_),
    .A(_2069_),
    .B(\audio_inst.i_jump.decay_value[16] ));
 sg13g2_nand2b_1 _4987_ (.Y(_1928_),
    .B(\audio_inst.i_jump.decay_value[17] ),
    .A_N(\audio_inst.i_jump.counter[17] ));
 sg13g2_nand3b_1 _4988_ (.B(_1927_),
    .C(_1928_),
    .Y(_1929_),
    .A_N(_1926_));
 sg13g2_a21oi_1 _4989_ (.A1(_1926_),
    .A2(_1928_),
    .Y(_1930_),
    .B1(net774));
 sg13g2_o21ai_1 _4990_ (.B1(_1930_),
    .Y(_1931_),
    .A1(_1924_),
    .A2(_1929_));
 sg13g2_nor2_1 _4991_ (.A(net777),
    .B(_1931_),
    .Y(_1932_));
 sg13g2_a21oi_1 _4992_ (.A1(_0652_),
    .A2(_1931_),
    .Y(_1933_),
    .B1(net481));
 sg13g2_nor2b_1 _4993_ (.A(_1932_),
    .B_N(_1933_),
    .Y(_0363_));
 sg13g2_nand2_2 _4994_ (.Y(_1934_),
    .A(_0641_),
    .B(_0653_));
 sg13g2_and3_1 _4995_ (.X(_1935_),
    .A(net646),
    .B(_0641_),
    .C(_0653_));
 sg13g2_nor3_2 _4996_ (.A(_2050_),
    .B(\audio_inst.i_jump.state[1] ),
    .C(_0652_),
    .Y(_1936_));
 sg13g2_nor2_1 _4997_ (.A(net646),
    .B(_1936_),
    .Y(_1937_));
 sg13g2_nor3_1 _4998_ (.A(_0429_),
    .B(_1935_),
    .C(net647),
    .Y(_0364_));
 sg13g2_a22oi_1 _4999_ (.Y(_1938_),
    .B1(_1936_),
    .B2(_0898_),
    .A2(_1934_),
    .A1(net533));
 sg13g2_nor2_1 _5000_ (.A(_0429_),
    .B(net891),
    .Y(_0365_));
 sg13g2_nor2_1 _5001_ (.A(_0021_),
    .B(_0878_),
    .Y(_1939_));
 sg13g2_xor2_1 _5002_ (.B(_0878_),
    .A(_0021_),
    .X(_1940_));
 sg13g2_a22oi_1 _5003_ (.Y(_1941_),
    .B1(_1936_),
    .B2(_1940_),
    .A2(_1934_),
    .A1(net531));
 sg13g2_nor2_1 _5004_ (.A(_0429_),
    .B(net878),
    .Y(_0366_));
 sg13g2_xnor2_1 _5005_ (.Y(_1942_),
    .A(net744),
    .B(_1939_));
 sg13g2_a22oi_1 _5006_ (.Y(_1943_),
    .B1(_1936_),
    .B2(_1942_),
    .A2(_1934_),
    .A1(net528));
 sg13g2_nor2_1 _5007_ (.A(_0429_),
    .B(net745),
    .Y(_0367_));
 sg13g2_xor2_1 _5008_ (.B(_0886_),
    .A(net700),
    .X(_1944_));
 sg13g2_a22oi_1 _5009_ (.Y(_1945_),
    .B1(_1936_),
    .B2(_1944_),
    .A2(_1934_),
    .A1(net525));
 sg13g2_nor2_1 _5010_ (.A(_0429_),
    .B(net701),
    .Y(_0368_));
 sg13g2_nor2b_1 _5011_ (.A(\gamepad_pmod.driver.pmod_latch_prev ),
    .B_N(net386),
    .Y(_1946_));
 sg13g2_nor2_1 _5012_ (.A(net598),
    .B(net514),
    .Y(_1947_));
 sg13g2_a22oi_1 _5013_ (.Y(_0369_),
    .B1(net503),
    .B2(_2052_),
    .A2(net515),
    .A1(_2005_));
 sg13g2_a22oi_1 _5014_ (.Y(_0370_),
    .B1(net503),
    .B2(_2053_),
    .A2(net515),
    .A1(_2004_));
 sg13g2_a22oi_1 _5015_ (.Y(_0371_),
    .B1(net502),
    .B2(_2054_),
    .A2(net514),
    .A1(_2003_));
 sg13g2_a22oi_1 _5016_ (.Y(_0372_),
    .B1(net502),
    .B2(_2055_),
    .A2(net515),
    .A1(_2002_));
 sg13g2_a22oi_1 _5017_ (.Y(_0373_),
    .B1(net503),
    .B2(_2056_),
    .A2(net515),
    .A1(_2001_));
 sg13g2_a22oi_1 _5018_ (.Y(_0374_),
    .B1(net503),
    .B2(_2057_),
    .A2(net515),
    .A1(_2000_));
 sg13g2_a22oi_1 _5019_ (.Y(_0375_),
    .B1(net502),
    .B2(_2058_),
    .A2(net514),
    .A1(_1999_));
 sg13g2_a22oi_1 _5020_ (.Y(_0376_),
    .B1(net502),
    .B2(_2059_),
    .A2(net514),
    .A1(_1998_));
 sg13g2_a22oi_1 _5021_ (.Y(_0377_),
    .B1(net502),
    .B2(_2060_),
    .A2(net514),
    .A1(_1997_));
 sg13g2_a22oi_1 _5022_ (.Y(_0378_),
    .B1(net502),
    .B2(_2061_),
    .A2(net514),
    .A1(_1996_));
 sg13g2_a22oi_1 _5023_ (.Y(_0379_),
    .B1(net502),
    .B2(_2062_),
    .A2(net514),
    .A1(_1995_));
 sg13g2_a22oi_1 _5024_ (.Y(_0380_),
    .B1(net502),
    .B2(_2063_),
    .A2(net514),
    .A1(_1994_));
 sg13g2_a21oi_1 _5025_ (.A1(_2182_),
    .A2(net630),
    .Y(_0381_),
    .B1(net597));
 sg13g2_o21ai_1 _5026_ (.B1(net620),
    .Y(_1948_),
    .A1(net777),
    .A2(net466));
 sg13g2_inv_1 _5027_ (.Y(_0382_),
    .A(_1948_));
 sg13g2_nand4_1 _5028_ (.B(net428),
    .C(net436),
    .A(net655),
    .Y(_1949_),
    .D(net642));
 sg13g2_nand4_1 _5029_ (.B(net439),
    .C(net654),
    .A(net411),
    .Y(_1950_),
    .D(net671));
 sg13g2_nand4_1 _5030_ (.B(net430),
    .C(net418),
    .A(net449),
    .Y(_1951_),
    .D(net468));
 sg13g2_nor3_2 _5031_ (.A(_1949_),
    .B(_1950_),
    .C(_1951_),
    .Y(_1952_));
 sg13g2_inv_1 _5032_ (.Y(_1953_),
    .A(_1952_));
 sg13g2_nand2_2 _5033_ (.Y(_1954_),
    .A(_2026_),
    .B(_0465_));
 sg13g2_nand2_1 _5034_ (.Y(_1955_),
    .A(net779),
    .B(net662));
 sg13g2_nor2_1 _5035_ (.A(net447),
    .B(\ai_controller_inst.restart_counter[6] ),
    .Y(_1956_));
 sg13g2_nand3_1 _5036_ (.B(net767),
    .C(_1956_),
    .A(net659),
    .Y(_1957_));
 sg13g2_nor4_1 _5037_ (.A(net751),
    .B(net690),
    .C(_1955_),
    .D(_1957_),
    .Y(_1958_));
 sg13g2_nand4_1 _5038_ (.B(_1952_),
    .C(_1954_),
    .A(_2135_),
    .Y(_1959_),
    .D(_1958_));
 sg13g2_nand2_1 _5039_ (.Y(_1960_),
    .A(net501),
    .B(_1952_));
 sg13g2_nor2b_1 _5040_ (.A(_1960_),
    .B_N(_1954_),
    .Y(_1961_));
 sg13g2_nand2_1 _5041_ (.Y(_1962_),
    .A(net610),
    .B(_1959_));
 sg13g2_inv_1 _5042_ (.Y(_1963_),
    .A(_1962_));
 sg13g2_nor2_1 _5043_ (.A(net690),
    .B(_1961_),
    .Y(_1964_));
 sg13g2_and4_1 _5044_ (.A(net690),
    .B(net501),
    .C(_1952_),
    .D(_1954_),
    .X(_1965_));
 sg13g2_nor3_1 _5045_ (.A(_1962_),
    .B(_1964_),
    .C(_1965_),
    .Y(_0383_));
 sg13g2_and2_1 _5046_ (.A(net751),
    .B(_1965_),
    .X(_1966_));
 sg13g2_o21ai_1 _5047_ (.B1(net611),
    .Y(_1967_),
    .A1(net751),
    .A2(_1965_));
 sg13g2_nor2_1 _5048_ (.A(_1966_),
    .B(_1967_),
    .Y(_0384_));
 sg13g2_nor2_1 _5049_ (.A(net662),
    .B(_1966_),
    .Y(_1968_));
 sg13g2_and2_1 _5050_ (.A(net662),
    .B(_1966_),
    .X(_1969_));
 sg13g2_nor3_1 _5051_ (.A(_1962_),
    .B(net663),
    .C(_1969_),
    .Y(_0385_));
 sg13g2_and2_1 _5052_ (.A(net779),
    .B(_1969_),
    .X(_1970_));
 sg13g2_o21ai_1 _5053_ (.B1(_1963_),
    .Y(_1971_),
    .A1(net779),
    .A2(_1969_));
 sg13g2_nor2_1 _5054_ (.A(_1970_),
    .B(_1971_),
    .Y(_0386_));
 sg13g2_and2_1 _5055_ (.A(net767),
    .B(_1970_),
    .X(_1972_));
 sg13g2_o21ai_1 _5056_ (.B1(_1963_),
    .Y(_1973_),
    .A1(net767),
    .A2(_1970_));
 sg13g2_nor2_1 _5057_ (.A(_1972_),
    .B(net768),
    .Y(_0387_));
 sg13g2_o21ai_1 _5058_ (.B1(_1963_),
    .Y(_1974_),
    .A1(net659),
    .A2(_1972_));
 sg13g2_a21oi_1 _5059_ (.A1(net659),
    .A2(_1972_),
    .Y(_0388_),
    .B1(_1974_));
 sg13g2_a21oi_1 _5060_ (.A1(\ai_controller_inst.restart_counter[5] ),
    .A2(_1972_),
    .Y(_1975_),
    .B1(net441));
 sg13g2_nand3_1 _5061_ (.B(\ai_controller_inst.restart_counter[5] ),
    .C(_1972_),
    .A(net441),
    .Y(_1976_));
 sg13g2_nand2_1 _5062_ (.Y(_1977_),
    .A(net610),
    .B(_1976_));
 sg13g2_nor2_1 _5063_ (.A(net442),
    .B(_1977_),
    .Y(_0389_));
 sg13g2_o21ai_1 _5064_ (.B1(net610),
    .Y(_1978_),
    .A1(_1993_),
    .A2(_1976_));
 sg13g2_a21oi_1 _5065_ (.A1(_1993_),
    .A2(_1976_),
    .Y(_0390_),
    .B1(_1978_));
 sg13g2_a21oi_1 _5066_ (.A1(net501),
    .A2(_1954_),
    .Y(_1979_),
    .B1(_1953_));
 sg13g2_nand2_1 _5067_ (.Y(_1980_),
    .A(_2058_),
    .B(_2063_));
 sg13g2_a22oi_1 _5068_ (.Y(_1981_),
    .B1(_1980_),
    .B2(_1953_),
    .A2(_1979_),
    .A1(net522));
 sg13g2_nor2_1 _5069_ (.A(net596),
    .B(_1981_),
    .Y(_0391_));
 sg13g2_nand2b_1 _5070_ (.Y(_1982_),
    .B(_0518_),
    .A_N(\ai_controller_inst.obstacle2_pos[6] ));
 sg13g2_nor2b_1 _5071_ (.A(_0478_),
    .B_N(_0477_),
    .Y(_1983_));
 sg13g2_a21oi_1 _5072_ (.A1(\ai_controller_inst.obstacle2_pos[7] ),
    .A2(_1982_),
    .Y(_1984_),
    .B1(_1983_));
 sg13g2_o21ai_1 _5073_ (.B1(_2030_),
    .Y(_1985_),
    .A1(_2031_),
    .A2(_0471_));
 sg13g2_a22oi_1 _5074_ (.Y(_1986_),
    .B1(_1985_),
    .B2(\ai_controller_inst.obstacle1_pos[7] ),
    .A2(_0483_),
    .A1(_0469_));
 sg13g2_nand2b_1 _5075_ (.Y(_1987_),
    .B(_1952_),
    .A_N(net802));
 sg13g2_o21ai_1 _5076_ (.B1(_1987_),
    .Y(_1988_),
    .A1(net468),
    .A2(net671));
 sg13g2_a22oi_1 _5077_ (.Y(_1989_),
    .B1(_1986_),
    .B2(_0468_),
    .A2(_1984_),
    .A1(_0490_));
 sg13g2_nor2_1 _5078_ (.A(_1954_),
    .B(_1989_),
    .Y(_1990_));
 sg13g2_o21ai_1 _5079_ (.B1(net614),
    .Y(_1991_),
    .A1(_1960_),
    .A2(_1990_));
 sg13g2_a21oi_1 _5080_ (.A1(_1960_),
    .A2(_1988_),
    .Y(_0392_),
    .B1(_1991_));
 sg13g2_a22oi_1 _5081_ (.Y(_1992_),
    .B1(_1979_),
    .B2(net800),
    .A2(_1953_),
    .A1(net655));
 sg13g2_a21oi_1 _5082_ (.A1(_1959_),
    .A2(_1992_),
    .Y(_0393_),
    .B1(net598));
 sg13g2_dfrbp_1 _5083_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net36),
    .D(net894),
    .Q_N(_2528_),
    .Q(\audio_inst.i_jump.state[1] ));
 sg13g2_dfrbp_1 _5084_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net158),
    .D(_0037_),
    .Q_N(_2527_),
    .Q(\audio_inst.i_jump.state[0] ));
 sg13g2_dfrbp_1 _5085_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net157),
    .D(_0038_),
    .Q_N(_2526_),
    .Q(\audio_inst.i_over.state[1] ));
 sg13g2_dfrbp_1 _5086_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net156),
    .D(_0039_),
    .Q_N(_2525_),
    .Q(\score_inst_5.num_r[0] ));
 sg13g2_dfrbp_1 _5087_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net155),
    .D(_0040_),
    .Q_N(_2524_),
    .Q(\score_inst_5.num_r[1] ));
 sg13g2_dfrbp_1 _5088_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net154),
    .D(_0041_),
    .Q_N(_2523_),
    .Q(\score_inst_5.num_r[2] ));
 sg13g2_dfrbp_1 _5089_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net153),
    .D(_0042_),
    .Q_N(_2522_),
    .Q(\score_inst_5.num_r[3] ));
 sg13g2_dfrbp_1 _5090_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net152),
    .D(_0043_),
    .Q_N(_0035_),
    .Q(\graphics_inst.hpos[0] ));
 sg13g2_dfrbp_1 _5091_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net151),
    .D(_0044_),
    .Q_N(_2521_),
    .Q(\graphics_inst.hpos[1] ));
 sg13g2_dfrbp_1 _5092_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net150),
    .D(_0045_),
    .Q_N(\score_inst_2.x_offset[2] ),
    .Q(\bg_render_inst.i_hpos[2] ));
 sg13g2_dfrbp_1 _5093_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net149),
    .D(_0046_),
    .Q_N(\dino_inst.x_offset[3] ),
    .Q(\bg_render_inst.i_hpos[3] ));
 sg13g2_dfrbp_1 _5094_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net148),
    .D(_0047_),
    .Q_N(\score_inst_1.x_offset[4] ),
    .Q(\bg_render_inst.i_hpos[4] ));
 sg13g2_dfrbp_1 _5095_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net147),
    .D(_0048_),
    .Q_N(_0029_),
    .Q(\bg_render_inst.i_hpos[5] ));
 sg13g2_dfrbp_1 _5096_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0049_),
    .Q_N(\score_inst_5.x_offset[6] ),
    .Q(\bg_render_inst.i_hpos[6] ));
 sg13g2_dfrbp_1 _5097_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net145),
    .D(_0050_),
    .Q_N(_2520_),
    .Q(\bg_render_inst.i_hpos[7] ));
 sg13g2_dfrbp_1 _5098_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net144),
    .D(_0051_),
    .Q_N(_0030_),
    .Q(\bg_render_inst.i_hpos[8] ));
 sg13g2_dfrbp_1 _5099_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net143),
    .D(_0052_),
    .Q_N(_0010_),
    .Q(\bg_render_inst.i_hpos[9] ));
 sg13g2_dfrbp_1 _5100_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net37),
    .D(net658),
    .Q_N(_2529_),
    .Q(\audio_inst.i_jump.decay_value[17] ));
 sg13g2_dfrbp_1 _5101_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net321),
    .D(net385),
    .Q_N(_2530_),
    .Q(\gamepad_pmod.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _5102_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net142),
    .D(net386),
    .Q_N(_2519_),
    .Q(\gamepad_pmod.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _5103_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net140),
    .D(net421),
    .Q_N(_2518_),
    .Q(\gamepad_pmod.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _5104_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net138),
    .D(net638),
    .Q_N(_2517_),
    .Q(\gamepad_pmod.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _5105_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net136),
    .D(net665),
    .Q_N(_2516_),
    .Q(\gamepad_pmod.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _5106_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net134),
    .D(_0057_),
    .Q_N(_2515_),
    .Q(\gamepad_pmod.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _5107_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net132),
    .D(net734),
    .Q_N(_2514_),
    .Q(\gamepad_pmod.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _5108_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net130),
    .D(net719),
    .Q_N(_2513_),
    .Q(\gamepad_pmod.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _5109_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net128),
    .D(net645),
    .Q_N(_2512_),
    .Q(\gamepad_pmod.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _5110_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net126),
    .D(net651),
    .Q_N(_2511_),
    .Q(\gamepad_pmod.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _5111_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net124),
    .D(net682),
    .Q_N(_2510_),
    .Q(\gamepad_pmod.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _5112_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net122),
    .D(net641),
    .Q_N(_2509_),
    .Q(\gamepad_pmod.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _5113_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net120),
    .D(net695),
    .Q_N(_2508_),
    .Q(\gamepad_pmod.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _5114_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net118),
    .D(net633),
    .Q_N(_2507_),
    .Q(\gamepad_pmod.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _5115_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net116),
    .D(_0066_),
    .Q_N(_2506_),
    .Q(\gamepad_pmod.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _5116_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net115),
    .D(_0067_),
    .Q_N(_2505_),
    .Q(\gamepad_pmod.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _5117_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net114),
    .D(_0068_),
    .Q_N(_2504_),
    .Q(\gamepad_pmod.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _5118_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net113),
    .D(_0069_),
    .Q_N(_2503_),
    .Q(\gamepad_pmod.driver.pmod_clk_sync[1] ));
 sg13g2_dfrbp_1 _5119_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net112),
    .D(_0070_),
    .Q_N(_2502_),
    .Q(\dino_inst.i_ypos[0] ));
 sg13g2_dfrbp_1 _5120_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net110),
    .D(_0071_),
    .Q_N(_2501_),
    .Q(\dino_inst.i_ypos[1] ));
 sg13g2_dfrbp_1 _5121_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net108),
    .D(_0072_),
    .Q_N(_2500_),
    .Q(\dino_inst.i_ypos[2] ));
 sg13g2_dfrbp_1 _5122_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net106),
    .D(_0073_),
    .Q_N(_2499_),
    .Q(\dino_inst.i_ypos[3] ));
 sg13g2_dfrbp_1 _5123_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net104),
    .D(_0074_),
    .Q_N(_2498_),
    .Q(\dino_inst.i_ypos[4] ));
 sg13g2_dfrbp_1 _5124_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net102),
    .D(_0075_),
    .Q_N(_2497_),
    .Q(\dino_inst.i_ypos[5] ));
 sg13g2_dfrbp_1 _5125_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net100),
    .D(_0076_),
    .Q_N(_2496_),
    .Q(\player_constroller_inst.u_player_physics.velocity[0] ));
 sg13g2_dfrbp_1 _5126_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net98),
    .D(net670),
    .Q_N(_2495_),
    .Q(\player_constroller_inst.u_player_physics.velocity[1] ));
 sg13g2_dfrbp_1 _5127_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net96),
    .D(net653),
    .Q_N(_2494_),
    .Q(\player_constroller_inst.u_player_physics.velocity[2] ));
 sg13g2_dfrbp_1 _5128_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net94),
    .D(_0079_),
    .Q_N(_2493_),
    .Q(\player_constroller_inst.u_player_physics.velocity[3] ));
 sg13g2_dfrbp_1 _5129_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net92),
    .D(_0080_),
    .Q_N(_2492_),
    .Q(\obstacles_inst.obstacle2_cross_gen_line_reg ));
 sg13g2_dfrbp_1 _5130_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net90),
    .D(_0081_),
    .Q_N(_2491_),
    .Q(\obstacles_inst.obstacle1_cross_gen_line_reg ));
 sg13g2_dfrbp_1 _5131_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net88),
    .D(net454),
    .Q_N(_2490_),
    .Q(\obs_rom_inst_2.i_obs_type[0] ));
 sg13g2_dfrbp_1 _5132_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net86),
    .D(_0083_),
    .Q_N(_2489_),
    .Q(\obs_rom_inst_2.i_obs_type[1] ));
 sg13g2_dfrbp_1 _5133_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net84),
    .D(net721),
    .Q_N(_0013_),
    .Q(\obs_rom_inst_2.i_obs_type[2] ));
 sg13g2_dfrbp_1 _5134_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net82),
    .D(net714),
    .Q_N(_2488_),
    .Q(\obs_rom_inst_1.i_obs_type[0] ));
 sg13g2_dfrbp_1 _5135_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net80),
    .D(_0086_),
    .Q_N(_2487_),
    .Q(\obs_rom_inst_1.i_obs_type[1] ));
 sg13g2_dfrbp_1 _5136_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net78),
    .D(net748),
    .Q_N(_0012_),
    .Q(\obs_rom_inst_1.i_obs_type[2] ));
 sg13g2_dfrbp_1 _5137_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net76),
    .D(net823),
    .Q_N(_0017_),
    .Q(\ai_controller_inst.obstacle2_pos[2] ));
 sg13g2_dfrbp_1 _5138_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net74),
    .D(_0089_),
    .Q_N(_2486_),
    .Q(\ai_controller_inst.obstacle2_pos[3] ));
 sg13g2_dfrbp_1 _5139_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net72),
    .D(_0090_),
    .Q_N(_2485_),
    .Q(\ai_controller_inst.obstacle2_pos[4] ));
 sg13g2_dfrbp_1 _5140_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net70),
    .D(_0091_),
    .Q_N(_2484_),
    .Q(\ai_controller_inst.obstacle2_pos[5] ));
 sg13g2_dfrbp_1 _5141_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net68),
    .D(_0092_),
    .Q_N(_2483_),
    .Q(\ai_controller_inst.obstacle2_pos[6] ));
 sg13g2_dfrbp_1 _5142_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net66),
    .D(_0093_),
    .Q_N(_2482_),
    .Q(\ai_controller_inst.obstacle2_pos[7] ));
 sg13g2_dfrbp_1 _5143_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net64),
    .D(_0094_),
    .Q_N(_2481_),
    .Q(\ai_controller_inst.obstacle2_pos[8] ));
 sg13g2_dfrbp_1 _5144_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net62),
    .D(_0095_),
    .Q_N(_2480_),
    .Q(\ai_controller_inst.obstacle2_pos[9] ));
 sg13g2_dfrbp_1 _5145_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net60),
    .D(net850),
    .Q_N(_0016_),
    .Q(\ai_controller_inst.obstacle1_pos[2] ));
 sg13g2_dfrbp_1 _5146_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net58),
    .D(net862),
    .Q_N(_2479_),
    .Q(\ai_controller_inst.obstacle1_pos[3] ));
 sg13g2_dfrbp_1 _5147_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net56),
    .D(_0098_),
    .Q_N(_2478_),
    .Q(\ai_controller_inst.obstacle1_pos[4] ));
 sg13g2_dfrbp_1 _5148_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net54),
    .D(net793),
    .Q_N(_2477_),
    .Q(\ai_controller_inst.obstacle1_pos[5] ));
 sg13g2_dfrbp_1 _5149_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net52),
    .D(_0100_),
    .Q_N(_2476_),
    .Q(\ai_controller_inst.obstacle1_pos[6] ));
 sg13g2_dfrbp_1 _5150_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net50),
    .D(_0101_),
    .Q_N(_2475_),
    .Q(\ai_controller_inst.obstacle1_pos[7] ));
 sg13g2_dfrbp_1 _5151_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net48),
    .D(_0102_),
    .Q_N(_2474_),
    .Q(\ai_controller_inst.obstacle1_pos[8] ));
 sg13g2_dfrbp_1 _5152_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net46),
    .D(net727),
    .Q_N(_2473_),
    .Q(\ai_controller_inst.obstacle1_pos[9] ));
 sg13g2_dfrbp_1 _5153_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net44),
    .D(net825),
    .Q_N(_0018_),
    .Q(\bg_object_inst.bg_object_pos[2] ));
 sg13g2_dfrbp_1 _5154_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net42),
    .D(_0105_),
    .Q_N(_2472_),
    .Q(\bg_object_inst.bg_object_pos[3] ));
 sg13g2_dfrbp_1 _5155_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net40),
    .D(net762),
    .Q_N(_2471_),
    .Q(\bg_object_inst.bg_object_pos[4] ));
 sg13g2_dfrbp_1 _5156_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net38),
    .D(_0107_),
    .Q_N(_2470_),
    .Q(\bg_object_inst.bg_object_pos[5] ));
 sg13g2_dfrbp_1 _5157_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net34),
    .D(_0108_),
    .Q_N(_2469_),
    .Q(\bg_object_inst.bg_object_pos[6] ));
 sg13g2_dfrbp_1 _5158_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net32),
    .D(net854),
    .Q_N(_2468_),
    .Q(\bg_object_inst.bg_object_pos[7] ));
 sg13g2_dfrbp_1 _5159_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net30),
    .D(_0110_),
    .Q_N(_2467_),
    .Q(\bg_object_inst.bg_object_pos[8] ));
 sg13g2_dfrbp_1 _5160_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net28),
    .D(net738),
    .Q_N(_2466_),
    .Q(\bg_object_inst.bg_object_pos[9] ));
 sg13g2_dfrbp_1 _5161_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net26),
    .D(_0112_),
    .Q_N(_2465_),
    .Q(\dino_inst.x_offset_r[5] ));
 sg13g2_dfrbp_1 _5162_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net25),
    .D(_0113_),
    .Q_N(_2464_),
    .Q(\dino_inst.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5163_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net24),
    .D(_0114_),
    .Q_N(_2463_),
    .Q(\dino_inst.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5164_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net23),
    .D(_0115_),
    .Q_N(_2462_),
    .Q(\dino_inst.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5165_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net22),
    .D(_0116_),
    .Q_N(_2461_),
    .Q(\dino_inst.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5166_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net21),
    .D(_0117_),
    .Q_N(_2460_),
    .Q(\audio_inst.i_jump.decay_value[16] ));
 sg13g2_dfrbp_1 _5167_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net19),
    .D(_0118_),
    .Q_N(_2459_),
    .Q(\obs_inst_2.o_rom_counter[0] ));
 sg13g2_dfrbp_1 _5168_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net18),
    .D(_0119_),
    .Q_N(_2458_),
    .Q(\obs_inst_2.o_rom_counter[1] ));
 sg13g2_dfrbp_1 _5169_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net383),
    .D(_0120_),
    .Q_N(_2457_),
    .Q(\obs_inst_2.o_rom_counter[2] ));
 sg13g2_dfrbp_1 _5170_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net382),
    .D(_0121_),
    .Q_N(_2456_),
    .Q(\obs_inst_2.o_rom_counter[3] ));
 sg13g2_dfrbp_1 _5171_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net381),
    .D(_0122_),
    .Q_N(_2455_),
    .Q(\obs_inst_2.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5172_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net380),
    .D(_0123_),
    .Q_N(_2454_),
    .Q(\obs_inst_2.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5173_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net379),
    .D(_0124_),
    .Q_N(_2453_),
    .Q(\obs_inst_2.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5174_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net378),
    .D(_0125_),
    .Q_N(_2452_),
    .Q(\obs_inst_2.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5175_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net377),
    .D(_0126_),
    .Q_N(_0034_),
    .Q(\audio_inst.i_jump.counter[0] ));
 sg13g2_dfrbp_1 _5176_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net375),
    .D(net832),
    .Q_N(_2451_),
    .Q(\audio_inst.i_jump.counter[1] ));
 sg13g2_dfrbp_1 _5177_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net373),
    .D(_0128_),
    .Q_N(_2450_),
    .Q(\audio_inst.i_jump.counter[2] ));
 sg13g2_dfrbp_1 _5178_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net371),
    .D(_0129_),
    .Q_N(_2449_),
    .Q(\audio_inst.i_jump.counter[3] ));
 sg13g2_dfrbp_1 _5179_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net369),
    .D(net806),
    .Q_N(_2448_),
    .Q(\audio_inst.i_jump.counter[4] ));
 sg13g2_dfrbp_1 _5180_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net367),
    .D(net788),
    .Q_N(_2447_),
    .Q(\audio_inst.i_jump.counter[5] ));
 sg13g2_dfrbp_1 _5181_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net365),
    .D(net686),
    .Q_N(_2446_),
    .Q(\audio_inst.i_jump.counter[6] ));
 sg13g2_dfrbp_1 _5182_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net363),
    .D(net635),
    .Q_N(_2445_),
    .Q(\audio_inst.i_jump.counter[7] ));
 sg13g2_dfrbp_1 _5183_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net361),
    .D(_0134_),
    .Q_N(_2444_),
    .Q(\audio_inst.i_jump.counter[8] ));
 sg13g2_dfrbp_1 _5184_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net359),
    .D(net770),
    .Q_N(_2443_),
    .Q(\audio_inst.i_jump.counter[9] ));
 sg13g2_dfrbp_1 _5185_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net357),
    .D(_0136_),
    .Q_N(_2442_),
    .Q(\audio_inst.i_jump.counter[10] ));
 sg13g2_dfrbp_1 _5186_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net355),
    .D(_0137_),
    .Q_N(_2441_),
    .Q(\audio_inst.i_jump.counter[11] ));
 sg13g2_dfrbp_1 _5187_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net353),
    .D(net916),
    .Q_N(_2440_),
    .Q(\audio_inst.i_jump.counter[12] ));
 sg13g2_dfrbp_1 _5188_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net351),
    .D(net743),
    .Q_N(_2439_),
    .Q(\audio_inst.i_jump.counter[13] ));
 sg13g2_dfrbp_1 _5189_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net349),
    .D(_0140_),
    .Q_N(_2438_),
    .Q(\audio_inst.i_jump.counter[14] ));
 sg13g2_dfrbp_1 _5190_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net347),
    .D(net776),
    .Q_N(_2437_),
    .Q(\audio_inst.i_jump.counter[15] ));
 sg13g2_dfrbp_1 _5191_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net345),
    .D(_0142_),
    .Q_N(_2436_),
    .Q(\audio_inst.i_jump.counter[16] ));
 sg13g2_dfrbp_1 _5192_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net343),
    .D(net755),
    .Q_N(_2435_),
    .Q(\audio_inst.i_jump.counter[17] ));
 sg13g2_dfrbp_1 _5193_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net341),
    .D(_0144_),
    .Q_N(_2434_),
    .Q(\audio_inst.i_jump.counter[18] ));
 sg13g2_dfrbp_1 _5194_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net339),
    .D(net460),
    .Q_N(_2433_),
    .Q(\audio_inst.i_over.decay_value[0] ));
 sg13g2_dfrbp_1 _5195_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net338),
    .D(net456),
    .Q_N(_2432_),
    .Q(\audio_inst.i_over.decay_value[1] ));
 sg13g2_dfrbp_1 _5196_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net337),
    .D(_0147_),
    .Q_N(_2431_),
    .Q(\audio_inst.i_over.decay_value[2] ));
 sg13g2_dfrbp_1 _5197_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net336),
    .D(_0148_),
    .Q_N(_2430_),
    .Q(\audio_inst.i_over.decay_value[3] ));
 sg13g2_dfrbp_1 _5198_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net335),
    .D(_0149_),
    .Q_N(_2429_),
    .Q(\audio_inst.i_over.decay_value[4] ));
 sg13g2_dfrbp_1 _5199_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net334),
    .D(_0150_),
    .Q_N(_2428_),
    .Q(\audio_inst.i_over.decay_value[5] ));
 sg13g2_dfrbp_1 _5200_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net333),
    .D(_0151_),
    .Q_N(_2427_),
    .Q(\audio_inst.i_over.decay_value[6] ));
 sg13g2_dfrbp_1 _5201_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net332),
    .D(_0152_),
    .Q_N(_2426_),
    .Q(\audio_inst.i_over.decay_value[7] ));
 sg13g2_dfrbp_1 _5202_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net331),
    .D(_0153_),
    .Q_N(_2425_),
    .Q(\audio_inst.i_over.decay_value[8] ));
 sg13g2_dfrbp_1 _5203_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net330),
    .D(_0154_),
    .Q_N(_2424_),
    .Q(\audio_inst.i_over.decay_value[9] ));
 sg13g2_dfrbp_1 _5204_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net329),
    .D(net764),
    .Q_N(_2423_),
    .Q(\audio_inst.i_over.decay_value[10] ));
 sg13g2_dfrbp_1 _5205_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net328),
    .D(net773),
    .Q_N(_2422_),
    .Q(\audio_inst.i_over.decay_value[11] ));
 sg13g2_dfrbp_1 _5206_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net327),
    .D(_0157_),
    .Q_N(_2421_),
    .Q(\audio_inst.i_over.decay_value[12] ));
 sg13g2_dfrbp_1 _5207_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net320),
    .D(_0158_),
    .Q_N(_2420_),
    .Q(\audio_inst.i_over.decay_value[13] ));
 sg13g2_dfrbp_1 _5208_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net319),
    .D(_0159_),
    .Q_N(_2419_),
    .Q(\audio_inst.i_over.decay_value[14] ));
 sg13g2_dfrbp_1 _5209_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net318),
    .D(_0160_),
    .Q_N(_2418_),
    .Q(\audio_inst.i_over.decay_value[15] ));
 sg13g2_dfrbp_1 _5210_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net317),
    .D(net753),
    .Q_N(_2417_),
    .Q(\audio_inst.i_jump.decay_value[14] ));
 sg13g2_dfrbp_1 _5211_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net315),
    .D(net445),
    .Q_N(_2416_),
    .Q(\audio_inst.i_jump.decay_value[15] ));
 sg13g2_dfrbp_1 _5212_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net313),
    .D(_0163_),
    .Q_N(_2415_),
    .Q(\audio_inst.i_jump.decay_value[0] ));
 sg13g2_dfrbp_1 _5213_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net312),
    .D(_0164_),
    .Q_N(_2414_),
    .Q(\audio_inst.i_jump.decay_value[1] ));
 sg13g2_dfrbp_1 _5214_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net311),
    .D(_0165_),
    .Q_N(_2413_),
    .Q(\audio_inst.i_jump.decay_value[2] ));
 sg13g2_dfrbp_1 _5215_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net310),
    .D(_0166_),
    .Q_N(_2412_),
    .Q(\audio_inst.i_jump.decay_value[3] ));
 sg13g2_dfrbp_1 _5216_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net309),
    .D(_0167_),
    .Q_N(_2411_),
    .Q(\audio_inst.i_jump.decay_value[4] ));
 sg13g2_dfrbp_1 _5217_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net308),
    .D(_0168_),
    .Q_N(_2410_),
    .Q(\audio_inst.i_jump.decay_value[5] ));
 sg13g2_dfrbp_1 _5218_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net307),
    .D(_0169_),
    .Q_N(_2409_),
    .Q(\audio_inst.i_jump.decay_value[6] ));
 sg13g2_dfrbp_1 _5219_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net306),
    .D(_0170_),
    .Q_N(_2408_),
    .Q(\audio_inst.i_jump.decay_value[7] ));
 sg13g2_dfrbp_1 _5220_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net305),
    .D(_0171_),
    .Q_N(_2407_),
    .Q(\audio_inst.i_jump.decay_value[8] ));
 sg13g2_dfrbp_1 _5221_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net304),
    .D(_0172_),
    .Q_N(_2406_),
    .Q(\audio_inst.i_jump.decay_value[9] ));
 sg13g2_dfrbp_1 _5222_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net303),
    .D(_0173_),
    .Q_N(_2405_),
    .Q(\audio_inst.i_jump.decay_value[10] ));
 sg13g2_dfrbp_1 _5223_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net302),
    .D(net698),
    .Q_N(_2404_),
    .Q(\audio_inst.i_jump.decay_value[11] ));
 sg13g2_dfrbp_1 _5224_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net301),
    .D(_0175_),
    .Q_N(_2403_),
    .Q(\audio_inst.i_jump.decay_value[12] ));
 sg13g2_dfrbp_1 _5225_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net300),
    .D(_0176_),
    .Q_N(_2402_),
    .Q(\audio_inst.i_jump.decay_value[13] ));
 sg13g2_dfrbp_1 _5226_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net299),
    .D(net434),
    .Q_N(_2401_),
    .Q(\audio_inst.i_over.state[0] ));
 sg13g2_dfrbp_1 _5227_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net298),
    .D(_0178_),
    .Q_N(_2400_),
    .Q(\score_inst_1.x_offset_r[4] ));
 sg13g2_dfrbp_1 _5228_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net297),
    .D(_0179_),
    .Q_N(_2399_),
    .Q(\score_inst_1.x_offset_r[5] ));
 sg13g2_dfrbp_1 _5229_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net296),
    .D(_0180_),
    .Q_N(_2398_),
    .Q(\score_inst_1.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5230_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net295),
    .D(_0181_),
    .Q_N(_2397_),
    .Q(\score_inst_1.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5231_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net294),
    .D(_0182_),
    .Q_N(_2396_),
    .Q(\score_inst_1.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5232_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net293),
    .D(_0183_),
    .Q_N(_2395_),
    .Q(\score_inst_1.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5233_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net292),
    .D(_0184_),
    .Q_N(_2394_),
    .Q(\score_inst_1.y_offset_r[5] ));
 sg13g2_dfrbp_1 _5234_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net291),
    .D(_0185_),
    .Q_N(_2393_),
    .Q(\score_inst_1.y_offset_r[6] ));
 sg13g2_dfrbp_1 _5235_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net290),
    .D(_0186_),
    .Q_N(_2392_),
    .Q(\score_inst_1.y_offset_r[7] ));
 sg13g2_dfrbp_1 _5236_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net289),
    .D(_0187_),
    .Q_N(_2391_),
    .Q(\score_inst_1.y_offset_r[8] ));
 sg13g2_dfrbp_1 _5237_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net288),
    .D(_0188_),
    .Q_N(_2390_),
    .Q(\score_inst_1.y_offset_r[9] ));
 sg13g2_dfrbp_1 _5238_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net287),
    .D(_0189_),
    .Q_N(_2389_),
    .Q(\score_inst_2.x_offset_r[3] ));
 sg13g2_dfrbp_1 _5239_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net286),
    .D(_0190_),
    .Q_N(_2388_),
    .Q(\score_inst_2.x_offset_r[4] ));
 sg13g2_dfrbp_1 _5240_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net285),
    .D(_0191_),
    .Q_N(_2387_),
    .Q(\score_inst_2.x_offset_r[5] ));
 sg13g2_dfrbp_1 _5241_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net284),
    .D(_0192_),
    .Q_N(_2386_),
    .Q(\score_inst_2.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5242_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net283),
    .D(_0193_),
    .Q_N(_2385_),
    .Q(\score_inst_2.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5243_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net282),
    .D(_0194_),
    .Q_N(_2384_),
    .Q(\score_inst_2.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5244_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net281),
    .D(_0195_),
    .Q_N(_2383_),
    .Q(\score_inst_2.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5245_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net280),
    .D(_0196_),
    .Q_N(_2382_),
    .Q(\score_inst_1.num_r[0] ));
 sg13g2_dfrbp_1 _5246_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net279),
    .D(_0197_),
    .Q_N(_2381_),
    .Q(\score_inst_1.num_r[1] ));
 sg13g2_dfrbp_1 _5247_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net278),
    .D(_0198_),
    .Q_N(_2380_),
    .Q(\score_inst_1.num_r[2] ));
 sg13g2_dfrbp_1 _5248_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net277),
    .D(_0199_),
    .Q_N(_2379_),
    .Q(\score_inst_1.num_r[3] ));
 sg13g2_dfrbp_1 _5249_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net276),
    .D(_0200_),
    .Q_N(_2378_),
    .Q(\dino_inst.o_rom_counter[1] ));
 sg13g2_dfrbp_1 _5250_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net275),
    .D(_0201_),
    .Q_N(_2377_),
    .Q(\dino_inst.o_rom_counter[2] ));
 sg13g2_dfrbp_1 _5251_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net274),
    .D(_0202_),
    .Q_N(_2376_),
    .Q(\score_inst_3.x_offset_r[5] ));
 sg13g2_dfrbp_1 _5252_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net273),
    .D(_0203_),
    .Q_N(_2375_),
    .Q(\score_inst_3.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5253_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net272),
    .D(_0204_),
    .Q_N(_2374_),
    .Q(\score_inst_3.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5254_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net271),
    .D(_0205_),
    .Q_N(_2373_),
    .Q(\score_inst_3.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5255_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net270),
    .D(_0206_),
    .Q_N(_2372_),
    .Q(\score_inst_3.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5256_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net269),
    .D(_0207_),
    .Q_N(_2371_),
    .Q(\score_inst_2.num_r[0] ));
 sg13g2_dfrbp_1 _5257_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net268),
    .D(_0208_),
    .Q_N(_2370_),
    .Q(\score_inst_2.num_r[1] ));
 sg13g2_dfrbp_1 _5258_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net267),
    .D(_0209_),
    .Q_N(_2369_),
    .Q(\score_inst_2.num_r[2] ));
 sg13g2_dfrbp_1 _5259_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net266),
    .D(_0210_),
    .Q_N(_2368_),
    .Q(\score_inst_2.num_r[3] ));
 sg13g2_dfrbp_1 _5260_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net265),
    .D(_0211_),
    .Q_N(_2367_),
    .Q(\score_inst_2.x_offset_r[2] ));
 sg13g2_dfrbp_1 _5261_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net264),
    .D(_0212_),
    .Q_N(_2366_),
    .Q(\score_inst_4.x_offset_r[3] ));
 sg13g2_dfrbp_1 _5262_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net263),
    .D(_0213_),
    .Q_N(_2365_),
    .Q(\score_inst_4.x_offset_r[4] ));
 sg13g2_dfrbp_1 _5263_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net262),
    .D(_0214_),
    .Q_N(_2364_),
    .Q(\score_inst_4.x_offset_r[5] ));
 sg13g2_dfrbp_1 _5264_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net261),
    .D(_0215_),
    .Q_N(_2363_),
    .Q(\score_inst_4.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5265_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net260),
    .D(_0216_),
    .Q_N(_2362_),
    .Q(\score_inst_4.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5266_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net259),
    .D(_0217_),
    .Q_N(_2361_),
    .Q(\score_inst_4.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5267_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net258),
    .D(_0218_),
    .Q_N(_2360_),
    .Q(\score_inst_4.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5268_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net257),
    .D(_0219_),
    .Q_N(_2359_),
    .Q(\score_inst_3.num_r[0] ));
 sg13g2_dfrbp_1 _5269_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net256),
    .D(_0220_),
    .Q_N(_2358_),
    .Q(\score_inst_3.num_r[1] ));
 sg13g2_dfrbp_1 _5270_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net255),
    .D(_0221_),
    .Q_N(_2357_),
    .Q(\score_inst_3.num_r[2] ));
 sg13g2_dfrbp_1 _5271_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net254),
    .D(_0222_),
    .Q_N(_2356_),
    .Q(\score_inst_3.num_r[3] ));
 sg13g2_dfrbp_1 _5272_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net253),
    .D(_0223_),
    .Q_N(_2355_),
    .Q(\dino_inst.o_rom_counter[0] ));
 sg13g2_dfrbp_1 _5273_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net252),
    .D(_0224_),
    .Q_N(_2354_),
    .Q(\score_inst_1.x_offset_r[3] ));
 sg13g2_dfrbp_1 _5274_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net251),
    .D(_0225_),
    .Q_N(_2353_),
    .Q(\score_inst_5.x_offset_r[4] ));
 sg13g2_dfrbp_1 _5275_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net250),
    .D(_0226_),
    .Q_N(_2352_),
    .Q(\score_inst_5.x_offset_r[5] ));
 sg13g2_dfrbp_1 _5276_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net249),
    .D(_0227_),
    .Q_N(_2351_),
    .Q(\score_inst_5.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5277_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net248),
    .D(_0228_),
    .Q_N(_2350_),
    .Q(\score_inst_5.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5278_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net247),
    .D(_0229_),
    .Q_N(_2349_),
    .Q(\score_inst_5.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5279_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net246),
    .D(net692),
    .Q_N(_2348_),
    .Q(\score_inst_5.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5280_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net245),
    .D(_0231_),
    .Q_N(_2347_),
    .Q(\score_inst_4.num_r[0] ));
 sg13g2_dfrbp_1 _5281_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net244),
    .D(_0232_),
    .Q_N(_2346_),
    .Q(\score_inst_4.num_r[1] ));
 sg13g2_dfrbp_1 _5282_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net243),
    .D(_0233_),
    .Q_N(_2345_),
    .Q(\score_inst_4.num_r[2] ));
 sg13g2_dfrbp_1 _5283_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net242),
    .D(_0234_),
    .Q_N(_2344_),
    .Q(\score_inst_4.num_r[3] ));
 sg13g2_dfrbp_1 _5284_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net241),
    .D(_0235_),
    .Q_N(_2343_),
    .Q(\dino_inst.o_rom_counter[3] ));
 sg13g2_dfrbp_1 _5285_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net240),
    .D(_0236_),
    .Q_N(_2342_),
    .Q(\dino_inst.o_rom_counter[4] ));
 sg13g2_dfrbp_1 _5286_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net239),
    .D(_0237_),
    .Q_N(_0014_),
    .Q(\dino_inst.o_rom_counter[5] ));
 sg13g2_dfrbp_1 _5287_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net238),
    .D(_0238_),
    .Q_N(_2341_),
    .Q(\dino_inst.y_offset_r[5] ));
 sg13g2_dfrbp_1 _5288_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net237),
    .D(_0239_),
    .Q_N(_2340_),
    .Q(\dino_inst.y_offset_r[6] ));
 sg13g2_dfrbp_1 _5289_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net236),
    .D(_0240_),
    .Q_N(_2339_),
    .Q(\dino_inst.y_offset_r[7] ));
 sg13g2_dfrbp_1 _5290_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net235),
    .D(_0241_),
    .Q_N(_2338_),
    .Q(\dino_inst.y_offset_r[8] ));
 sg13g2_dfrbp_1 _5291_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net234),
    .D(_0242_),
    .Q_N(_2337_),
    .Q(\dino_inst.y_offset_r[9] ));
 sg13g2_dfrbp_1 _5292_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net233),
    .D(_0243_),
    .Q_N(_2336_),
    .Q(\bg_object_rom_inst.i_rom_counter[0] ));
 sg13g2_dfrbp_1 _5293_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net232),
    .D(_0244_),
    .Q_N(_2335_),
    .Q(\bg_object_rom_inst.i_rom_counter[1] ));
 sg13g2_dfrbp_1 _5294_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net231),
    .D(_0245_),
    .Q_N(_2334_),
    .Q(\bg_object_rom_inst.i_rom_counter[2] ));
 sg13g2_dfrbp_1 _5295_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net230),
    .D(_0246_),
    .Q_N(_2333_),
    .Q(\bg_render_inst.x_offset_r[5] ));
 sg13g2_dfrbp_1 _5296_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net229),
    .D(_0247_),
    .Q_N(_2332_),
    .Q(\bg_render_inst.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5297_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net228),
    .D(_0248_),
    .Q_N(_2331_),
    .Q(\bg_render_inst.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5298_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net227),
    .D(_0249_),
    .Q_N(_2330_),
    .Q(\bg_render_inst.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5299_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net226),
    .D(_0250_),
    .Q_N(_2329_),
    .Q(\bg_render_inst.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5300_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net225),
    .D(_0251_),
    .Q_N(_2328_),
    .Q(\obs_inst_1.o_rom_counter[4] ));
 sg13g2_dfrbp_1 _5301_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net224),
    .D(_0252_),
    .Q_N(_2327_),
    .Q(\obs_inst_1.o_rom_counter[5] ));
 sg13g2_dfrbp_1 _5302_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net223),
    .D(_0253_),
    .Q_N(_2326_),
    .Q(\obs_inst_1.o_rom_counter[6] ));
 sg13g2_dfrbp_1 _5303_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net222),
    .D(_0254_),
    .Q_N(_2325_),
    .Q(\obs_inst_1.o_rom_counter[7] ));
 sg13g2_dfrbp_1 _5304_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net221),
    .D(_0255_),
    .Q_N(_2324_),
    .Q(\obs_inst_1.y_offset_r[6] ));
 sg13g2_dfrbp_1 _5305_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net220),
    .D(_0256_),
    .Q_N(_2323_),
    .Q(\obs_inst_1.y_offset_r[7] ));
 sg13g2_dfrbp_1 _5306_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net219),
    .D(_0257_),
    .Q_N(_2322_),
    .Q(\obs_inst_1.y_offset_r[8] ));
 sg13g2_dfrbp_1 _5307_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net218),
    .D(_0258_),
    .Q_N(_2321_),
    .Q(\obs_inst_1.y_offset_r[9] ));
 sg13g2_dfrbp_1 _5308_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net217),
    .D(_0259_),
    .Q_N(_2320_),
    .Q(\lfsr_inst.r_lfsr[1] ));
 sg13g2_dfrbp_1 _5309_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net216),
    .D(_0260_),
    .Q_N(_2319_),
    .Q(\lfsr_inst.r_lfsr[2] ));
 sg13g2_dfrbp_1 _5310_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net215),
    .D(_0261_),
    .Q_N(_2318_),
    .Q(\lfsr_inst.r_lfsr[3] ));
 sg13g2_dfrbp_1 _5311_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net214),
    .D(_0262_),
    .Q_N(_2317_),
    .Q(\lfsr_inst.r_lfsr[4] ));
 sg13g2_dfrbp_1 _5312_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net213),
    .D(_0263_),
    .Q_N(_2316_),
    .Q(\lfsr_inst.r_lfsr[5] ));
 sg13g2_dfrbp_1 _5313_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net212),
    .D(_0264_),
    .Q_N(_2315_),
    .Q(\lfsr_inst.r_lfsr[6] ));
 sg13g2_dfrbp_1 _5314_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net211),
    .D(_0265_),
    .Q_N(_2314_),
    .Q(\lfsr_inst.r_lfsr[7] ));
 sg13g2_dfrbp_1 _5315_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net210),
    .D(_0266_),
    .Q_N(_2313_),
    .Q(\lfsr_inst.r_lfsr[8] ));
 sg13g2_dfrbp_1 _5316_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net209),
    .D(_0267_),
    .Q_N(_2312_),
    .Q(\lfsr_inst.r_lfsr[9] ));
 sg13g2_dfrbp_1 _5317_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net208),
    .D(_0268_),
    .Q_N(_2311_),
    .Q(\lfsr_inst.r_lfsr[10] ));
 sg13g2_dfrbp_1 _5318_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net207),
    .D(_0269_),
    .Q_N(_2310_),
    .Q(\lfsr_inst.r_lfsr[11] ));
 sg13g2_dfrbp_1 _5319_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net206),
    .D(_0270_),
    .Q_N(_2309_),
    .Q(\lfsr_inst.r_lfsr[12] ));
 sg13g2_dfrbp_1 _5320_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net205),
    .D(_0271_),
    .Q_N(_2308_),
    .Q(\lfsr_inst.r_lfsr[13] ));
 sg13g2_dfrbp_1 _5321_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net204),
    .D(_0272_),
    .Q_N(_2307_),
    .Q(\lfsr_inst.r_lfsr[14] ));
 sg13g2_dfrbp_1 _5322_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net203),
    .D(_0273_),
    .Q_N(_2306_),
    .Q(\lfsr_inst.r_lfsr[15] ));
 sg13g2_dfrbp_1 _5323_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net202),
    .D(_0274_),
    .Q_N(_2305_),
    .Q(\obs_inst_1.o_rom_counter[0] ));
 sg13g2_dfrbp_1 _5324_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net201),
    .D(_0275_),
    .Q_N(_2304_),
    .Q(\obs_inst_1.o_rom_counter[1] ));
 sg13g2_dfrbp_1 _5325_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net200),
    .D(_0276_),
    .Q_N(_2303_),
    .Q(\obs_inst_1.o_rom_counter[2] ));
 sg13g2_dfrbp_1 _5326_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net199),
    .D(_0277_),
    .Q_N(_2302_),
    .Q(\obs_inst_1.o_rom_counter[3] ));
 sg13g2_dfrbp_1 _5327_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net198),
    .D(_0278_),
    .Q_N(_2301_),
    .Q(\obs_inst_1.x_offset_r[6] ));
 sg13g2_dfrbp_1 _5328_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net197),
    .D(_0279_),
    .Q_N(_2300_),
    .Q(\obs_inst_1.x_offset_r[7] ));
 sg13g2_dfrbp_1 _5329_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net196),
    .D(_0280_),
    .Q_N(_2299_),
    .Q(\obs_inst_1.x_offset_r[8] ));
 sg13g2_dfrbp_1 _5330_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net195),
    .D(_0281_),
    .Q_N(_2298_),
    .Q(\obs_inst_1.x_offset_r[9] ));
 sg13g2_dfrbp_1 _5331_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net194),
    .D(_0282_),
    .Q_N(_2297_),
    .Q(\bg_object_rom_inst.i_rom_counter[3] ));
 sg13g2_dfrbp_1 _5332_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net193),
    .D(_0283_),
    .Q_N(_0025_),
    .Q(\bg_object_rom_inst.i_rom_counter[4] ));
 sg13g2_dfrbp_1 _5333_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net192),
    .D(_0284_),
    .Q_N(_0024_),
    .Q(\bg_object_rom_inst.i_rom_counter[5] ));
 sg13g2_dfrbp_1 _5334_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net191),
    .D(_0285_),
    .Q_N(_2296_),
    .Q(\bg_render_inst.y_offset_r[5] ));
 sg13g2_dfrbp_1 _5335_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net190),
    .D(_0286_),
    .Q_N(_2295_),
    .Q(\bg_render_inst.y_offset_r[6] ));
 sg13g2_dfrbp_1 _5336_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net189),
    .D(_0287_),
    .Q_N(_2294_),
    .Q(\bg_render_inst.y_offset_r[7] ));
 sg13g2_dfrbp_1 _5337_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net188),
    .D(_0288_),
    .Q_N(_2293_),
    .Q(\bg_render_inst.y_offset_r[8] ));
 sg13g2_dfrbp_1 _5338_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net187),
    .D(_0289_),
    .Q_N(_2292_),
    .Q(\bg_render_inst.y_offset_r[9] ));
 sg13g2_dfrbp_1 _5339_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net186),
    .D(net393),
    .Q_N(_0033_),
    .Q(\graphics_inst.hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _5340_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net184),
    .D(_0291_),
    .Q_N(_2291_),
    .Q(\graphics_inst.hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _5341_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net182),
    .D(_0292_),
    .Q_N(\bg_render_inst.y_offset[2] ),
    .Q(\bg_line_inst.i_vpos[2] ));
 sg13g2_dfrbp_1 _5342_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net180),
    .D(_0293_),
    .Q_N(\obs_inst_1.y_offset[3] ),
    .Q(\bg_line_inst.i_vpos[3] ));
 sg13g2_dfrbp_1 _5343_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net178),
    .D(_0294_),
    .Q_N(_2290_),
    .Q(\bg_line_inst.i_vpos[4] ));
 sg13g2_dfrbp_1 _5344_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net176),
    .D(_0295_),
    .Q_N(_0011_),
    .Q(\bg_line_inst.i_vpos[5] ));
 sg13g2_dfrbp_1 _5345_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net174),
    .D(_0296_),
    .Q_N(_0031_),
    .Q(\bg_line_inst.i_vpos[6] ));
 sg13g2_dfrbp_1 _5346_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net172),
    .D(_0297_),
    .Q_N(_2289_),
    .Q(\bg_line_inst.i_vpos[7] ));
 sg13g2_dfrbp_1 _5347_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net170),
    .D(_0298_),
    .Q_N(_0032_),
    .Q(\bg_line_inst.i_vpos[8] ));
 sg13g2_dfrbp_1 _5348_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net168),
    .D(_0299_),
    .Q_N(_2288_),
    .Q(\bg_line_inst.i_vpos[9] ));
 sg13g2_dfrbp_1 _5349_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net166),
    .D(_0300_),
    .Q_N(_2287_),
    .Q(\graphics_inst.display_on_r_r ));
 sg13g2_dfrbp_1 _5350_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net165),
    .D(_0301_),
    .Q_N(_2286_),
    .Q(\graphics_inst.display_on_r ));
 sg13g2_dfrbp_1 _5351_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net164),
    .D(_0302_),
    .Q_N(_2285_),
    .Q(\graphics_inst.o_vsync ));
 sg13g2_dfrbp_1 _5352_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net163),
    .D(_0303_),
    .Q_N(_2284_),
    .Q(\graphics_inst.hsync_r_r ));
 sg13g2_dfrbp_1 _5353_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net162),
    .D(_0304_),
    .Q_N(_2283_),
    .Q(\graphics_inst.vsync_r ));
 sg13g2_dfrbp_1 _5354_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net161),
    .D(_0305_),
    .Q_N(_2282_),
    .Q(\graphics_inst.hsync_r ));
 sg13g2_dfrbp_1 _5355_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net160),
    .D(_0306_),
    .Q_N(_2281_),
    .Q(\graphics_inst.B_r[0] ));
 sg13g2_dfrbp_1 _5356_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net159),
    .D(_0307_),
    .Q_N(_2280_),
    .Q(\graphics_inst.B_r[1] ));
 sg13g2_dfrbp_1 _5357_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net141),
    .D(_0308_),
    .Q_N(_2279_),
    .Q(\graphics_inst.G_r[0] ));
 sg13g2_dfrbp_1 _5358_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net139),
    .D(_0309_),
    .Q_N(_2278_),
    .Q(\graphics_inst.G_r[1] ));
 sg13g2_dfrbp_1 _5359_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net137),
    .D(_0310_),
    .Q_N(_2277_),
    .Q(\graphics_inst.R_r[1] ));
 sg13g2_dfrbp_1 _5360_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net135),
    .D(_0311_),
    .Q_N(_2276_),
    .Q(\graphics_inst.game_tick_r ));
 sg13g2_dfrbp_1 _5361_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net133),
    .D(_0312_),
    .Q_N(_2275_),
    .Q(\ai_controller_inst.crash ));
 sg13g2_dfrbp_1 _5362_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net129),
    .D(_0313_),
    .Q_N(_2274_),
    .Q(\gamepad_pmod.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _5363_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net127),
    .D(_0314_),
    .Q_N(_2273_),
    .Q(\gamepad_pmod.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _5364_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net125),
    .D(_0315_),
    .Q_N(_2272_),
    .Q(\graphics_inst.frame_counter[0] ));
 sg13g2_dfrbp_1 _5365_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net121),
    .D(_0316_),
    .Q_N(_2271_),
    .Q(\graphics_inst.frame_counter[1] ));
 sg13g2_dfrbp_1 _5366_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net117),
    .D(_0317_),
    .Q_N(_2270_),
    .Q(\score[16] ));
 sg13g2_dfrbp_1 _5367_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net109),
    .D(_0318_),
    .Q_N(_2269_),
    .Q(\score[17] ));
 sg13g2_dfrbp_1 _5368_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net105),
    .D(_0319_),
    .Q_N(_2268_),
    .Q(\score[18] ));
 sg13g2_dfrbp_1 _5369_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net101),
    .D(_0320_),
    .Q_N(_2267_),
    .Q(\score[19] ));
 sg13g2_dfrbp_1 _5370_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net97),
    .D(_0321_),
    .Q_N(_2266_),
    .Q(\score[12] ));
 sg13g2_dfrbp_1 _5371_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net93),
    .D(_0322_),
    .Q_N(_2265_),
    .Q(\score[13] ));
 sg13g2_dfrbp_1 _5372_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net89),
    .D(_0323_),
    .Q_N(_2264_),
    .Q(\graphics_inst.color_decoder_inst.rgb_scheme ));
 sg13g2_dfrbp_1 _5373_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net85),
    .D(_0324_),
    .Q_N(_2263_),
    .Q(\score[15] ));
 sg13g2_dfrbp_1 _5374_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net81),
    .D(_0325_),
    .Q_N(_2262_),
    .Q(\score[8] ));
 sg13g2_dfrbp_1 _5375_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net77),
    .D(_0326_),
    .Q_N(_2261_),
    .Q(\score[9] ));
 sg13g2_dfrbp_1 _5376_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net73),
    .D(_0327_),
    .Q_N(_0023_),
    .Q(\graphics_inst.color_decoder_inst.invert ));
 sg13g2_dfrbp_1 _5377_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net69),
    .D(_0328_),
    .Q_N(_2260_),
    .Q(\score[11] ));
 sg13g2_dfrbp_1 _5378_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net65),
    .D(_0329_),
    .Q_N(_2259_),
    .Q(\score[4] ));
 sg13g2_dfrbp_1 _5379_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net61),
    .D(_0330_),
    .Q_N(_2258_),
    .Q(\score[5] ));
 sg13g2_dfrbp_1 _5380_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net57),
    .D(_0331_),
    .Q_N(_2257_),
    .Q(\score[6] ));
 sg13g2_dfrbp_1 _5381_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net53),
    .D(_0332_),
    .Q_N(_2256_),
    .Q(\score[7] ));
 sg13g2_dfrbp_1 _5382_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net49),
    .D(_0333_),
    .Q_N(_2255_),
    .Q(\score[0] ));
 sg13g2_dfrbp_1 _5383_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net45),
    .D(_0334_),
    .Q_N(_2254_),
    .Q(\score[1] ));
 sg13g2_dfrbp_1 _5384_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net41),
    .D(_0335_),
    .Q_N(_2253_),
    .Q(\score[2] ));
 sg13g2_dfrbp_1 _5385_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net322),
    .D(_0336_),
    .Q_N(_2531_),
    .Q(\score[3] ));
 sg13g2_dfrbp_1 _5386_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net323),
    .D(_0000_),
    .Q_N(_2532_),
    .Q(\player_constroller_inst.game_state[0] ));
 sg13g2_dfrbp_1 _5387_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net324),
    .D(net796),
    .Q_N(_0015_),
    .Q(\player_constroller_inst.game_state[1] ));
 sg13g2_dfrbp_1 _5388_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net325),
    .D(net844),
    .Q_N(_2533_),
    .Q(\player_constroller_inst.game_state[2] ));
 sg13g2_dfrbp_1 _5389_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net326),
    .D(net840),
    .Q_N(_2534_),
    .Q(\player_constroller_inst.game_state[3] ));
 sg13g2_dfrbp_1 _5390_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net75),
    .D(_0004_),
    .Q_N(_2535_),
    .Q(\player_constroller_inst.game_over ));
 sg13g2_dfrbp_1 _5391_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net35),
    .D(_0005_),
    .Q_N(_2252_),
    .Q(\player_constroller_inst.game_state[5] ));
 sg13g2_dfrbp_1 _5392_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net31),
    .D(net467),
    .Q_N(_2251_),
    .Q(\audio_inst.game_over_sound ));
 sg13g2_dfrbp_1 _5393_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net27),
    .D(_0338_),
    .Q_N(_0028_),
    .Q(\audio_inst.i_over.stage_index[0] ));
 sg13g2_dfrbp_1 _5394_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net376),
    .D(_0339_),
    .Q_N(_0027_),
    .Q(\audio_inst.i_over.stage_index[1] ));
 sg13g2_dfrbp_1 _5395_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net372),
    .D(_0340_),
    .Q_N(_0008_),
    .Q(\audio_inst.i_over.stage_index[2] ));
 sg13g2_dfrbp_1 _5396_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net368),
    .D(_0341_),
    .Q_N(_0009_),
    .Q(\audio_inst.i_over.stage_index[3] ));
 sg13g2_dfrbp_1 _5397_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net364),
    .D(net783),
    .Q_N(_0026_),
    .Q(\audio_inst.i_over.stage_index[4] ));
 sg13g2_dfrbp_1 _5398_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net360),
    .D(net786),
    .Q_N(_2250_),
    .Q(\audio_inst.i_over.counter[0] ));
 sg13g2_dfrbp_1 _5399_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net356),
    .D(_0344_),
    .Q_N(_2249_),
    .Q(\audio_inst.i_over.counter[1] ));
 sg13g2_dfrbp_1 _5400_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net352),
    .D(_0345_),
    .Q_N(_2248_),
    .Q(\audio_inst.i_over.counter[2] ));
 sg13g2_dfrbp_1 _5401_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net348),
    .D(_0346_),
    .Q_N(_2247_),
    .Q(\audio_inst.i_over.counter[3] ));
 sg13g2_dfrbp_1 _5402_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net344),
    .D(_0347_),
    .Q_N(_2246_),
    .Q(\audio_inst.i_over.counter[4] ));
 sg13g2_dfrbp_1 _5403_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net340),
    .D(_0348_),
    .Q_N(_2245_),
    .Q(\audio_inst.i_over.counter[5] ));
 sg13g2_dfrbp_1 _5404_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net314),
    .D(_0349_),
    .Q_N(_2244_),
    .Q(\audio_inst.i_over.counter[6] ));
 sg13g2_dfrbp_1 _5405_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net183),
    .D(_0350_),
    .Q_N(_2243_),
    .Q(\audio_inst.i_over.counter[7] ));
 sg13g2_dfrbp_1 _5406_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net179),
    .D(_0351_),
    .Q_N(_2242_),
    .Q(\audio_inst.i_over.counter[8] ));
 sg13g2_dfrbp_1 _5407_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net175),
    .D(_0352_),
    .Q_N(_2241_),
    .Q(\audio_inst.i_over.counter[9] ));
 sg13g2_dfrbp_1 _5408_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net171),
    .D(_0353_),
    .Q_N(_2240_),
    .Q(\audio_inst.i_over.counter[10] ));
 sg13g2_dfrbp_1 _5409_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net167),
    .D(_0354_),
    .Q_N(_2239_),
    .Q(\audio_inst.i_over.counter[11] ));
 sg13g2_dfrbp_1 _5410_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net123),
    .D(_0355_),
    .Q_N(_2238_),
    .Q(\audio_inst.i_over.counter[12] ));
 sg13g2_dfrbp_1 _5411_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net111),
    .D(_0356_),
    .Q_N(_2237_),
    .Q(\audio_inst.i_over.counter[13] ));
 sg13g2_dfrbp_1 _5412_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net103),
    .D(_0357_),
    .Q_N(_2236_),
    .Q(\audio_inst.i_over.counter[14] ));
 sg13g2_dfrbp_1 _5413_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net95),
    .D(_0358_),
    .Q_N(_2235_),
    .Q(\audio_inst.i_over.counter[15] ));
 sg13g2_dfrbp_1 _5414_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net87),
    .D(_0359_),
    .Q_N(_2234_),
    .Q(\audio_inst.i_over.counter[16] ));
 sg13g2_dfrbp_1 _5415_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net79),
    .D(_0360_),
    .Q_N(_2233_),
    .Q(\audio_inst.i_over.counter[17] ));
 sg13g2_dfrbp_1 _5416_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net71),
    .D(_0361_),
    .Q_N(_0007_),
    .Q(\audio_inst.i_over.counter[18] ));
 sg13g2_dfrbp_1 _5417_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net63),
    .D(_0362_),
    .Q_N(_2232_),
    .Q(\audio_inst.i_over.active ));
 sg13g2_dfrbp_1 _5418_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net55),
    .D(net778),
    .Q_N(_2231_),
    .Q(\audio_inst.i_jump.wave_out ));
 sg13g2_dfrbp_1 _5419_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net47),
    .D(net648),
    .Q_N(_0022_),
    .Q(\audio_inst.i_jump.stage_index[0] ));
 sg13g2_dfrbp_1 _5420_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net39),
    .D(_0365_),
    .Q_N(_0006_),
    .Q(\audio_inst.i_jump.stage_index[1] ));
 sg13g2_dfrbp_1 _5421_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net29),
    .D(_0366_),
    .Q_N(_0021_),
    .Q(\audio_inst.i_jump.stage_index[2] ));
 sg13g2_dfrbp_1 _5422_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net374),
    .D(_0367_),
    .Q_N(_0020_),
    .Q(\audio_inst.i_jump.stage_index[3] ));
 sg13g2_dfrbp_1 _5423_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net366),
    .D(_0368_),
    .Q_N(_0019_),
    .Q(\audio_inst.i_jump.stage_index[4] ));
 sg13g2_dfrbp_1 _5424_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net358),
    .D(net450),
    .Q_N(_2230_),
    .Q(\gamepad_pmod.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _5425_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net350),
    .D(net431),
    .Q_N(_2229_),
    .Q(\gamepad_pmod.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _5426_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net342),
    .D(net419),
    .Q_N(_2228_),
    .Q(\gamepad_pmod.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _5427_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net185),
    .D(net627),
    .Q_N(_2227_),
    .Q(\gamepad_pmod.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _5428_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net177),
    .D(net412),
    .Q_N(_2226_),
    .Q(\gamepad_pmod.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _5429_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net169),
    .D(net440),
    .Q_N(_2225_),
    .Q(\gamepad_pmod.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _5430_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net119),
    .D(_0375_),
    .Q_N(_2224_),
    .Q(\gamepad_pmod.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _5431_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net99),
    .D(_0376_),
    .Q_N(_2223_),
    .Q(\gamepad_pmod.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _5432_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net83),
    .D(net656),
    .Q_N(_2222_),
    .Q(\gamepad_pmod.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _5433_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net67),
    .D(net429),
    .Q_N(_2221_),
    .Q(\gamepad_pmod.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _5434_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net51),
    .D(net437),
    .Q_N(_2220_),
    .Q(\gamepad_pmod.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _5435_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net33),
    .D(net643),
    .Q_N(_2219_),
    .Q(\gamepad_pmod.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _5436_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net370),
    .D(net631),
    .Q_N(_2218_),
    .Q(\audio_inst.i_jump.active ));
 sg13g2_dfrbp_1 _5437_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net354),
    .D(_0382_),
    .Q_N(_2217_),
    .Q(\audio_inst.sound ));
 sg13g2_dfrbp_1 _5438_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net346),
    .D(_0383_),
    .Q_N(_2216_),
    .Q(\ai_controller_inst.restart_counter[0] ));
 sg13g2_dfrbp_1 _5439_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net181),
    .D(_0384_),
    .Q_N(_2215_),
    .Q(\ai_controller_inst.restart_counter[1] ));
 sg13g2_dfrbp_1 _5440_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net131),
    .D(_0385_),
    .Q_N(_2214_),
    .Q(\ai_controller_inst.restart_counter[2] ));
 sg13g2_dfrbp_1 _5441_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net91),
    .D(_0386_),
    .Q_N(_2213_),
    .Q(\ai_controller_inst.restart_counter[3] ));
 sg13g2_dfrbp_1 _5442_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net59),
    .D(_0387_),
    .Q_N(_2212_),
    .Q(\ai_controller_inst.restart_counter[4] ));
 sg13g2_dfrbp_1 _5443_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net20),
    .D(net660),
    .Q_N(_2211_),
    .Q(\ai_controller_inst.restart_counter[5] ));
 sg13g2_dfrbp_1 _5444_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net316),
    .D(net443),
    .Q_N(_2210_),
    .Q(\ai_controller_inst.restart_counter[6] ));
 sg13g2_dfrbp_1 _5445_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net107),
    .D(net448),
    .Q_N(_2209_),
    .Q(\ai_controller_inst.restart_counter[7] ));
 sg13g2_dfrbp_1 _5446_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net43),
    .D(_0391_),
    .Q_N(_2208_),
    .Q(\ai_controller_inst.button_down ));
 sg13g2_dfrbp_1 _5447_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net173),
    .D(_0392_),
    .Q_N(_2207_),
    .Q(\ai_controller_inst.button_up ));
 sg13g2_dfrbp_1 _5448_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net362),
    .D(net801),
    .Q_N(_2206_),
    .Q(\ai_controller_inst.button_start ));
 sg13g2_tiehi _5167__19 (.L_HI(net19));
 sg13g2_tiehi _5443__20 (.L_HI(net20));
 sg13g2_tiehi _5166__21 (.L_HI(net21));
 sg13g2_tiehi _5165__22 (.L_HI(net22));
 sg13g2_tiehi _5164__23 (.L_HI(net23));
 sg13g2_tiehi _5163__24 (.L_HI(net24));
 sg13g2_tiehi _5162__25 (.L_HI(net25));
 sg13g2_tiehi _5161__26 (.L_HI(net26));
 sg13g2_tiehi _5393__27 (.L_HI(net27));
 sg13g2_tiehi _5160__28 (.L_HI(net28));
 sg13g2_tiehi _5421__29 (.L_HI(net29));
 sg13g2_tiehi _5159__30 (.L_HI(net30));
 sg13g2_tiehi _5392__31 (.L_HI(net31));
 sg13g2_tiehi _5158__32 (.L_HI(net32));
 sg13g2_tiehi _5435__33 (.L_HI(net33));
 sg13g2_tiehi _5157__34 (.L_HI(net34));
 sg13g2_tiehi _5391__35 (.L_HI(net35));
 sg13g2_tiehi _5083__36 (.L_HI(net36));
 sg13g2_tiehi _5100__37 (.L_HI(net37));
 sg13g2_tiehi _5156__38 (.L_HI(net38));
 sg13g2_tiehi _5420__39 (.L_HI(net39));
 sg13g2_tiehi _5155__40 (.L_HI(net40));
 sg13g2_tiehi _5384__41 (.L_HI(net41));
 sg13g2_tiehi _5154__42 (.L_HI(net42));
 sg13g2_tiehi _5446__43 (.L_HI(net43));
 sg13g2_tiehi _5153__44 (.L_HI(net44));
 sg13g2_tiehi _5383__45 (.L_HI(net45));
 sg13g2_tiehi _5152__46 (.L_HI(net46));
 sg13g2_tiehi _5419__47 (.L_HI(net47));
 sg13g2_tiehi _5151__48 (.L_HI(net48));
 sg13g2_tiehi _5382__49 (.L_HI(net49));
 sg13g2_tiehi _5150__50 (.L_HI(net50));
 sg13g2_tiehi _5434__51 (.L_HI(net51));
 sg13g2_tiehi _5149__52 (.L_HI(net52));
 sg13g2_tiehi _5381__53 (.L_HI(net53));
 sg13g2_tiehi _5148__54 (.L_HI(net54));
 sg13g2_tiehi _5418__55 (.L_HI(net55));
 sg13g2_tiehi _5147__56 (.L_HI(net56));
 sg13g2_tiehi _5380__57 (.L_HI(net57));
 sg13g2_tiehi _5146__58 (.L_HI(net58));
 sg13g2_tiehi _5442__59 (.L_HI(net59));
 sg13g2_tiehi _5145__60 (.L_HI(net60));
 sg13g2_tiehi _5379__61 (.L_HI(net61));
 sg13g2_tiehi _5144__62 (.L_HI(net62));
 sg13g2_tiehi _5417__63 (.L_HI(net63));
 sg13g2_tiehi _5143__64 (.L_HI(net64));
 sg13g2_tiehi _5378__65 (.L_HI(net65));
 sg13g2_tiehi _5142__66 (.L_HI(net66));
 sg13g2_tiehi _5433__67 (.L_HI(net67));
 sg13g2_tiehi _5141__68 (.L_HI(net68));
 sg13g2_tiehi _5377__69 (.L_HI(net69));
 sg13g2_tiehi _5140__70 (.L_HI(net70));
 sg13g2_tiehi _5416__71 (.L_HI(net71));
 sg13g2_tiehi _5139__72 (.L_HI(net72));
 sg13g2_tiehi _5376__73 (.L_HI(net73));
 sg13g2_tiehi _5138__74 (.L_HI(net74));
 sg13g2_tiehi _5390__75 (.L_HI(net75));
 sg13g2_tiehi _5137__76 (.L_HI(net76));
 sg13g2_tiehi _5375__77 (.L_HI(net77));
 sg13g2_tiehi _5136__78 (.L_HI(net78));
 sg13g2_tiehi _5415__79 (.L_HI(net79));
 sg13g2_tiehi _5135__80 (.L_HI(net80));
 sg13g2_tiehi _5374__81 (.L_HI(net81));
 sg13g2_tiehi _5134__82 (.L_HI(net82));
 sg13g2_tiehi _5432__83 (.L_HI(net83));
 sg13g2_tiehi _5133__84 (.L_HI(net84));
 sg13g2_tiehi _5373__85 (.L_HI(net85));
 sg13g2_tiehi _5132__86 (.L_HI(net86));
 sg13g2_tiehi _5414__87 (.L_HI(net87));
 sg13g2_tiehi _5131__88 (.L_HI(net88));
 sg13g2_tiehi _5372__89 (.L_HI(net89));
 sg13g2_tiehi _5130__90 (.L_HI(net90));
 sg13g2_tiehi _5441__91 (.L_HI(net91));
 sg13g2_tiehi _5129__92 (.L_HI(net92));
 sg13g2_tiehi _5371__93 (.L_HI(net93));
 sg13g2_tiehi _5128__94 (.L_HI(net94));
 sg13g2_tiehi _5413__95 (.L_HI(net95));
 sg13g2_tiehi _5127__96 (.L_HI(net96));
 sg13g2_tiehi _5370__97 (.L_HI(net97));
 sg13g2_tiehi _5126__98 (.L_HI(net98));
 sg13g2_tiehi _5431__99 (.L_HI(net99));
 sg13g2_tiehi _5125__100 (.L_HI(net100));
 sg13g2_tiehi _5369__101 (.L_HI(net101));
 sg13g2_tiehi _5124__102 (.L_HI(net102));
 sg13g2_tiehi _5412__103 (.L_HI(net103));
 sg13g2_tiehi _5123__104 (.L_HI(net104));
 sg13g2_tiehi _5368__105 (.L_HI(net105));
 sg13g2_tiehi _5122__106 (.L_HI(net106));
 sg13g2_tiehi _5445__107 (.L_HI(net107));
 sg13g2_tiehi _5121__108 (.L_HI(net108));
 sg13g2_tiehi _5367__109 (.L_HI(net109));
 sg13g2_tiehi _5120__110 (.L_HI(net110));
 sg13g2_tiehi _5411__111 (.L_HI(net111));
 sg13g2_tiehi _5119__112 (.L_HI(net112));
 sg13g2_tiehi _5118__113 (.L_HI(net113));
 sg13g2_tiehi _5117__114 (.L_HI(net114));
 sg13g2_tiehi _5116__115 (.L_HI(net115));
 sg13g2_tiehi _5115__116 (.L_HI(net116));
 sg13g2_tiehi _5366__117 (.L_HI(net117));
 sg13g2_tiehi _5114__118 (.L_HI(net118));
 sg13g2_tiehi _5430__119 (.L_HI(net119));
 sg13g2_tiehi _5113__120 (.L_HI(net120));
 sg13g2_tiehi _5365__121 (.L_HI(net121));
 sg13g2_tiehi _5112__122 (.L_HI(net122));
 sg13g2_tiehi _5410__123 (.L_HI(net123));
 sg13g2_tiehi _5111__124 (.L_HI(net124));
 sg13g2_tiehi _5364__125 (.L_HI(net125));
 sg13g2_tiehi _5110__126 (.L_HI(net126));
 sg13g2_tiehi _5363__127 (.L_HI(net127));
 sg13g2_tiehi _5109__128 (.L_HI(net128));
 sg13g2_tiehi _5362__129 (.L_HI(net129));
 sg13g2_tiehi _5108__130 (.L_HI(net130));
 sg13g2_tiehi _5440__131 (.L_HI(net131));
 sg13g2_tiehi _5107__132 (.L_HI(net132));
 sg13g2_tiehi _5361__133 (.L_HI(net133));
 sg13g2_tiehi _5106__134 (.L_HI(net134));
 sg13g2_tiehi _5360__135 (.L_HI(net135));
 sg13g2_tiehi _5105__136 (.L_HI(net136));
 sg13g2_tiehi _5359__137 (.L_HI(net137));
 sg13g2_tiehi _5104__138 (.L_HI(net138));
 sg13g2_tiehi _5358__139 (.L_HI(net139));
 sg13g2_tiehi _5103__140 (.L_HI(net140));
 sg13g2_tiehi _5357__141 (.L_HI(net141));
 sg13g2_tiehi _5102__142 (.L_HI(net142));
 sg13g2_tiehi _5099__143 (.L_HI(net143));
 sg13g2_tiehi _5098__144 (.L_HI(net144));
 sg13g2_tiehi _5097__145 (.L_HI(net145));
 sg13g2_tiehi _5096__146 (.L_HI(net146));
 sg13g2_tiehi _5095__147 (.L_HI(net147));
 sg13g2_tiehi _5094__148 (.L_HI(net148));
 sg13g2_tiehi _5093__149 (.L_HI(net149));
 sg13g2_tiehi _5092__150 (.L_HI(net150));
 sg13g2_tiehi _5091__151 (.L_HI(net151));
 sg13g2_tiehi _5090__152 (.L_HI(net152));
 sg13g2_tiehi _5089__153 (.L_HI(net153));
 sg13g2_tiehi _5088__154 (.L_HI(net154));
 sg13g2_tiehi _5087__155 (.L_HI(net155));
 sg13g2_tiehi _5086__156 (.L_HI(net156));
 sg13g2_tiehi _5085__157 (.L_HI(net157));
 sg13g2_tiehi _5084__158 (.L_HI(net158));
 sg13g2_tiehi _5356__159 (.L_HI(net159));
 sg13g2_tiehi _5355__160 (.L_HI(net160));
 sg13g2_tiehi _5354__161 (.L_HI(net161));
 sg13g2_tiehi _5353__162 (.L_HI(net162));
 sg13g2_tiehi _5352__163 (.L_HI(net163));
 sg13g2_tiehi _5351__164 (.L_HI(net164));
 sg13g2_tiehi _5350__165 (.L_HI(net165));
 sg13g2_tiehi _5349__166 (.L_HI(net166));
 sg13g2_tiehi _5409__167 (.L_HI(net167));
 sg13g2_tiehi _5348__168 (.L_HI(net168));
 sg13g2_tiehi _5429__169 (.L_HI(net169));
 sg13g2_tiehi _5347__170 (.L_HI(net170));
 sg13g2_tiehi _5408__171 (.L_HI(net171));
 sg13g2_tiehi _5346__172 (.L_HI(net172));
 sg13g2_tiehi _5447__173 (.L_HI(net173));
 sg13g2_tiehi _5345__174 (.L_HI(net174));
 sg13g2_tiehi _5407__175 (.L_HI(net175));
 sg13g2_tiehi _5344__176 (.L_HI(net176));
 sg13g2_tiehi _5428__177 (.L_HI(net177));
 sg13g2_tiehi _5343__178 (.L_HI(net178));
 sg13g2_tiehi _5406__179 (.L_HI(net179));
 sg13g2_tiehi _5342__180 (.L_HI(net180));
 sg13g2_tiehi _5439__181 (.L_HI(net181));
 sg13g2_tiehi _5341__182 (.L_HI(net182));
 sg13g2_tiehi _5405__183 (.L_HI(net183));
 sg13g2_tiehi _5340__184 (.L_HI(net184));
 sg13g2_tiehi _5427__185 (.L_HI(net185));
 sg13g2_tiehi _5339__186 (.L_HI(net186));
 sg13g2_tiehi _5338__187 (.L_HI(net187));
 sg13g2_tiehi _5337__188 (.L_HI(net188));
 sg13g2_tiehi _5336__189 (.L_HI(net189));
 sg13g2_tiehi _5335__190 (.L_HI(net190));
 sg13g2_tiehi _5334__191 (.L_HI(net191));
 sg13g2_tiehi _5333__192 (.L_HI(net192));
 sg13g2_tiehi _5332__193 (.L_HI(net193));
 sg13g2_tiehi _5331__194 (.L_HI(net194));
 sg13g2_tiehi _5330__195 (.L_HI(net195));
 sg13g2_tiehi _5329__196 (.L_HI(net196));
 sg13g2_tiehi _5328__197 (.L_HI(net197));
 sg13g2_tiehi _5327__198 (.L_HI(net198));
 sg13g2_tiehi _5326__199 (.L_HI(net199));
 sg13g2_tiehi _5325__200 (.L_HI(net200));
 sg13g2_tiehi _5324__201 (.L_HI(net201));
 sg13g2_tiehi _5323__202 (.L_HI(net202));
 sg13g2_tiehi _5322__203 (.L_HI(net203));
 sg13g2_tiehi _5321__204 (.L_HI(net204));
 sg13g2_tiehi _5320__205 (.L_HI(net205));
 sg13g2_tiehi _5319__206 (.L_HI(net206));
 sg13g2_tiehi _5318__207 (.L_HI(net207));
 sg13g2_tiehi _5317__208 (.L_HI(net208));
 sg13g2_tiehi _5316__209 (.L_HI(net209));
 sg13g2_tiehi _5315__210 (.L_HI(net210));
 sg13g2_tiehi _5314__211 (.L_HI(net211));
 sg13g2_tiehi _5313__212 (.L_HI(net212));
 sg13g2_tiehi _5312__213 (.L_HI(net213));
 sg13g2_tiehi _5311__214 (.L_HI(net214));
 sg13g2_tiehi _5310__215 (.L_HI(net215));
 sg13g2_tiehi _5309__216 (.L_HI(net216));
 sg13g2_tiehi _5308__217 (.L_HI(net217));
 sg13g2_tiehi _5307__218 (.L_HI(net218));
 sg13g2_tiehi _5306__219 (.L_HI(net219));
 sg13g2_tiehi _5305__220 (.L_HI(net220));
 sg13g2_tiehi _5304__221 (.L_HI(net221));
 sg13g2_tiehi _5303__222 (.L_HI(net222));
 sg13g2_tiehi _5302__223 (.L_HI(net223));
 sg13g2_tiehi _5301__224 (.L_HI(net224));
 sg13g2_tiehi _5300__225 (.L_HI(net225));
 sg13g2_tiehi _5299__226 (.L_HI(net226));
 sg13g2_tiehi _5298__227 (.L_HI(net227));
 sg13g2_tiehi _5297__228 (.L_HI(net228));
 sg13g2_tiehi _5296__229 (.L_HI(net229));
 sg13g2_tiehi _5295__230 (.L_HI(net230));
 sg13g2_tiehi _5294__231 (.L_HI(net231));
 sg13g2_tiehi _5293__232 (.L_HI(net232));
 sg13g2_tiehi _5292__233 (.L_HI(net233));
 sg13g2_tiehi _5291__234 (.L_HI(net234));
 sg13g2_tiehi _5290__235 (.L_HI(net235));
 sg13g2_tiehi _5289__236 (.L_HI(net236));
 sg13g2_tiehi _5288__237 (.L_HI(net237));
 sg13g2_tiehi _5287__238 (.L_HI(net238));
 sg13g2_tiehi _5286__239 (.L_HI(net239));
 sg13g2_tiehi _5285__240 (.L_HI(net240));
 sg13g2_tiehi _5284__241 (.L_HI(net241));
 sg13g2_tiehi _5283__242 (.L_HI(net242));
 sg13g2_tiehi _5282__243 (.L_HI(net243));
 sg13g2_tiehi _5281__244 (.L_HI(net244));
 sg13g2_tiehi _5280__245 (.L_HI(net245));
 sg13g2_tiehi _5279__246 (.L_HI(net246));
 sg13g2_tiehi _5278__247 (.L_HI(net247));
 sg13g2_tiehi _5277__248 (.L_HI(net248));
 sg13g2_tiehi _5276__249 (.L_HI(net249));
 sg13g2_tiehi _5275__250 (.L_HI(net250));
 sg13g2_tiehi _5274__251 (.L_HI(net251));
 sg13g2_tiehi _5273__252 (.L_HI(net252));
 sg13g2_tiehi _5272__253 (.L_HI(net253));
 sg13g2_tiehi _5271__254 (.L_HI(net254));
 sg13g2_tiehi _5270__255 (.L_HI(net255));
 sg13g2_tiehi _5269__256 (.L_HI(net256));
 sg13g2_tiehi _5268__257 (.L_HI(net257));
 sg13g2_tiehi _5267__258 (.L_HI(net258));
 sg13g2_tiehi _5266__259 (.L_HI(net259));
 sg13g2_tiehi _5265__260 (.L_HI(net260));
 sg13g2_tiehi _5264__261 (.L_HI(net261));
 sg13g2_tiehi _5263__262 (.L_HI(net262));
 sg13g2_tiehi _5262__263 (.L_HI(net263));
 sg13g2_tiehi _5261__264 (.L_HI(net264));
 sg13g2_tiehi _5260__265 (.L_HI(net265));
 sg13g2_tiehi _5259__266 (.L_HI(net266));
 sg13g2_tiehi _5258__267 (.L_HI(net267));
 sg13g2_tiehi _5257__268 (.L_HI(net268));
 sg13g2_tiehi _5256__269 (.L_HI(net269));
 sg13g2_tiehi _5255__270 (.L_HI(net270));
 sg13g2_tiehi _5254__271 (.L_HI(net271));
 sg13g2_tiehi _5253__272 (.L_HI(net272));
 sg13g2_tiehi _5252__273 (.L_HI(net273));
 sg13g2_tiehi _5251__274 (.L_HI(net274));
 sg13g2_tiehi _5250__275 (.L_HI(net275));
 sg13g2_tiehi _5249__276 (.L_HI(net276));
 sg13g2_tiehi _5248__277 (.L_HI(net277));
 sg13g2_tiehi _5247__278 (.L_HI(net278));
 sg13g2_tiehi _5246__279 (.L_HI(net279));
 sg13g2_tiehi _5245__280 (.L_HI(net280));
 sg13g2_tiehi _5244__281 (.L_HI(net281));
 sg13g2_tiehi _5243__282 (.L_HI(net282));
 sg13g2_tiehi _5242__283 (.L_HI(net283));
 sg13g2_tiehi _5241__284 (.L_HI(net284));
 sg13g2_tiehi _5240__285 (.L_HI(net285));
 sg13g2_tiehi _5239__286 (.L_HI(net286));
 sg13g2_tiehi _5238__287 (.L_HI(net287));
 sg13g2_tiehi _5237__288 (.L_HI(net288));
 sg13g2_tiehi _5236__289 (.L_HI(net289));
 sg13g2_tiehi _5235__290 (.L_HI(net290));
 sg13g2_tiehi _5234__291 (.L_HI(net291));
 sg13g2_tiehi _5233__292 (.L_HI(net292));
 sg13g2_tiehi _5232__293 (.L_HI(net293));
 sg13g2_tiehi _5231__294 (.L_HI(net294));
 sg13g2_tiehi _5230__295 (.L_HI(net295));
 sg13g2_tiehi _5229__296 (.L_HI(net296));
 sg13g2_tiehi _5228__297 (.L_HI(net297));
 sg13g2_tiehi _5227__298 (.L_HI(net298));
 sg13g2_tiehi _5226__299 (.L_HI(net299));
 sg13g2_tiehi _5225__300 (.L_HI(net300));
 sg13g2_tiehi _5224__301 (.L_HI(net301));
 sg13g2_tiehi _5223__302 (.L_HI(net302));
 sg13g2_tiehi _5222__303 (.L_HI(net303));
 sg13g2_tiehi _5221__304 (.L_HI(net304));
 sg13g2_tiehi _5220__305 (.L_HI(net305));
 sg13g2_tiehi _5219__306 (.L_HI(net306));
 sg13g2_tiehi _5218__307 (.L_HI(net307));
 sg13g2_tiehi _5217__308 (.L_HI(net308));
 sg13g2_tiehi _5216__309 (.L_HI(net309));
 sg13g2_tiehi _5215__310 (.L_HI(net310));
 sg13g2_tiehi _5214__311 (.L_HI(net311));
 sg13g2_tiehi _5213__312 (.L_HI(net312));
 sg13g2_tiehi _5212__313 (.L_HI(net313));
 sg13g2_tiehi _5404__314 (.L_HI(net314));
 sg13g2_tiehi _5211__315 (.L_HI(net315));
 sg13g2_tiehi _5444__316 (.L_HI(net316));
 sg13g2_tiehi _5210__317 (.L_HI(net317));
 sg13g2_tiehi _5209__318 (.L_HI(net318));
 sg13g2_tiehi _5208__319 (.L_HI(net319));
 sg13g2_tiehi _5207__320 (.L_HI(net320));
 sg13g2_tiehi _5101__321 (.L_HI(net321));
 sg13g2_tiehi _5385__322 (.L_HI(net322));
 sg13g2_tiehi _5386__323 (.L_HI(net323));
 sg13g2_tiehi _5387__324 (.L_HI(net324));
 sg13g2_tiehi _5388__325 (.L_HI(net325));
 sg13g2_tiehi _5389__326 (.L_HI(net326));
 sg13g2_tiehi _5206__327 (.L_HI(net327));
 sg13g2_tiehi _5205__328 (.L_HI(net328));
 sg13g2_tiehi _5204__329 (.L_HI(net329));
 sg13g2_tiehi _5203__330 (.L_HI(net330));
 sg13g2_tiehi _5202__331 (.L_HI(net331));
 sg13g2_tiehi _5201__332 (.L_HI(net332));
 sg13g2_tiehi _5200__333 (.L_HI(net333));
 sg13g2_tiehi _5199__334 (.L_HI(net334));
 sg13g2_tiehi _5198__335 (.L_HI(net335));
 sg13g2_tiehi _5197__336 (.L_HI(net336));
 sg13g2_tiehi _5196__337 (.L_HI(net337));
 sg13g2_tiehi _5195__338 (.L_HI(net338));
 sg13g2_tiehi _5194__339 (.L_HI(net339));
 sg13g2_tiehi _5403__340 (.L_HI(net340));
 sg13g2_tiehi _5193__341 (.L_HI(net341));
 sg13g2_tiehi _5426__342 (.L_HI(net342));
 sg13g2_tiehi _5192__343 (.L_HI(net343));
 sg13g2_tiehi _5402__344 (.L_HI(net344));
 sg13g2_tiehi _5191__345 (.L_HI(net345));
 sg13g2_tiehi _5438__346 (.L_HI(net346));
 sg13g2_tiehi _5190__347 (.L_HI(net347));
 sg13g2_tiehi _5401__348 (.L_HI(net348));
 sg13g2_tiehi _5189__349 (.L_HI(net349));
 sg13g2_tiehi _5425__350 (.L_HI(net350));
 sg13g2_tiehi _5188__351 (.L_HI(net351));
 sg13g2_tiehi _5400__352 (.L_HI(net352));
 sg13g2_tiehi _5187__353 (.L_HI(net353));
 sg13g2_tiehi _5437__354 (.L_HI(net354));
 sg13g2_tiehi _5186__355 (.L_HI(net355));
 sg13g2_tiehi _5399__356 (.L_HI(net356));
 sg13g2_tiehi _5185__357 (.L_HI(net357));
 sg13g2_tiehi _5424__358 (.L_HI(net358));
 sg13g2_tiehi _5184__359 (.L_HI(net359));
 sg13g2_tiehi _5398__360 (.L_HI(net360));
 sg13g2_tiehi _5183__361 (.L_HI(net361));
 sg13g2_tiehi _5448__362 (.L_HI(net362));
 sg13g2_tiehi _5182__363 (.L_HI(net363));
 sg13g2_tiehi _5397__364 (.L_HI(net364));
 sg13g2_tiehi _5181__365 (.L_HI(net365));
 sg13g2_tiehi _5423__366 (.L_HI(net366));
 sg13g2_tiehi _5180__367 (.L_HI(net367));
 sg13g2_tiehi _5396__368 (.L_HI(net368));
 sg13g2_tiehi _5179__369 (.L_HI(net369));
 sg13g2_tiehi _5436__370 (.L_HI(net370));
 sg13g2_tiehi _5178__371 (.L_HI(net371));
 sg13g2_tiehi _5395__372 (.L_HI(net372));
 sg13g2_tiehi _5177__373 (.L_HI(net373));
 sg13g2_tiehi _5422__374 (.L_HI(net374));
 sg13g2_tiehi _5176__375 (.L_HI(net375));
 sg13g2_tiehi _5394__376 (.L_HI(net376));
 sg13g2_tiehi _5175__377 (.L_HI(net377));
 sg13g2_tiehi _5174__378 (.L_HI(net378));
 sg13g2_tiehi _5173__379 (.L_HI(net379));
 sg13g2_tiehi _5172__380 (.L_HI(net380));
 sg13g2_tiehi _5171__381 (.L_HI(net381));
 sg13g2_tiehi _5170__382 (.L_HI(net382));
 sg13g2_tiehi _5169__383 (.L_HI(net383));
 sg13g2_tiehi tt_um_uwasic_dinogame_384 (.L_HI(net384));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_uwasic_dinogame_5 (.L_LO(net5));
 sg13g2_tielo tt_um_uwasic_dinogame_6 (.L_LO(net6));
 sg13g2_tielo tt_um_uwasic_dinogame_7 (.L_LO(net7));
 sg13g2_tielo tt_um_uwasic_dinogame_8 (.L_LO(net8));
 sg13g2_tielo tt_um_uwasic_dinogame_9 (.L_LO(net9));
 sg13g2_tielo tt_um_uwasic_dinogame_10 (.L_LO(net10));
 sg13g2_tielo tt_um_uwasic_dinogame_11 (.L_LO(net11));
 sg13g2_tielo tt_um_uwasic_dinogame_12 (.L_LO(net12));
 sg13g2_tielo tt_um_uwasic_dinogame_13 (.L_LO(net13));
 sg13g2_tielo tt_um_uwasic_dinogame_14 (.L_LO(net14));
 sg13g2_tielo tt_um_uwasic_dinogame_15 (.L_LO(net15));
 sg13g2_tielo tt_um_uwasic_dinogame_16 (.L_LO(net16));
 sg13g2_tielo tt_um_uwasic_dinogame_17 (.L_LO(net17));
 sg13g2_tiehi _5168__18 (.L_HI(net18));
 sg13g2_buf_1 _5830_ (.A(\audio_inst.sound ),
    .X(uio_out[7]));
 sg13g2_buf_1 _5831_ (.A(uo_out[4]),
    .X(uo_out[2]));
 sg13g2_buf_1 _5832_ (.A(\graphics_inst.o_vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _5833_ (.A(\graphics_inst.hsync_r_r ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_0656_),
    .X(net470));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(_1836_));
 sg13g2_buf_2 fanout472 (.A(_1836_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_0728_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_0642_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(net481),
    .X(net478));
 sg13g2_buf_1 fanout479 (.A(net481),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(net481),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_0430_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net485),
    .X(net482));
 sg13g2_buf_1 fanout483 (.A(net485),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_1 fanout485 (.A(_0727_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net487),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_0467_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(net491),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(_0467_));
 sg13g2_buf_2 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_1 fanout493 (.A(_0437_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_0492_),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(_0474_));
 sg13g2_buf_1 fanout496 (.A(_0474_),
    .X(net496));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(_2137_));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(_0473_));
 sg13g2_buf_2 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_2136_),
    .X(net500));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(_2135_));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(_1947_));
 sg13g2_buf_2 fanout503 (.A(_1947_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_1411_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_1404_),
    .X(net505));
 sg13g2_buf_1 fanout506 (.A(_1404_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_1213_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_1213_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_1212_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_1212_),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_0436_));
 sg13g2_buf_2 fanout512 (.A(_0436_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_2186_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_1946_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_1946_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_1518_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_0435_),
    .X(net517));
 sg13g2_buf_1 fanout518 (.A(_0435_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_2099_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_2007_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net883),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net525),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(net525),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(\audio_inst.i_jump.stage_index[4] ),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(\audio_inst.i_jump.stage_index[3] ),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net531),
    .X(net529));
 sg13g2_buf_1 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(net877),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(\audio_inst.i_jump.stage_index[1] ));
 sg13g2_buf_2 fanout533 (.A(net890),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(\audio_inst.i_jump.stage_index[0] ),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(net538),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(net852),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net540),
    .X(net539));
 sg13g2_buf_1 fanout540 (.A(_0008_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net856),
    .X(net543));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(net874));
 sg13g2_buf_1 fanout545 (.A(\audio_inst.i_over.stage_index[1] ),
    .X(net545));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(\audio_inst.i_over.stage_index[0] ));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net843),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(\bg_line_inst.i_vpos[7] ),
    .X(net550));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(\bg_line_inst.i_vpos[6] ));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(\bg_line_inst.i_vpos[5] ),
    .X(net553));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(net816));
 sg13g2_buf_2 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(\bg_line_inst.i_vpos[3] ),
    .X(net556));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(net432));
 sg13g2_buf_2 fanout558 (.A(\bg_object_rom_inst.i_rom_counter[5] ),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(\obs_inst_1.o_rom_counter[0] ),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(\obs_inst_1.o_rom_counter[7] ),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(\obs_inst_1.o_rom_counter[6] ),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(\obs_inst_1.o_rom_counter[5] ),
    .X(net564));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(net566));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(\obs_inst_1.o_rom_counter[4] ));
 sg13g2_buf_2 fanout567 (.A(\dino_inst.o_rom_counter[4] ),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(\dino_inst.o_rom_counter[3] ),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(\dino_inst.o_rom_counter[0] ),
    .X(net569));
 sg13g2_buf_1 fanout570 (.A(\dino_inst.o_rom_counter[0] ),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(\obs_inst_2.o_rom_counter[0] ),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net797),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_1 fanout574 (.A(\obs_rom_inst_2.i_obs_type[0] ),
    .X(net574));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net898));
 sg13g2_buf_2 fanout576 (.A(net892),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(\bg_render_inst.i_hpos[9] ),
    .X(net577));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(net579));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(\bg_render_inst.i_hpos[8] ));
 sg13g2_buf_2 fanout581 (.A(net583),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(\bg_render_inst.i_hpos[7] ));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(\bg_render_inst.i_hpos[6] ));
 sg13g2_buf_2 fanout587 (.A(net811),
    .X(net587));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(net589));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(\bg_render_inst.i_hpos[5] ));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(net886));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(net886));
 sg13g2_buf_2 fanout592 (.A(net594),
    .X(net592));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(net594));
 sg13g2_buf_2 fanout594 (.A(\bg_render_inst.i_hpos[3] ),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(\bg_render_inst.i_hpos[2] ));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(net606));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(net599));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(net599));
 sg13g2_buf_2 fanout599 (.A(net606),
    .X(net599));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(net602));
 sg13g2_buf_1 fanout601 (.A(net602),
    .X(net601));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(net606));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(_2051_));
 sg13g2_buf_4 fanout607 (.X(net607),
    .A(net608));
 sg13g2_buf_2 fanout608 (.A(net616),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(net616),
    .X(net609));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(net615));
 sg13g2_buf_1 fanout611 (.A(net615),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net614),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net616),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(rst_n),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net624),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(net624),
    .X(net620));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(net623));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(net623));
 sg13g2_buf_2 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(rst_n),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(ena),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(ena),
    .X(net626));
 sg13g2_buf_2 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[5]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_tielo tt_um_uwasic_dinogame_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_45_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_50_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_1_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_3_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_43_clk));
 sg13g2_inv_8 clkload9 (.A(clknet_leaf_51_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_38_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_40_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_18_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_23_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_25_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gamepad_pmod.driver.pmod_clk_sync[1] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gamepad_pmod.driver.pmod_latch_sync[1] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0035_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold4 (.A(\dino_inst.x_offset[3] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0034_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0657_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold7 (.A(\lfsr_inst.r_lfsr[11] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0033_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0290_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold10 (.A(\gamepad_pmod.driver.pmod_data_sync[0] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold11 (.A(\graphics_inst.vsync_r ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold12 (.A(\bg_render_inst.y_offset[2] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold13 (.A(\obs_inst_1.y_offset[3] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold14 (.A(\graphics_inst.hsync_r ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold15 (.A(\gamepad_pmod.driver.pmod_latch_sync[0] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold16 (.A(\lfsr_inst.r_lfsr[13] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold17 (.A(\lfsr_inst.r_lfsr[9] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold18 (.A(\gamepad_pmod.driver.pmod_clk_sync[0] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold19 (.A(\score[2] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold20 (.A(\lfsr_inst.r_lfsr[14] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold21 (.A(\score[3] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold22 (.A(\score[0] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0007_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold24 (.A(_1881_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold25 (.A(\graphics_inst.display_on_r ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold26 (.A(\score[12] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold27 (.A(\gamepad_pmod.decoder.data_reg[4] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0373_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold29 (.A(\score[13] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold30 (.A(\lfsr_inst.r_lfsr[10] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0028_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold32 (.A(_1838_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold33 (.A(\lfsr_inst.r_lfsr[12] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold34 (.A(\gamepad_pmod.decoder.data_reg[2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0371_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold36 (.A(\gamepad_pmod.driver.pmod_data_sync[1] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0054_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold38 (.A(\score[16] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold39 (.A(\lfsr_inst.r_lfsr[1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold40 (.A(\audio_inst.i_jump.decay_value[2] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold41 (.A(\audio_inst.i_jump.decay_value[1] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold42 (.A(\score[1] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold43 (.A(\graphics_inst.color_decoder_inst.invert ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold44 (.A(\gamepad_pmod.decoder.data_reg[9] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0378_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold46 (.A(\gamepad_pmod.decoder.data_reg[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0370_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold48 (.A(\bg_line_inst.i_vpos[2] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold49 (.A(\audio_inst.i_over.active ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0177_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold51 (.A(\score[15] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold52 (.A(\gamepad_pmod.decoder.data_reg[10] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0379_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold54 (.A(\audio_inst.i_jump.decay_value[16] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold55 (.A(\gamepad_pmod.decoder.data_reg[5] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0374_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ai_controller_inst.restart_counter[6] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1975_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0389_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold60 (.A(\audio_inst.i_jump.decay_value[15] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0162_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold62 (.A(\audio_inst.i_over.decay_value[7] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold63 (.A(\ai_controller_inst.restart_counter[7] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0390_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold65 (.A(\gamepad_pmod.decoder.data_reg[0] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0369_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold67 (.A(\audio_inst.i_jump.decay_value[7] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold68 (.A(\score[6] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold69 (.A(\obs_rom_inst_2.i_obs_type[0] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0082_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold71 (.A(\audio_inst.i_over.decay_value[1] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0146_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold73 (.A(\graphics_inst.frame_counter[1] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold74 (.A(\audio_inst.i_jump.decay_value[5] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold75 (.A(\audio_inst.i_over.decay_value[0] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0145_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold77 (.A(\score[19] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ai_controller_inst.crash ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold79 (.A(\score[4] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold80 (.A(\audio_inst.i_jump.decay_value[12] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold81 (.A(\audio_inst.i_jump.counter[3] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold82 (.A(\audio_inst.game_over_sound ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0337_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold84 (.A(\gamepad_pmod.decoder.data_reg[3] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0372_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold86 (.A(\score[9] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold87 (.A(\audio_inst.i_jump.active ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold88 (.A(_2198_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0381_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold90 (.A(\gamepad_pmod.driver.shift_reg[11] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0065_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold92 (.A(\audio_inst.i_jump.counter[7] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0133_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold94 (.A(\player_constroller_inst.game_state[0] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold95 (.A(\gamepad_pmod.driver.shift_reg[1] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0055_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold97 (.A(\audio_inst.i_jump.counter[14] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold98 (.A(\gamepad_pmod.driver.shift_reg[9] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0063_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold100 (.A(\gamepad_pmod.decoder.data_reg[11] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0380_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold102 (.A(\gamepad_pmod.driver.shift_reg[6] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0060_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold104 (.A(\audio_inst.i_jump.stage_index[0] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold105 (.A(_1937_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0364_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold107 (.A(\score[7] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold108 (.A(\gamepad_pmod.driver.shift_reg[7] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0061_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold110 (.A(\player_constroller_inst.u_player_physics.velocity[2] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0078_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold112 (.A(\gamepad_pmod.decoder.data_reg[6] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold113 (.A(\gamepad_pmod.decoder.data_reg[8] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0377_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold115 (.A(\audio_inst.i_jump.decay_value[17] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0053_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold117 (.A(\ai_controller_inst.restart_counter[5] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0388_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold119 (.A(\audio_inst.i_jump.decay_value[13] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ai_controller_inst.restart_counter[2] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold121 (.A(_1968_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold122 (.A(\gamepad_pmod.driver.shift_reg[2] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0056_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold124 (.A(\audio_inst.i_jump.decay_value[3] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold125 (.A(\score_inst_2.x_offset[2] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold126 (.A(\score[11] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold127 (.A(\player_constroller_inst.u_player_physics.velocity[1] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0077_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold129 (.A(\gamepad_pmod.decoder.data_reg[7] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold130 (.A(\graphics_inst.hvsync_gen.vpos[0] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold131 (.A(\score[5] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold132 (.A(_1771_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold133 (.A(\audio_inst.i_jump.decay_value[0] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold134 (.A(\audio_inst.i_over.counter[2] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold135 (.A(\audio_inst.i_jump.decay_value[8] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold136 (.A(\audio_inst.i_jump.counter[16] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold137 (.A(\audio_inst.i_over.decay_value[13] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold138 (.A(\audio_inst.i_over.decay_value[12] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold139 (.A(\gamepad_pmod.driver.shift_reg[8] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0062_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold141 (.A(\gamepad_pmod.driver.shift_reg[3] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold142 (.A(\score[8] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold143 (.A(\audio_inst.i_jump.counter[6] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0132_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold145 (.A(\audio_inst.i_over.decay_value[8] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold146 (.A(\audio_inst.i_over.decay_value[5] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold147 (.A(\audio_inst.i_jump.decay_value[9] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ai_controller_inst.restart_counter[0] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0010_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0230_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold151 (.A(\audio_inst.i_over.decay_value[14] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold152 (.A(\gamepad_pmod.driver.shift_reg[10] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0064_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold154 (.A(\audio_inst.i_over.decay_value[3] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold155 (.A(\audio_inst.i_jump.decay_value[11] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0174_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold157 (.A(\player_constroller_inst.u_player_physics.velocity[0] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0019_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold159 (.A(_1945_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold160 (.A(\audio_inst.i_jump.decay_value[6] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold161 (.A(\score[7] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold162 (.A(_1729_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold163 (.A(_1740_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold164 (.A(\audio_inst.i_jump.decay_value[4] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold165 (.A(\audio_inst.i_jump.decay_value[10] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold166 (.A(\audio_inst.i_over.counter[16] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold167 (.A(\audio_inst.i_over.decay_value[4] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold168 (.A(\audio_inst.i_jump.counter[11] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold169 (.A(\obstacles_inst.obstacle1_cross_gen_line_reg ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0486_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold171 (.A(\lfsr_inst.r_lfsr[6] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0085_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold173 (.A(\score[18] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold174 (.A(\audio_inst.i_over.decay_value[6] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0032_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold176 (.A(\gamepad_pmod.driver.shift_reg[5] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0059_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold178 (.A(\obs_rom_inst_2.i_obs_type[2] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0084_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold180 (.A(\score[0] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold181 (.A(_1736_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold182 (.A(\player_constroller_inst.game_over ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold183 (.A(_2189_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold184 (.A(\ai_controller_inst.obstacle1_pos[9] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0103_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold186 (.A(\audio_inst.i_over.counter[7] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold187 (.A(_1859_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold188 (.A(\audio_inst.i_over.counter[5] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1855_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold190 (.A(\audio_inst.i_over.decay_value[2] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold191 (.A(\gamepad_pmod.driver.shift_reg[4] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0058_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold193 (.A(\lfsr_inst.r_lfsr[15] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold194 (.A(\lfsr_inst.r_lfsr[7] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold195 (.A(\bg_object_inst.bg_object_pos[9] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0111_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold197 (.A(\audio_inst.i_over.counter[3] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold198 (.A(\audio_inst.i_over.counter[1] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold199 (.A(_1848_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold200 (.A(\audio_inst.i_jump.counter[13] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0139_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0020_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold203 (.A(_1943_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold204 (.A(\audio_inst.i_over.decay_value[15] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold205 (.A(\lfsr_inst.r_lfsr[8] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0087_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold207 (.A(\audio_inst.i_over.decay_value[9] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold208 (.A(\score[17] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold209 (.A(\ai_controller_inst.restart_counter[1] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold210 (.A(\audio_inst.i_jump.decay_value[14] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0161_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold212 (.A(\audio_inst.i_jump.counter[17] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0143_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold214 (.A(\dino_inst.i_ypos[2] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold215 (.A(\player_constroller_inst.game_state[5] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold216 (.A(_2179_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0011_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold218 (.A(\lfsr_inst.r_lfsr[3] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold219 (.A(\bg_object_inst.bg_object_pos[4] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0106_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold221 (.A(\audio_inst.i_over.decay_value[10] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0155_),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold223 (.A(\audio_inst.i_over.counter[17] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold224 (.A(\obstacles_inst.obstacle2_cross_gen_line_reg ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold225 (.A(\ai_controller_inst.restart_counter[4] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold226 (.A(_1973_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold227 (.A(\audio_inst.i_jump.counter[9] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0135_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold229 (.A(\graphics_inst.color_decoder_inst.rgb_scheme ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold230 (.A(\audio_inst.i_over.decay_value[11] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0156_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold232 (.A(\audio_inst.i_jump.counter[18] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold233 (.A(\audio_inst.i_jump.counter[15] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0141_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold235 (.A(\audio_inst.i_jump.wave_out ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0363_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold237 (.A(\ai_controller_inst.restart_counter[3] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold238 (.A(\audio_inst.i_jump.counter[2] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold239 (.A(\graphics_inst.hvsync_gen.vpos[1] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0026_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0342_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold242 (.A(\lfsr_inst.r_lfsr[5] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold243 (.A(\audio_inst.i_over.counter[0] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0343_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold245 (.A(\audio_inst.i_jump.counter[5] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0131_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold247 (.A(\obs_rom_inst_2.i_obs_type[1] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold248 (.A(\score[8] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold249 (.A(_1761_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold250 (.A(\ai_controller_inst.obstacle1_pos[5] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0099_),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold252 (.A(\dino_inst.i_ypos[0] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold253 (.A(\player_constroller_inst.game_state[1] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0001_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold255 (.A(\obs_rom_inst_1.i_obs_type[1] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold256 (.A(\audio_inst.i_jump.state[0] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold257 (.A(_2199_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold258 (.A(\ai_controller_inst.button_start ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0393_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold260 (.A(\ai_controller_inst.button_up ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold261 (.A(\ai_controller_inst.obstacle2_pos[9] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold262 (.A(\audio_inst.i_over.counter[8] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold263 (.A(\audio_inst.i_jump.counter[4] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0130_),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold265 (.A(\audio_inst.i_over.counter[9] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold266 (.A(\graphics_inst.frame_counter[0] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold267 (.A(\audio_inst.i_over.counter[6] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold268 (.A(\audio_inst.i_jump.counter[10] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0029_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold270 (.A(\audio_inst.i_jump.counter[8] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold271 (.A(\lfsr_inst.r_lfsr[4] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold272 (.A(\audio_inst.i_jump.counter[12] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold273 (.A(\ai_controller_inst.obstacle1_pos[4] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold274 (.A(\bg_line_inst.i_vpos[4] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold275 (.A(\graphics_inst.hpos[0] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0397_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0409_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold278 (.A(\ai_controller_inst.obstacle1_pos[7] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0549_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold280 (.A(\ai_controller_inst.obstacle2_pos[2] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0088_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold282 (.A(\bg_object_inst.bg_object_pos[2] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0104_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold284 (.A(\dino_inst.i_ypos[3] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold285 (.A(\ai_controller_inst.obstacle2_pos[4] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold286 (.A(\bg_object_inst.bg_object_pos[5] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0570_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold288 (.A(\score_inst_5.x_offset[6] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold289 (.A(\audio_inst.i_jump.counter[1] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0127_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold291 (.A(\dino_inst.i_ypos[0] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold292 (.A(\ai_controller_inst.obstacle2_pos[6] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0522_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold294 (.A(\bg_object_inst.bg_object_pos[6] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0573_),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold296 (.A(\player_constroller_inst.game_state[3] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold297 (.A(_2180_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0003_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold299 (.A(\player_constroller_inst.u_player_physics.velocity[3] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0462_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold301 (.A(\graphics_inst.game_tick_r ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0002_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold303 (.A(\score_inst_1.x_offset[4] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold304 (.A(\audio_inst.i_over.counter[12] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold305 (.A(_1869_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold306 (.A(\dino_inst.i_ypos[4] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0016_),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0096_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold309 (.A(\audio_inst.i_over.counter[4] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold310 (.A(\audio_inst.i_over.stage_index[3] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold311 (.A(\bg_object_inst.bg_object_pos[7] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0109_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0031_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold314 (.A(\audio_inst.i_over.stage_index[2] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold315 (.A(\lfsr_inst.r_lfsr[2] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold316 (.A(\audio_inst.i_over.counter[13] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold317 (.A(\bg_line_inst.i_vpos[9] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold318 (.A(\dino_inst.i_ypos[1] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold319 (.A(\ai_controller_inst.obstacle1_pos[3] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0097_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold321 (.A(\audio_inst.i_over.counter[11] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold322 (.A(_1867_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold323 (.A(\ai_controller_inst.obstacle2_pos[3] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold324 (.A(\graphics_inst.hpos[1] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold325 (.A(\audio_inst.i_over.state[1] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0396_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold327 (.A(\bg_object_inst.bg_object_pos[3] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold328 (.A(\audio_inst.i_over.counter[10] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold329 (.A(\ai_controller_inst.obstacle1_pos[6] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold330 (.A(\bg_line_inst.i_vpos[6] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold331 (.A(net551),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold332 (.A(\audio_inst.i_over.stage_index[1] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0011_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold334 (.A(\ai_controller_inst.obstacle2_pos[5] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold335 (.A(\audio_inst.i_jump.stage_index[2] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold336 (.A(_1941_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold337 (.A(\bg_object_inst.bg_object_pos[8] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold338 (.A(\audio_inst.i_over.counter[14] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold339 (.A(\bg_render_inst.i_hpos[2] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold340 (.A(\bg_line_inst.i_vpos[8] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold341 (.A(\ai_controller_inst.button_down ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0030_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold343 (.A(\ai_controller_inst.obstacle1_pos[8] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold344 (.A(\bg_render_inst.i_hpos[4] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold345 (.A(\ai_controller_inst.obstacle2_pos[8] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0529_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold347 (.A(\ai_controller_inst.obstacle2_pos[7] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold348 (.A(\audio_inst.i_jump.stage_index[1] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold349 (.A(_1938_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0010_),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold351 (.A(\audio_inst.i_jump.state[1] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0036_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold353 (.A(\graphics_inst.hvsync_gen.vpos[0] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold354 (.A(\ai_controller_inst.obstacle1_pos[2] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold355 (.A(\audio_inst.i_over.counter[15] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold356 (.A(\dino_inst.i_ypos[5] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold357 (.A(\bg_object_inst.bg_object_pos[3] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold358 (.A(\bg_line_inst.i_vpos[9] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0032_),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold360 (.A(\audio_inst.i_jump.counter[10] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold361 (.A(\audio_inst.i_jump.counter[1] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold362 (.A(\audio_inst.i_jump.counter[2] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0661_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold364 (.A(\ai_controller_inst.obstacle2_pos[7] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0528_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold366 (.A(\ai_controller_inst.obstacle1_pos[6] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold367 (.A(\audio_inst.i_over.counter[11] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold368 (.A(_1870_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold369 (.A(\audio_inst.i_jump.counter[13] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold370 (.A(\dino_inst.i_ypos[5] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold371 (.A(\ai_controller_inst.obstacle2_pos[2] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold372 (.A(\audio_inst.i_over.counter[0] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold373 (.A(\audio_inst.i_jump.counter[10] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0138_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0026_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold376 (.A(\ai_controller_inst.obstacle2_pos[2] ),
    .X(net918));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_fill_1 FILLER_0_56 ();
 sg13g2_fill_2 FILLER_0_74 ();
 sg13g2_fill_1 FILLER_0_76 ();
 sg13g2_fill_2 FILLER_0_85 ();
 sg13g2_fill_1 FILLER_0_87 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_fill_1 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_4 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_176 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_fill_1 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_fill_1 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_fill_1 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_4 FILLER_0_287 ();
 sg13g2_fill_1 FILLER_0_291 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_fill_2 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_85 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_fill_2 FILLER_1_140 ();
 sg13g2_fill_1 FILLER_1_168 ();
 sg13g2_fill_2 FILLER_1_203 ();
 sg13g2_fill_2 FILLER_1_249 ();
 sg13g2_fill_2 FILLER_1_277 ();
 sg13g2_fill_1 FILLER_1_279 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_4 FILLER_2_28 ();
 sg13g2_fill_2 FILLER_2_32 ();
 sg13g2_fill_1 FILLER_2_60 ();
 sg13g2_fill_2 FILLER_2_125 ();
 sg13g2_fill_1 FILLER_2_127 ();
 sg13g2_fill_2 FILLER_2_154 ();
 sg13g2_fill_1 FILLER_2_156 ();
 sg13g2_fill_2 FILLER_2_183 ();
 sg13g2_fill_1 FILLER_2_191 ();
 sg13g2_fill_1 FILLER_2_207 ();
 sg13g2_fill_1 FILLER_2_270 ();
 sg13g2_fill_2 FILLER_2_302 ();
 sg13g2_fill_2 FILLER_2_310 ();
 sg13g2_fill_1 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_4 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_118 ();
 sg13g2_decap_4 FILLER_3_125 ();
 sg13g2_fill_1 FILLER_3_129 ();
 sg13g2_fill_1 FILLER_3_156 ();
 sg13g2_fill_2 FILLER_3_169 ();
 sg13g2_fill_2 FILLER_3_192 ();
 sg13g2_fill_1 FILLER_3_194 ();
 sg13g2_fill_2 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_244 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_30 ();
 sg13g2_fill_2 FILLER_4_70 ();
 sg13g2_fill_2 FILLER_4_86 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_128 ();
 sg13g2_fill_2 FILLER_4_213 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_fill_2 FILLER_4_235 ();
 sg13g2_fill_1 FILLER_4_271 ();
 sg13g2_fill_2 FILLER_4_290 ();
 sg13g2_fill_1 FILLER_4_292 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_fill_1 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_65 ();
 sg13g2_fill_1 FILLER_5_72 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_fill_1 FILLER_5_91 ();
 sg13g2_fill_2 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_fill_2 FILLER_5_130 ();
 sg13g2_fill_1 FILLER_5_132 ();
 sg13g2_fill_2 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_209 ();
 sg13g2_decap_4 FILLER_5_216 ();
 sg13g2_fill_2 FILLER_5_220 ();
 sg13g2_fill_2 FILLER_5_253 ();
 sg13g2_fill_1 FILLER_5_255 ();
 sg13g2_fill_1 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_4 FILLER_5_294 ();
 sg13g2_fill_1 FILLER_5_298 ();
 sg13g2_fill_2 FILLER_5_309 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_fill_2 FILLER_5_330 ();
 sg13g2_fill_2 FILLER_5_337 ();
 sg13g2_fill_1 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_4 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_25 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_180 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_fill_2 FILLER_6_207 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_decap_8 FILLER_6_240 ();
 sg13g2_fill_1 FILLER_6_247 ();
 sg13g2_fill_2 FILLER_6_282 ();
 sg13g2_decap_8 FILLER_6_295 ();
 sg13g2_fill_2 FILLER_6_306 ();
 sg13g2_fill_1 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_18 ();
 sg13g2_fill_2 FILLER_7_77 ();
 sg13g2_fill_2 FILLER_7_174 ();
 sg13g2_decap_4 FILLER_7_193 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_229 ();
 sg13g2_fill_2 FILLER_7_236 ();
 sg13g2_fill_1 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_257 ();
 sg13g2_fill_2 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_271 ();
 sg13g2_fill_1 FILLER_7_276 ();
 sg13g2_fill_1 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_28 ();
 sg13g2_fill_2 FILLER_8_65 ();
 sg13g2_fill_2 FILLER_8_89 ();
 sg13g2_fill_1 FILLER_8_100 ();
 sg13g2_fill_2 FILLER_8_140 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_fill_2 FILLER_8_152 ();
 sg13g2_fill_1 FILLER_8_154 ();
 sg13g2_fill_2 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_fill_1 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_1 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_297 ();
 sg13g2_fill_2 FILLER_8_304 ();
 sg13g2_fill_1 FILLER_8_306 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_fill_2 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_59 ();
 sg13g2_fill_2 FILLER_9_123 ();
 sg13g2_fill_1 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_135 ();
 sg13g2_decap_4 FILLER_9_150 ();
 sg13g2_fill_1 FILLER_9_168 ();
 sg13g2_fill_2 FILLER_9_204 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_fill_2 FILLER_9_231 ();
 sg13g2_decap_4 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_297 ();
 sg13g2_fill_2 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_2 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_28 ();
 sg13g2_fill_2 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_85 ();
 sg13g2_fill_2 FILLER_10_121 ();
 sg13g2_fill_1 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_129 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_171 ();
 sg13g2_fill_2 FILLER_10_206 ();
 sg13g2_fill_1 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_219 ();
 sg13g2_fill_2 FILLER_10_236 ();
 sg13g2_fill_1 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_decap_4 FILLER_10_393 ();
 sg13g2_fill_1 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_33 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_142 ();
 sg13g2_decap_4 FILLER_11_199 ();
 sg13g2_fill_2 FILLER_11_241 ();
 sg13g2_fill_1 FILLER_11_243 ();
 sg13g2_fill_2 FILLER_11_254 ();
 sg13g2_fill_1 FILLER_11_256 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_270 ();
 sg13g2_fill_2 FILLER_11_303 ();
 sg13g2_fill_2 FILLER_11_362 ();
 sg13g2_fill_1 FILLER_11_364 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_4 ();
 sg13g2_fill_2 FILLER_12_78 ();
 sg13g2_fill_2 FILLER_12_124 ();
 sg13g2_decap_4 FILLER_12_140 ();
 sg13g2_fill_2 FILLER_12_149 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_205 ();
 sg13g2_fill_2 FILLER_12_221 ();
 sg13g2_fill_2 FILLER_12_250 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_4 FILLER_12_324 ();
 sg13g2_fill_2 FILLER_12_354 ();
 sg13g2_fill_1 FILLER_12_356 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_113 ();
 sg13g2_fill_2 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_195 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_235 ();
 sg13g2_decap_4 FILLER_13_250 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_4 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_fill_2 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_324 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_351 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_1 FILLER_14_17 ();
 sg13g2_decap_8 FILLER_14_40 ();
 sg13g2_fill_1 FILLER_14_47 ();
 sg13g2_fill_2 FILLER_14_60 ();
 sg13g2_fill_2 FILLER_14_66 ();
 sg13g2_decap_8 FILLER_14_86 ();
 sg13g2_fill_2 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_decap_4 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_156 ();
 sg13g2_fill_2 FILLER_14_188 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_decap_4 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_decap_8 FILLER_14_281 ();
 sg13g2_fill_2 FILLER_14_288 ();
 sg13g2_fill_2 FILLER_14_325 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_36 ();
 sg13g2_decap_4 FILLER_15_43 ();
 sg13g2_fill_2 FILLER_15_58 ();
 sg13g2_fill_2 FILLER_15_69 ();
 sg13g2_fill_1 FILLER_15_71 ();
 sg13g2_decap_4 FILLER_15_100 ();
 sg13g2_fill_1 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_114 ();
 sg13g2_decap_8 FILLER_15_121 ();
 sg13g2_fill_2 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_156 ();
 sg13g2_decap_8 FILLER_15_222 ();
 sg13g2_decap_8 FILLER_15_229 ();
 sg13g2_fill_1 FILLER_15_236 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_decap_4 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_360 ();
 sg13g2_fill_2 FILLER_16_22 ();
 sg13g2_fill_1 FILLER_16_24 ();
 sg13g2_fill_2 FILLER_16_76 ();
 sg13g2_fill_1 FILLER_16_78 ();
 sg13g2_fill_2 FILLER_16_123 ();
 sg13g2_fill_1 FILLER_16_133 ();
 sg13g2_decap_4 FILLER_16_137 ();
 sg13g2_decap_4 FILLER_16_145 ();
 sg13g2_fill_1 FILLER_16_149 ();
 sg13g2_fill_2 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_fill_1 FILLER_16_254 ();
 sg13g2_fill_2 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_145 ();
 sg13g2_decap_4 FILLER_17_152 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_fill_2 FILLER_17_184 ();
 sg13g2_decap_4 FILLER_17_253 ();
 sg13g2_fill_2 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_51 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_decap_8 FILLER_18_174 ();
 sg13g2_decap_8 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_261 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_fill_2 FILLER_18_301 ();
 sg13g2_fill_1 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_fill_2 FILLER_18_335 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_11 ();
 sg13g2_fill_2 FILLER_19_27 ();
 sg13g2_fill_1 FILLER_19_29 ();
 sg13g2_fill_2 FILLER_19_46 ();
 sg13g2_fill_2 FILLER_19_61 ();
 sg13g2_fill_2 FILLER_19_120 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_decap_4 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_185 ();
 sg13g2_decap_8 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_fill_2 FILLER_19_232 ();
 sg13g2_decap_4 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_289 ();
 sg13g2_decap_4 FILLER_19_296 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_decap_4 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_375 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_115 ();
 sg13g2_fill_2 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_fill_1 FILLER_20_159 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_12 ();
 sg13g2_fill_1 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_38 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_199 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_decap_4 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_247 ();
 sg13g2_fill_2 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_353 ();
 sg13g2_fill_2 FILLER_21_381 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_2 FILLER_22_12 ();
 sg13g2_fill_1 FILLER_22_29 ();
 sg13g2_fill_2 FILLER_22_44 ();
 sg13g2_fill_1 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_111 ();
 sg13g2_fill_2 FILLER_22_129 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_fill_1 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_195 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_decap_8 FILLER_22_281 ();
 sg13g2_fill_2 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_290 ();
 sg13g2_fill_2 FILLER_22_299 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_27 ();
 sg13g2_fill_1 FILLER_23_29 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_249 ();
 sg13g2_fill_2 FILLER_23_260 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_fill_2 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_11 ();
 sg13g2_fill_2 FILLER_24_50 ();
 sg13g2_fill_2 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_178 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_4 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_24 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_fill_2 FILLER_25_270 ();
 sg13g2_fill_2 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_fill_2 FILLER_26_26 ();
 sg13g2_fill_2 FILLER_26_45 ();
 sg13g2_fill_1 FILLER_26_47 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_decap_4 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_4 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_229 ();
 sg13g2_decap_4 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_16 ();
 sg13g2_fill_1 FILLER_27_32 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_fill_1 FILLER_27_198 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_decap_4 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_252 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_301 ();
 sg13g2_fill_2 FILLER_27_370 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_117 ();
 sg13g2_fill_2 FILLER_28_136 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_8 FILLER_28_212 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_decap_8 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_243 ();
 sg13g2_decap_4 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_254 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_decap_4 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_decap_4 FILLER_28_289 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_333 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_decap_4 FILLER_29_222 ();
 sg13g2_fill_2 FILLER_29_226 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_19 ();
 sg13g2_fill_1 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_166 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_211 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_276 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_38 ();
 sg13g2_fill_2 FILLER_31_45 ();
 sg13g2_fill_2 FILLER_31_55 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_decap_4 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_59 ();
 sg13g2_decap_8 FILLER_32_64 ();
 sg13g2_decap_4 FILLER_32_71 ();
 sg13g2_fill_2 FILLER_32_75 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_90 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_decap_4 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_decap_4 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_decap_4 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_372 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_decap_4 FILLER_33_78 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_124 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_222 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_2 FILLER_33_286 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_34_26 ();
 sg13g2_fill_2 FILLER_34_32 ();
 sg13g2_decap_8 FILLER_34_104 ();
 sg13g2_decap_4 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_2 FILLER_34_156 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_360 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_50 ();
 sg13g2_fill_2 FILLER_35_110 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_decap_4 FILLER_35_153 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_239 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_319 ();
 sg13g2_decap_8 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_4 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_fill_2 FILLER_36_20 ();
 sg13g2_fill_1 FILLER_36_22 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_fill_2 FILLER_36_138 ();
 sg13g2_fill_2 FILLER_36_158 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_204 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_367 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_15 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_fill_1 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_164 ();
 sg13g2_fill_1 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_180 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_201 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_213 ();
 sg13g2_decap_4 FILLER_37_220 ();
 sg13g2_decap_4 FILLER_37_245 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_271 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_decap_4 FILLER_37_280 ();
 sg13g2_fill_1 FILLER_37_284 ();
 sg13g2_fill_2 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_150 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_decap_4 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_fill_1 FILLER_39_88 ();
 sg13g2_fill_2 FILLER_39_135 ();
 sg13g2_fill_1 FILLER_39_137 ();
 sg13g2_decap_8 FILLER_39_152 ();
 sg13g2_decap_8 FILLER_39_159 ();
 sg13g2_decap_8 FILLER_39_166 ();
 sg13g2_decap_4 FILLER_39_182 ();
 sg13g2_fill_1 FILLER_39_191 ();
 sg13g2_fill_2 FILLER_39_231 ();
 sg13g2_fill_1 FILLER_39_233 ();
 sg13g2_decap_4 FILLER_39_248 ();
 sg13g2_fill_2 FILLER_39_252 ();
 sg13g2_fill_2 FILLER_39_263 ();
 sg13g2_fill_1 FILLER_39_265 ();
 sg13g2_decap_8 FILLER_39_292 ();
 sg13g2_decap_8 FILLER_39_299 ();
 sg13g2_decap_8 FILLER_39_306 ();
 sg13g2_decap_8 FILLER_39_313 ();
 sg13g2_decap_8 FILLER_39_320 ();
 sg13g2_decap_8 FILLER_39_327 ();
 sg13g2_decap_4 FILLER_39_334 ();
 sg13g2_fill_2 FILLER_39_338 ();
 sg13g2_decap_8 FILLER_39_344 ();
 sg13g2_fill_2 FILLER_39_356 ();
 sg13g2_fill_1 FILLER_39_358 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_4 FILLER_40_28 ();
 sg13g2_fill_2 FILLER_40_32 ();
 sg13g2_fill_1 FILLER_40_51 ();
 sg13g2_fill_1 FILLER_40_87 ();
 sg13g2_fill_1 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_142 ();
 sg13g2_fill_1 FILLER_40_144 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_205 ();
 sg13g2_fill_1 FILLER_40_212 ();
 sg13g2_fill_1 FILLER_40_222 ();
 sg13g2_decap_4 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_345 ();
 sg13g2_decap_4 FILLER_40_352 ();
 sg13g2_fill_2 FILLER_40_356 ();
 sg13g2_decap_8 FILLER_40_375 ();
 sg13g2_fill_2 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_393 ();
 sg13g2_fill_2 FILLER_40_400 ();
 sg13g2_fill_1 FILLER_40_402 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_4 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_46 ();
 sg13g2_decap_4 FILLER_41_52 ();
 sg13g2_decap_8 FILLER_41_109 ();
 sg13g2_decap_8 FILLER_41_116 ();
 sg13g2_fill_2 FILLER_41_123 ();
 sg13g2_fill_1 FILLER_41_125 ();
 sg13g2_decap_4 FILLER_41_131 ();
 sg13g2_fill_2 FILLER_41_135 ();
 sg13g2_fill_1 FILLER_41_198 ();
 sg13g2_decap_8 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_228 ();
 sg13g2_fill_1 FILLER_41_230 ();
 sg13g2_fill_1 FILLER_41_261 ();
 sg13g2_fill_2 FILLER_41_288 ();
 sg13g2_fill_2 FILLER_41_302 ();
 sg13g2_decap_4 FILLER_41_360 ();
 sg13g2_fill_1 FILLER_41_364 ();
 sg13g2_fill_2 FILLER_41_368 ();
 sg13g2_fill_1 FILLER_41_373 ();
 sg13g2_decap_8 FILLER_41_377 ();
 sg13g2_decap_8 FILLER_41_384 ();
 sg13g2_decap_8 FILLER_41_401 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_28 ();
 sg13g2_fill_1 FILLER_42_30 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_115 ();
 sg13g2_decap_8 FILLER_42_125 ();
 sg13g2_fill_1 FILLER_42_132 ();
 sg13g2_fill_2 FILLER_42_147 ();
 sg13g2_fill_2 FILLER_42_153 ();
 sg13g2_fill_1 FILLER_42_155 ();
 sg13g2_decap_8 FILLER_42_174 ();
 sg13g2_decap_8 FILLER_42_181 ();
 sg13g2_decap_8 FILLER_42_188 ();
 sg13g2_decap_8 FILLER_42_195 ();
 sg13g2_decap_4 FILLER_42_202 ();
 sg13g2_decap_4 FILLER_42_227 ();
 sg13g2_fill_1 FILLER_42_257 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_277 ();
 sg13g2_decap_8 FILLER_42_282 ();
 sg13g2_decap_4 FILLER_42_294 ();
 sg13g2_fill_2 FILLER_42_298 ();
 sg13g2_fill_2 FILLER_42_304 ();
 sg13g2_fill_1 FILLER_42_306 ();
 sg13g2_fill_2 FILLER_42_369 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_53 ();
 sg13g2_decap_8 FILLER_43_60 ();
 sg13g2_decap_8 FILLER_43_67 ();
 sg13g2_fill_1 FILLER_43_74 ();
 sg13g2_fill_1 FILLER_43_89 ();
 sg13g2_decap_4 FILLER_43_136 ();
 sg13g2_fill_1 FILLER_43_140 ();
 sg13g2_decap_4 FILLER_43_167 ();
 sg13g2_fill_1 FILLER_43_171 ();
 sg13g2_fill_1 FILLER_43_201 ();
 sg13g2_fill_2 FILLER_43_239 ();
 sg13g2_fill_1 FILLER_43_241 ();
 sg13g2_fill_2 FILLER_43_251 ();
 sg13g2_fill_1 FILLER_43_253 ();
 sg13g2_decap_8 FILLER_43_276 ();
 sg13g2_decap_8 FILLER_43_283 ();
 sg13g2_fill_2 FILLER_43_290 ();
 sg13g2_fill_1 FILLER_43_292 ();
 sg13g2_decap_4 FILLER_43_310 ();
 sg13g2_fill_1 FILLER_43_314 ();
 sg13g2_decap_8 FILLER_43_323 ();
 sg13g2_fill_2 FILLER_43_330 ();
 sg13g2_fill_1 FILLER_43_362 ();
 sg13g2_fill_2 FILLER_43_384 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_14 ();
 sg13g2_fill_1 FILLER_44_46 ();
 sg13g2_fill_2 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_58 ();
 sg13g2_decap_4 FILLER_44_67 ();
 sg13g2_fill_2 FILLER_44_79 ();
 sg13g2_decap_8 FILLER_44_89 ();
 sg13g2_decap_8 FILLER_44_96 ();
 sg13g2_fill_2 FILLER_44_103 ();
 sg13g2_decap_4 FILLER_44_109 ();
 sg13g2_fill_2 FILLER_44_164 ();
 sg13g2_decap_4 FILLER_44_171 ();
 sg13g2_fill_2 FILLER_44_215 ();
 sg13g2_decap_4 FILLER_44_232 ();
 sg13g2_fill_2 FILLER_44_267 ();
 sg13g2_fill_1 FILLER_44_269 ();
 sg13g2_fill_1 FILLER_44_287 ();
 sg13g2_decap_4 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_323 ();
 sg13g2_decap_4 FILLER_44_330 ();
 sg13g2_fill_1 FILLER_44_339 ();
 sg13g2_fill_1 FILLER_44_374 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_14 ();
 sg13g2_fill_1 FILLER_45_47 ();
 sg13g2_fill_2 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_72 ();
 sg13g2_fill_1 FILLER_45_79 ();
 sg13g2_fill_2 FILLER_45_106 ();
 sg13g2_fill_1 FILLER_45_108 ();
 sg13g2_decap_4 FILLER_45_122 ();
 sg13g2_fill_2 FILLER_45_136 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_fill_2 FILLER_45_165 ();
 sg13g2_fill_1 FILLER_45_167 ();
 sg13g2_fill_2 FILLER_45_178 ();
 sg13g2_fill_1 FILLER_45_180 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_fill_1 FILLER_45_314 ();
 sg13g2_fill_2 FILLER_45_324 ();
 sg13g2_fill_1 FILLER_45_326 ();
 sg13g2_decap_4 FILLER_45_336 ();
 sg13g2_fill_1 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_356 ();
 sg13g2_decap_8 FILLER_45_365 ();
 sg13g2_decap_8 FILLER_45_372 ();
 sg13g2_fill_1 FILLER_45_379 ();
 sg13g2_fill_1 FILLER_45_390 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_fill_1 FILLER_46_43 ();
 sg13g2_fill_2 FILLER_46_70 ();
 sg13g2_decap_4 FILLER_46_107 ();
 sg13g2_fill_1 FILLER_46_111 ();
 sg13g2_fill_2 FILLER_46_148 ();
 sg13g2_decap_8 FILLER_46_158 ();
 sg13g2_decap_4 FILLER_46_165 ();
 sg13g2_fill_2 FILLER_46_169 ();
 sg13g2_decap_8 FILLER_46_198 ();
 sg13g2_decap_8 FILLER_46_205 ();
 sg13g2_fill_2 FILLER_46_212 ();
 sg13g2_fill_1 FILLER_46_223 ();
 sg13g2_fill_2 FILLER_46_238 ();
 sg13g2_fill_1 FILLER_46_240 ();
 sg13g2_fill_1 FILLER_46_252 ();
 sg13g2_fill_2 FILLER_46_300 ();
 sg13g2_fill_1 FILLER_46_324 ();
 sg13g2_fill_1 FILLER_46_337 ();
 sg13g2_decap_8 FILLER_46_356 ();
 sg13g2_decap_8 FILLER_46_363 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_fill_1 FILLER_46_376 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_40 ();
 sg13g2_fill_1 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_64 ();
 sg13g2_fill_2 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_107 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_4 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_170 ();
 sg13g2_decap_8 FILLER_47_177 ();
 sg13g2_decap_8 FILLER_47_184 ();
 sg13g2_decap_4 FILLER_47_191 ();
 sg13g2_fill_2 FILLER_47_195 ();
 sg13g2_decap_4 FILLER_47_201 ();
 sg13g2_fill_2 FILLER_47_205 ();
 sg13g2_fill_1 FILLER_47_215 ();
 sg13g2_fill_1 FILLER_47_233 ();
 sg13g2_fill_2 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_275 ();
 sg13g2_decap_8 FILLER_47_282 ();
 sg13g2_fill_2 FILLER_47_289 ();
 sg13g2_fill_2 FILLER_47_328 ();
 sg13g2_fill_1 FILLER_47_330 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_11 ();
 sg13g2_fill_1 FILLER_48_20 ();
 sg13g2_fill_2 FILLER_48_37 ();
 sg13g2_fill_1 FILLER_48_39 ();
 sg13g2_fill_2 FILLER_48_63 ();
 sg13g2_fill_1 FILLER_48_90 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_decap_4 FILLER_48_123 ();
 sg13g2_fill_2 FILLER_48_140 ();
 sg13g2_fill_2 FILLER_48_146 ();
 sg13g2_decap_4 FILLER_48_187 ();
 sg13g2_fill_2 FILLER_48_191 ();
 sg13g2_fill_1 FILLER_48_232 ();
 sg13g2_fill_2 FILLER_48_250 ();
 sg13g2_fill_1 FILLER_48_252 ();
 sg13g2_fill_2 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_290 ();
 sg13g2_decap_8 FILLER_48_295 ();
 sg13g2_fill_1 FILLER_48_307 ();
 sg13g2_fill_2 FILLER_48_317 ();
 sg13g2_fill_1 FILLER_48_319 ();
 sg13g2_fill_1 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_8 ();
 sg13g2_fill_1 FILLER_49_34 ();
 sg13g2_fill_1 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_68 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_fill_1 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_109 ();
 sg13g2_fill_1 FILLER_49_111 ();
 sg13g2_fill_2 FILLER_49_116 ();
 sg13g2_fill_1 FILLER_49_118 ();
 sg13g2_fill_2 FILLER_49_133 ();
 sg13g2_fill_2 FILLER_49_169 ();
 sg13g2_fill_2 FILLER_49_197 ();
 sg13g2_fill_1 FILLER_49_199 ();
 sg13g2_fill_2 FILLER_49_219 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_fill_1 FILLER_49_239 ();
 sg13g2_fill_1 FILLER_49_244 ();
 sg13g2_fill_1 FILLER_49_279 ();
 sg13g2_decap_8 FILLER_49_306 ();
 sg13g2_decap_8 FILLER_49_313 ();
 sg13g2_decap_8 FILLER_49_320 ();
 sg13g2_decap_4 FILLER_49_327 ();
 sg13g2_decap_8 FILLER_49_345 ();
 sg13g2_decap_8 FILLER_49_352 ();
 sg13g2_fill_2 FILLER_49_364 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_fill_1 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_27 ();
 sg13g2_fill_1 FILLER_50_29 ();
 sg13g2_fill_1 FILLER_50_48 ();
 sg13g2_fill_1 FILLER_50_54 ();
 sg13g2_fill_2 FILLER_50_66 ();
 sg13g2_fill_1 FILLER_50_68 ();
 sg13g2_fill_2 FILLER_50_99 ();
 sg13g2_fill_2 FILLER_50_127 ();
 sg13g2_fill_2 FILLER_50_156 ();
 sg13g2_fill_1 FILLER_50_158 ();
 sg13g2_fill_1 FILLER_50_167 ();
 sg13g2_fill_1 FILLER_50_176 ();
 sg13g2_fill_2 FILLER_50_211 ();
 sg13g2_fill_1 FILLER_50_213 ();
 sg13g2_decap_4 FILLER_50_227 ();
 sg13g2_fill_1 FILLER_50_231 ();
 sg13g2_fill_1 FILLER_50_298 ();
 sg13g2_decap_8 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_313 ();
 sg13g2_decap_8 FILLER_50_326 ();
 sg13g2_decap_8 FILLER_50_333 ();
 sg13g2_fill_2 FILLER_50_340 ();
 sg13g2_fill_1 FILLER_50_342 ();
 sg13g2_fill_1 FILLER_50_347 ();
 sg13g2_fill_2 FILLER_50_361 ();
 sg13g2_fill_2 FILLER_50_381 ();
 sg13g2_fill_1 FILLER_50_383 ();
 sg13g2_fill_1 FILLER_50_396 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_2 FILLER_51_72 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_fill_2 FILLER_51_87 ();
 sg13g2_fill_1 FILLER_51_89 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_4 FILLER_51_119 ();
 sg13g2_fill_1 FILLER_51_123 ();
 sg13g2_fill_1 FILLER_51_153 ();
 sg13g2_fill_2 FILLER_51_166 ();
 sg13g2_fill_1 FILLER_51_173 ();
 sg13g2_fill_2 FILLER_51_184 ();
 sg13g2_fill_1 FILLER_51_186 ();
 sg13g2_decap_8 FILLER_51_191 ();
 sg13g2_decap_8 FILLER_51_198 ();
 sg13g2_decap_8 FILLER_51_205 ();
 sg13g2_fill_2 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_decap_8 FILLER_51_231 ();
 sg13g2_decap_4 FILLER_51_238 ();
 sg13g2_fill_1 FILLER_51_242 ();
 sg13g2_decap_4 FILLER_51_247 ();
 sg13g2_fill_1 FILLER_51_251 ();
 sg13g2_fill_2 FILLER_51_260 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_fill_1 FILLER_51_286 ();
 sg13g2_fill_2 FILLER_51_329 ();
 sg13g2_fill_2 FILLER_51_384 ();
 sg13g2_fill_1 FILLER_51_386 ();
 sg13g2_fill_2 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_52_11 ();
 sg13g2_fill_2 FILLER_52_17 ();
 sg13g2_fill_1 FILLER_52_33 ();
 sg13g2_decap_4 FILLER_52_79 ();
 sg13g2_fill_1 FILLER_52_83 ();
 sg13g2_decap_4 FILLER_52_94 ();
 sg13g2_fill_2 FILLER_52_98 ();
 sg13g2_fill_1 FILLER_52_135 ();
 sg13g2_decap_8 FILLER_52_198 ();
 sg13g2_fill_2 FILLER_52_205 ();
 sg13g2_fill_1 FILLER_52_207 ();
 sg13g2_fill_2 FILLER_52_217 ();
 sg13g2_fill_1 FILLER_52_219 ();
 sg13g2_decap_4 FILLER_52_226 ();
 sg13g2_fill_2 FILLER_52_264 ();
 sg13g2_fill_1 FILLER_52_301 ();
 sg13g2_fill_1 FILLER_52_316 ();
 sg13g2_fill_1 FILLER_52_348 ();
 sg13g2_fill_1 FILLER_52_363 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_20 ();
 sg13g2_fill_1 FILLER_53_22 ();
 sg13g2_fill_2 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_37 ();
 sg13g2_fill_1 FILLER_53_130 ();
 sg13g2_fill_2 FILLER_53_160 ();
 sg13g2_fill_1 FILLER_53_171 ();
 sg13g2_fill_1 FILLER_53_216 ();
 sg13g2_decap_4 FILLER_53_248 ();
 sg13g2_fill_1 FILLER_53_278 ();
 sg13g2_fill_2 FILLER_53_319 ();
 sg13g2_fill_1 FILLER_53_361 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_11 ();
 sg13g2_fill_1 FILLER_54_28 ();
 sg13g2_fill_1 FILLER_54_50 ();
 sg13g2_decap_4 FILLER_54_68 ();
 sg13g2_fill_2 FILLER_54_97 ();
 sg13g2_fill_1 FILLER_54_99 ();
 sg13g2_fill_1 FILLER_54_126 ();
 sg13g2_fill_1 FILLER_54_142 ();
 sg13g2_decap_4 FILLER_54_208 ();
 sg13g2_fill_2 FILLER_54_212 ();
 sg13g2_fill_2 FILLER_54_221 ();
 sg13g2_fill_1 FILLER_54_238 ();
 sg13g2_decap_8 FILLER_54_247 ();
 sg13g2_decap_8 FILLER_54_254 ();
 sg13g2_fill_2 FILLER_54_261 ();
 sg13g2_fill_2 FILLER_54_279 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_fill_2 FILLER_54_351 ();
 sg13g2_fill_2 FILLER_54_380 ();
 sg13g2_fill_2 FILLER_54_386 ();
 sg13g2_fill_2 FILLER_54_406 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_2 ();
 sg13g2_fill_1 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_33 ();
 sg13g2_fill_2 FILLER_55_43 ();
 sg13g2_fill_1 FILLER_55_45 ();
 sg13g2_fill_1 FILLER_55_77 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_1 FILLER_55_140 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_2 FILLER_55_199 ();
 sg13g2_decap_4 FILLER_55_254 ();
 sg13g2_fill_1 FILLER_55_258 ();
 sg13g2_fill_1 FILLER_55_307 ();
 sg13g2_fill_1 FILLER_55_322 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_fill_1 FILLER_56_28 ();
 sg13g2_fill_2 FILLER_56_34 ();
 sg13g2_decap_8 FILLER_56_48 ();
 sg13g2_fill_1 FILLER_56_55 ();
 sg13g2_decap_4 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_69 ();
 sg13g2_fill_1 FILLER_56_77 ();
 sg13g2_fill_1 FILLER_56_113 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_decap_8 FILLER_56_176 ();
 sg13g2_fill_2 FILLER_56_209 ();
 sg13g2_fill_1 FILLER_56_211 ();
 sg13g2_decap_4 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_251 ();
 sg13g2_decap_4 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_266 ();
 sg13g2_fill_2 FILLER_56_300 ();
 sg13g2_fill_2 FILLER_56_364 ();
 sg13g2_fill_2 FILLER_57_53 ();
 sg13g2_decap_8 FILLER_57_69 ();
 sg13g2_fill_2 FILLER_57_76 ();
 sg13g2_decap_4 FILLER_57_85 ();
 sg13g2_fill_1 FILLER_57_102 ();
 sg13g2_fill_1 FILLER_57_135 ();
 sg13g2_fill_1 FILLER_57_155 ();
 sg13g2_fill_1 FILLER_57_164 ();
 sg13g2_decap_8 FILLER_57_179 ();
 sg13g2_decap_4 FILLER_57_190 ();
 sg13g2_decap_8 FILLER_57_198 ();
 sg13g2_fill_2 FILLER_57_205 ();
 sg13g2_fill_2 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_234 ();
 sg13g2_fill_1 FILLER_57_241 ();
 sg13g2_fill_1 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_279 ();
 sg13g2_fill_1 FILLER_57_332 ();
 sg13g2_fill_1 FILLER_57_338 ();
 sg13g2_fill_1 FILLER_57_370 ();
 sg13g2_fill_2 FILLER_57_377 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_16 ();
 sg13g2_fill_2 FILLER_58_26 ();
 sg13g2_fill_2 FILLER_58_33 ();
 sg13g2_fill_2 FILLER_58_44 ();
 sg13g2_fill_2 FILLER_58_61 ();
 sg13g2_fill_2 FILLER_58_72 ();
 sg13g2_fill_1 FILLER_58_74 ();
 sg13g2_decap_8 FILLER_58_93 ();
 sg13g2_decap_4 FILLER_58_100 ();
 sg13g2_fill_1 FILLER_58_108 ();
 sg13g2_fill_1 FILLER_58_139 ();
 sg13g2_fill_2 FILLER_58_162 ();
 sg13g2_fill_2 FILLER_58_198 ();
 sg13g2_fill_1 FILLER_58_200 ();
 sg13g2_fill_1 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_226 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_262 ();
 sg13g2_fill_1 FILLER_58_264 ();
 sg13g2_decap_4 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_366 ();
 sg13g2_fill_1 FILLER_58_386 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_69 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_2 FILLER_59_177 ();
 sg13g2_decap_8 FILLER_59_205 ();
 sg13g2_decap_8 FILLER_59_216 ();
 sg13g2_decap_4 FILLER_59_223 ();
 sg13g2_fill_1 FILLER_59_236 ();
 sg13g2_decap_8 FILLER_59_309 ();
 sg13g2_fill_1 FILLER_59_324 ();
 sg13g2_fill_2 FILLER_59_334 ();
 sg13g2_fill_2 FILLER_59_362 ();
 sg13g2_fill_1 FILLER_59_377 ();
 sg13g2_fill_2 FILLER_59_383 ();
 sg13g2_fill_1 FILLER_59_385 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_fill_2 FILLER_60_30 ();
 sg13g2_fill_1 FILLER_60_32 ();
 sg13g2_fill_2 FILLER_60_53 ();
 sg13g2_decap_4 FILLER_60_65 ();
 sg13g2_fill_1 FILLER_60_69 ();
 sg13g2_fill_2 FILLER_60_79 ();
 sg13g2_fill_1 FILLER_60_81 ();
 sg13g2_fill_2 FILLER_60_119 ();
 sg13g2_fill_1 FILLER_60_121 ();
 sg13g2_fill_2 FILLER_60_158 ();
 sg13g2_fill_1 FILLER_60_185 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_fill_1 FILLER_60_193 ();
 sg13g2_fill_1 FILLER_60_220 ();
 sg13g2_fill_2 FILLER_60_229 ();
 sg13g2_fill_1 FILLER_60_244 ();
 sg13g2_fill_2 FILLER_60_287 ();
 sg13g2_fill_1 FILLER_60_309 ();
 sg13g2_decap_4 FILLER_60_323 ();
 sg13g2_fill_2 FILLER_60_336 ();
 sg13g2_decap_4 FILLER_60_364 ();
 sg13g2_fill_1 FILLER_60_368 ();
 sg13g2_fill_2 FILLER_60_387 ();
 sg13g2_decap_4 FILLER_60_405 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_12 ();
 sg13g2_fill_2 FILLER_61_23 ();
 sg13g2_fill_2 FILLER_61_34 ();
 sg13g2_fill_2 FILLER_61_41 ();
 sg13g2_decap_8 FILLER_61_52 ();
 sg13g2_decap_4 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_68 ();
 sg13g2_fill_1 FILLER_61_70 ();
 sg13g2_fill_2 FILLER_61_130 ();
 sg13g2_fill_1 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_188 ();
 sg13g2_decap_8 FILLER_61_194 ();
 sg13g2_fill_2 FILLER_61_201 ();
 sg13g2_fill_1 FILLER_61_203 ();
 sg13g2_decap_4 FILLER_61_208 ();
 sg13g2_fill_1 FILLER_61_225 ();
 sg13g2_fill_1 FILLER_61_293 ();
 sg13g2_decap_8 FILLER_61_359 ();
 sg13g2_decap_8 FILLER_61_366 ();
 sg13g2_decap_8 FILLER_61_373 ();
 sg13g2_fill_1 FILLER_61_380 ();
 sg13g2_decap_8 FILLER_61_402 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_4 FILLER_62_54 ();
 sg13g2_fill_1 FILLER_62_99 ();
 sg13g2_decap_8 FILLER_62_146 ();
 sg13g2_decap_4 FILLER_62_153 ();
 sg13g2_fill_2 FILLER_62_157 ();
 sg13g2_decap_8 FILLER_62_172 ();
 sg13g2_decap_4 FILLER_62_179 ();
 sg13g2_decap_8 FILLER_62_187 ();
 sg13g2_fill_1 FILLER_62_220 ();
 sg13g2_fill_2 FILLER_62_229 ();
 sg13g2_fill_1 FILLER_62_236 ();
 sg13g2_fill_2 FILLER_62_267 ();
 sg13g2_fill_2 FILLER_62_278 ();
 sg13g2_fill_1 FILLER_62_280 ();
 sg13g2_decap_4 FILLER_62_355 ();
 sg13g2_fill_2 FILLER_62_359 ();
 sg13g2_fill_1 FILLER_62_373 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_4 FILLER_62_385 ();
 sg13g2_fill_1 FILLER_62_389 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_decap_8 FILLER_62_402 ();
 sg13g2_decap_4 FILLER_63_47 ();
 sg13g2_fill_2 FILLER_63_64 ();
 sg13g2_decap_8 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_99 ();
 sg13g2_fill_2 FILLER_63_109 ();
 sg13g2_decap_4 FILLER_63_149 ();
 sg13g2_decap_8 FILLER_63_158 ();
 sg13g2_decap_4 FILLER_63_165 ();
 sg13g2_fill_1 FILLER_63_169 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_fill_2 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_209 ();
 sg13g2_decap_4 FILLER_63_220 ();
 sg13g2_fill_1 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_229 ();
 sg13g2_fill_2 FILLER_63_243 ();
 sg13g2_fill_2 FILLER_63_317 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_fill_2 FILLER_63_358 ();
 sg13g2_fill_1 FILLER_63_360 ();
 sg13g2_fill_1 FILLER_63_386 ();
 sg13g2_decap_4 FILLER_63_404 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_4 ();
 sg13g2_fill_2 FILLER_64_23 ();
 sg13g2_fill_2 FILLER_64_74 ();
 sg13g2_fill_1 FILLER_64_138 ();
 sg13g2_fill_1 FILLER_64_144 ();
 sg13g2_decap_8 FILLER_64_150 ();
 sg13g2_decap_4 FILLER_64_157 ();
 sg13g2_decap_8 FILLER_64_166 ();
 sg13g2_decap_8 FILLER_64_199 ();
 sg13g2_decap_8 FILLER_64_206 ();
 sg13g2_fill_2 FILLER_64_213 ();
 sg13g2_fill_1 FILLER_64_232 ();
 sg13g2_fill_1 FILLER_64_256 ();
 sg13g2_fill_2 FILLER_64_288 ();
 sg13g2_fill_2 FILLER_64_331 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_65 ();
 sg13g2_fill_1 FILLER_65_80 ();
 sg13g2_decap_4 FILLER_65_84 ();
 sg13g2_fill_2 FILLER_65_88 ();
 sg13g2_fill_1 FILLER_65_126 ();
 sg13g2_decap_4 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_203 ();
 sg13g2_fill_2 FILLER_65_221 ();
 sg13g2_fill_1 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_240 ();
 sg13g2_fill_1 FILLER_65_281 ();
 sg13g2_fill_2 FILLER_65_286 ();
 sg13g2_fill_1 FILLER_65_288 ();
 sg13g2_fill_2 FILLER_65_293 ();
 sg13g2_fill_2 FILLER_65_300 ();
 sg13g2_fill_1 FILLER_65_302 ();
 sg13g2_fill_1 FILLER_65_307 ();
 sg13g2_fill_1 FILLER_65_312 ();
 sg13g2_decap_8 FILLER_65_330 ();
 sg13g2_fill_2 FILLER_65_337 ();
 sg13g2_fill_1 FILLER_65_339 ();
 sg13g2_fill_1 FILLER_65_348 ();
 sg13g2_fill_1 FILLER_65_357 ();
 sg13g2_fill_2 FILLER_65_391 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_decap_8 FILLER_66_116 ();
 sg13g2_decap_4 FILLER_66_123 ();
 sg13g2_decap_8 FILLER_66_153 ();
 sg13g2_decap_8 FILLER_66_164 ();
 sg13g2_decap_8 FILLER_66_171 ();
 sg13g2_fill_2 FILLER_66_178 ();
 sg13g2_fill_1 FILLER_66_192 ();
 sg13g2_decap_4 FILLER_66_198 ();
 sg13g2_fill_2 FILLER_66_211 ();
 sg13g2_fill_2 FILLER_66_222 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_229 ();
 sg13g2_fill_2 FILLER_66_236 ();
 sg13g2_fill_2 FILLER_66_242 ();
 sg13g2_fill_1 FILLER_66_244 ();
 sg13g2_fill_2 FILLER_66_255 ();
 sg13g2_fill_2 FILLER_66_267 ();
 sg13g2_fill_2 FILLER_66_273 ();
 sg13g2_fill_1 FILLER_66_311 ();
 sg13g2_fill_2 FILLER_66_369 ();
 sg13g2_fill_1 FILLER_66_371 ();
 sg13g2_fill_1 FILLER_66_378 ();
 sg13g2_decap_4 FILLER_67_43 ();
 sg13g2_fill_1 FILLER_67_51 ();
 sg13g2_fill_2 FILLER_67_59 ();
 sg13g2_fill_2 FILLER_67_104 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_4 FILLER_67_126 ();
 sg13g2_fill_1 FILLER_67_130 ();
 sg13g2_decap_4 FILLER_67_163 ();
 sg13g2_fill_2 FILLER_67_167 ();
 sg13g2_decap_8 FILLER_67_174 ();
 sg13g2_decap_8 FILLER_67_181 ();
 sg13g2_decap_4 FILLER_67_188 ();
 sg13g2_fill_1 FILLER_67_192 ();
 sg13g2_fill_1 FILLER_67_207 ();
 sg13g2_decap_8 FILLER_67_227 ();
 sg13g2_fill_1 FILLER_67_234 ();
 sg13g2_fill_2 FILLER_67_247 ();
 sg13g2_fill_1 FILLER_67_249 ();
 sg13g2_decap_4 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_304 ();
 sg13g2_fill_2 FILLER_67_315 ();
 sg13g2_fill_2 FILLER_67_329 ();
 sg13g2_decap_8 FILLER_67_340 ();
 sg13g2_decap_8 FILLER_67_347 ();
 sg13g2_decap_8 FILLER_67_354 ();
 sg13g2_fill_1 FILLER_67_361 ();
 sg13g2_fill_1 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_fill_2 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_71 ();
 sg13g2_fill_1 FILLER_68_106 ();
 sg13g2_fill_1 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_4 FILLER_68_175 ();
 sg13g2_fill_1 FILLER_68_184 ();
 sg13g2_decap_4 FILLER_68_231 ();
 sg13g2_fill_2 FILLER_68_267 ();
 sg13g2_fill_1 FILLER_68_269 ();
 sg13g2_fill_1 FILLER_68_289 ();
 sg13g2_fill_1 FILLER_68_354 ();
 sg13g2_decap_8 FILLER_68_363 ();
 sg13g2_decap_8 FILLER_68_370 ();
 sg13g2_fill_2 FILLER_68_377 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_45 ();
 sg13g2_fill_1 FILLER_69_70 ();
 sg13g2_fill_2 FILLER_69_75 ();
 sg13g2_decap_4 FILLER_69_159 ();
 sg13g2_fill_2 FILLER_69_163 ();
 sg13g2_fill_2 FILLER_69_191 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_2 FILLER_69_204 ();
 sg13g2_fill_2 FILLER_69_224 ();
 sg13g2_fill_1 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_303 ();
 sg13g2_fill_2 FILLER_69_341 ();
 sg13g2_fill_1 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_370 ();
 sg13g2_fill_2 FILLER_69_377 ();
 sg13g2_fill_1 FILLER_69_379 ();
 sg13g2_fill_1 FILLER_69_394 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_4 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_25 ();
 sg13g2_decap_8 FILLER_70_52 ();
 sg13g2_fill_1 FILLER_70_59 ();
 sg13g2_fill_1 FILLER_70_74 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_decap_8 FILLER_70_132 ();
 sg13g2_fill_1 FILLER_70_139 ();
 sg13g2_decap_8 FILLER_70_144 ();
 sg13g2_decap_8 FILLER_70_151 ();
 sg13g2_fill_2 FILLER_70_158 ();
 sg13g2_fill_2 FILLER_70_182 ();
 sg13g2_fill_1 FILLER_70_184 ();
 sg13g2_decap_4 FILLER_70_211 ();
 sg13g2_fill_1 FILLER_70_215 ();
 sg13g2_fill_1 FILLER_70_234 ();
 sg13g2_fill_1 FILLER_70_250 ();
 sg13g2_decap_4 FILLER_70_264 ();
 sg13g2_fill_2 FILLER_70_307 ();
 sg13g2_decap_4 FILLER_70_317 ();
 sg13g2_fill_1 FILLER_70_321 ();
 sg13g2_fill_2 FILLER_70_345 ();
 sg13g2_fill_1 FILLER_70_347 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_decap_8 FILLER_71_4 ();
 sg13g2_decap_8 FILLER_71_16 ();
 sg13g2_fill_2 FILLER_71_23 ();
 sg13g2_decap_4 FILLER_71_45 ();
 sg13g2_fill_1 FILLER_71_49 ();
 sg13g2_fill_1 FILLER_71_86 ();
 sg13g2_fill_1 FILLER_71_103 ();
 sg13g2_decap_8 FILLER_71_131 ();
 sg13g2_decap_8 FILLER_71_138 ();
 sg13g2_decap_8 FILLER_71_145 ();
 sg13g2_fill_2 FILLER_71_178 ();
 sg13g2_fill_1 FILLER_71_180 ();
 sg13g2_decap_4 FILLER_71_201 ();
 sg13g2_fill_2 FILLER_71_205 ();
 sg13g2_fill_2 FILLER_71_210 ();
 sg13g2_fill_1 FILLER_71_222 ();
 sg13g2_fill_2 FILLER_71_228 ();
 sg13g2_fill_2 FILLER_71_235 ();
 sg13g2_fill_2 FILLER_71_247 ();
 sg13g2_fill_2 FILLER_71_290 ();
 sg13g2_fill_1 FILLER_71_292 ();
 sg13g2_fill_2 FILLER_71_309 ();
 sg13g2_fill_2 FILLER_71_332 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_72_54 ();
 sg13g2_decap_4 FILLER_72_157 ();
 sg13g2_fill_1 FILLER_72_161 ();
 sg13g2_fill_1 FILLER_72_201 ();
 sg13g2_fill_2 FILLER_72_213 ();
 sg13g2_decap_8 FILLER_72_261 ();
 sg13g2_fill_1 FILLER_72_268 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_2 FILLER_72_295 ();
 sg13g2_fill_1 FILLER_72_297 ();
 sg13g2_fill_2 FILLER_72_318 ();
 sg13g2_fill_2 FILLER_72_337 ();
 sg13g2_fill_1 FILLER_72_344 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_fill_2 FILLER_73_77 ();
 sg13g2_fill_1 FILLER_73_79 ();
 sg13g2_fill_1 FILLER_73_112 ();
 sg13g2_fill_2 FILLER_73_193 ();
 sg13g2_fill_1 FILLER_73_195 ();
 sg13g2_fill_2 FILLER_73_227 ();
 sg13g2_fill_1 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_355 ();
 sg13g2_fill_1 FILLER_73_365 ();
 sg13g2_fill_1 FILLER_73_376 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_fill_2 FILLER_74_68 ();
 sg13g2_fill_2 FILLER_74_80 ();
 sg13g2_fill_2 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_93 ();
 sg13g2_fill_1 FILLER_74_103 ();
 sg13g2_fill_2 FILLER_74_135 ();
 sg13g2_fill_2 FILLER_74_207 ();
 sg13g2_decap_8 FILLER_74_234 ();
 sg13g2_decap_4 FILLER_74_241 ();
 sg13g2_fill_1 FILLER_74_245 ();
 sg13g2_fill_2 FILLER_74_272 ();
 sg13g2_fill_1 FILLER_74_283 ();
 sg13g2_fill_2 FILLER_74_366 ();
 sg13g2_decap_8 FILLER_74_375 ();
 sg13g2_decap_4 FILLER_74_382 ();
 sg13g2_fill_1 FILLER_74_386 ();
 sg13g2_decap_4 FILLER_74_390 ();
 sg13g2_fill_1 FILLER_74_394 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_19 ();
 sg13g2_fill_1 FILLER_75_21 ();
 sg13g2_fill_1 FILLER_75_40 ();
 sg13g2_fill_1 FILLER_75_76 ();
 sg13g2_fill_1 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_104 ();
 sg13g2_fill_1 FILLER_75_106 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_137 ();
 sg13g2_decap_4 FILLER_75_144 ();
 sg13g2_fill_2 FILLER_75_148 ();
 sg13g2_decap_4 FILLER_75_158 ();
 sg13g2_fill_2 FILLER_75_197 ();
 sg13g2_fill_1 FILLER_75_199 ();
 sg13g2_fill_2 FILLER_75_205 ();
 sg13g2_decap_8 FILLER_75_222 ();
 sg13g2_decap_8 FILLER_75_229 ();
 sg13g2_decap_8 FILLER_75_236 ();
 sg13g2_fill_2 FILLER_75_243 ();
 sg13g2_fill_1 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_277 ();
 sg13g2_fill_2 FILLER_75_284 ();
 sg13g2_fill_1 FILLER_75_286 ();
 sg13g2_fill_1 FILLER_75_310 ();
 sg13g2_decap_8 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_fill_2 FILLER_75_375 ();
 sg13g2_fill_1 FILLER_75_377 ();
 sg13g2_fill_2 FILLER_75_387 ();
 sg13g2_fill_1 FILLER_75_389 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_fill_2 FILLER_76_26 ();
 sg13g2_fill_1 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_42 ();
 sg13g2_fill_2 FILLER_76_66 ();
 sg13g2_fill_1 FILLER_76_68 ();
 sg13g2_fill_1 FILLER_76_88 ();
 sg13g2_decap_8 FILLER_76_144 ();
 sg13g2_decap_4 FILLER_76_151 ();
 sg13g2_decap_4 FILLER_76_160 ();
 sg13g2_fill_2 FILLER_76_164 ();
 sg13g2_decap_8 FILLER_76_200 ();
 sg13g2_decap_8 FILLER_76_207 ();
 sg13g2_decap_4 FILLER_76_214 ();
 sg13g2_fill_2 FILLER_76_218 ();
 sg13g2_decap_8 FILLER_76_225 ();
 sg13g2_decap_8 FILLER_76_240 ();
 sg13g2_fill_1 FILLER_76_247 ();
 sg13g2_decap_8 FILLER_76_270 ();
 sg13g2_decap_8 FILLER_76_277 ();
 sg13g2_decap_8 FILLER_76_284 ();
 sg13g2_fill_2 FILLER_76_291 ();
 sg13g2_fill_1 FILLER_76_293 ();
 sg13g2_fill_2 FILLER_76_350 ();
 sg13g2_fill_1 FILLER_76_352 ();
 sg13g2_fill_2 FILLER_76_362 ();
 sg13g2_fill_1 FILLER_76_364 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_2 ();
 sg13g2_fill_2 FILLER_77_69 ();
 sg13g2_fill_1 FILLER_77_97 ();
 sg13g2_fill_2 FILLER_77_103 ();
 sg13g2_fill_2 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_173 ();
 sg13g2_fill_2 FILLER_77_214 ();
 sg13g2_fill_2 FILLER_77_247 ();
 sg13g2_fill_1 FILLER_77_249 ();
 sg13g2_fill_2 FILLER_77_276 ();
 sg13g2_fill_1 FILLER_77_283 ();
 sg13g2_fill_2 FILLER_77_336 ();
 sg13g2_fill_1 FILLER_77_338 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_30 ();
 sg13g2_fill_2 FILLER_78_124 ();
 sg13g2_fill_1 FILLER_78_192 ();
 sg13g2_fill_1 FILLER_78_274 ();
 sg13g2_fill_2 FILLER_78_301 ();
 sg13g2_fill_1 FILLER_78_303 ();
 sg13g2_fill_2 FILLER_78_318 ();
 sg13g2_fill_1 FILLER_78_320 ();
 sg13g2_fill_1 FILLER_78_367 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_41 ();
 sg13g2_fill_1 FILLER_79_43 ();
 sg13g2_fill_2 FILLER_79_83 ();
 sg13g2_fill_1 FILLER_79_85 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_fill_2 FILLER_79_133 ();
 sg13g2_fill_1 FILLER_79_135 ();
 sg13g2_fill_2 FILLER_79_149 ();
 sg13g2_fill_1 FILLER_79_156 ();
 sg13g2_fill_1 FILLER_79_191 ();
 sg13g2_decap_4 FILLER_79_252 ();
 sg13g2_fill_1 FILLER_79_256 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_18 ();
 sg13g2_fill_2 FILLER_80_44 ();
 sg13g2_fill_2 FILLER_80_84 ();
 sg13g2_fill_2 FILLER_80_91 ();
 sg13g2_fill_1 FILLER_80_102 ();
 sg13g2_fill_2 FILLER_80_140 ();
 sg13g2_fill_1 FILLER_80_142 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_8 FILLER_80_184 ();
 sg13g2_decap_8 FILLER_80_191 ();
 sg13g2_decap_8 FILLER_80_198 ();
 sg13g2_fill_2 FILLER_80_205 ();
 sg13g2_fill_1 FILLER_80_207 ();
 sg13g2_decap_8 FILLER_80_216 ();
 sg13g2_decap_8 FILLER_80_223 ();
 sg13g2_fill_2 FILLER_80_230 ();
 sg13g2_fill_1 FILLER_80_232 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_8 FILLER_80_249 ();
 sg13g2_decap_8 FILLER_80_256 ();
 sg13g2_decap_4 FILLER_80_263 ();
 sg13g2_fill_1 FILLER_80_267 ();
 sg13g2_fill_2 FILLER_80_310 ();
 sg13g2_fill_2 FILLER_80_325 ();
 sg13g2_fill_1 FILLER_80_327 ();
 sg13g2_fill_1 FILLER_80_333 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_370 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net384;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
endmodule

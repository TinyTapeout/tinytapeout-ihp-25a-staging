module tt_um_stochastic_addmultiply_CL123abc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire SN_Bit_1;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire clknet_leaf_0_clk;
 wire \add_avg[0] ;
 wire \add_avg[1] ;
 wire \add_avg[2] ;
 wire \add_avg[3] ;
 wire \add_avg[4] ;
 wire \add_avg[5] ;
 wire \add_avg[6] ;
 wire \add_avg[7] ;
 wire \add_avg[8] ;
 wire add_bit_out;
 wire \add_output.bitseq[0] ;
 wire \add_output.bitseq[1] ;
 wire \add_output.bitseq[2] ;
 wire \add_output.bitseq[3] ;
 wire \add_output.bitseq[4] ;
 wire \add_output.bitseq[5] ;
 wire \add_output.bitseq[6] ;
 wire \add_output.bitseq[7] ;
 wire \add_output.bitseq[8] ;
 wire \add_output.counter[0] ;
 wire \add_output.counter[1] ;
 wire \add_output.counter[2] ;
 wire \add_output.counter[3] ;
 wire \add_up_counter.clk_counter[0] ;
 wire \add_up_counter.clk_counter[10] ;
 wire \add_up_counter.clk_counter[11] ;
 wire \add_up_counter.clk_counter[12] ;
 wire \add_up_counter.clk_counter[13] ;
 wire \add_up_counter.clk_counter[14] ;
 wire \add_up_counter.clk_counter[15] ;
 wire \add_up_counter.clk_counter[16] ;
 wire \add_up_counter.clk_counter[17] ;
 wire \add_up_counter.clk_counter[1] ;
 wire \add_up_counter.clk_counter[2] ;
 wire \add_up_counter.clk_counter[3] ;
 wire \add_up_counter.clk_counter[4] ;
 wire \add_up_counter.clk_counter[5] ;
 wire \add_up_counter.clk_counter[6] ;
 wire \add_up_counter.clk_counter[7] ;
 wire \add_up_counter.clk_counter[8] ;
 wire \add_up_counter.clk_counter[9] ;
 wire \add_up_counter.prob_counter[0] ;
 wire \add_up_counter.prob_counter[10] ;
 wire \add_up_counter.prob_counter[11] ;
 wire \add_up_counter.prob_counter[12] ;
 wire \add_up_counter.prob_counter[13] ;
 wire \add_up_counter.prob_counter[14] ;
 wire \add_up_counter.prob_counter[15] ;
 wire \add_up_counter.prob_counter[16] ;
 wire \add_up_counter.prob_counter[1] ;
 wire \add_up_counter.prob_counter[2] ;
 wire \add_up_counter.prob_counter[3] ;
 wire \add_up_counter.prob_counter[4] ;
 wire \add_up_counter.prob_counter[5] ;
 wire \add_up_counter.prob_counter[6] ;
 wire \add_up_counter.prob_counter[7] ;
 wire \add_up_counter.prob_counter[8] ;
 wire \add_up_counter.prob_counter[9] ;
 wire \global_SN_gen.Input_1[0] ;
 wire \global_SN_gen.Input_1[1] ;
 wire \global_SN_gen.Input_1[2] ;
 wire \global_SN_gen.Input_1[3] ;
 wire \global_SN_gen.Input_1[4] ;
 wire \global_SN_gen.Input_1[5] ;
 wire \global_SN_gen.Input_1[6] ;
 wire \global_SN_gen.Input_1[7] ;
 wire \global_SN_gen.Input_1[8] ;
 wire \global_SN_gen.Input_2[0] ;
 wire \global_SN_gen.Input_2[1] ;
 wire \global_SN_gen.Input_2[2] ;
 wire \global_SN_gen.Input_2[3] ;
 wire \global_SN_gen.Input_2[4] ;
 wire \global_SN_gen.Input_2[5] ;
 wire \global_SN_gen.Input_2[6] ;
 wire \global_SN_gen.Input_2[7] ;
 wire \global_SN_gen.Input_2[8] ;
 wire \global_SN_gen.lfsr[0] ;
 wire \global_SN_gen.lfsr[10] ;
 wire \global_SN_gen.lfsr[11] ;
 wire \global_SN_gen.lfsr[12] ;
 wire \global_SN_gen.lfsr[13] ;
 wire \global_SN_gen.lfsr[14] ;
 wire \global_SN_gen.lfsr[15] ;
 wire \global_SN_gen.lfsr[16] ;
 wire \global_SN_gen.lfsr[17] ;
 wire \global_SN_gen.lfsr[18] ;
 wire \global_SN_gen.lfsr[19] ;
 wire \global_SN_gen.lfsr[1] ;
 wire \global_SN_gen.lfsr[20] ;
 wire \global_SN_gen.lfsr[21] ;
 wire \global_SN_gen.lfsr[22] ;
 wire \global_SN_gen.lfsr[23] ;
 wire \global_SN_gen.lfsr[24] ;
 wire \global_SN_gen.lfsr[25] ;
 wire \global_SN_gen.lfsr[26] ;
 wire \global_SN_gen.lfsr[27] ;
 wire \global_SN_gen.lfsr[28] ;
 wire \global_SN_gen.lfsr[29] ;
 wire \global_SN_gen.lfsr[2] ;
 wire \global_SN_gen.lfsr[30] ;
 wire \global_SN_gen.lfsr[3] ;
 wire \global_SN_gen.lfsr[4] ;
 wire \global_SN_gen.lfsr[5] ;
 wire \global_SN_gen.lfsr[6] ;
 wire \global_SN_gen.lfsr[7] ;
 wire \global_SN_gen.lfsr[8] ;
 wire \global_SN_gen.lfsr[9] ;
 wire \global_input.adjustment[0] ;
 wire \global_input.adjustment[1] ;
 wire \global_input.adjustment[2] ;
 wire \global_input.adjustment[3] ;
 wire \global_input.adjustment[4] ;
 wire \global_input.loop ;
 wire \global_input.output_bitcounter_1[0] ;
 wire \global_input.output_bitcounter_1[1] ;
 wire \global_input.output_bitcounter_1[2] ;
 wire \global_input.output_bitcounter_1[3] ;
 wire \global_input.output_bitcounter_1[4] ;
 wire \global_input.output_bitcounter_1[5] ;
 wire \global_input.output_bitcounter_1[6] ;
 wire \global_input.output_bitcounter_1[7] ;
 wire \global_input.output_bitcounter_1[8] ;
 wire \global_input.output_bitcounter_2[0] ;
 wire \global_input.output_bitcounter_2[1] ;
 wire \global_input.output_bitcounter_2[2] ;
 wire \global_input.output_bitcounter_2[3] ;
 wire \global_input.output_bitcounter_2[4] ;
 wire \global_input.output_bitcounter_2[5] ;
 wire \global_input.output_bitcounter_2[6] ;
 wire \global_input.output_bitcounter_2[7] ;
 wire \global_input.output_bitcounter_2[8] ;
 wire \global_input.output_case[0] ;
 wire \global_input.output_case[1] ;
 wire \global_input.output_case[2] ;
 wire \global_input.output_case[3] ;
 wire \mul_avg[0] ;
 wire \mul_avg[1] ;
 wire \mul_avg[2] ;
 wire \mul_avg[3] ;
 wire \mul_avg[4] ;
 wire \mul_avg[5] ;
 wire \mul_avg[6] ;
 wire \mul_avg[7] ;
 wire \mul_avg[8] ;
 wire mul_bit_out;
 wire \mul_output.bitseq[0] ;
 wire \mul_output.bitseq[1] ;
 wire \mul_output.bitseq[2] ;
 wire \mul_output.bitseq[3] ;
 wire \mul_output.bitseq[4] ;
 wire \mul_output.bitseq[5] ;
 wire \mul_output.bitseq[6] ;
 wire \mul_output.bitseq[7] ;
 wire \mul_output.bitseq[8] ;
 wire \mul_output.counter[0] ;
 wire \mul_output.counter[1] ;
 wire \mul_output.counter[2] ;
 wire \mul_output.counter[3] ;
 wire \mul_up_counter.prob_counter[0] ;
 wire \mul_up_counter.prob_counter[10] ;
 wire \mul_up_counter.prob_counter[11] ;
 wire \mul_up_counter.prob_counter[12] ;
 wire \mul_up_counter.prob_counter[13] ;
 wire \mul_up_counter.prob_counter[14] ;
 wire \mul_up_counter.prob_counter[15] ;
 wire \mul_up_counter.prob_counter[16] ;
 wire \mul_up_counter.prob_counter[1] ;
 wire \mul_up_counter.prob_counter[2] ;
 wire \mul_up_counter.prob_counter[3] ;
 wire \mul_up_counter.prob_counter[4] ;
 wire \mul_up_counter.prob_counter[5] ;
 wire \mul_up_counter.prob_counter[6] ;
 wire \mul_up_counter.prob_counter[7] ;
 wire \mul_up_counter.prob_counter[8] ;
 wire \mul_up_counter.prob_counter[9] ;
 wire \smul.SN_Bit_Q ;
 wire \smul_avg[0] ;
 wire \smul_avg[1] ;
 wire \smul_avg[2] ;
 wire \smul_avg[3] ;
 wire \smul_avg[4] ;
 wire \smul_avg[5] ;
 wire \smul_avg[6] ;
 wire \smul_avg[7] ;
 wire \smul_avg[8] ;
 wire smul_bit_out;
 wire \smul_output.bitseq[0] ;
 wire \smul_output.bitseq[1] ;
 wire \smul_output.bitseq[2] ;
 wire \smul_output.bitseq[3] ;
 wire \smul_output.bitseq[4] ;
 wire \smul_output.bitseq[5] ;
 wire \smul_output.bitseq[6] ;
 wire \smul_output.bitseq[7] ;
 wire \smul_output.bitseq[8] ;
 wire \smul_output.counter[0] ;
 wire \smul_output.counter[1] ;
 wire \smul_output.counter[2] ;
 wire \smul_output.counter[3] ;
 wire \smul_up_counter.prob_counter[0] ;
 wire \smul_up_counter.prob_counter[10] ;
 wire \smul_up_counter.prob_counter[11] ;
 wire \smul_up_counter.prob_counter[12] ;
 wire \smul_up_counter.prob_counter[13] ;
 wire \smul_up_counter.prob_counter[14] ;
 wire \smul_up_counter.prob_counter[15] ;
 wire \smul_up_counter.prob_counter[16] ;
 wire \smul_up_counter.prob_counter[1] ;
 wire \smul_up_counter.prob_counter[2] ;
 wire \smul_up_counter.prob_counter[3] ;
 wire \smul_up_counter.prob_counter[4] ;
 wire \smul_up_counter.prob_counter[5] ;
 wire \smul_up_counter.prob_counter[6] ;
 wire \smul_up_counter.prob_counter[7] ;
 wire \smul_up_counter.prob_counter[8] ;
 wire \smul_up_counter.prob_counter[9] ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;

 sg13g2_inv_1 _1071_ (.Y(_0414_),
    .A(net115));
 sg13g2_inv_1 _1072_ (.Y(_0588_),
    .A(net135));
 sg13g2_inv_1 _1073_ (.Y(_0589_),
    .A(net390));
 sg13g2_inv_1 _1074_ (.Y(_0590_),
    .A(net413));
 sg13g2_inv_1 _1075_ (.Y(_0591_),
    .A(net398));
 sg13g2_inv_1 _1076_ (.Y(_0592_),
    .A(net412));
 sg13g2_inv_1 _1077_ (.Y(_0593_),
    .A(net393));
 sg13g2_inv_1 _1078_ (.Y(_0594_),
    .A(net414));
 sg13g2_inv_1 _1079_ (.Y(_0595_),
    .A(net404));
 sg13g2_inv_1 _1080_ (.Y(_0596_),
    .A(net397));
 sg13g2_inv_1 _1081_ (.Y(_0597_),
    .A(net80));
 sg13g2_inv_1 _1082_ (.Y(_0401_),
    .A(net124));
 sg13g2_inv_1 _1083_ (.Y(_0598_),
    .A(net216));
 sg13g2_inv_1 _1084_ (.Y(_0599_),
    .A(net358));
 sg13g2_inv_1 _1085_ (.Y(_0600_),
    .A(net377));
 sg13g2_inv_1 _1086_ (.Y(_0601_),
    .A(net370));
 sg13g2_inv_1 _1087_ (.Y(_0602_),
    .A(net366));
 sg13g2_inv_2 _1088_ (.Y(_0603_),
    .A(net356));
 sg13g2_inv_2 _1089_ (.Y(_0604_),
    .A(net374));
 sg13g2_inv_1 _1090_ (.Y(_0605_),
    .A(net379));
 sg13g2_inv_1 _1091_ (.Y(_0606_),
    .A(net364));
 sg13g2_inv_1 _1092_ (.Y(_0607_),
    .A(net406));
 sg13g2_inv_1 _1093_ (.Y(_0608_),
    .A(net180));
 sg13g2_inv_1 _1094_ (.Y(_0609_),
    .A(net360));
 sg13g2_inv_1 _1095_ (.Y(_0610_),
    .A(net229));
 sg13g2_inv_1 _1096_ (.Y(_0611_),
    .A(net244));
 sg13g2_inv_1 _1097_ (.Y(_0612_),
    .A(net264));
 sg13g2_inv_1 _1098_ (.Y(_0613_),
    .A(net355));
 sg13g2_inv_1 _1099_ (.Y(_0614_),
    .A(\global_SN_gen.lfsr[16] ));
 sg13g2_inv_1 _1100_ (.Y(_0225_),
    .A(net30));
 sg13g2_inv_1 _1101_ (.Y(_0223_),
    .A(net29));
 sg13g2_inv_2 _1102_ (.Y(_0221_),
    .A(net49));
 sg13g2_inv_1 _1103_ (.Y(_0615_),
    .A(\global_SN_gen.lfsr[3] ));
 sg13g2_inv_1 _1104_ (.Y(_0212_),
    .A(net41));
 sg13g2_inv_1 _1105_ (.Y(_0616_),
    .A(net309));
 sg13g2_inv_1 _1106_ (.Y(_0617_),
    .A(\global_input.output_case[2] ));
 sg13g2_inv_1 _1107_ (.Y(_0618_),
    .A(net415));
 sg13g2_inv_1 _1108_ (.Y(_0619_),
    .A(net155));
 sg13g2_inv_1 _1109_ (.Y(_0620_),
    .A(\global_SN_gen.Input_2[6] ));
 sg13g2_inv_1 _1110_ (.Y(_0621_),
    .A(\global_SN_gen.Input_2[5] ));
 sg13g2_inv_1 _1111_ (.Y(_0622_),
    .A(\global_SN_gen.Input_2[4] ));
 sg13g2_inv_1 _1112_ (.Y(_0623_),
    .A(net363));
 sg13g2_inv_1 _1113_ (.Y(_0624_),
    .A(net402));
 sg13g2_inv_1 _1114_ (.Y(_0625_),
    .A(net387));
 sg13g2_inv_1 _1115_ (.Y(_0626_),
    .A(net385));
 sg13g2_inv_1 _1116_ (.Y(_0627_),
    .A(net408));
 sg13g2_inv_1 _1117_ (.Y(_0628_),
    .A(net395));
 sg13g2_inv_1 _1118_ (.Y(_0629_),
    .A(net389));
 sg13g2_inv_1 _1119_ (.Y(_0630_),
    .A(net407));
 sg13g2_inv_1 _1120_ (.Y(_0631_),
    .A(\global_input.adjustment[4] ));
 sg13g2_inv_1 _1121_ (.Y(_0632_),
    .A(net250));
 sg13g2_inv_1 _1122_ (.Y(_0633_),
    .A(net87));
 sg13g2_inv_1 _1123_ (.Y(_0289_),
    .A(net152));
 sg13g2_inv_1 _1124_ (.Y(_0634_),
    .A(net105));
 sg13g2_inv_1 _1125_ (.Y(_0635_),
    .A(\global_SN_gen.lfsr[18] ));
 sg13g2_inv_1 _1126_ (.Y(_0636_),
    .A(\global_SN_gen.lfsr[17] ));
 sg13g2_inv_1 _1127_ (.Y(_0637_),
    .A(\global_SN_gen.lfsr[15] ));
 sg13g2_inv_1 _1128_ (.Y(_0638_),
    .A(\global_SN_gen.lfsr[14] ));
 sg13g2_inv_1 _1129_ (.Y(_0639_),
    .A(\add_up_counter.clk_counter[3] ));
 sg13g2_inv_1 _1130_ (.Y(_0640_),
    .A(net203));
 sg13g2_inv_1 _1131_ (.Y(_0641_),
    .A(\add_up_counter.clk_counter[16] ));
 sg13g2_inv_1 _1132_ (.Y(_0642_),
    .A(\smul.SN_Bit_Q ));
 sg13g2_inv_1 _1133_ (.Y(_0060_),
    .A(net319));
 sg13g2_and2_1 _1134_ (.A(net249),
    .B(net115),
    .X(_0643_));
 sg13g2_nand2_1 _1135_ (.Y(_0644_),
    .A(net214),
    .B(_0643_));
 sg13g2_nor2_1 _1136_ (.A(\add_output.counter[2] ),
    .B(\add_output.counter[1] ),
    .Y(_0645_));
 sg13g2_and3_1 _1137_ (.X(_0646_),
    .A(\add_output.counter[3] ),
    .B(\add_output.counter[0] ),
    .C(_0645_));
 sg13g2_nand3_1 _1138_ (.B(\add_output.counter[0] ),
    .C(_0645_),
    .A(\add_output.counter[3] ),
    .Y(_0647_));
 sg13g2_xor2_1 _1139_ (.B(_0644_),
    .A(net369),
    .X(_0648_));
 sg13g2_nor2_1 _1140_ (.A(net299),
    .B(_0648_),
    .Y(_0417_));
 sg13g2_xor2_1 _1141_ (.B(_0643_),
    .A(net214),
    .X(_0416_));
 sg13g2_nor2_1 _1142_ (.A(net249),
    .B(net115),
    .Y(_0649_));
 sg13g2_nor3_1 _1143_ (.A(_0643_),
    .B(net299),
    .C(_0649_),
    .Y(_0415_));
 sg13g2_nor4_2 _1144_ (.A(\add_up_counter.clk_counter[5] ),
    .B(\add_up_counter.clk_counter[4] ),
    .C(\add_up_counter.clk_counter[7] ),
    .Y(_0650_),
    .D(\add_up_counter.clk_counter[6] ));
 sg13g2_nor4_1 _1145_ (.A(\add_up_counter.clk_counter[1] ),
    .B(\add_up_counter.clk_counter[0] ),
    .C(\add_up_counter.clk_counter[3] ),
    .D(\add_up_counter.clk_counter[2] ),
    .Y(_0651_));
 sg13g2_and2_1 _1146_ (.A(_0650_),
    .B(_0651_),
    .X(_0652_));
 sg13g2_nor4_2 _1147_ (.A(\add_up_counter.clk_counter[9] ),
    .B(\add_up_counter.clk_counter[8] ),
    .C(\add_up_counter.clk_counter[11] ),
    .Y(_0653_),
    .D(\add_up_counter.clk_counter[10] ));
 sg13g2_nor4_2 _1148_ (.A(\add_up_counter.clk_counter[13] ),
    .B(\add_up_counter.clk_counter[12] ),
    .C(\add_up_counter.clk_counter[15] ),
    .Y(_0654_),
    .D(\add_up_counter.clk_counter[14] ));
 sg13g2_and4_1 _1149_ (.A(\add_up_counter.clk_counter[17] ),
    .B(_0652_),
    .C(_0653_),
    .D(_0654_),
    .X(_0655_));
 sg13g2_and2_1 _1150_ (.A(_0641_),
    .B(_0655_),
    .X(_0656_));
 sg13g2_nand2_1 _1151_ (.Y(_0657_),
    .A(_0641_),
    .B(_0655_));
 sg13g2_nor2_1 _1152_ (.A(net132),
    .B(net293),
    .Y(_0658_));
 sg13g2_a21oi_1 _1153_ (.A1(_0588_),
    .A2(net293),
    .Y(_0413_),
    .B1(_0658_));
 sg13g2_nand2_1 _1154_ (.Y(_0659_),
    .A(net101),
    .B(net285));
 sg13g2_o21ai_1 _1155_ (.B1(_0659_),
    .Y(_0412_),
    .A1(_0589_),
    .A2(net285));
 sg13g2_nand2_1 _1156_ (.Y(_0660_),
    .A(net145),
    .B(net285));
 sg13g2_o21ai_1 _1157_ (.B1(_0660_),
    .Y(_0411_),
    .A1(_0590_),
    .A2(net285));
 sg13g2_nand2_1 _1158_ (.Y(_0661_),
    .A(net66),
    .B(net284));
 sg13g2_o21ai_1 _1159_ (.B1(_0661_),
    .Y(_0410_),
    .A1(_0591_),
    .A2(net284));
 sg13g2_nand2_1 _1160_ (.Y(_0662_),
    .A(net82),
    .B(net284));
 sg13g2_o21ai_1 _1161_ (.B1(_0662_),
    .Y(_0409_),
    .A1(_0592_),
    .A2(net284));
 sg13g2_nor2_1 _1162_ (.A(net189),
    .B(net293),
    .Y(_0663_));
 sg13g2_a21oi_1 _1163_ (.A1(_0593_),
    .A2(net291),
    .Y(_0408_),
    .B1(_0663_));
 sg13g2_nand2_1 _1164_ (.Y(_0664_),
    .A(net72),
    .B(net284));
 sg13g2_o21ai_1 _1165_ (.B1(_0664_),
    .Y(_0407_),
    .A1(_0594_),
    .A2(net284));
 sg13g2_nand2_1 _1166_ (.Y(_0665_),
    .A(net68),
    .B(net284));
 sg13g2_o21ai_1 _1167_ (.B1(_0665_),
    .Y(_0406_),
    .A1(_0595_),
    .A2(net284));
 sg13g2_nand2_1 _1168_ (.Y(_0666_),
    .A(net80),
    .B(net285));
 sg13g2_o21ai_1 _1169_ (.B1(_0666_),
    .Y(_0405_),
    .A1(_0596_),
    .A2(net285));
 sg13g2_and2_1 _1170_ (.A(net263),
    .B(net124),
    .X(_0667_));
 sg13g2_nand2_1 _1171_ (.Y(_0668_),
    .A(net210),
    .B(_0667_));
 sg13g2_nor2_1 _1172_ (.A(\mul_output.counter[2] ),
    .B(\mul_output.counter[1] ),
    .Y(_0669_));
 sg13g2_and3_1 _1173_ (.X(_0670_),
    .A(net420),
    .B(\mul_output.counter[0] ),
    .C(_0669_));
 sg13g2_nand3_1 _1174_ (.B(\mul_output.counter[0] ),
    .C(_0669_),
    .A(\mul_output.counter[3] ),
    .Y(_0671_));
 sg13g2_xor2_1 _1175_ (.B(_0668_),
    .A(net373),
    .X(_0672_));
 sg13g2_nor2_1 _1176_ (.A(net297),
    .B(_0672_),
    .Y(_0404_));
 sg13g2_xor2_1 _1177_ (.B(_0667_),
    .A(net210),
    .X(_0403_));
 sg13g2_nor2_1 _1178_ (.A(net263),
    .B(net124),
    .Y(_0673_));
 sg13g2_nor3_1 _1179_ (.A(_0667_),
    .B(net297),
    .C(_0673_),
    .Y(_0402_));
 sg13g2_nor2b_1 _1180_ (.A(\global_SN_gen.lfsr[19] ),
    .B_N(\global_SN_gen.Input_1[7] ),
    .Y(_0674_));
 sg13g2_a21o_1 _1181_ (.A2(_0635_),
    .A1(\global_SN_gen.Input_1[6] ),
    .B1(_0674_),
    .X(_0675_));
 sg13g2_nand2b_1 _1182_ (.Y(_0676_),
    .B(\global_SN_gen.lfsr[18] ),
    .A_N(\global_SN_gen.Input_1[6] ));
 sg13g2_nand2b_1 _1183_ (.Y(_0677_),
    .B(\global_SN_gen.lfsr[19] ),
    .A_N(\global_SN_gen.Input_1[7] ));
 sg13g2_nand2b_1 _1184_ (.Y(_0678_),
    .B(\global_SN_gen.lfsr[17] ),
    .A_N(\global_SN_gen.Input_1[5] ));
 sg13g2_nand3_1 _1185_ (.B(_0677_),
    .C(_0678_),
    .A(_0676_),
    .Y(_0679_));
 sg13g2_nor2_1 _1186_ (.A(_0675_),
    .B(_0679_),
    .Y(_0680_));
 sg13g2_nor2_1 _1187_ (.A(_0614_),
    .B(\global_SN_gen.Input_1[4] ),
    .Y(_0681_));
 sg13g2_nand2b_1 _1188_ (.Y(_0682_),
    .B(\global_SN_gen.Input_1[4] ),
    .A_N(\global_SN_gen.lfsr[16] ));
 sg13g2_o21ai_1 _1189_ (.B1(_0682_),
    .Y(_0683_),
    .A1(_0623_),
    .A2(\global_SN_gen.lfsr[17] ));
 sg13g2_nor4_1 _1190_ (.A(_0675_),
    .B(_0679_),
    .C(_0681_),
    .D(_0683_),
    .Y(_0684_));
 sg13g2_nor2b_1 _1191_ (.A(\global_SN_gen.lfsr[15] ),
    .B_N(\global_SN_gen.Input_1[3] ),
    .Y(_0685_));
 sg13g2_nor2b_1 _1192_ (.A(\global_SN_gen.lfsr[14] ),
    .B_N(\global_SN_gen.Input_1[2] ),
    .Y(_0686_));
 sg13g2_nor2b_1 _1193_ (.A(\global_SN_gen.Input_1[2] ),
    .B_N(\global_SN_gen.lfsr[14] ),
    .Y(_0687_));
 sg13g2_nor2b_1 _1194_ (.A(\global_SN_gen.Input_1[3] ),
    .B_N(\global_SN_gen.lfsr[15] ),
    .Y(_0688_));
 sg13g2_nand2b_1 _1195_ (.Y(_0689_),
    .B(\global_SN_gen.lfsr[15] ),
    .A_N(\global_SN_gen.Input_1[3] ));
 sg13g2_or4_1 _1196_ (.A(_0685_),
    .B(_0686_),
    .C(_0687_),
    .D(_0688_),
    .X(_0690_));
 sg13g2_nand2b_1 _1197_ (.Y(_0691_),
    .B(\global_SN_gen.lfsr[12] ),
    .A_N(\global_SN_gen.Input_1[0] ));
 sg13g2_nand2b_1 _1198_ (.Y(_0692_),
    .B(\global_SN_gen.lfsr[13] ),
    .A_N(\global_SN_gen.Input_1[1] ));
 sg13g2_nand2_1 _1199_ (.Y(_0693_),
    .A(_0691_),
    .B(_0692_));
 sg13g2_nor2b_1 _1200_ (.A(\global_SN_gen.lfsr[13] ),
    .B_N(\global_SN_gen.Input_1[1] ),
    .Y(_0694_));
 sg13g2_a21oi_1 _1201_ (.A1(_0691_),
    .A2(_0692_),
    .Y(_0695_),
    .B1(_0694_));
 sg13g2_o21ai_1 _1202_ (.B1(_0689_),
    .Y(_0696_),
    .A1(_0685_),
    .A2(_0686_));
 sg13g2_o21ai_1 _1203_ (.B1(_0696_),
    .Y(_0697_),
    .A1(_0690_),
    .A2(_0695_));
 sg13g2_nor2b_1 _1204_ (.A(\global_SN_gen.lfsr[20] ),
    .B_N(\global_SN_gen.Input_1[8] ),
    .Y(_0698_));
 sg13g2_a21o_1 _1205_ (.A2(_0677_),
    .A1(_0675_),
    .B1(_0698_),
    .X(_0699_));
 sg13g2_a221oi_1 _1206_ (.B2(_0697_),
    .C1(_0699_),
    .B1(_0684_),
    .A1(_0680_),
    .Y(_0700_),
    .A2(_0683_));
 sg13g2_nor2b_1 _1207_ (.A(\global_SN_gen.Input_1[8] ),
    .B_N(\global_SN_gen.lfsr[20] ),
    .Y(_0701_));
 sg13g2_nand2b_1 _1208_ (.Y(_0702_),
    .B(\global_SN_gen.Input_1[0] ),
    .A_N(\global_SN_gen.lfsr[12] ));
 sg13g2_nand2b_1 _1209_ (.Y(_0703_),
    .B(_0702_),
    .A_N(_0694_));
 sg13g2_nor4_1 _1210_ (.A(_0690_),
    .B(_0693_),
    .C(_0698_),
    .D(_0703_),
    .Y(_0704_));
 sg13g2_a21o_1 _1211_ (.A2(_0704_),
    .A1(_0684_),
    .B1(_0701_),
    .X(_0705_));
 sg13g2_o21ai_1 _1212_ (.B1(_0642_),
    .Y(_0706_),
    .A1(_0700_),
    .A2(_0705_));
 sg13g2_or3_1 _1213_ (.A(_0642_),
    .B(_0700_),
    .C(_0705_),
    .X(_0707_));
 sg13g2_nand3_1 _1214_ (.B(_0706_),
    .C(_0707_),
    .A(net287),
    .Y(_0708_));
 sg13g2_a21oi_2 _1215_ (.B1(net292),
    .Y(_0709_),
    .A2(_0707_),
    .A1(_0706_));
 sg13g2_nand2_1 _1216_ (.Y(_0710_),
    .A(net355),
    .B(net248));
 sg13g2_nand3_1 _1217_ (.B(\smul_up_counter.prob_counter[1] ),
    .C(\smul_up_counter.prob_counter[0] ),
    .A(net264),
    .Y(_0711_));
 sg13g2_and4_1 _1218_ (.A(\smul_up_counter.prob_counter[3] ),
    .B(\smul_up_counter.prob_counter[2] ),
    .C(\smul_up_counter.prob_counter[1] ),
    .D(\smul_up_counter.prob_counter[0] ),
    .X(_0712_));
 sg13g2_and2_1 _1219_ (.A(net229),
    .B(_0712_),
    .X(_0713_));
 sg13g2_and4_2 _1220_ (.A(\smul_up_counter.prob_counter[6] ),
    .B(\smul_up_counter.prob_counter[5] ),
    .C(\smul_up_counter.prob_counter[4] ),
    .D(_0712_),
    .X(_0714_));
 sg13g2_nand3_1 _1221_ (.B(\smul_up_counter.prob_counter[7] ),
    .C(_0714_),
    .A(net364),
    .Y(_0715_));
 sg13g2_nor2_1 _1222_ (.A(_0605_),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_nand4_1 _1223_ (.B(\smul_up_counter.prob_counter[8] ),
    .C(\smul_up_counter.prob_counter[7] ),
    .A(net379),
    .Y(_0717_),
    .D(_0714_));
 sg13g2_nand2_1 _1224_ (.Y(_0718_),
    .A(net374),
    .B(_0716_));
 sg13g2_nor4_2 _1225_ (.A(_0602_),
    .B(_0603_),
    .C(_0604_),
    .Y(_0719_),
    .D(_0717_));
 sg13g2_nand2_1 _1226_ (.Y(_0720_),
    .A(net370),
    .B(_0719_));
 sg13g2_nand4_1 _1227_ (.B(\smul_up_counter.prob_counter[14] ),
    .C(\smul_up_counter.prob_counter[13] ),
    .A(net358),
    .Y(_0721_),
    .D(_0719_));
 sg13g2_xor2_1 _1228_ (.B(_0721_),
    .A(_0046_),
    .X(_0722_));
 sg13g2_nand3_1 _1229_ (.B(\smul_up_counter.prob_counter[10] ),
    .C(_0716_),
    .A(net356),
    .Y(_0723_));
 sg13g2_nand2_1 _1230_ (.Y(_0724_),
    .A(net277),
    .B(_0722_));
 sg13g2_o21ai_1 _1231_ (.B1(_0724_),
    .Y(_0400_),
    .A1(_0598_),
    .A2(net279));
 sg13g2_o21ai_1 _1232_ (.B1(_0599_),
    .Y(_0725_),
    .A1(_0600_),
    .A2(_0720_));
 sg13g2_nand3_1 _1233_ (.B(_0721_),
    .C(_0725_),
    .A(net277),
    .Y(_0726_));
 sg13g2_o21ai_1 _1234_ (.B1(_0726_),
    .Y(_0399_),
    .A1(_0599_),
    .A2(net279));
 sg13g2_xnor2_1 _1235_ (.Y(_0727_),
    .A(net377),
    .B(_0720_));
 sg13g2_nand2_1 _1236_ (.Y(_0728_),
    .A(net277),
    .B(_0727_));
 sg13g2_o21ai_1 _1237_ (.B1(_0728_),
    .Y(_0398_),
    .A1(_0600_),
    .A2(net279));
 sg13g2_or2_1 _1238_ (.X(_0729_),
    .B(_0719_),
    .A(net370));
 sg13g2_nand3_1 _1239_ (.B(_0720_),
    .C(_0729_),
    .A(net277),
    .Y(_0730_));
 sg13g2_o21ai_1 _1240_ (.B1(_0730_),
    .Y(_0397_),
    .A1(_0601_),
    .A2(net279));
 sg13g2_nand2_1 _1241_ (.Y(_0731_),
    .A(_0602_),
    .B(_0723_));
 sg13g2_nand3b_1 _1242_ (.B(_0731_),
    .C(net276),
    .Y(_0732_),
    .A_N(_0719_));
 sg13g2_o21ai_1 _1243_ (.B1(_0732_),
    .Y(_0396_),
    .A1(_0602_),
    .A2(_0708_));
 sg13g2_nand2_1 _1244_ (.Y(_0733_),
    .A(_0603_),
    .B(_0718_));
 sg13g2_nand3_1 _1245_ (.B(_0723_),
    .C(_0733_),
    .A(net276),
    .Y(_0734_));
 sg13g2_o21ai_1 _1246_ (.B1(_0734_),
    .Y(_0395_),
    .A1(_0603_),
    .A2(net278));
 sg13g2_nand2_1 _1247_ (.Y(_0735_),
    .A(_0604_),
    .B(_0717_));
 sg13g2_nand3_1 _1248_ (.B(_0718_),
    .C(_0735_),
    .A(_0709_),
    .Y(_0736_));
 sg13g2_o21ai_1 _1249_ (.B1(_0736_),
    .Y(_0394_),
    .A1(_0604_),
    .A2(net278));
 sg13g2_nand2_1 _1250_ (.Y(_0737_),
    .A(_0605_),
    .B(_0715_));
 sg13g2_nand3_1 _1251_ (.B(_0717_),
    .C(_0737_),
    .A(net276),
    .Y(_0738_));
 sg13g2_o21ai_1 _1252_ (.B1(_0738_),
    .Y(_0393_),
    .A1(_0605_),
    .A2(net278));
 sg13g2_a21o_1 _1253_ (.A2(_0714_),
    .A1(\smul_up_counter.prob_counter[7] ),
    .B1(net364),
    .X(_0739_));
 sg13g2_nand3_1 _1254_ (.B(_0715_),
    .C(_0739_),
    .A(net276),
    .Y(_0740_));
 sg13g2_o21ai_1 _1255_ (.B1(_0740_),
    .Y(_0392_),
    .A1(_0606_),
    .A2(net278));
 sg13g2_nor2_1 _1256_ (.A(_0607_),
    .B(net278),
    .Y(_0741_));
 sg13g2_xnor2_1 _1257_ (.Y(_0742_),
    .A(_0607_),
    .B(_0714_));
 sg13g2_a21o_1 _1258_ (.A2(_0742_),
    .A1(net276),
    .B1(_0741_),
    .X(_0391_));
 sg13g2_a21oi_1 _1259_ (.A1(\smul_up_counter.prob_counter[5] ),
    .A2(_0713_),
    .Y(_0743_),
    .B1(net180));
 sg13g2_nor2_1 _1260_ (.A(_0714_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nand2_1 _1261_ (.Y(_0745_),
    .A(net276),
    .B(_0744_));
 sg13g2_o21ai_1 _1262_ (.B1(_0745_),
    .Y(_0390_),
    .A1(_0608_),
    .A2(net278));
 sg13g2_xnor2_1 _1263_ (.Y(_0746_),
    .A(_0609_),
    .B(_0713_));
 sg13g2_nand2_1 _1264_ (.Y(_0747_),
    .A(net276),
    .B(_0746_));
 sg13g2_o21ai_1 _1265_ (.B1(_0747_),
    .Y(_0389_),
    .A1(_0609_),
    .A2(net278));
 sg13g2_or2_1 _1266_ (.X(_0748_),
    .B(_0712_),
    .A(net229));
 sg13g2_nand3b_1 _1267_ (.B(_0748_),
    .C(net276),
    .Y(_0749_),
    .A_N(_0713_));
 sg13g2_o21ai_1 _1268_ (.B1(_0749_),
    .Y(_0388_),
    .A1(_0610_),
    .A2(net278));
 sg13g2_nand2_1 _1269_ (.Y(_0750_),
    .A(_0611_),
    .B(_0711_));
 sg13g2_nand3b_1 _1270_ (.B(_0750_),
    .C(net277),
    .Y(_0751_),
    .A_N(_0712_));
 sg13g2_o21ai_1 _1271_ (.B1(_0751_),
    .Y(_0387_),
    .A1(_0611_),
    .A2(net279));
 sg13g2_nand2_1 _1272_ (.Y(_0752_),
    .A(_0612_),
    .B(_0710_));
 sg13g2_nand3_1 _1273_ (.B(_0711_),
    .C(_0752_),
    .A(net277),
    .Y(_0753_));
 sg13g2_o21ai_1 _1274_ (.B1(_0753_),
    .Y(_0386_),
    .A1(_0612_),
    .A2(net279));
 sg13g2_or2_1 _1275_ (.X(_0754_),
    .B(net248),
    .A(net355));
 sg13g2_nand3_1 _1276_ (.B(_0710_),
    .C(_0754_),
    .A(net277),
    .Y(_0755_));
 sg13g2_o21ai_1 _1277_ (.B1(_0755_),
    .Y(_0385_),
    .A1(_0613_),
    .A2(net279));
 sg13g2_nor2_1 _1278_ (.A(net248),
    .B(net277),
    .Y(_0756_));
 sg13g2_a21oi_1 _1279_ (.A1(net248),
    .A2(net279),
    .Y(_0384_),
    .B1(_0756_));
 sg13g2_xnor2_1 _1280_ (.Y(_0210_),
    .A(net54),
    .B(net43));
 sg13g2_mux2_1 _1281_ (.A0(net1),
    .A1(net191),
    .S(net312),
    .X(_0383_));
 sg13g2_mux2_1 _1282_ (.A0(net191),
    .A1(net186),
    .S(net312),
    .X(_0382_));
 sg13g2_mux2_1 _1283_ (.A0(net186),
    .A1(net111),
    .S(net311),
    .X(_0381_));
 sg13g2_mux2_1 _1284_ (.A0(net111),
    .A1(\global_input.output_bitcounter_1[5] ),
    .S(net311),
    .X(_0380_));
 sg13g2_mux2_1 _1285_ (.A0(net235),
    .A1(net218),
    .S(net311),
    .X(_0379_));
 sg13g2_mux2_1 _1286_ (.A0(net218),
    .A1(net107),
    .S(net309),
    .X(_0378_));
 sg13g2_mux2_1 _1287_ (.A0(net107),
    .A1(net170),
    .S(net309),
    .X(_0377_));
 sg13g2_mux2_1 _1288_ (.A0(net170),
    .A1(net171),
    .S(net309),
    .X(_0376_));
 sg13g2_mux2_1 _1289_ (.A0(net171),
    .A1(\global_input.output_bitcounter_1[0] ),
    .S(net309),
    .X(_0375_));
 sg13g2_nand3_1 _1290_ (.B(net308),
    .C(net293),
    .A(net310),
    .Y(_0757_));
 sg13g2_nand4_1 _1291_ (.B(net415),
    .C(net308),
    .A(net309),
    .Y(_0758_),
    .D(net292));
 sg13g2_nor2_1 _1292_ (.A(_0617_),
    .B(_0758_),
    .Y(_0759_));
 sg13g2_and4_1 _1293_ (.A(\global_input.output_case[3] ),
    .B(_0617_),
    .C(_0618_),
    .D(net308),
    .X(_0760_));
 sg13g2_nand3_1 _1294_ (.B(net292),
    .C(_0760_),
    .A(net309),
    .Y(_0761_));
 sg13g2_xor2_1 _1295_ (.B(_0759_),
    .A(net403),
    .X(_0762_));
 sg13g2_and2_1 _1296_ (.A(_0761_),
    .B(_0762_),
    .X(_0374_));
 sg13g2_xnor2_1 _1297_ (.Y(_0373_),
    .A(net252),
    .B(_0758_));
 sg13g2_nand2_1 _1298_ (.Y(_0763_),
    .A(_0618_),
    .B(_0757_));
 sg13g2_and3_1 _1299_ (.X(_0372_),
    .A(_0758_),
    .B(_0761_),
    .C(_0763_));
 sg13g2_a21o_1 _1300_ (.A2(net292),
    .A1(net309),
    .B1(net308),
    .X(_0764_));
 sg13g2_and2_1 _1301_ (.A(_0757_),
    .B(_0764_),
    .X(_0371_));
 sg13g2_mux2_1 _1302_ (.A0(net2),
    .A1(net158),
    .S(net311),
    .X(_0370_));
 sg13g2_mux2_1 _1303_ (.A0(net158),
    .A1(net188),
    .S(net311),
    .X(_0369_));
 sg13g2_mux2_1 _1304_ (.A0(net188),
    .A1(net175),
    .S(net312),
    .X(_0368_));
 sg13g2_mux2_1 _1305_ (.A0(net175),
    .A1(net173),
    .S(net311),
    .X(_0367_));
 sg13g2_mux2_1 _1306_ (.A0(net173),
    .A1(net167),
    .S(net311),
    .X(_0366_));
 sg13g2_mux2_1 _1307_ (.A0(net167),
    .A1(net138),
    .S(net310),
    .X(_0365_));
 sg13g2_mux2_1 _1308_ (.A0(net138),
    .A1(net169),
    .S(net310),
    .X(_0364_));
 sg13g2_mux2_1 _1309_ (.A0(net169),
    .A1(net162),
    .S(net310),
    .X(_0363_));
 sg13g2_mux2_1 _1310_ (.A0(\global_input.output_bitcounter_2[1] ),
    .A1(net153),
    .S(net310),
    .X(_0362_));
 sg13g2_nand2b_1 _1311_ (.Y(_0765_),
    .B(\add_up_counter.clk_counter[3] ),
    .A_N(\global_input.adjustment[3] ));
 sg13g2_nand2b_1 _1312_ (.Y(_0766_),
    .B(\add_up_counter.clk_counter[0] ),
    .A_N(\global_input.adjustment[0] ));
 sg13g2_nor2b_1 _1313_ (.A(\add_up_counter.clk_counter[0] ),
    .B_N(\global_input.adjustment[0] ),
    .Y(_0767_));
 sg13g2_xor2_1 _1314_ (.B(\add_up_counter.clk_counter[1] ),
    .A(\global_input.adjustment[1] ),
    .X(_0768_));
 sg13g2_o21ai_1 _1315_ (.B1(_0766_),
    .Y(_0769_),
    .A1(_0631_),
    .A2(\add_up_counter.clk_counter[4] ));
 sg13g2_nor4_1 _1316_ (.A(net311),
    .B(_0767_),
    .C(_0768_),
    .D(_0769_),
    .Y(_0770_));
 sg13g2_xnor2_1 _1317_ (.Y(_0771_),
    .A(\global_input.adjustment[2] ),
    .B(\add_up_counter.clk_counter[2] ));
 sg13g2_a22oi_1 _1318_ (.Y(_0772_),
    .B1(\global_input.adjustment[3] ),
    .B2(_0639_),
    .A2(\add_up_counter.clk_counter[4] ),
    .A1(_0631_));
 sg13g2_nand4_1 _1319_ (.B(_0770_),
    .C(_0771_),
    .A(_0765_),
    .Y(_0773_),
    .D(_0772_));
 sg13g2_mux2_1 _1320_ (.A0(net158),
    .A1(\global_SN_gen.Input_2[8] ),
    .S(net281),
    .X(_0361_));
 sg13g2_nor2_1 _1321_ (.A(\global_input.output_bitcounter_2[7] ),
    .B(net282),
    .Y(_0774_));
 sg13g2_a21oi_1 _1322_ (.A1(_0619_),
    .A2(net281),
    .Y(_0360_),
    .B1(_0774_));
 sg13g2_nor2_1 _1323_ (.A(net175),
    .B(net281),
    .Y(_0775_));
 sg13g2_a21oi_1 _1324_ (.A1(_0620_),
    .A2(net281),
    .Y(_0359_),
    .B1(_0775_));
 sg13g2_nor2_1 _1325_ (.A(net173),
    .B(net281),
    .Y(_0776_));
 sg13g2_a21oi_1 _1326_ (.A1(_0621_),
    .A2(net281),
    .Y(_0358_),
    .B1(_0776_));
 sg13g2_nor2_1 _1327_ (.A(net167),
    .B(net281),
    .Y(_0777_));
 sg13g2_a21oi_1 _1328_ (.A1(_0622_),
    .A2(net281),
    .Y(_0357_),
    .B1(_0777_));
 sg13g2_mux2_1 _1329_ (.A0(net138),
    .A1(\global_SN_gen.Input_2[3] ),
    .S(net283),
    .X(_0356_));
 sg13g2_mux2_1 _1330_ (.A0(net169),
    .A1(net179),
    .S(net283),
    .X(_0355_));
 sg13g2_mux2_1 _1331_ (.A0(net162),
    .A1(\global_SN_gen.Input_2[1] ),
    .S(net280),
    .X(_0354_));
 sg13g2_mux2_1 _1332_ (.A0(net153),
    .A1(net184),
    .S(net280),
    .X(_0353_));
 sg13g2_nand2b_1 _1333_ (.Y(_0778_),
    .B(\global_SN_gen.Input_1[6] ),
    .A_N(\global_SN_gen.lfsr[6] ));
 sg13g2_nand2b_1 _1334_ (.Y(_0779_),
    .B(\global_SN_gen.Input_1[7] ),
    .A_N(\global_SN_gen.lfsr[7] ));
 sg13g2_nand2_1 _1335_ (.Y(_0780_),
    .A(_0778_),
    .B(_0779_));
 sg13g2_nor2b_1 _1336_ (.A(\global_SN_gen.Input_1[6] ),
    .B_N(\global_SN_gen.lfsr[6] ),
    .Y(_0781_));
 sg13g2_nor2b_1 _1337_ (.A(\global_SN_gen.Input_1[7] ),
    .B_N(\global_SN_gen.lfsr[7] ),
    .Y(_0782_));
 sg13g2_nor2b_1 _1338_ (.A(\global_SN_gen.Input_1[5] ),
    .B_N(\global_SN_gen.lfsr[5] ),
    .Y(_0783_));
 sg13g2_or3_1 _1339_ (.A(_0781_),
    .B(_0782_),
    .C(_0783_),
    .X(_0784_));
 sg13g2_nor2_1 _1340_ (.A(_0780_),
    .B(_0784_),
    .Y(_0785_));
 sg13g2_nand2b_1 _1341_ (.Y(_0786_),
    .B(\global_SN_gen.Input_1[4] ),
    .A_N(\global_SN_gen.lfsr[4] ));
 sg13g2_o21ai_1 _1342_ (.B1(_0786_),
    .Y(_0787_),
    .A1(\global_SN_gen.lfsr[5] ),
    .A2(_0623_));
 sg13g2_nor2b_1 _1343_ (.A(\global_SN_gen.Input_1[4] ),
    .B_N(\global_SN_gen.lfsr[4] ),
    .Y(_0788_));
 sg13g2_nor4_2 _1344_ (.A(_0780_),
    .B(_0784_),
    .C(_0787_),
    .Y(_0789_),
    .D(_0788_));
 sg13g2_nor2b_1 _1345_ (.A(\global_SN_gen.lfsr[2] ),
    .B_N(\global_SN_gen.Input_1[2] ),
    .Y(_0790_));
 sg13g2_nor2b_1 _1346_ (.A(\global_SN_gen.lfsr[3] ),
    .B_N(\global_SN_gen.Input_1[3] ),
    .Y(_0791_));
 sg13g2_nor2b_1 _1347_ (.A(\global_SN_gen.Input_1[2] ),
    .B_N(\global_SN_gen.lfsr[2] ),
    .Y(_0792_));
 sg13g2_nor2b_1 _1348_ (.A(\global_SN_gen.Input_1[3] ),
    .B_N(\global_SN_gen.lfsr[3] ),
    .Y(_0793_));
 sg13g2_nand2b_1 _1349_ (.Y(_0794_),
    .B(\global_SN_gen.lfsr[3] ),
    .A_N(\global_SN_gen.Input_1[3] ));
 sg13g2_or4_1 _1350_ (.A(_0790_),
    .B(_0791_),
    .C(_0792_),
    .D(_0793_),
    .X(_0795_));
 sg13g2_nor2b_1 _1351_ (.A(\global_SN_gen.lfsr[1] ),
    .B_N(\global_SN_gen.Input_1[1] ),
    .Y(_0796_));
 sg13g2_nand2b_1 _1352_ (.Y(_0797_),
    .B(\global_SN_gen.lfsr[0] ),
    .A_N(\global_SN_gen.Input_1[0] ));
 sg13g2_xnor2_1 _1353_ (.Y(_0798_),
    .A(\global_SN_gen.Input_1[1] ),
    .B(\global_SN_gen.lfsr[1] ));
 sg13g2_a21oi_1 _1354_ (.A1(_0797_),
    .A2(_0798_),
    .Y(_0799_),
    .B1(_0796_));
 sg13g2_o21ai_1 _1355_ (.B1(_0794_),
    .Y(_0800_),
    .A1(_0790_),
    .A2(_0791_));
 sg13g2_o21ai_1 _1356_ (.B1(_0800_),
    .Y(_0801_),
    .A1(_0795_),
    .A2(_0799_));
 sg13g2_a21oi_1 _1357_ (.A1(_0778_),
    .A2(_0779_),
    .Y(_0802_),
    .B1(_0782_));
 sg13g2_a21o_1 _1358_ (.A2(\global_SN_gen.Input_1[8] ),
    .A1(_0221_),
    .B1(_0802_),
    .X(_0803_));
 sg13g2_a221oi_1 _1359_ (.B2(_0801_),
    .C1(_0803_),
    .B1(_0789_),
    .A1(_0785_),
    .Y(_0804_),
    .A2(_0787_));
 sg13g2_a221oi_1 _1360_ (.B2(_0212_),
    .C1(_0795_),
    .B1(\global_SN_gen.Input_1[0] ),
    .A1(_0221_),
    .Y(_0805_),
    .A2(\global_SN_gen.Input_1[8] ));
 sg13g2_and4_1 _1361_ (.A(_0789_),
    .B(_0797_),
    .C(_0798_),
    .D(_0805_),
    .X(_0806_));
 sg13g2_nor2_1 _1362_ (.A(_0221_),
    .B(net409),
    .Y(_0807_));
 sg13g2_nor3_2 _1363_ (.A(_0804_),
    .B(_0806_),
    .C(_0807_),
    .Y(SN_Bit_1));
 sg13g2_nor4_1 _1364_ (.A(_0615_),
    .B(_0804_),
    .C(_0806_),
    .D(_0807_),
    .Y(_0808_));
 sg13g2_nand2b_1 _1365_ (.Y(_0809_),
    .B(\global_SN_gen.Input_2[8] ),
    .A_N(\global_SN_gen.lfsr[20] ));
 sg13g2_nand2b_1 _1366_ (.Y(_0810_),
    .B(\global_SN_gen.lfsr[13] ),
    .A_N(\global_SN_gen.Input_2[1] ));
 sg13g2_nor2b_1 _1367_ (.A(\global_SN_gen.lfsr[12] ),
    .B_N(\global_SN_gen.Input_2[0] ),
    .Y(_0811_));
 sg13g2_nor2b_1 _1368_ (.A(\global_SN_gen.lfsr[13] ),
    .B_N(\global_SN_gen.Input_2[1] ),
    .Y(_0812_));
 sg13g2_a221oi_1 _1369_ (.B2(_0811_),
    .C1(_0812_),
    .B1(_0810_),
    .A1(\global_SN_gen.Input_2[2] ),
    .Y(_0813_),
    .A2(_0638_));
 sg13g2_nand2b_1 _1370_ (.Y(_0814_),
    .B(\global_SN_gen.lfsr[15] ),
    .A_N(\global_SN_gen.Input_2[3] ));
 sg13g2_o21ai_1 _1371_ (.B1(_0814_),
    .Y(_0815_),
    .A1(\global_SN_gen.Input_2[2] ),
    .A2(_0638_));
 sg13g2_a22oi_1 _1372_ (.Y(_0816_),
    .B1(\global_SN_gen.Input_2[3] ),
    .B2(_0637_),
    .A2(\global_SN_gen.Input_2[4] ),
    .A1(_0614_));
 sg13g2_o21ai_1 _1373_ (.B1(_0816_),
    .Y(_0817_),
    .A1(_0813_),
    .A2(_0815_));
 sg13g2_a22oi_1 _1374_ (.Y(_0818_),
    .B1(\global_SN_gen.lfsr[17] ),
    .B2(_0621_),
    .A2(_0622_),
    .A1(\global_SN_gen.lfsr[16] ));
 sg13g2_a22oi_1 _1375_ (.Y(_0819_),
    .B1(\global_SN_gen.lfsr[18] ),
    .B2(_0620_),
    .A2(\global_SN_gen.lfsr[19] ),
    .A1(_0619_));
 sg13g2_nor2b_1 _1376_ (.A(\global_SN_gen.lfsr[19] ),
    .B_N(\global_SN_gen.Input_2[7] ),
    .Y(_0820_));
 sg13g2_a221oi_1 _1377_ (.B2(\global_SN_gen.Input_2[5] ),
    .C1(_0820_),
    .B1(_0636_),
    .A1(\global_SN_gen.Input_2[6] ),
    .Y(_0821_),
    .A2(_0635_));
 sg13g2_nand2_1 _1378_ (.Y(_0822_),
    .A(_0819_),
    .B(_0821_));
 sg13g2_a21oi_1 _1379_ (.A1(_0817_),
    .A2(_0818_),
    .Y(_0823_),
    .B1(_0822_));
 sg13g2_nand2b_1 _1380_ (.Y(_0824_),
    .B(\global_SN_gen.lfsr[20] ),
    .A_N(\global_SN_gen.Input_2[8] ));
 sg13g2_o21ai_1 _1381_ (.B1(_0824_),
    .Y(_0825_),
    .A1(_0819_),
    .A2(_0820_));
 sg13g2_o21ai_1 _1382_ (.B1(_0809_),
    .Y(_0826_),
    .A1(_0823_),
    .A2(_0825_));
 sg13g2_a221oi_1 _1383_ (.B2(_0615_),
    .C1(_0808_),
    .B1(_0826_),
    .A1(_0641_),
    .Y(_0827_),
    .A2(_0655_));
 sg13g2_nand2_1 _1384_ (.Y(_0828_),
    .A(net84),
    .B(net275));
 sg13g2_nand3_1 _1385_ (.B(net419),
    .C(\add_up_counter.prob_counter[0] ),
    .A(net140),
    .Y(_0829_));
 sg13g2_and4_2 _1386_ (.A(net151),
    .B(net140),
    .C(net419),
    .D(\add_up_counter.prob_counter[0] ),
    .X(_0830_));
 sg13g2_nand3_1 _1387_ (.B(\add_up_counter.prob_counter[4] ),
    .C(_0830_),
    .A(net208),
    .Y(_0831_));
 sg13g2_and4_2 _1388_ (.A(net182),
    .B(net208),
    .C(net418),
    .D(_0830_),
    .X(_0832_));
 sg13g2_nand3_1 _1389_ (.B(net247),
    .C(_0832_),
    .A(net136),
    .Y(_0833_));
 sg13g2_and4_2 _1390_ (.A(net193),
    .B(\add_up_counter.prob_counter[8] ),
    .C(net247),
    .D(_0832_),
    .X(_0834_));
 sg13g2_and4_1 _1391_ (.A(\add_up_counter.prob_counter[12] ),
    .B(\add_up_counter.prob_counter[11] ),
    .C(\add_up_counter.prob_counter[10] ),
    .D(_0834_),
    .X(_0835_));
 sg13g2_and2_1 _1392_ (.A(\add_up_counter.prob_counter[13] ),
    .B(_0835_),
    .X(_0836_));
 sg13g2_and3_1 _1393_ (.X(_0837_),
    .A(net221),
    .B(\add_up_counter.prob_counter[14] ),
    .C(_0836_));
 sg13g2_or2_1 _1394_ (.X(_0838_),
    .B(net275),
    .A(net291));
 sg13g2_and3_1 _1395_ (.X(_0839_),
    .A(net197),
    .B(net417),
    .C(_0834_));
 sg13g2_xor2_1 _1396_ (.B(_0837_),
    .A(_0048_),
    .X(_0840_));
 sg13g2_o21ai_1 _1397_ (.B1(_0828_),
    .Y(_0352_),
    .A1(net268),
    .A2(_0840_));
 sg13g2_a21oi_1 _1398_ (.A1(net219),
    .A2(_0836_),
    .Y(_0841_),
    .B1(net201));
 sg13g2_nor4_1 _1399_ (.A(net291),
    .B(net275),
    .C(_0837_),
    .D(_0841_),
    .Y(_0842_));
 sg13g2_a21o_1 _1400_ (.A2(net275),
    .A1(net201),
    .B1(_0842_),
    .X(_0351_));
 sg13g2_nand2_1 _1401_ (.Y(_0843_),
    .A(net219),
    .B(net275));
 sg13g2_xnor2_1 _1402_ (.Y(_0844_),
    .A(net219),
    .B(_0836_));
 sg13g2_o21ai_1 _1403_ (.B1(_0843_),
    .Y(_0350_),
    .A1(net268),
    .A2(_0844_));
 sg13g2_nand2_1 _1404_ (.Y(_0845_),
    .A(net224),
    .B(net275));
 sg13g2_xnor2_1 _1405_ (.Y(_0846_),
    .A(net224),
    .B(_0835_));
 sg13g2_o21ai_1 _1406_ (.B1(_0845_),
    .Y(_0349_),
    .A1(_0838_),
    .A2(_0846_));
 sg13g2_nand2_1 _1407_ (.Y(_0847_),
    .A(net240),
    .B(net274));
 sg13g2_xnor2_1 _1408_ (.Y(_0848_),
    .A(net240),
    .B(_0839_));
 sg13g2_o21ai_1 _1409_ (.B1(_0847_),
    .Y(_0348_),
    .A1(net267),
    .A2(_0848_));
 sg13g2_nand2_1 _1410_ (.Y(_0849_),
    .A(net197),
    .B(net274));
 sg13g2_a21oi_1 _1411_ (.A1(\add_up_counter.prob_counter[10] ),
    .A2(_0834_),
    .Y(_0850_),
    .B1(net197));
 sg13g2_or2_1 _1412_ (.X(_0851_),
    .B(_0850_),
    .A(_0839_));
 sg13g2_o21ai_1 _1413_ (.B1(_0849_),
    .Y(_0347_),
    .A1(net267),
    .A2(_0851_));
 sg13g2_nand2_1 _1414_ (.Y(_0852_),
    .A(net256),
    .B(net274));
 sg13g2_xnor2_1 _1415_ (.Y(_0853_),
    .A(net256),
    .B(_0834_));
 sg13g2_o21ai_1 _1416_ (.B1(_0852_),
    .Y(_0346_),
    .A1(net267),
    .A2(_0853_));
 sg13g2_nand2_1 _1417_ (.Y(_0854_),
    .A(net193),
    .B(net274));
 sg13g2_xor2_1 _1418_ (.B(_0833_),
    .A(net193),
    .X(_0855_));
 sg13g2_o21ai_1 _1419_ (.B1(_0854_),
    .Y(_0345_),
    .A1(net268),
    .A2(_0855_));
 sg13g2_nand2_1 _1420_ (.Y(_0856_),
    .A(net136),
    .B(net273));
 sg13g2_a21o_1 _1421_ (.A2(_0832_),
    .A1(net239),
    .B1(net136),
    .X(_0857_));
 sg13g2_nand2_1 _1422_ (.Y(_0858_),
    .A(_0833_),
    .B(_0857_));
 sg13g2_o21ai_1 _1423_ (.B1(_0856_),
    .Y(_0344_),
    .A1(net268),
    .A2(_0858_));
 sg13g2_nand2_1 _1424_ (.Y(_0859_),
    .A(net239),
    .B(net274));
 sg13g2_xnor2_1 _1425_ (.Y(_0860_),
    .A(net239),
    .B(_0832_));
 sg13g2_o21ai_1 _1426_ (.B1(_0859_),
    .Y(_0343_),
    .A1(net268),
    .A2(_0860_));
 sg13g2_nand2_1 _1427_ (.Y(_0861_),
    .A(net182),
    .B(net273));
 sg13g2_xor2_1 _1428_ (.B(_0831_),
    .A(net182),
    .X(_0862_));
 sg13g2_o21ai_1 _1429_ (.B1(_0861_),
    .Y(_0342_),
    .A1(net267),
    .A2(_0862_));
 sg13g2_nand2_1 _1430_ (.Y(_0863_),
    .A(net208),
    .B(net273));
 sg13g2_a21o_1 _1431_ (.A2(_0830_),
    .A1(\add_up_counter.prob_counter[4] ),
    .B1(net208),
    .X(_0864_));
 sg13g2_nand2_1 _1432_ (.Y(_0865_),
    .A(_0831_),
    .B(_0864_));
 sg13g2_o21ai_1 _1433_ (.B1(_0863_),
    .Y(_0341_),
    .A1(net267),
    .A2(_0865_));
 sg13g2_nand2_1 _1434_ (.Y(_0866_),
    .A(net243),
    .B(net273));
 sg13g2_xnor2_1 _1435_ (.Y(_0867_),
    .A(net243),
    .B(_0830_));
 sg13g2_o21ai_1 _1436_ (.B1(_0866_),
    .Y(_0340_),
    .A1(net267),
    .A2(_0867_));
 sg13g2_nand2_1 _1437_ (.Y(_0418_),
    .A(net151),
    .B(net273));
 sg13g2_xor2_1 _1438_ (.B(_0829_),
    .A(net151),
    .X(_0419_));
 sg13g2_o21ai_1 _1439_ (.B1(_0418_),
    .Y(_0339_),
    .A1(net268),
    .A2(_0419_));
 sg13g2_nand2_1 _1440_ (.Y(_0420_),
    .A(net140),
    .B(net273));
 sg13g2_a21o_1 _1441_ (.A2(\add_up_counter.prob_counter[0] ),
    .A1(\add_up_counter.prob_counter[1] ),
    .B1(net140),
    .X(_0421_));
 sg13g2_nand2_1 _1442_ (.Y(_0422_),
    .A(_0829_),
    .B(_0421_));
 sg13g2_o21ai_1 _1443_ (.B1(_0420_),
    .Y(_0338_),
    .A1(net268),
    .A2(_0422_));
 sg13g2_nand2_1 _1444_ (.Y(_0423_),
    .A(net261),
    .B(net273));
 sg13g2_xnor2_1 _1445_ (.Y(_0424_),
    .A(net261),
    .B(\add_up_counter.prob_counter[0] ));
 sg13g2_o21ai_1 _1446_ (.B1(_0423_),
    .Y(_0337_),
    .A1(net267),
    .A2(_0424_));
 sg13g2_nand2_1 _1447_ (.Y(_0425_),
    .A(net371),
    .B(net273));
 sg13g2_o21ai_1 _1448_ (.B1(_0425_),
    .Y(_0336_),
    .A1(net371),
    .A2(net267));
 sg13g2_mux2_1 _1449_ (.A0(net191),
    .A1(\global_SN_gen.Input_1[8] ),
    .S(net282),
    .X(_0335_));
 sg13g2_mux2_1 _1450_ (.A0(net186),
    .A1(\global_SN_gen.Input_1[7] ),
    .S(net282),
    .X(_0334_));
 sg13g2_mux2_1 _1451_ (.A0(net111),
    .A1(net205),
    .S(net282),
    .X(_0333_));
 sg13g2_nor2_1 _1452_ (.A(net235),
    .B(net282),
    .Y(_0426_));
 sg13g2_a21oi_1 _1453_ (.A1(_0623_),
    .A2(net282),
    .Y(_0332_),
    .B1(_0426_));
 sg13g2_mux2_1 _1454_ (.A0(net218),
    .A1(net260),
    .S(net280),
    .X(_0331_));
 sg13g2_mux2_1 _1455_ (.A0(net107),
    .A1(\global_SN_gen.Input_1[3] ),
    .S(net280),
    .X(_0330_));
 sg13g2_mux2_1 _1456_ (.A0(net170),
    .A1(net178),
    .S(net280),
    .X(_0329_));
 sg13g2_mux2_1 _1457_ (.A0(net171),
    .A1(net185),
    .S(net280),
    .X(_0328_));
 sg13g2_mux2_1 _1458_ (.A0(net212),
    .A1(\global_SN_gen.Input_1[0] ),
    .S(net280),
    .X(_0327_));
 sg13g2_nor2_1 _1459_ (.A(net381),
    .B(net152),
    .Y(_0427_));
 sg13g2_nor2_1 _1460_ (.A(\smul_output.counter[2] ),
    .B(\smul_output.counter[1] ),
    .Y(_0428_));
 sg13g2_nor4_2 _1461_ (.A(net142),
    .B(\smul_output.counter[2] ),
    .C(\smul_output.counter[1] ),
    .Y(_0429_),
    .D(net152));
 sg13g2_and3_2 _1462_ (.X(_0430_),
    .A(\smul_output.counter[3] ),
    .B(\smul_output.counter[0] ),
    .C(_0428_));
 sg13g2_nand3_1 _1463_ (.B(\smul_output.counter[0] ),
    .C(_0428_),
    .A(\smul_output.counter[3] ),
    .Y(_0431_));
 sg13g2_o21ai_1 _1464_ (.B1(net294),
    .Y(_0432_),
    .A1(net104),
    .A2(net307));
 sg13g2_a21oi_1 _1465_ (.A1(_0633_),
    .A2(net307),
    .Y(_0326_),
    .B1(_0432_));
 sg13g2_nand2_1 _1466_ (.Y(_0433_),
    .A(SN_Bit_1),
    .B(_0826_));
 sg13g2_nor2_1 _1467_ (.A(SN_Bit_1),
    .B(_0826_),
    .Y(_0434_));
 sg13g2_or2_1 _1468_ (.X(_0435_),
    .B(_0826_),
    .A(SN_Bit_1));
 sg13g2_a21o_1 _1469_ (.A2(_0826_),
    .A1(SN_Bit_1),
    .B1(net291),
    .X(_0436_));
 sg13g2_nor2_1 _1470_ (.A(net271),
    .B(net269),
    .Y(_0437_));
 sg13g2_nor3_1 _1471_ (.A(_0588_),
    .B(net272),
    .C(net270),
    .Y(_0438_));
 sg13g2_nor2_1 _1472_ (.A(_0589_),
    .B(_0590_),
    .Y(_0439_));
 sg13g2_nand3_1 _1473_ (.B(\mul_up_counter.prob_counter[1] ),
    .C(\mul_up_counter.prob_counter[0] ),
    .A(net389),
    .Y(_0440_));
 sg13g2_and4_2 _1474_ (.A(\mul_up_counter.prob_counter[3] ),
    .B(\mul_up_counter.prob_counter[2] ),
    .C(\mul_up_counter.prob_counter[1] ),
    .D(\mul_up_counter.prob_counter[0] ),
    .X(_0441_));
 sg13g2_nand3_1 _1475_ (.B(\mul_up_counter.prob_counter[4] ),
    .C(_0441_),
    .A(net385),
    .Y(_0442_));
 sg13g2_and4_2 _1476_ (.A(\mul_up_counter.prob_counter[6] ),
    .B(\mul_up_counter.prob_counter[5] ),
    .C(\mul_up_counter.prob_counter[4] ),
    .D(_0441_),
    .X(_0443_));
 sg13g2_nand3_1 _1477_ (.B(\mul_up_counter.prob_counter[7] ),
    .C(_0443_),
    .A(\mul_up_counter.prob_counter[8] ),
    .Y(_0444_));
 sg13g2_nor2_1 _1478_ (.A(_0595_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_a21oi_1 _1479_ (.A1(_0433_),
    .A2(_0435_),
    .Y(_0446_),
    .B1(net291));
 sg13g2_nor4_2 _1480_ (.A(_0593_),
    .B(_0594_),
    .C(_0595_),
    .Y(_0447_),
    .D(_0444_));
 sg13g2_and3_2 _1481_ (.X(_0448_),
    .A(\mul_up_counter.prob_counter[13] ),
    .B(\mul_up_counter.prob_counter[12] ),
    .C(_0447_));
 sg13g2_nand2_1 _1482_ (.Y(_0449_),
    .A(_0439_),
    .B(_0448_));
 sg13g2_xor2_1 _1483_ (.B(_0449_),
    .A(net368),
    .X(_0450_));
 sg13g2_a21o_1 _1484_ (.A2(_0450_),
    .A1(net266),
    .B1(_0438_),
    .X(_0325_));
 sg13g2_nor3_1 _1485_ (.A(_0589_),
    .B(net272),
    .C(net270),
    .Y(_0451_));
 sg13g2_a21o_1 _1486_ (.A2(_0448_),
    .A1(\mul_up_counter.prob_counter[14] ),
    .B1(net390),
    .X(_0452_));
 sg13g2_a221oi_1 _1487_ (.B2(_0448_),
    .C1(net291),
    .B1(_0439_),
    .A1(_0433_),
    .Y(_0453_),
    .A2(_0435_));
 sg13g2_a21o_1 _1488_ (.A2(_0453_),
    .A1(net391),
    .B1(_0451_),
    .X(_0324_));
 sg13g2_nor3_1 _1489_ (.A(_0590_),
    .B(_0434_),
    .C(_0436_),
    .Y(_0454_));
 sg13g2_xnor2_1 _1490_ (.Y(_0455_),
    .A(_0590_),
    .B(_0448_));
 sg13g2_a21o_1 _1491_ (.A2(_0455_),
    .A1(net266),
    .B1(_0454_),
    .X(_0323_));
 sg13g2_nor3_1 _1492_ (.A(_0591_),
    .B(net272),
    .C(net270),
    .Y(_0456_));
 sg13g2_a21oi_1 _1493_ (.A1(\mul_up_counter.prob_counter[12] ),
    .A2(_0447_),
    .Y(_0457_),
    .B1(net398));
 sg13g2_nor2_1 _1494_ (.A(_0448_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_a21o_1 _1495_ (.A2(_0458_),
    .A1(net266),
    .B1(_0456_),
    .X(_0322_));
 sg13g2_nor3_1 _1496_ (.A(_0592_),
    .B(net271),
    .C(net269),
    .Y(_0459_));
 sg13g2_xnor2_1 _1497_ (.Y(_0460_),
    .A(_0592_),
    .B(_0447_));
 sg13g2_a21o_1 _1498_ (.A2(_0460_),
    .A1(net265),
    .B1(_0459_),
    .X(_0321_));
 sg13g2_nor3_1 _1499_ (.A(_0593_),
    .B(net272),
    .C(net270),
    .Y(_0461_));
 sg13g2_a21oi_1 _1500_ (.A1(\mul_up_counter.prob_counter[10] ),
    .A2(_0445_),
    .Y(_0462_),
    .B1(net393));
 sg13g2_nor2_1 _1501_ (.A(_0447_),
    .B(net394),
    .Y(_0463_));
 sg13g2_a21o_1 _1502_ (.A2(_0463_),
    .A1(net266),
    .B1(_0461_),
    .X(_0320_));
 sg13g2_nor3_1 _1503_ (.A(_0594_),
    .B(net272),
    .C(net270),
    .Y(_0464_));
 sg13g2_xnor2_1 _1504_ (.Y(_0465_),
    .A(_0594_),
    .B(_0445_));
 sg13g2_a21o_1 _1505_ (.A2(_0465_),
    .A1(net266),
    .B1(_0464_),
    .X(_0319_));
 sg13g2_nor3_1 _1506_ (.A(_0595_),
    .B(net272),
    .C(net270),
    .Y(_0466_));
 sg13g2_xnor2_1 _1507_ (.Y(_0467_),
    .A(net404),
    .B(_0444_));
 sg13g2_a21o_1 _1508_ (.A2(_0467_),
    .A1(net266),
    .B1(_0466_),
    .X(_0318_));
 sg13g2_nor3_1 _1509_ (.A(_0596_),
    .B(_0434_),
    .C(_0436_),
    .Y(_0468_));
 sg13g2_a21o_1 _1510_ (.A2(_0443_),
    .A1(\mul_up_counter.prob_counter[7] ),
    .B1(\mul_up_counter.prob_counter[8] ),
    .X(_0469_));
 sg13g2_and2_1 _1511_ (.A(_0444_),
    .B(_0469_),
    .X(_0470_));
 sg13g2_a21o_1 _1512_ (.A2(_0470_),
    .A1(net266),
    .B1(_0468_),
    .X(_0317_));
 sg13g2_nor3_1 _1513_ (.A(_0624_),
    .B(net272),
    .C(net270),
    .Y(_0471_));
 sg13g2_xnor2_1 _1514_ (.Y(_0472_),
    .A(_0624_),
    .B(_0443_));
 sg13g2_a21o_1 _1515_ (.A2(_0472_),
    .A1(_0446_),
    .B1(_0471_),
    .X(_0316_));
 sg13g2_nor3_1 _1516_ (.A(_0625_),
    .B(net271),
    .C(net269),
    .Y(_0473_));
 sg13g2_xnor2_1 _1517_ (.Y(_0474_),
    .A(net387),
    .B(_0442_));
 sg13g2_a21o_1 _1518_ (.A2(_0474_),
    .A1(net265),
    .B1(_0473_),
    .X(_0315_));
 sg13g2_nor3_1 _1519_ (.A(_0626_),
    .B(net271),
    .C(net269),
    .Y(_0475_));
 sg13g2_a21o_1 _1520_ (.A2(_0441_),
    .A1(\mul_up_counter.prob_counter[4] ),
    .B1(\mul_up_counter.prob_counter[5] ),
    .X(_0476_));
 sg13g2_and2_1 _1521_ (.A(_0442_),
    .B(_0476_),
    .X(_0477_));
 sg13g2_a21o_1 _1522_ (.A2(_0477_),
    .A1(net265),
    .B1(_0475_),
    .X(_0314_));
 sg13g2_nor3_1 _1523_ (.A(_0627_),
    .B(net271),
    .C(net269),
    .Y(_0478_));
 sg13g2_xnor2_1 _1524_ (.Y(_0479_),
    .A(_0627_),
    .B(_0441_));
 sg13g2_a21o_1 _1525_ (.A2(_0479_),
    .A1(net265),
    .B1(_0478_),
    .X(_0313_));
 sg13g2_nor3_1 _1526_ (.A(_0628_),
    .B(net271),
    .C(net269),
    .Y(_0480_));
 sg13g2_xnor2_1 _1527_ (.Y(_0481_),
    .A(net395),
    .B(_0440_));
 sg13g2_a21o_1 _1528_ (.A2(_0481_),
    .A1(net265),
    .B1(_0480_),
    .X(_0312_));
 sg13g2_nor3_1 _1529_ (.A(_0629_),
    .B(net271),
    .C(net269),
    .Y(_0482_));
 sg13g2_a21o_1 _1530_ (.A2(\mul_up_counter.prob_counter[0] ),
    .A1(\mul_up_counter.prob_counter[1] ),
    .B1(\mul_up_counter.prob_counter[2] ),
    .X(_0483_));
 sg13g2_and2_1 _1531_ (.A(_0440_),
    .B(_0483_),
    .X(_0484_));
 sg13g2_a21o_1 _1532_ (.A2(_0484_),
    .A1(net265),
    .B1(_0482_),
    .X(_0311_));
 sg13g2_nor3_1 _1533_ (.A(_0630_),
    .B(net271),
    .C(net269),
    .Y(_0485_));
 sg13g2_xor2_1 _1534_ (.B(net382),
    .A(net407),
    .X(_0486_));
 sg13g2_a21o_1 _1535_ (.A2(_0486_),
    .A1(net265),
    .B1(_0485_),
    .X(_0310_));
 sg13g2_mux2_1 _1536_ (.A0(net265),
    .A1(_0437_),
    .S(net382),
    .X(_0309_));
 sg13g2_nor4_1 _1537_ (.A(\add_output.counter[3] ),
    .B(\add_output.counter[2] ),
    .C(\add_output.counter[1] ),
    .D(\add_output.counter[0] ),
    .Y(_0487_));
 sg13g2_o21ai_1 _1538_ (.B1(net298),
    .Y(_0488_),
    .A1(\add_output.bitseq[0] ),
    .A2(net305));
 sg13g2_a21oi_1 _1539_ (.A1(_0634_),
    .A2(net305),
    .Y(_0308_),
    .B1(_0488_));
 sg13g2_nor4_1 _1540_ (.A(\mul_output.counter[3] ),
    .B(\mul_output.counter[2] ),
    .C(\mul_output.counter[1] ),
    .D(\mul_output.counter[0] ),
    .Y(_0489_));
 sg13g2_o21ai_1 _1541_ (.B1(net296),
    .Y(_0490_),
    .A1(net103),
    .A2(net301));
 sg13g2_a21oi_1 _1542_ (.A1(_0597_),
    .A2(net301),
    .Y(_0307_),
    .B1(_0490_));
 sg13g2_o21ai_1 _1543_ (.B1(\global_input.output_case[3] ),
    .Y(_0491_),
    .A1(\global_input.output_case[2] ),
    .A2(\global_input.output_case[1] ));
 sg13g2_nand2_1 _1544_ (.Y(_0492_),
    .A(_0616_),
    .B(_0491_));
 sg13g2_nor3_1 _1545_ (.A(\add_up_counter.clk_counter[16] ),
    .B(\add_up_counter.clk_counter[17] ),
    .C(_0492_),
    .Y(_0493_));
 sg13g2_nand4_1 _1546_ (.B(_0653_),
    .C(_0654_),
    .A(_0652_),
    .Y(_0494_),
    .D(_0493_));
 sg13g2_nor2_1 _1547_ (.A(\global_input.output_case[3] ),
    .B(_0617_),
    .Y(_0495_));
 sg13g2_nand3_1 _1548_ (.B(net308),
    .C(_0495_),
    .A(_0618_),
    .Y(_0496_));
 sg13g2_or2_1 _1549_ (.X(_0497_),
    .B(\global_input.output_case[2] ),
    .A(\global_input.output_case[3] ));
 sg13g2_nor2_1 _1550_ (.A(_0618_),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_nand2_1 _1551_ (.Y(_0499_),
    .A(\global_input.output_case[0] ),
    .B(_0498_));
 sg13g2_nand2_1 _1552_ (.Y(_0500_),
    .A(_0496_),
    .B(_0499_));
 sg13g2_nand2_1 _1553_ (.Y(_0501_),
    .A(\global_input.output_case[1] ),
    .B(_0495_));
 sg13g2_a21oi_1 _1554_ (.A1(_0497_),
    .A2(_0501_),
    .Y(_0502_),
    .B1(net308));
 sg13g2_nor2b_1 _1555_ (.A(_0500_),
    .B_N(_0501_),
    .Y(_0503_));
 sg13g2_nor4_2 _1556_ (.A(_0760_),
    .B(_0494_),
    .C(_0500_),
    .Y(_0504_),
    .D(_0502_));
 sg13g2_a21o_1 _1557_ (.A2(_0494_),
    .A1(net160),
    .B1(_0504_),
    .X(_0306_));
 sg13g2_a21o_1 _1558_ (.A2(_0494_),
    .A1(net133),
    .B1(_0504_),
    .X(_0305_));
 sg13g2_nor3_1 _1559_ (.A(_0618_),
    .B(net308),
    .C(_0497_),
    .Y(_0505_));
 sg13g2_nor3_1 _1560_ (.A(_0760_),
    .B(_0494_),
    .C(_0505_),
    .Y(_0506_));
 sg13g2_a22oi_1 _1561_ (.Y(_0304_),
    .B1(_0496_),
    .B2(_0506_),
    .A2(_0494_),
    .A1(_0632_));
 sg13g2_nand2_1 _1562_ (.Y(_0507_),
    .A(net117),
    .B(_0494_));
 sg13g2_o21ai_1 _1563_ (.B1(_0507_),
    .Y(_0303_),
    .A1(_0494_),
    .A2(_0503_));
 sg13g2_mux2_1 _1564_ (.A0(net308),
    .A1(net149),
    .S(_0494_),
    .X(_0302_));
 sg13g2_nand2_1 _1565_ (.Y(_0508_),
    .A(net70),
    .B(net288));
 sg13g2_o21ai_1 _1566_ (.B1(_0508_),
    .Y(_0301_),
    .A1(_0598_),
    .A2(net287));
 sg13g2_nand2_1 _1567_ (.Y(_0509_),
    .A(net76),
    .B(net287));
 sg13g2_o21ai_1 _1568_ (.B1(_0509_),
    .Y(_0300_),
    .A1(_0599_),
    .A2(net287));
 sg13g2_nand2_1 _1569_ (.Y(_0510_),
    .A(net64),
    .B(net287));
 sg13g2_o21ai_1 _1570_ (.B1(_0510_),
    .Y(_0299_),
    .A1(_0600_),
    .A2(net287));
 sg13g2_nand2_1 _1571_ (.Y(_0511_),
    .A(net78),
    .B(net287));
 sg13g2_o21ai_1 _1572_ (.B1(_0511_),
    .Y(_0298_),
    .A1(_0601_),
    .A2(net287));
 sg13g2_nand2_1 _1573_ (.Y(_0512_),
    .A(net74),
    .B(net289));
 sg13g2_o21ai_1 _1574_ (.B1(_0512_),
    .Y(_0297_),
    .A1(_0602_),
    .A2(net289));
 sg13g2_nor2_1 _1575_ (.A(net122),
    .B(net292),
    .Y(_0513_));
 sg13g2_a21oi_1 _1576_ (.A1(_0603_),
    .A2(net292),
    .Y(_0296_),
    .B1(_0513_));
 sg13g2_nand2_1 _1577_ (.Y(_0514_),
    .A(net62),
    .B(net288));
 sg13g2_o21ai_1 _1578_ (.B1(_0514_),
    .Y(_0295_),
    .A1(_0604_),
    .A2(net288));
 sg13g2_nand2_1 _1579_ (.Y(_0515_),
    .A(net60),
    .B(net288));
 sg13g2_o21ai_1 _1580_ (.B1(_0515_),
    .Y(_0294_),
    .A1(_0605_),
    .A2(net288));
 sg13g2_nand2_1 _1581_ (.Y(_0516_),
    .A(net87),
    .B(net288));
 sg13g2_o21ai_1 _1582_ (.B1(_0516_),
    .Y(_0293_),
    .A1(_0606_),
    .A2(net288));
 sg13g2_and2_1 _1583_ (.A(net381),
    .B(net152),
    .X(_0517_));
 sg13g2_and2_1 _1584_ (.A(net254),
    .B(_0517_),
    .X(_0518_));
 sg13g2_a21oi_1 _1585_ (.A1(net142),
    .A2(_0518_),
    .Y(_0519_),
    .B1(net295));
 sg13g2_o21ai_1 _1586_ (.B1(_0519_),
    .Y(_0520_),
    .A1(net142),
    .A2(_0518_));
 sg13g2_inv_1 _1587_ (.Y(_0292_),
    .A(_0520_));
 sg13g2_xor2_1 _1588_ (.B(_0517_),
    .A(net254),
    .X(_0291_));
 sg13g2_nor3_1 _1589_ (.A(_0427_),
    .B(net143),
    .C(_0517_),
    .Y(_0290_));
 sg13g2_mux2_1 _1590_ (.A0(net84),
    .A1(net125),
    .S(net286),
    .X(_0288_));
 sg13g2_mux2_1 _1591_ (.A0(net201),
    .A1(\add_avg[7] ),
    .S(net286),
    .X(_0287_));
 sg13g2_mux2_1 _1592_ (.A0(net219),
    .A1(net246),
    .S(net286),
    .X(_0286_));
 sg13g2_mux2_1 _1593_ (.A0(net224),
    .A1(net232),
    .S(net286),
    .X(_0285_));
 sg13g2_mux2_1 _1594_ (.A0(\add_up_counter.prob_counter[12] ),
    .A1(net230),
    .S(net286),
    .X(_0284_));
 sg13g2_mux2_1 _1595_ (.A0(net197),
    .A1(net228),
    .S(net286),
    .X(_0283_));
 sg13g2_mux2_1 _1596_ (.A0(\add_up_counter.prob_counter[10] ),
    .A1(net222),
    .S(net286),
    .X(_0282_));
 sg13g2_mux2_1 _1597_ (.A0(net193),
    .A1(net196),
    .S(net286),
    .X(_0281_));
 sg13g2_nand2_1 _1598_ (.Y(_0521_),
    .A(net136),
    .B(net291));
 sg13g2_o21ai_1 _1599_ (.B1(_0521_),
    .Y(_0280_),
    .A1(_0634_),
    .A2(net291));
 sg13g2_nand2_1 _1600_ (.Y(_0522_),
    .A(net116),
    .B(net296));
 sg13g2_a22oi_1 _1601_ (.Y(_0523_),
    .B1(net301),
    .B2(net68),
    .A2(net421),
    .A1(net103));
 sg13g2_o21ai_1 _1602_ (.B1(_0523_),
    .Y(_0028_),
    .A1(net300),
    .A2(_0522_));
 sg13g2_nand2_1 _1603_ (.Y(_0524_),
    .A(net89),
    .B(net296));
 sg13g2_a22oi_1 _1604_ (.Y(_0525_),
    .B1(net300),
    .B2(net72),
    .A2(net297),
    .A1(\mul_output.bitseq[1] ));
 sg13g2_o21ai_1 _1605_ (.B1(_0525_),
    .Y(_0029_),
    .A1(net300),
    .A2(_0524_));
 sg13g2_nand2_1 _1606_ (.Y(_0526_),
    .A(net55),
    .B(net296));
 sg13g2_a22oi_1 _1607_ (.Y(_0527_),
    .B1(net300),
    .B2(\mul_avg[3] ),
    .A2(net297),
    .A1(\mul_output.bitseq[2] ));
 sg13g2_o21ai_1 _1608_ (.B1(_0527_),
    .Y(_0030_),
    .A1(net300),
    .A2(_0526_));
 sg13g2_nand2_1 _1609_ (.Y(_0528_),
    .A(net86),
    .B(net296));
 sg13g2_a22oi_1 _1610_ (.Y(_0529_),
    .B1(net300),
    .B2(net82),
    .A2(net297),
    .A1(net55));
 sg13g2_o21ai_1 _1611_ (.B1(_0529_),
    .Y(_0031_),
    .A1(net300),
    .A2(_0528_));
 sg13g2_nand2_1 _1612_ (.Y(_0530_),
    .A(net233),
    .B(_0671_));
 sg13g2_a22oi_1 _1613_ (.Y(_0531_),
    .B1(net300),
    .B2(net66),
    .A2(net297),
    .A1(net86));
 sg13g2_o21ai_1 _1614_ (.B1(_0531_),
    .Y(_0032_),
    .A1(net302),
    .A2(net234));
 sg13g2_nand2_1 _1615_ (.Y(_0532_),
    .A(net93),
    .B(net296));
 sg13g2_a22oi_1 _1616_ (.Y(_0533_),
    .B1(net301),
    .B2(\mul_avg[6] ),
    .A2(_0670_),
    .A1(\mul_output.bitseq[5] ));
 sg13g2_o21ai_1 _1617_ (.B1(_0533_),
    .Y(_0033_),
    .A1(net302),
    .A2(_0532_));
 sg13g2_nand2_1 _1618_ (.Y(_0534_),
    .A(net91),
    .B(net296));
 sg13g2_a22oi_1 _1619_ (.Y(_0535_),
    .B1(net301),
    .B2(\mul_avg[7] ),
    .A2(net297),
    .A1(\mul_output.bitseq[6] ));
 sg13g2_o21ai_1 _1620_ (.B1(_0535_),
    .Y(_0034_),
    .A1(net301),
    .A2(_0534_));
 sg13g2_nand2_1 _1621_ (.Y(_0536_),
    .A(net52),
    .B(net296));
 sg13g2_a22oi_1 _1622_ (.Y(_0537_),
    .B1(net301),
    .B2(net132),
    .A2(net297),
    .A1(net91));
 sg13g2_o21ai_1 _1623_ (.B1(_0537_),
    .Y(_0035_),
    .A1(net301),
    .A2(_0536_));
 sg13g2_and2_1 _1624_ (.A(net52),
    .B(_0670_),
    .X(_0036_));
 sg13g2_nand2_1 _1625_ (.Y(_0538_),
    .A(net97),
    .B(net298));
 sg13g2_a22oi_1 _1626_ (.Y(_0539_),
    .B1(net305),
    .B2(\add_avg[1] ),
    .A2(net299),
    .A1(\add_output.bitseq[0] ));
 sg13g2_o21ai_1 _1627_ (.B1(_0539_),
    .Y(_0018_),
    .A1(net303),
    .A2(_0538_));
 sg13g2_nand2_1 _1628_ (.Y(_0540_),
    .A(net109),
    .B(net298));
 sg13g2_a22oi_1 _1629_ (.Y(_0541_),
    .B1(net303),
    .B2(\add_avg[2] ),
    .A2(_0646_),
    .A1(net97));
 sg13g2_o21ai_1 _1630_ (.B1(_0541_),
    .Y(_0019_),
    .A1(net303),
    .A2(_0540_));
 sg13g2_nand2_1 _1631_ (.Y(_0542_),
    .A(net95),
    .B(net298));
 sg13g2_a22oi_1 _1632_ (.Y(_0543_),
    .B1(net303),
    .B2(\add_avg[3] ),
    .A2(net299),
    .A1(\add_output.bitseq[2] ));
 sg13g2_o21ai_1 _1633_ (.B1(_0543_),
    .Y(_0020_),
    .A1(net303),
    .A2(_0542_));
 sg13g2_nand2_1 _1634_ (.Y(_0544_),
    .A(net119),
    .B(net298));
 sg13g2_a22oi_1 _1635_ (.Y(_0545_),
    .B1(net303),
    .B2(\add_avg[4] ),
    .A2(_0646_),
    .A1(net95));
 sg13g2_o21ai_1 _1636_ (.B1(_0545_),
    .Y(_0021_),
    .A1(net303),
    .A2(_0544_));
 sg13g2_nand2_1 _1637_ (.Y(_0546_),
    .A(net164),
    .B(_0647_));
 sg13g2_a22oi_1 _1638_ (.Y(_0547_),
    .B1(net304),
    .B2(\add_avg[5] ),
    .A2(_0646_),
    .A1(net119));
 sg13g2_o21ai_1 _1639_ (.B1(_0547_),
    .Y(_0022_),
    .A1(net303),
    .A2(net165));
 sg13g2_nand2_1 _1640_ (.Y(_0548_),
    .A(net128),
    .B(net298));
 sg13g2_a22oi_1 _1641_ (.Y(_0549_),
    .B1(net305),
    .B2(\add_avg[6] ),
    .A2(net299),
    .A1(\add_output.bitseq[5] ));
 sg13g2_o21ai_1 _1642_ (.B1(_0549_),
    .Y(_0023_),
    .A1(net304),
    .A2(_0548_));
 sg13g2_nand2_1 _1643_ (.Y(_0550_),
    .A(net99),
    .B(net298));
 sg13g2_a22oi_1 _1644_ (.Y(_0551_),
    .B1(net305),
    .B2(\add_avg[7] ),
    .A2(net299),
    .A1(\add_output.bitseq[6] ));
 sg13g2_o21ai_1 _1645_ (.B1(_0551_),
    .Y(_0024_),
    .A1(net304),
    .A2(_0550_));
 sg13g2_nand2_1 _1646_ (.Y(_0552_),
    .A(net58),
    .B(net298));
 sg13g2_a22oi_1 _1647_ (.Y(_0553_),
    .B1(net304),
    .B2(net125),
    .A2(net299),
    .A1(net99));
 sg13g2_o21ai_1 _1648_ (.B1(_0553_),
    .Y(_0025_),
    .A1(net304),
    .A2(_0552_));
 sg13g2_and2_1 _1649_ (.A(net58),
    .B(net299),
    .X(_0026_));
 sg13g2_nand2_1 _1650_ (.Y(_0554_),
    .A(net137),
    .B(net294));
 sg13g2_a22oi_1 _1651_ (.Y(_0555_),
    .B1(net295),
    .B2(net104),
    .A2(net307),
    .A1(net60));
 sg13g2_o21ai_1 _1652_ (.B1(_0555_),
    .Y(_0037_),
    .A1(net307),
    .A2(_0554_));
 sg13g2_nand2_1 _1653_ (.Y(_0556_),
    .A(net130),
    .B(_0431_));
 sg13g2_a22oi_1 _1654_ (.Y(_0557_),
    .B1(_0430_),
    .B2(\smul_output.bitseq[1] ),
    .A2(_0429_),
    .A1(net62));
 sg13g2_o21ai_1 _1655_ (.B1(_0557_),
    .Y(_0038_),
    .A1(net307),
    .A2(_0556_));
 sg13g2_nand2_1 _1656_ (.Y(_0558_),
    .A(net199),
    .B(net294));
 sg13g2_a22oi_1 _1657_ (.Y(_0559_),
    .B1(net143),
    .B2(net130),
    .A2(_0429_),
    .A1(net122));
 sg13g2_o21ai_1 _1658_ (.B1(_0559_),
    .Y(_0039_),
    .A1(_0429_),
    .A2(_0558_));
 sg13g2_nand2_1 _1659_ (.Y(_0560_),
    .A(net147),
    .B(net294));
 sg13g2_a22oi_1 _1660_ (.Y(_0561_),
    .B1(net295),
    .B2(\smul_output.bitseq[3] ),
    .A2(net307),
    .A1(net74));
 sg13g2_o21ai_1 _1661_ (.B1(_0561_),
    .Y(_0040_),
    .A1(net307),
    .A2(_0560_));
 sg13g2_nand2_1 _1662_ (.Y(_0562_),
    .A(net157),
    .B(net294));
 sg13g2_a22oi_1 _1663_ (.Y(_0563_),
    .B1(net295),
    .B2(net147),
    .A2(net306),
    .A1(net78));
 sg13g2_o21ai_1 _1664_ (.B1(_0563_),
    .Y(_0041_),
    .A1(net306),
    .A2(_0562_));
 sg13g2_nand2_1 _1665_ (.Y(_0564_),
    .A(net126),
    .B(net294));
 sg13g2_a22oi_1 _1666_ (.Y(_0565_),
    .B1(net295),
    .B2(\smul_output.bitseq[5] ),
    .A2(net306),
    .A1(net64));
 sg13g2_o21ai_1 _1667_ (.B1(_0565_),
    .Y(_0042_),
    .A1(net306),
    .A2(_0564_));
 sg13g2_nand2_1 _1668_ (.Y(_0566_),
    .A(net113),
    .B(net294));
 sg13g2_a22oi_1 _1669_ (.Y(_0567_),
    .B1(net295),
    .B2(\smul_output.bitseq[6] ),
    .A2(net306),
    .A1(net76));
 sg13g2_o21ai_1 _1670_ (.B1(_0567_),
    .Y(_0043_),
    .A1(net306),
    .A2(_0566_));
 sg13g2_nand2_1 _1671_ (.Y(_0568_),
    .A(net59),
    .B(net294));
 sg13g2_a22oi_1 _1672_ (.Y(_0569_),
    .B1(net295),
    .B2(net113),
    .A2(net306),
    .A1(net70));
 sg13g2_o21ai_1 _1673_ (.B1(_0569_),
    .Y(_0044_),
    .A1(net306),
    .A2(_0568_));
 sg13g2_and2_1 _1674_ (.A(net59),
    .B(net144),
    .X(_0045_));
 sg13g2_nor2_1 _1675_ (.A(net372),
    .B(net292),
    .Y(_0000_));
 sg13g2_xor2_1 _1676_ (.B(net372),
    .A(net376),
    .X(_0009_));
 sg13g2_nand3_1 _1677_ (.B(net372),
    .C(net411),
    .A(net376),
    .Y(_0570_));
 sg13g2_a21o_1 _1678_ (.A2(net372),
    .A1(net376),
    .B1(net411),
    .X(_0571_));
 sg13g2_and2_1 _1679_ (.A(_0570_),
    .B(_0571_),
    .X(_0010_));
 sg13g2_and4_2 _1680_ (.A(\add_up_counter.clk_counter[1] ),
    .B(\add_up_counter.clk_counter[0] ),
    .C(net361),
    .D(\add_up_counter.clk_counter[2] ),
    .X(_0572_));
 sg13g2_xnor2_1 _1681_ (.Y(_0011_),
    .A(net361),
    .B(_0570_));
 sg13g2_xor2_1 _1682_ (.B(_0572_),
    .A(net383),
    .X(_0012_));
 sg13g2_nand3_1 _1683_ (.B(\add_up_counter.clk_counter[4] ),
    .C(_0572_),
    .A(net400),
    .Y(_0573_));
 sg13g2_a21o_1 _1684_ (.A2(_0572_),
    .A1(net383),
    .B1(net400),
    .X(_0574_));
 sg13g2_and2_1 _1685_ (.A(_0573_),
    .B(_0574_),
    .X(_0013_));
 sg13g2_nand4_1 _1686_ (.B(\add_up_counter.clk_counter[4] ),
    .C(net226),
    .A(\add_up_counter.clk_counter[5] ),
    .Y(_0575_),
    .D(_0572_));
 sg13g2_xnor2_1 _1687_ (.Y(_0014_),
    .A(net226),
    .B(_0573_));
 sg13g2_nor2_2 _1688_ (.A(_0640_),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_xnor2_1 _1689_ (.Y(_0015_),
    .A(net203),
    .B(_0575_));
 sg13g2_xor2_1 _1690_ (.B(_0576_),
    .A(net351),
    .X(_0016_));
 sg13g2_nand3_1 _1691_ (.B(net351),
    .C(_0576_),
    .A(net392),
    .Y(_0577_));
 sg13g2_a21o_1 _1692_ (.A2(_0576_),
    .A1(net351),
    .B1(net392),
    .X(_0578_));
 sg13g2_and2_1 _1693_ (.A(_0577_),
    .B(_0578_),
    .X(_0017_));
 sg13g2_and4_2 _1694_ (.A(\add_up_counter.clk_counter[9] ),
    .B(\add_up_counter.clk_counter[8] ),
    .C(net194),
    .D(_0576_),
    .X(_0579_));
 sg13g2_xnor2_1 _1695_ (.Y(_0001_),
    .A(net194),
    .B(_0577_));
 sg13g2_xor2_1 _1696_ (.B(_0579_),
    .A(net258),
    .X(_0002_));
 sg13g2_nand3_1 _1697_ (.B(net405),
    .C(_0579_),
    .A(net258),
    .Y(_0580_));
 sg13g2_a21o_1 _1698_ (.A2(_0579_),
    .A1(net258),
    .B1(net405),
    .X(_0581_));
 sg13g2_and2_1 _1699_ (.A(_0580_),
    .B(_0581_),
    .X(_0003_));
 sg13g2_and4_2 _1700_ (.A(net258),
    .B(net206),
    .C(\add_up_counter.clk_counter[12] ),
    .D(_0579_),
    .X(_0582_));
 sg13g2_xnor2_1 _1701_ (.Y(_0004_),
    .A(net206),
    .B(_0580_));
 sg13g2_xor2_1 _1702_ (.B(_0582_),
    .A(net353),
    .X(_0005_));
 sg13g2_a21oi_1 _1703_ (.A1(\add_up_counter.clk_counter[14] ),
    .A2(_0582_),
    .Y(_0583_),
    .B1(net236));
 sg13g2_nand3_1 _1704_ (.B(\add_up_counter.clk_counter[14] ),
    .C(_0582_),
    .A(net236),
    .Y(_0584_));
 sg13g2_nor2b_1 _1705_ (.A(net237),
    .B_N(_0584_),
    .Y(_0006_));
 sg13g2_nand4_1 _1706_ (.B(net353),
    .C(net241),
    .A(net236),
    .Y(_0585_),
    .D(_0582_));
 sg13g2_xnor2_1 _1707_ (.Y(_0007_),
    .A(net241),
    .B(_0584_));
 sg13g2_nand2_1 _1708_ (.Y(_0586_),
    .A(net378),
    .B(net289));
 sg13g2_mux2_1 _1709_ (.A0(net378),
    .A1(_0586_),
    .S(_0585_),
    .X(_0587_));
 sg13g2_inv_1 _1710_ (.Y(_0008_),
    .A(_0587_));
 sg13g2_o21ai_1 _1711_ (.B1(net280),
    .Y(_0027_),
    .A1(_0616_),
    .A2(net292));
 sg13g2_inv_1 _1712_ (.Y(_0061_),
    .A(net318));
 sg13g2_inv_1 _1713_ (.Y(_0062_),
    .A(net313));
 sg13g2_inv_1 _1714_ (.Y(_0063_),
    .A(net313));
 sg13g2_inv_1 _1715_ (.Y(_0064_),
    .A(net313));
 sg13g2_inv_1 _1716_ (.Y(_0065_),
    .A(net313));
 sg13g2_inv_1 _1717_ (.Y(_0066_),
    .A(net319));
 sg13g2_inv_1 _1718_ (.Y(_0067_),
    .A(net319));
 sg13g2_inv_1 _1719_ (.Y(_0068_),
    .A(net319));
 sg13g2_inv_1 _1720_ (.Y(_0069_),
    .A(net335));
 sg13g2_inv_1 _1721_ (.Y(_0070_),
    .A(net335));
 sg13g2_inv_1 _1722_ (.Y(_0071_),
    .A(net335));
 sg13g2_inv_1 _1723_ (.Y(_0072_),
    .A(net335));
 sg13g2_inv_1 _1724_ (.Y(_0073_),
    .A(net335));
 sg13g2_inv_1 _1725_ (.Y(_0074_),
    .A(net335));
 sg13g2_inv_1 _1726_ (.Y(_0075_),
    .A(net334));
 sg13g2_inv_1 _1727_ (.Y(_0076_),
    .A(net334));
 sg13g2_inv_1 _1728_ (.Y(_0077_),
    .A(net331));
 sg13g2_inv_1 _1729_ (.Y(_0078_),
    .A(net331));
 sg13g2_inv_1 _1730_ (.Y(_0079_),
    .A(net330));
 sg13g2_inv_1 _1731_ (.Y(_0080_),
    .A(net332));
 sg13g2_inv_1 _1732_ (.Y(_0081_),
    .A(net332));
 sg13g2_inv_1 _1733_ (.Y(_0082_),
    .A(net323));
 sg13g2_inv_1 _1734_ (.Y(_0083_),
    .A(net322));
 sg13g2_inv_1 _1735_ (.Y(_0084_),
    .A(net323));
 sg13g2_inv_1 _1736_ (.Y(_0085_),
    .A(net322));
 sg13g2_inv_1 _1737_ (.Y(_0086_),
    .A(net323));
 sg13g2_inv_1 _1738_ (.Y(_0087_),
    .A(net323));
 sg13g2_inv_1 _1739_ (.Y(_0088_),
    .A(net325));
 sg13g2_inv_1 _1740_ (.Y(_0089_),
    .A(net323));
 sg13g2_inv_1 _1741_ (.Y(_0090_),
    .A(net329));
 sg13g2_inv_1 _1742_ (.Y(_0091_),
    .A(net345));
 sg13g2_inv_1 _1743_ (.Y(_0092_),
    .A(net345));
 sg13g2_inv_1 _1744_ (.Y(_0093_),
    .A(net340));
 sg13g2_inv_1 _1745_ (.Y(_0094_),
    .A(net345));
 sg13g2_inv_1 _1746_ (.Y(_0095_),
    .A(net345));
 sg13g2_inv_1 _1747_ (.Y(_0096_),
    .A(net337));
 sg13g2_inv_1 _1748_ (.Y(_0097_),
    .A(net313));
 sg13g2_inv_1 _1749_ (.Y(_0098_),
    .A(net314));
 sg13g2_inv_1 _1750_ (.Y(_0099_),
    .A(net314));
 sg13g2_inv_1 _1751_ (.Y(_0100_),
    .A(net313));
 sg13g2_inv_1 _1752_ (.Y(_0101_),
    .A(net316));
 sg13g2_inv_1 _1753_ (.Y(_0102_),
    .A(net316));
 sg13g2_inv_1 _1754_ (.Y(_0103_),
    .A(net316));
 sg13g2_inv_1 _1755_ (.Y(_0104_),
    .A(net316));
 sg13g2_inv_1 _1756_ (.Y(_0105_),
    .A(net315));
 sg13g2_inv_1 _1757_ (.Y(_0106_),
    .A(net337));
 sg13g2_inv_1 _1758_ (.Y(_0107_),
    .A(net337));
 sg13g2_inv_1 _1759_ (.Y(_0108_),
    .A(net336));
 sg13g2_inv_1 _1760_ (.Y(_0109_),
    .A(net336));
 sg13g2_inv_1 _1761_ (.Y(_0110_),
    .A(net333));
 sg13g2_inv_1 _1762_ (.Y(_0111_),
    .A(net333));
 sg13g2_inv_1 _1763_ (.Y(_0112_),
    .A(net332));
 sg13g2_inv_1 _1764_ (.Y(_0113_),
    .A(net332));
 sg13g2_inv_1 _1765_ (.Y(_0114_),
    .A(net332));
 sg13g2_inv_1 _1766_ (.Y(_0115_),
    .A(net332));
 sg13g2_inv_1 _1767_ (.Y(_0116_),
    .A(net322));
 sg13g2_inv_1 _1768_ (.Y(_0117_),
    .A(net322));
 sg13g2_inv_1 _1769_ (.Y(_0118_),
    .A(net315));
 sg13g2_inv_1 _1770_ (.Y(_0119_),
    .A(net315));
 sg13g2_inv_1 _1771_ (.Y(_0120_),
    .A(net315));
 sg13g2_inv_1 _1772_ (.Y(_0121_),
    .A(net315));
 sg13g2_inv_1 _1773_ (.Y(_0122_),
    .A(net315));
 sg13g2_inv_1 _1774_ (.Y(_0123_),
    .A(net316));
 sg13g2_inv_1 _1775_ (.Y(_0124_),
    .A(net319));
 sg13g2_inv_1 _1776_ (.Y(_0125_),
    .A(net316));
 sg13g2_inv_1 _1777_ (.Y(_0126_),
    .A(net316));
 sg13g2_inv_1 _1778_ (.Y(_0127_),
    .A(net316));
 sg13g2_inv_1 _1779_ (.Y(_0128_),
    .A(net322));
 sg13g2_inv_1 _1780_ (.Y(_0129_),
    .A(net322));
 sg13g2_inv_1 _1781_ (.Y(_0130_),
    .A(net328));
 sg13g2_inv_1 _1782_ (.Y(_0131_),
    .A(net328));
 sg13g2_inv_1 _1783_ (.Y(_0132_),
    .A(net319));
 sg13g2_inv_1 _1784_ (.Y(_0133_),
    .A(net336));
 sg13g2_inv_1 _1785_ (.Y(_0134_),
    .A(net345));
 sg13g2_inv_1 _1786_ (.Y(_0135_),
    .A(net344));
 sg13g2_inv_1 _1787_ (.Y(_0136_),
    .A(net345));
 sg13g2_inv_1 _1788_ (.Y(_0137_),
    .A(net344));
 sg13g2_inv_1 _1789_ (.Y(_0138_),
    .A(net344));
 sg13g2_inv_1 _1790_ (.Y(_0139_),
    .A(net344));
 sg13g2_inv_1 _1791_ (.Y(_0140_),
    .A(net344));
 sg13g2_inv_1 _1792_ (.Y(_0141_),
    .A(net344));
 sg13g2_inv_1 _1793_ (.Y(_0142_),
    .A(net337));
 sg13g2_inv_1 _1794_ (.Y(_0143_),
    .A(net337));
 sg13g2_inv_1 _1795_ (.Y(_0144_),
    .A(net337));
 sg13g2_inv_1 _1796_ (.Y(_0145_),
    .A(net337));
 sg13g2_inv_1 _1797_ (.Y(_0146_),
    .A(net336));
 sg13g2_inv_1 _1798_ (.Y(_0147_),
    .A(net336));
 sg13g2_inv_1 _1799_ (.Y(_0148_),
    .A(net336));
 sg13g2_inv_1 _1800_ (.Y(_0149_),
    .A(net336));
 sg13g2_inv_1 _1801_ (.Y(_0150_),
    .A(net333));
 sg13g2_inv_1 _1802_ (.Y(_0151_),
    .A(net336));
 sg13g2_inv_1 _1803_ (.Y(_0152_),
    .A(net326));
 sg13g2_inv_1 _1804_ (.Y(_0153_),
    .A(net326));
 sg13g2_inv_1 _1805_ (.Y(_0154_),
    .A(net325));
 sg13g2_inv_1 _1806_ (.Y(_0155_),
    .A(net340));
 sg13g2_inv_1 _1807_ (.Y(_0156_),
    .A(net340));
 sg13g2_inv_1 _1808_ (.Y(_0157_),
    .A(net346));
 sg13g2_inv_1 _1809_ (.Y(_0158_),
    .A(net346));
 sg13g2_inv_1 _1810_ (.Y(_0159_),
    .A(net348));
 sg13g2_inv_1 _1811_ (.Y(_0160_),
    .A(net348));
 sg13g2_inv_1 _1812_ (.Y(_0161_),
    .A(net340));
 sg13g2_inv_1 _1813_ (.Y(_0162_),
    .A(net317));
 sg13g2_inv_1 _1814_ (.Y(_0163_),
    .A(net317));
 sg13g2_inv_1 _1815_ (.Y(_0164_),
    .A(net317));
 sg13g2_inv_1 _1816_ (.Y(_0165_),
    .A(net317));
 sg13g2_inv_1 _1817_ (.Y(_0166_),
    .A(net317));
 sg13g2_inv_1 _1818_ (.Y(_0167_),
    .A(net317));
 sg13g2_inv_1 _1819_ (.Y(_0168_),
    .A(net317));
 sg13g2_inv_1 _1820_ (.Y(_0169_),
    .A(net317));
 sg13g2_inv_1 _1821_ (.Y(_0170_),
    .A(net318));
 sg13g2_inv_1 _1822_ (.Y(_0171_),
    .A(net318));
 sg13g2_inv_1 _1823_ (.Y(_0172_),
    .A(net318));
 sg13g2_inv_1 _1824_ (.Y(_0173_),
    .A(net313));
 sg13g2_inv_1 _1825_ (.Y(_0174_),
    .A(net313));
 sg13g2_inv_1 _1826_ (.Y(_0175_),
    .A(net318));
 sg13g2_inv_1 _1827_ (.Y(_0176_),
    .A(net320));
 sg13g2_inv_1 _1828_ (.Y(_0177_),
    .A(net320));
 sg13g2_inv_1 _1829_ (.Y(_0178_),
    .A(net319));
 sg13g2_inv_1 _1830_ (.Y(_0179_),
    .A(net326));
 sg13g2_inv_1 _1831_ (.Y(_0180_),
    .A(net341));
 sg13g2_inv_1 _1832_ (.Y(_0181_),
    .A(net341));
 sg13g2_inv_1 _1833_ (.Y(_0182_),
    .A(net341));
 sg13g2_inv_1 _1834_ (.Y(_0183_),
    .A(net341));
 sg13g2_inv_1 _1835_ (.Y(_0184_),
    .A(net347));
 sg13g2_inv_1 _1836_ (.Y(_0185_),
    .A(net347));
 sg13g2_inv_1 _1837_ (.Y(_0186_),
    .A(net346));
 sg13g2_inv_1 _1838_ (.Y(_0187_),
    .A(net347));
 sg13g2_inv_1 _1839_ (.Y(_0188_),
    .A(net326));
 sg13g2_inv_1 _1840_ (.Y(_0189_),
    .A(net341));
 sg13g2_inv_1 _1841_ (.Y(_0190_),
    .A(net341));
 sg13g2_inv_1 _1842_ (.Y(_0191_),
    .A(net342));
 sg13g2_inv_1 _1843_ (.Y(_0192_),
    .A(net346));
 sg13g2_inv_1 _1844_ (.Y(_0193_),
    .A(net346));
 sg13g2_inv_1 _1845_ (.Y(_0194_),
    .A(net347));
 sg13g2_inv_1 _1846_ (.Y(_0195_),
    .A(net347));
 sg13g2_inv_1 _1847_ (.Y(_0196_),
    .A(net347));
 sg13g2_inv_1 _1848_ (.Y(_0197_),
    .A(net340));
 sg13g2_inv_1 _1849_ (.Y(_0198_),
    .A(net333));
 sg13g2_inv_1 _1850_ (.Y(_0199_),
    .A(net332));
 sg13g2_inv_1 _1851_ (.Y(_0200_),
    .A(net332));
 sg13g2_inv_1 _1852_ (.Y(_0201_),
    .A(net325));
 sg13g2_inv_1 _1853_ (.Y(_0202_),
    .A(net325));
 sg13g2_inv_1 _1854_ (.Y(_0203_),
    .A(net325));
 sg13g2_inv_1 _1855_ (.Y(_0204_),
    .A(net340));
 sg13g2_inv_1 _1856_ (.Y(_0205_),
    .A(net343));
 sg13g2_inv_1 _1857_ (.Y(_0206_),
    .A(net345));
 sg13g2_inv_1 _1858_ (.Y(_0207_),
    .A(net344));
 sg13g2_inv_1 _1859_ (.Y(_0208_),
    .A(net344));
 sg13g2_inv_1 _1860_ (.Y(_0209_),
    .A(net347));
 sg13g2_inv_1 _1861_ (.Y(_0211_),
    .A(net328));
 sg13g2_inv_1 _1862_ (.Y(_0213_),
    .A(net326));
 sg13g2_inv_1 _1863_ (.Y(_0214_),
    .A(net340));
 sg13g2_inv_1 _1864_ (.Y(_0215_),
    .A(net340));
 sg13g2_inv_1 _1865_ (.Y(_0216_),
    .A(net343));
 sg13g2_inv_1 _1866_ (.Y(_0217_),
    .A(net343));
 sg13g2_inv_1 _1867_ (.Y(_0218_),
    .A(net342));
 sg13g2_inv_1 _1868_ (.Y(_0219_),
    .A(net342));
 sg13g2_inv_1 _1869_ (.Y(_0220_),
    .A(net342));
 sg13g2_inv_1 _1870_ (.Y(_0222_),
    .A(net326));
 sg13g2_inv_1 _1871_ (.Y(_0224_),
    .A(net326));
 sg13g2_inv_1 _1872_ (.Y(_0226_),
    .A(net328));
 sg13g2_inv_1 _1873_ (.Y(_0227_),
    .A(net326));
 sg13g2_inv_1 _1874_ (.Y(_0228_),
    .A(net328));
 sg13g2_inv_1 _1875_ (.Y(_0229_),
    .A(net341));
 sg13g2_inv_1 _1876_ (.Y(_0230_),
    .A(net341));
 sg13g2_inv_1 _1877_ (.Y(_0231_),
    .A(net342));
 sg13g2_inv_1 _1878_ (.Y(_0232_),
    .A(net342));
 sg13g2_inv_1 _1879_ (.Y(_0233_),
    .A(net346));
 sg13g2_inv_1 _1880_ (.Y(_0234_),
    .A(net346));
 sg13g2_inv_1 _1881_ (.Y(_0235_),
    .A(net346));
 sg13g2_inv_1 _1882_ (.Y(_0236_),
    .A(net327));
 sg13g2_inv_1 _1883_ (.Y(_0237_),
    .A(net327));
 sg13g2_inv_1 _1884_ (.Y(_0238_),
    .A(net327));
 sg13g2_inv_1 _1885_ (.Y(_0239_),
    .A(net324));
 sg13g2_inv_1 _1886_ (.Y(_0240_),
    .A(net324));
 sg13g2_inv_1 _1887_ (.Y(_0241_),
    .A(net324));
 sg13g2_inv_1 _1888_ (.Y(_0242_),
    .A(net327));
 sg13g2_inv_1 _1889_ (.Y(_0243_),
    .A(net327));
 sg13g2_inv_1 _1890_ (.Y(_0244_),
    .A(net327));
 sg13g2_inv_1 _1891_ (.Y(_0245_),
    .A(net327));
 sg13g2_inv_1 _1892_ (.Y(_0246_),
    .A(net330));
 sg13g2_inv_1 _1893_ (.Y(_0247_),
    .A(net330));
 sg13g2_inv_1 _1894_ (.Y(_0248_),
    .A(net330));
 sg13g2_inv_1 _1895_ (.Y(_0249_),
    .A(net331));
 sg13g2_inv_1 _1896_ (.Y(_0250_),
    .A(net330));
 sg13g2_inv_1 _1897_ (.Y(_0251_),
    .A(net334));
 sg13g2_inv_1 _1898_ (.Y(_0252_),
    .A(net334));
 sg13g2_inv_1 _1899_ (.Y(_0253_),
    .A(net334));
 sg13g2_inv_1 _1900_ (.Y(_0254_),
    .A(net338));
 sg13g2_inv_1 _1901_ (.Y(_0255_),
    .A(net334));
 sg13g2_inv_1 _1902_ (.Y(_0256_),
    .A(net334));
 sg13g2_inv_1 _1903_ (.Y(_0257_),
    .A(net334));
 sg13g2_inv_1 _1904_ (.Y(_0258_),
    .A(net335));
 sg13g2_inv_1 _1905_ (.Y(_0259_),
    .A(net331));
 sg13g2_inv_1 _1906_ (.Y(_0260_),
    .A(net330));
 sg13g2_inv_1 _1907_ (.Y(_0261_),
    .A(net330));
 sg13g2_inv_1 _1908_ (.Y(_0262_),
    .A(net330));
 sg13g2_inv_1 _1909_ (.Y(_0263_),
    .A(net329));
 sg13g2_inv_1 _1910_ (.Y(_0264_),
    .A(net324));
 sg13g2_inv_1 _1911_ (.Y(_0265_),
    .A(net324));
 sg13g2_inv_1 _1912_ (.Y(_0266_),
    .A(net324));
 sg13g2_inv_1 _1913_ (.Y(_0267_),
    .A(net319));
 sg13g2_inv_1 _1914_ (.Y(_0268_),
    .A(net324));
 sg13g2_inv_1 _1915_ (.Y(_0269_),
    .A(net322));
 sg13g2_inv_1 _1916_ (.Y(_0270_),
    .A(net323));
 sg13g2_inv_1 _1917_ (.Y(_0271_),
    .A(net323));
 sg13g2_inv_1 _1918_ (.Y(_0272_),
    .A(net322));
 sg13g2_inv_1 _1919_ (.Y(_0273_),
    .A(net325));
 sg13g2_inv_1 _1920_ (.Y(_0274_),
    .A(net325));
 sg13g2_inv_1 _1921_ (.Y(_0275_),
    .A(net325));
 sg13g2_inv_1 _1922_ (.Y(_0276_),
    .A(net314));
 sg13g2_inv_1 _1923_ (.Y(_0277_),
    .A(net315));
 sg13g2_inv_1 _1924_ (.Y(_0278_),
    .A(net315));
 sg13g2_inv_1 _1925_ (.Y(_0279_),
    .A(net314));
 sg13g2_dfrbp_1 _1926_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0060_),
    .D(_0280_),
    .Q_N(_1069_),
    .Q(\add_avg[0] ));
 sg13g2_dfrbp_1 _1927_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0061_),
    .D(_0281_),
    .Q_N(_1068_),
    .Q(\add_avg[1] ));
 sg13g2_dfrbp_1 _1928_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0062_),
    .D(net223),
    .Q_N(_1067_),
    .Q(\add_avg[2] ));
 sg13g2_dfrbp_1 _1929_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0063_),
    .D(_0283_),
    .Q_N(_1066_),
    .Q(\add_avg[3] ));
 sg13g2_dfrbp_1 _1930_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0064_),
    .D(net231),
    .Q_N(_1065_),
    .Q(\add_avg[4] ));
 sg13g2_dfrbp_1 _1931_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0065_),
    .D(_0285_),
    .Q_N(_1064_),
    .Q(\add_avg[5] ));
 sg13g2_dfrbp_1 _1932_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0066_),
    .D(_0286_),
    .Q_N(_1063_),
    .Q(\add_avg[6] ));
 sg13g2_dfrbp_1 _1933_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0067_),
    .D(net202),
    .Q_N(_1062_),
    .Q(\add_avg[7] ));
 sg13g2_dfrbp_1 _1934_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0068_),
    .D(_0288_),
    .Q_N(_1061_),
    .Q(\add_avg[8] ));
 sg13g2_dfrbp_1 _1935_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0069_),
    .D(_0289_),
    .Q_N(_1060_),
    .Q(\smul_output.counter[0] ));
 sg13g2_dfrbp_1 _1936_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0070_),
    .D(_0290_),
    .Q_N(_1059_),
    .Q(\smul_output.counter[1] ));
 sg13g2_dfrbp_1 _1937_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0071_),
    .D(net255),
    .Q_N(_1058_),
    .Q(\smul_output.counter[2] ));
 sg13g2_dfrbp_1 _1938_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0072_),
    .D(_0292_),
    .Q_N(_1057_),
    .Q(\smul_output.counter[3] ));
 sg13g2_dfrbp_1 _1939_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0073_),
    .D(net88),
    .Q_N(_1056_),
    .Q(\smul_avg[0] ));
 sg13g2_dfrbp_1 _1940_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0074_),
    .D(net61),
    .Q_N(_1055_),
    .Q(\smul_avg[1] ));
 sg13g2_dfrbp_1 _1941_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0075_),
    .D(net63),
    .Q_N(_1054_),
    .Q(\smul_avg[2] ));
 sg13g2_dfrbp_1 _1942_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0076_),
    .D(net123),
    .Q_N(_1053_),
    .Q(\smul_avg[3] ));
 sg13g2_dfrbp_1 _1943_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0077_),
    .D(net75),
    .Q_N(_1052_),
    .Q(\smul_avg[4] ));
 sg13g2_dfrbp_1 _1944_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0078_),
    .D(net79),
    .Q_N(_1051_),
    .Q(\smul_avg[5] ));
 sg13g2_dfrbp_1 _1945_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0079_),
    .D(net65),
    .Q_N(_1050_),
    .Q(\smul_avg[6] ));
 sg13g2_dfrbp_1 _1946_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0080_),
    .D(net77),
    .Q_N(_1049_),
    .Q(\smul_avg[7] ));
 sg13g2_dfrbp_1 _1947_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0081_),
    .D(net71),
    .Q_N(_1048_),
    .Q(\smul_avg[8] ));
 sg13g2_dfrbp_1 _1948_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0082_),
    .D(_0028_),
    .Q_N(_1047_),
    .Q(\mul_output.bitseq[0] ));
 sg13g2_dfrbp_1 _1949_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0083_),
    .D(net90),
    .Q_N(_1046_),
    .Q(\mul_output.bitseq[1] ));
 sg13g2_dfrbp_1 _1950_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0084_),
    .D(net56),
    .Q_N(_1045_),
    .Q(\mul_output.bitseq[2] ));
 sg13g2_dfrbp_1 _1951_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0085_),
    .D(_0031_),
    .Q_N(_1044_),
    .Q(\mul_output.bitseq[3] ));
 sg13g2_dfrbp_1 _1952_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0086_),
    .D(_0032_),
    .Q_N(_1043_),
    .Q(\mul_output.bitseq[4] ));
 sg13g2_dfrbp_1 _1953_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0087_),
    .D(net94),
    .Q_N(_1042_),
    .Q(\mul_output.bitseq[5] ));
 sg13g2_dfrbp_1 _1954_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0088_),
    .D(net92),
    .Q_N(_1041_),
    .Q(\mul_output.bitseq[6] ));
 sg13g2_dfrbp_1 _1955_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0089_),
    .D(_0035_),
    .Q_N(_1040_),
    .Q(\mul_output.bitseq[7] ));
 sg13g2_dfrbp_1 _1956_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0090_),
    .D(net53),
    .Q_N(_1039_),
    .Q(\mul_output.bitseq[8] ));
 sg13g2_dfrbp_1 _1957_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0091_),
    .D(net150),
    .Q_N(\global_input.adjustment[0] ),
    .Q(_0049_));
 sg13g2_dfrbp_1 _1958_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0092_),
    .D(net118),
    .Q_N(_1038_),
    .Q(\global_input.adjustment[1] ));
 sg13g2_dfrbp_1 _1959_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0093_),
    .D(net251),
    .Q_N(_1037_),
    .Q(\global_input.adjustment[2] ));
 sg13g2_dfrbp_1 _1960_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0094_),
    .D(net134),
    .Q_N(\global_input.adjustment[3] ),
    .Q(_0050_));
 sg13g2_dfrbp_1 _1961_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0095_),
    .D(net161),
    .Q_N(_1036_),
    .Q(\global_input.adjustment[4] ));
 sg13g2_dfrbp_1 _1962_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0096_),
    .D(_0307_),
    .Q_N(_1035_),
    .Q(mul_bit_out));
 sg13g2_dfrbp_1 _1963_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0097_),
    .D(net98),
    .Q_N(_1034_),
    .Q(\add_output.bitseq[0] ));
 sg13g2_dfrbp_1 _1964_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0098_),
    .D(net110),
    .Q_N(_1033_),
    .Q(\add_output.bitseq[1] ));
 sg13g2_dfrbp_1 _1965_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0099_),
    .D(net96),
    .Q_N(_1032_),
    .Q(\add_output.bitseq[2] ));
 sg13g2_dfrbp_1 _1966_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0100_),
    .D(net120),
    .Q_N(_1031_),
    .Q(\add_output.bitseq[3] ));
 sg13g2_dfrbp_1 _1967_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0101_),
    .D(net166),
    .Q_N(_1030_),
    .Q(\add_output.bitseq[4] ));
 sg13g2_dfrbp_1 _1968_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0102_),
    .D(net129),
    .Q_N(_1029_),
    .Q(\add_output.bitseq[5] ));
 sg13g2_dfrbp_1 _1969_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0103_),
    .D(net100),
    .Q_N(_1028_),
    .Q(\add_output.bitseq[6] ));
 sg13g2_dfrbp_1 _1970_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0104_),
    .D(_0025_),
    .Q_N(_1027_),
    .Q(\add_output.bitseq[7] ));
 sg13g2_dfrbp_1 _1971_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0105_),
    .D(_0026_),
    .Q_N(_1026_),
    .Q(\add_output.bitseq[8] ));
 sg13g2_dfrbp_1 _1972_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0106_),
    .D(net106),
    .Q_N(_1025_),
    .Q(add_bit_out));
 sg13g2_dfrbp_1 _1973_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0107_),
    .D(_0037_),
    .Q_N(_1024_),
    .Q(\smul_output.bitseq[0] ));
 sg13g2_dfrbp_1 _1974_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0108_),
    .D(net131),
    .Q_N(_1023_),
    .Q(\smul_output.bitseq[1] ));
 sg13g2_dfrbp_1 _1975_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0109_),
    .D(net200),
    .Q_N(_1022_),
    .Q(\smul_output.bitseq[2] ));
 sg13g2_dfrbp_1 _1976_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0110_),
    .D(net148),
    .Q_N(_1021_),
    .Q(\smul_output.bitseq[3] ));
 sg13g2_dfrbp_1 _1977_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0111_),
    .D(_0041_),
    .Q_N(_1020_),
    .Q(\smul_output.bitseq[4] ));
 sg13g2_dfrbp_1 _1978_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0112_),
    .D(net127),
    .Q_N(_1019_),
    .Q(\smul_output.bitseq[5] ));
 sg13g2_dfrbp_1 _1979_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0113_),
    .D(net114),
    .Q_N(_1018_),
    .Q(\smul_output.bitseq[6] ));
 sg13g2_dfrbp_1 _1980_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0114_),
    .D(_0044_),
    .Q_N(_1017_),
    .Q(\smul_output.bitseq[7] ));
 sg13g2_dfrbp_1 _1981_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0115_),
    .D(_0045_),
    .Q_N(_1016_),
    .Q(\smul_output.bitseq[8] ));
 sg13g2_dfrbp_1 _1982_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0116_),
    .D(_0309_),
    .Q_N(_1015_),
    .Q(\mul_up_counter.prob_counter[0] ));
 sg13g2_dfrbp_1 _1983_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0117_),
    .D(_0310_),
    .Q_N(_1014_),
    .Q(\mul_up_counter.prob_counter[1] ));
 sg13g2_dfrbp_1 _1984_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0118_),
    .D(_0311_),
    .Q_N(_1013_),
    .Q(\mul_up_counter.prob_counter[2] ));
 sg13g2_dfrbp_1 _1985_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0119_),
    .D(net396),
    .Q_N(_1012_),
    .Q(\mul_up_counter.prob_counter[3] ));
 sg13g2_dfrbp_1 _1986_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0120_),
    .D(_0313_),
    .Q_N(_1011_),
    .Q(\mul_up_counter.prob_counter[4] ));
 sg13g2_dfrbp_1 _1987_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0121_),
    .D(net386),
    .Q_N(_1010_),
    .Q(\mul_up_counter.prob_counter[5] ));
 sg13g2_dfrbp_1 _1988_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0122_),
    .D(net388),
    .Q_N(_1009_),
    .Q(\mul_up_counter.prob_counter[6] ));
 sg13g2_dfrbp_1 _1989_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0123_),
    .D(_0316_),
    .Q_N(_1008_),
    .Q(\mul_up_counter.prob_counter[7] ));
 sg13g2_dfrbp_1 _1990_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0124_),
    .D(_0317_),
    .Q_N(_1007_),
    .Q(\mul_up_counter.prob_counter[8] ));
 sg13g2_dfrbp_1 _1991_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0125_),
    .D(_0318_),
    .Q_N(_1006_),
    .Q(\mul_up_counter.prob_counter[9] ));
 sg13g2_dfrbp_1 _1992_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0126_),
    .D(_0319_),
    .Q_N(_1005_),
    .Q(\mul_up_counter.prob_counter[10] ));
 sg13g2_dfrbp_1 _1993_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0127_),
    .D(_0320_),
    .Q_N(_1004_),
    .Q(\mul_up_counter.prob_counter[11] ));
 sg13g2_dfrbp_1 _1994_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0128_),
    .D(_0321_),
    .Q_N(_1003_),
    .Q(\mul_up_counter.prob_counter[12] ));
 sg13g2_dfrbp_1 _1995_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0129_),
    .D(net399),
    .Q_N(_1002_),
    .Q(\mul_up_counter.prob_counter[13] ));
 sg13g2_dfrbp_1 _1996_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0130_),
    .D(_0323_),
    .Q_N(_1001_),
    .Q(\mul_up_counter.prob_counter[14] ));
 sg13g2_dfrbp_1 _1997_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0131_),
    .D(_0324_),
    .Q_N(_1000_),
    .Q(\mul_up_counter.prob_counter[15] ));
 sg13g2_dfrbp_1 _1998_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0132_),
    .D(_0325_),
    .Q_N(_0047_),
    .Q(\mul_up_counter.prob_counter[16] ));
 sg13g2_dfrbp_1 _1999_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0133_),
    .D(_0326_),
    .Q_N(_0999_),
    .Q(smul_bit_out));
 sg13g2_dfrbp_1 _2000_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0134_),
    .D(_0000_),
    .Q_N(_0998_),
    .Q(\add_up_counter.clk_counter[0] ));
 sg13g2_dfrbp_1 _2001_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0135_),
    .D(_0009_),
    .Q_N(_0997_),
    .Q(\add_up_counter.clk_counter[1] ));
 sg13g2_dfrbp_1 _2002_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0136_),
    .D(_0010_),
    .Q_N(_0996_),
    .Q(\add_up_counter.clk_counter[2] ));
 sg13g2_dfrbp_1 _2003_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0137_),
    .D(net362),
    .Q_N(_0995_),
    .Q(\add_up_counter.clk_counter[3] ));
 sg13g2_dfrbp_1 _2004_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0138_),
    .D(net384),
    .Q_N(_0994_),
    .Q(\add_up_counter.clk_counter[4] ));
 sg13g2_dfrbp_1 _2005_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0139_),
    .D(net401),
    .Q_N(_0993_),
    .Q(\add_up_counter.clk_counter[5] ));
 sg13g2_dfrbp_1 _2006_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0140_),
    .D(net227),
    .Q_N(_0992_),
    .Q(\add_up_counter.clk_counter[6] ));
 sg13g2_dfrbp_1 _2007_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0141_),
    .D(net204),
    .Q_N(_0991_),
    .Q(\add_up_counter.clk_counter[7] ));
 sg13g2_dfrbp_1 _2008_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0142_),
    .D(net352),
    .Q_N(_0990_),
    .Q(\add_up_counter.clk_counter[8] ));
 sg13g2_dfrbp_1 _2009_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0143_),
    .D(_0017_),
    .Q_N(_0989_),
    .Q(\add_up_counter.clk_counter[9] ));
 sg13g2_dfrbp_1 _2010_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0144_),
    .D(net195),
    .Q_N(_0988_),
    .Q(\add_up_counter.clk_counter[10] ));
 sg13g2_dfrbp_1 _2011_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0145_),
    .D(net259),
    .Q_N(_0987_),
    .Q(\add_up_counter.clk_counter[11] ));
 sg13g2_dfrbp_1 _2012_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0146_),
    .D(_0003_),
    .Q_N(_0986_),
    .Q(\add_up_counter.clk_counter[12] ));
 sg13g2_dfrbp_1 _2013_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0147_),
    .D(net207),
    .Q_N(_0985_),
    .Q(\add_up_counter.clk_counter[13] ));
 sg13g2_dfrbp_1 _2014_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0148_),
    .D(net354),
    .Q_N(_0984_),
    .Q(\add_up_counter.clk_counter[14] ));
 sg13g2_dfrbp_1 _2015_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0149_),
    .D(net238),
    .Q_N(_0983_),
    .Q(\add_up_counter.clk_counter[15] ));
 sg13g2_dfrbp_1 _2016_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0150_),
    .D(net242),
    .Q_N(_0982_),
    .Q(\add_up_counter.clk_counter[16] ));
 sg13g2_dfrbp_1 _2017_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0151_),
    .D(_0008_),
    .Q_N(_0981_),
    .Q(\add_up_counter.clk_counter[17] ));
 sg13g2_dfrbp_1 _2018_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0152_),
    .D(net213),
    .Q_N(_0980_),
    .Q(\global_SN_gen.Input_1[0] ));
 sg13g2_dfrbp_1 _2019_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0153_),
    .D(_0328_),
    .Q_N(_0979_),
    .Q(\global_SN_gen.Input_1[1] ));
 sg13g2_dfrbp_1 _2020_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0154_),
    .D(_0329_),
    .Q_N(_0978_),
    .Q(\global_SN_gen.Input_1[2] ));
 sg13g2_dfrbp_1 _2021_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0155_),
    .D(net108),
    .Q_N(_0977_),
    .Q(\global_SN_gen.Input_1[3] ));
 sg13g2_dfrbp_1 _2022_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0156_),
    .D(_0331_),
    .Q_N(_0976_),
    .Q(\global_SN_gen.Input_1[4] ));
 sg13g2_dfrbp_1 _2023_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0157_),
    .D(_0332_),
    .Q_N(_0975_),
    .Q(\global_SN_gen.Input_1[5] ));
 sg13g2_dfrbp_1 _2024_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0158_),
    .D(_0333_),
    .Q_N(_0974_),
    .Q(\global_SN_gen.Input_1[6] ));
 sg13g2_dfrbp_1 _2025_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0159_),
    .D(net187),
    .Q_N(_0973_),
    .Q(\global_SN_gen.Input_1[7] ));
 sg13g2_dfrbp_1 _2026_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0160_),
    .D(net192),
    .Q_N(_0972_),
    .Q(\global_SN_gen.Input_1[8] ));
 sg13g2_dfrbp_1 _2027_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0161_),
    .D(_0027_),
    .Q_N(_0971_),
    .Q(\global_input.loop ));
 sg13g2_dfrbp_1 _2028_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0162_),
    .D(_0336_),
    .Q_N(_0970_),
    .Q(\add_up_counter.prob_counter[0] ));
 sg13g2_dfrbp_1 _2029_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0163_),
    .D(net262),
    .Q_N(_0969_),
    .Q(\add_up_counter.prob_counter[1] ));
 sg13g2_dfrbp_1 _2030_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0164_),
    .D(net141),
    .Q_N(_0968_),
    .Q(\add_up_counter.prob_counter[2] ));
 sg13g2_dfrbp_1 _2031_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0165_),
    .D(_0339_),
    .Q_N(_0967_),
    .Q(\add_up_counter.prob_counter[3] ));
 sg13g2_dfrbp_1 _2032_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0166_),
    .D(_0340_),
    .Q_N(_0966_),
    .Q(\add_up_counter.prob_counter[4] ));
 sg13g2_dfrbp_1 _2033_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0167_),
    .D(net209),
    .Q_N(_0965_),
    .Q(\add_up_counter.prob_counter[5] ));
 sg13g2_dfrbp_1 _2034_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0168_),
    .D(net183),
    .Q_N(_0964_),
    .Q(\add_up_counter.prob_counter[6] ));
 sg13g2_dfrbp_1 _2035_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0169_),
    .D(_0343_),
    .Q_N(_0963_),
    .Q(\add_up_counter.prob_counter[7] ));
 sg13g2_dfrbp_1 _2036_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0170_),
    .D(_0344_),
    .Q_N(_0962_),
    .Q(\add_up_counter.prob_counter[8] ));
 sg13g2_dfrbp_1 _2037_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0171_),
    .D(_0345_),
    .Q_N(_0961_),
    .Q(\add_up_counter.prob_counter[9] ));
 sg13g2_dfrbp_1 _2038_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0172_),
    .D(net257),
    .Q_N(_0960_),
    .Q(\add_up_counter.prob_counter[10] ));
 sg13g2_dfrbp_1 _2039_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_0173_),
    .D(net198),
    .Q_N(_0959_),
    .Q(\add_up_counter.prob_counter[11] ));
 sg13g2_dfrbp_1 _2040_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0174_),
    .D(_0348_),
    .Q_N(_0958_),
    .Q(\add_up_counter.prob_counter[12] ));
 sg13g2_dfrbp_1 _2041_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0175_),
    .D(net225),
    .Q_N(_0957_),
    .Q(\add_up_counter.prob_counter[13] ));
 sg13g2_dfrbp_1 _2042_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0176_),
    .D(net220),
    .Q_N(_0956_),
    .Q(\add_up_counter.prob_counter[14] ));
 sg13g2_dfrbp_1 _2043_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0177_),
    .D(_0351_),
    .Q_N(_0955_),
    .Q(\add_up_counter.prob_counter[15] ));
 sg13g2_dfrbp_1 _2044_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0178_),
    .D(net85),
    .Q_N(_0048_),
    .Q(\add_up_counter.prob_counter[16] ));
 sg13g2_dfrbp_1 _2045_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0179_),
    .D(_0353_),
    .Q_N(_0954_),
    .Q(\global_SN_gen.Input_2[0] ));
 sg13g2_dfrbp_1 _2046_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0180_),
    .D(net163),
    .Q_N(_0953_),
    .Q(\global_SN_gen.Input_2[1] ));
 sg13g2_dfrbp_1 _2047_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0181_),
    .D(_0355_),
    .Q_N(_0952_),
    .Q(\global_SN_gen.Input_2[2] ));
 sg13g2_dfrbp_1 _2048_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0182_),
    .D(net139),
    .Q_N(_0951_),
    .Q(\global_SN_gen.Input_2[3] ));
 sg13g2_dfrbp_1 _2049_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0183_),
    .D(net168),
    .Q_N(_0950_),
    .Q(\global_SN_gen.Input_2[4] ));
 sg13g2_dfrbp_1 _2050_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0184_),
    .D(net174),
    .Q_N(_0949_),
    .Q(\global_SN_gen.Input_2[5] ));
 sg13g2_dfrbp_1 _2051_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0185_),
    .D(net176),
    .Q_N(_0948_),
    .Q(\global_SN_gen.Input_2[6] ));
 sg13g2_dfrbp_1 _2052_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0186_),
    .D(net156),
    .Q_N(_0947_),
    .Q(\global_SN_gen.Input_2[7] ));
 sg13g2_dfrbp_1 _2053_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0187_),
    .D(net159),
    .Q_N(_0946_),
    .Q(\global_SN_gen.Input_2[8] ));
 sg13g2_dfrbp_1 _2054_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0188_),
    .D(net154),
    .Q_N(_0945_),
    .Q(\global_input.output_bitcounter_2[0] ));
 sg13g2_dfrbp_1 _2055_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0189_),
    .D(_0363_),
    .Q_N(_0944_),
    .Q(\global_input.output_bitcounter_2[1] ));
 sg13g2_dfrbp_1 _2056_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0190_),
    .D(_0364_),
    .Q_N(_0943_),
    .Q(\global_input.output_bitcounter_2[2] ));
 sg13g2_dfrbp_1 _2057_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0191_),
    .D(_0365_),
    .Q_N(_0942_),
    .Q(\global_input.output_bitcounter_2[3] ));
 sg13g2_dfrbp_1 _2058_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0192_),
    .D(_0366_),
    .Q_N(_0941_),
    .Q(\global_input.output_bitcounter_2[4] ));
 sg13g2_dfrbp_1 _2059_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0193_),
    .D(_0367_),
    .Q_N(_0940_),
    .Q(\global_input.output_bitcounter_2[5] ));
 sg13g2_dfrbp_1 _2060_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0194_),
    .D(_0368_),
    .Q_N(_0939_),
    .Q(\global_input.output_bitcounter_2[6] ));
 sg13g2_dfrbp_1 _2061_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0195_),
    .D(_0369_),
    .Q_N(_0938_),
    .Q(\global_input.output_bitcounter_2[7] ));
 sg13g2_dfrbp_1 _2062_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0196_),
    .D(_0370_),
    .Q_N(_0937_),
    .Q(\global_input.output_bitcounter_2[8] ));
 sg13g2_dfrbp_1 _2063_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0197_),
    .D(_0371_),
    .Q_N(_0936_),
    .Q(\global_input.output_case[0] ));
 sg13g2_dfrbp_1 _2064_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0198_),
    .D(_0372_),
    .Q_N(_0935_),
    .Q(\global_input.output_case[1] ));
 sg13g2_dfrbp_1 _2065_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0199_),
    .D(net253),
    .Q_N(_0934_),
    .Q(\global_input.output_case[2] ));
 sg13g2_dfrbp_1 _2066_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0200_),
    .D(_0374_),
    .Q_N(_0933_),
    .Q(\global_input.output_case[3] ));
 sg13g2_dfrbp_1 _2067_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0201_),
    .D(net172),
    .Q_N(_0932_),
    .Q(\global_input.output_bitcounter_1[0] ));
 sg13g2_dfrbp_1 _2068_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0202_),
    .D(_0376_),
    .Q_N(_0931_),
    .Q(\global_input.output_bitcounter_1[1] ));
 sg13g2_dfrbp_1 _2069_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0203_),
    .D(_0377_),
    .Q_N(_0930_),
    .Q(\global_input.output_bitcounter_1[2] ));
 sg13g2_dfrbp_1 _2070_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0204_),
    .D(_0378_),
    .Q_N(_0929_),
    .Q(\global_input.output_bitcounter_1[3] ));
 sg13g2_dfrbp_1 _2071_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0205_),
    .D(_0379_),
    .Q_N(_0928_),
    .Q(\global_input.output_bitcounter_1[4] ));
 sg13g2_dfrbp_1 _2072_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0206_),
    .D(net112),
    .Q_N(_0927_),
    .Q(\global_input.output_bitcounter_1[5] ));
 sg13g2_dfrbp_1 _2073_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0207_),
    .D(_0381_),
    .Q_N(_0926_),
    .Q(\global_input.output_bitcounter_1[6] ));
 sg13g2_dfrbp_1 _2074_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0208_),
    .D(_0382_),
    .Q_N(_0925_),
    .Q(\global_input.output_bitcounter_1[7] ));
 sg13g2_dfrbp_1 _2075_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0209_),
    .D(_0383_),
    .Q_N(_0924_),
    .Q(\global_input.output_bitcounter_1[8] ));
 sg13g2_dfrbp_1 _2076_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0211_),
    .D(_0210_),
    .Q_N(\global_SN_gen.lfsr[0] ),
    .Q(_0051_));
 sg13g2_dfrbp_1 _2077_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0213_),
    .D(_0212_),
    .Q_N(\global_SN_gen.lfsr[1] ),
    .Q(_0052_));
 sg13g2_dfrbp_1 _2078_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0214_),
    .D(net42),
    .Q_N(_0923_),
    .Q(\global_SN_gen.lfsr[2] ));
 sg13g2_dfrbp_1 _2079_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0215_),
    .D(net47),
    .Q_N(_0922_),
    .Q(\global_SN_gen.lfsr[3] ));
 sg13g2_dfrbp_1 _2080_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0216_),
    .D(net24),
    .Q_N(\global_SN_gen.lfsr[4] ),
    .Q(_0053_));
 sg13g2_dfrbp_1 _2081_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0217_),
    .D(net34),
    .Q_N(_0921_),
    .Q(\global_SN_gen.lfsr[5] ));
 sg13g2_dfrbp_1 _2082_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0218_),
    .D(net28),
    .Q_N(\global_SN_gen.lfsr[6] ),
    .Q(_0054_));
 sg13g2_dfrbp_1 _2083_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0219_),
    .D(net33),
    .Q_N(_0920_),
    .Q(\global_SN_gen.lfsr[7] ));
 sg13g2_dfrbp_1 _2084_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0220_),
    .D(net27),
    .Q_N(\global_SN_gen.lfsr[8] ),
    .Q(_0055_));
 sg13g2_dfrbp_1 _2085_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0222_),
    .D(_0221_),
    .Q_N(\global_SN_gen.lfsr[9] ),
    .Q(_0056_));
 sg13g2_dfrbp_1 _2086_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0224_),
    .D(_0223_),
    .Q_N(\global_SN_gen.lfsr[10] ),
    .Q(_0057_));
 sg13g2_dfrbp_1 _2087_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0226_),
    .D(_0225_),
    .Q_N(\global_SN_gen.lfsr[11] ),
    .Q(_0058_));
 sg13g2_dfrbp_1 _2088_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0227_),
    .D(net25),
    .Q_N(_0919_),
    .Q(\global_SN_gen.lfsr[12] ));
 sg13g2_dfrbp_1 _2089_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0228_),
    .D(net44),
    .Q_N(_0918_),
    .Q(\global_SN_gen.lfsr[13] ));
 sg13g2_dfrbp_1 _2090_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0229_),
    .D(net51),
    .Q_N(_0917_),
    .Q(\global_SN_gen.lfsr[14] ));
 sg13g2_dfrbp_1 _2091_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0230_),
    .D(net45),
    .Q_N(_0916_),
    .Q(\global_SN_gen.lfsr[15] ));
 sg13g2_dfrbp_1 _2092_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0231_),
    .D(net57),
    .Q_N(_0915_),
    .Q(\global_SN_gen.lfsr[16] ));
 sg13g2_dfrbp_1 _2093_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0232_),
    .D(net26),
    .Q_N(\global_SN_gen.lfsr[17] ),
    .Q(_0059_));
 sg13g2_dfrbp_1 _2094_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0233_),
    .D(net50),
    .Q_N(_0914_),
    .Q(\global_SN_gen.lfsr[18] ));
 sg13g2_dfrbp_1 _2095_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0234_),
    .D(net46),
    .Q_N(_0913_),
    .Q(\global_SN_gen.lfsr[19] ));
 sg13g2_dfrbp_1 _2096_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0235_),
    .D(net48),
    .Q_N(_0912_),
    .Q(\global_SN_gen.lfsr[20] ));
 sg13g2_dfrbp_1 _2097_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0236_),
    .D(net121),
    .Q_N(_0911_),
    .Q(\global_SN_gen.lfsr[21] ));
 sg13g2_dfrbp_1 _2098_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0237_),
    .D(net38),
    .Q_N(_0910_),
    .Q(\global_SN_gen.lfsr[22] ));
 sg13g2_dfrbp_1 _2099_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0238_),
    .D(net39),
    .Q_N(_0909_),
    .Q(\global_SN_gen.lfsr[23] ));
 sg13g2_dfrbp_1 _2100_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0239_),
    .D(net32),
    .Q_N(_0908_),
    .Q(\global_SN_gen.lfsr[24] ));
 sg13g2_dfrbp_1 _2101_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0240_),
    .D(net37),
    .Q_N(_0907_),
    .Q(\global_SN_gen.lfsr[25] ));
 sg13g2_dfrbp_1 _2102_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0241_),
    .D(net35),
    .Q_N(_0906_),
    .Q(\global_SN_gen.lfsr[26] ));
 sg13g2_dfrbp_1 _2103_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0242_),
    .D(net40),
    .Q_N(_0905_),
    .Q(\global_SN_gen.lfsr[27] ));
 sg13g2_dfrbp_1 _2104_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0243_),
    .D(net43),
    .Q_N(_0904_),
    .Q(\global_SN_gen.lfsr[28] ));
 sg13g2_dfrbp_1 _2105_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0244_),
    .D(net31),
    .Q_N(_0903_),
    .Q(\global_SN_gen.lfsr[29] ));
 sg13g2_dfrbp_1 _2106_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0245_),
    .D(net36),
    .Q_N(_0902_),
    .Q(\global_SN_gen.lfsr[30] ));
 sg13g2_dfrbp_1 _2107_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0246_),
    .D(_0384_),
    .Q_N(_0901_),
    .Q(\smul_up_counter.prob_counter[0] ));
 sg13g2_dfrbp_1 _2108_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0247_),
    .D(_0385_),
    .Q_N(_0900_),
    .Q(\smul_up_counter.prob_counter[1] ));
 sg13g2_dfrbp_1 _2109_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0248_),
    .D(net350),
    .Q_N(_0899_),
    .Q(\smul_up_counter.prob_counter[2] ));
 sg13g2_dfrbp_1 _2110_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0249_),
    .D(net245),
    .Q_N(_0898_),
    .Q(\smul_up_counter.prob_counter[3] ));
 sg13g2_dfrbp_1 _2111_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0250_),
    .D(_0388_),
    .Q_N(_0897_),
    .Q(\smul_up_counter.prob_counter[4] ));
 sg13g2_dfrbp_1 _2112_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0251_),
    .D(_0389_),
    .Q_N(_0896_),
    .Q(\smul_up_counter.prob_counter[5] ));
 sg13g2_dfrbp_1 _2113_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0252_),
    .D(net181),
    .Q_N(_0895_),
    .Q(\smul_up_counter.prob_counter[6] ));
 sg13g2_dfrbp_1 _2114_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0253_),
    .D(_0391_),
    .Q_N(_0894_),
    .Q(\smul_up_counter.prob_counter[7] ));
 sg13g2_dfrbp_1 _2115_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0254_),
    .D(net365),
    .Q_N(_0893_),
    .Q(\smul_up_counter.prob_counter[8] ));
 sg13g2_dfrbp_1 _2116_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0255_),
    .D(net380),
    .Q_N(_0892_),
    .Q(\smul_up_counter.prob_counter[9] ));
 sg13g2_dfrbp_1 _2117_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0256_),
    .D(net375),
    .Q_N(_0891_),
    .Q(\smul_up_counter.prob_counter[10] ));
 sg13g2_dfrbp_1 _2118_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0257_),
    .D(net357),
    .Q_N(_0890_),
    .Q(\smul_up_counter.prob_counter[11] ));
 sg13g2_dfrbp_1 _2119_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0258_),
    .D(net367),
    .Q_N(_0889_),
    .Q(\smul_up_counter.prob_counter[12] ));
 sg13g2_dfrbp_1 _2120_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0259_),
    .D(_0397_),
    .Q_N(_0888_),
    .Q(\smul_up_counter.prob_counter[13] ));
 sg13g2_dfrbp_1 _2121_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0260_),
    .D(_0398_),
    .Q_N(_0887_),
    .Q(\smul_up_counter.prob_counter[14] ));
 sg13g2_dfrbp_1 _2122_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0261_),
    .D(net359),
    .Q_N(_0886_),
    .Q(\smul_up_counter.prob_counter[15] ));
 sg13g2_dfrbp_1 _2123_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0262_),
    .D(net217),
    .Q_N(_0046_),
    .Q(\smul_up_counter.prob_counter[16] ));
 sg13g2_dfrbp_1 _2124_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net23),
    .D(net410),
    .Q_N(_0885_),
    .Q(\smul.SN_Bit_Q ));
 sg13g2_dfrbp_1 _2125_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0263_),
    .D(_0401_),
    .Q_N(_0884_),
    .Q(\mul_output.counter[0] ));
 sg13g2_dfrbp_1 _2126_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0264_),
    .D(_0402_),
    .Q_N(_0883_),
    .Q(\mul_output.counter[1] ));
 sg13g2_dfrbp_1 _2127_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0265_),
    .D(net211),
    .Q_N(_0882_),
    .Q(\mul_output.counter[2] ));
 sg13g2_dfrbp_1 _2128_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0266_),
    .D(_0404_),
    .Q_N(_0881_),
    .Q(\mul_output.counter[3] ));
 sg13g2_dfrbp_1 _2129_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0267_),
    .D(net81),
    .Q_N(_0880_),
    .Q(\mul_avg[0] ));
 sg13g2_dfrbp_1 _2130_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0268_),
    .D(net69),
    .Q_N(_0879_),
    .Q(\mul_avg[1] ));
 sg13g2_dfrbp_1 _2131_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0269_),
    .D(net73),
    .Q_N(_0878_),
    .Q(\mul_avg[2] ));
 sg13g2_dfrbp_1 _2132_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0270_),
    .D(net190),
    .Q_N(_0877_),
    .Q(\mul_avg[3] ));
 sg13g2_dfrbp_1 _2133_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0271_),
    .D(net83),
    .Q_N(_0876_),
    .Q(\mul_avg[4] ));
 sg13g2_dfrbp_1 _2134_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0272_),
    .D(net67),
    .Q_N(_0875_),
    .Q(\mul_avg[5] ));
 sg13g2_dfrbp_1 _2135_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0273_),
    .D(net146),
    .Q_N(_0874_),
    .Q(\mul_avg[6] ));
 sg13g2_dfrbp_1 _2136_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0274_),
    .D(net102),
    .Q_N(_0873_),
    .Q(\mul_avg[7] ));
 sg13g2_dfrbp_1 _2137_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0275_),
    .D(_0413_),
    .Q_N(_0872_),
    .Q(\mul_avg[8] ));
 sg13g2_dfrbp_1 _2138_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_0276_),
    .D(_0414_),
    .Q_N(_0871_),
    .Q(\add_output.counter[0] ));
 sg13g2_dfrbp_1 _2139_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0277_),
    .D(_0415_),
    .Q_N(_0870_),
    .Q(\add_output.counter[1] ));
 sg13g2_dfrbp_1 _2140_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0278_),
    .D(net215),
    .Q_N(_0869_),
    .Q(\add_output.counter[2] ));
 sg13g2_dfrbp_1 _2141_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0279_),
    .D(_0417_),
    .Q_N(_0868_),
    .Q(\add_output.counter[3] ));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_4 (.L_LO(net4));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_5 (.L_LO(net5));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_6 (.L_LO(net6));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_7 (.L_LO(net7));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_8 (.L_LO(net8));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_9 (.L_LO(net9));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_10 (.L_LO(net10));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_11 (.L_LO(net11));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_12 (.L_LO(net12));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_13 (.L_LO(net13));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_14 (.L_LO(net14));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_15 (.L_LO(net15));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_16 (.L_LO(net16));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_17 (.L_LO(net17));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_18 (.L_LO(net18));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_19 (.L_LO(net19));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_20 (.L_LO(net20));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_21 (.L_LO(net21));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_22 (.L_LO(net22));
 sg13g2_tiehi _2124__23 (.L_HI(net23));
 sg13g2_buf_2 _2163_ (.A(mul_bit_out),
    .X(uo_out[0]));
 sg13g2_buf_2 _2164_ (.A(add_bit_out),
    .X(uo_out[1]));
 sg13g2_buf_1 _2165_ (.A(smul_bit_out),
    .X(uo_out[2]));
 sg13g2_buf_1 _2166_ (.A(\add_up_counter.clk_counter[17] ),
    .X(uo_out[3]));
 sg13g2_buf_2 fanout265 (.A(net266),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_0446_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(net268),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_0838_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_0436_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net272),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_0434_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_0827_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_0709_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_0709_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_0708_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_0708_),
    .X(net279));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(net283));
 sg13g2_buf_2 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(net283),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_0773_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(net290),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(net290),
    .X(net285));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(net290));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net290),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_0657_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net293),
    .X(net291));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(net293));
 sg13g2_buf_2 fanout293 (.A(_0656_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_0431_),
    .X(net294));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(_0430_));
 sg13g2_buf_2 fanout296 (.A(_0671_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_0670_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_0647_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_0646_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net302),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301));
 sg13g2_buf_1 fanout302 (.A(_0489_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net305),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net305),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_0487_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net307),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_0429_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(net416),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net310));
 sg13g2_buf_4 fanout310 (.X(net310),
    .A(net312));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(net312));
 sg13g2_buf_2 fanout312 (.A(net177),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(net321),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(net321),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net321),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net320),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_1 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(net349),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(net323),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(net329),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net328),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_1 fanout329 (.A(net349),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(net339),
    .X(net330));
 sg13g2_buf_1 fanout331 (.A(net339),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(net339),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(net335),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(net338),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net338),
    .X(net336));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(net338));
 sg13g2_buf_1 fanout338 (.A(net339),
    .X(net338));
 sg13g2_buf_1 fanout339 (.A(net349),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(net343),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net343),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net349),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(net348),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(net347),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_1 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(rst_n),
    .X(net349));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_stochastic_addmultiply_CL123abc_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_22_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_6_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0922_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold2 (.A(\global_SN_gen.lfsr[11] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0915_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0920_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0921_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold6 (.A(\global_SN_gen.lfsr[9] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold7 (.A(\global_SN_gen.lfsr[10] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold8 (.A(\global_SN_gen.lfsr[28] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold9 (.A(\global_SN_gen.lfsr[23] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold10 (.A(\global_SN_gen.lfsr[6] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold11 (.A(\global_SN_gen.lfsr[4] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold12 (.A(\global_SN_gen.lfsr[25] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold13 (.A(\global_SN_gen.lfsr[29] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold14 (.A(\global_SN_gen.lfsr[24] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold15 (.A(\global_SN_gen.lfsr[21] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold16 (.A(\global_SN_gen.lfsr[22] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold17 (.A(\global_SN_gen.lfsr[26] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold18 (.A(\global_SN_gen.lfsr[0] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold19 (.A(\global_SN_gen.lfsr[1] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold20 (.A(\global_SN_gen.lfsr[27] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold21 (.A(\global_SN_gen.lfsr[12] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold22 (.A(\global_SN_gen.lfsr[14] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold23 (.A(\global_SN_gen.lfsr[18] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold24 (.A(\global_SN_gen.lfsr[2] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold25 (.A(\global_SN_gen.lfsr[19] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold26 (.A(\global_SN_gen.lfsr[8] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold27 (.A(\global_SN_gen.lfsr[17] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold28 (.A(\global_SN_gen.lfsr[13] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mul_output.bitseq[8] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0036_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold31 (.A(\global_SN_gen.lfsr[30] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mul_output.bitseq[3] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0030_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold34 (.A(\global_SN_gen.lfsr[15] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold35 (.A(\add_output.bitseq[8] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold36 (.A(\smul_output.bitseq[8] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold37 (.A(\smul_avg[1] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0294_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold39 (.A(\smul_avg[2] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0295_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold41 (.A(\smul_avg[6] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0299_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mul_avg[5] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0410_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mul_avg[1] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0406_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold47 (.A(\smul_avg[8] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0301_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mul_avg[2] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0407_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold51 (.A(\smul_avg[4] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0297_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold53 (.A(\smul_avg[7] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0300_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold55 (.A(\smul_avg[5] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0298_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mul_avg[0] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0405_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mul_avg[4] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0409_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold61 (.A(\add_up_counter.prob_counter[16] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0352_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mul_output.bitseq[4] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold64 (.A(\smul_avg[0] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0293_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mul_output.bitseq[2] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0029_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mul_output.bitseq[7] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0034_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mul_output.bitseq[6] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0033_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold72 (.A(\add_output.bitseq[3] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0020_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold74 (.A(\add_output.bitseq[1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0018_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold76 (.A(\add_output.bitseq[7] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0024_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mul_avg[7] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0412_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mul_output.bitseq[0] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold81 (.A(\smul_output.bitseq[0] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold82 (.A(\add_avg[0] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0308_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold84 (.A(\global_input.output_bitcounter_1[3] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0330_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold86 (.A(\add_output.bitseq[2] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0019_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold88 (.A(\global_input.output_bitcounter_1[6] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0380_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold90 (.A(\smul_output.bitseq[7] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0043_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold92 (.A(\add_output.counter[0] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mul_output.bitseq[1] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold94 (.A(\global_input.adjustment[1] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0303_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold96 (.A(\add_output.bitseq[4] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0021_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold98 (.A(\global_SN_gen.lfsr[20] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold99 (.A(\smul_avg[3] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0296_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mul_output.counter[0] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold102 (.A(\add_avg[8] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold103 (.A(\smul_output.bitseq[6] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0042_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold105 (.A(\add_output.bitseq[6] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0023_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold107 (.A(\smul_output.bitseq[2] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0038_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mul_avg[8] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0050_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0305_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mul_up_counter.prob_counter[16] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold113 (.A(\add_up_counter.prob_counter[8] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold114 (.A(\smul_output.bitseq[1] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold115 (.A(\global_input.output_bitcounter_2[3] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0356_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold117 (.A(\add_up_counter.prob_counter[2] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0338_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold119 (.A(\smul_output.counter[3] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0430_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold121 (.A(net295),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mul_avg[6] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0411_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold124 (.A(\smul_output.bitseq[4] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0040_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0049_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0302_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold128 (.A(\add_up_counter.prob_counter[3] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold129 (.A(\smul_output.counter[0] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold130 (.A(\global_input.output_bitcounter_2[0] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0362_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold132 (.A(\global_SN_gen.Input_2[7] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0360_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold134 (.A(\smul_output.bitseq[5] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold135 (.A(\global_input.output_bitcounter_2[8] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0361_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold137 (.A(\global_input.adjustment[4] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0306_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold139 (.A(\global_input.output_bitcounter_2[1] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0354_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold141 (.A(\add_output.bitseq[5] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0546_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0022_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold144 (.A(\global_input.output_bitcounter_2[4] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0357_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold146 (.A(\global_input.output_bitcounter_2[2] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold147 (.A(\global_input.output_bitcounter_1[2] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold148 (.A(\global_input.output_bitcounter_1[1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0375_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold150 (.A(\global_input.output_bitcounter_2[5] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0358_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold152 (.A(\global_input.output_bitcounter_2[6] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0359_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold154 (.A(\global_input.loop ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold155 (.A(\global_SN_gen.Input_1[2] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold156 (.A(\global_SN_gen.Input_2[2] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold157 (.A(\smul_up_counter.prob_counter[6] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0390_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold159 (.A(\add_up_counter.prob_counter[6] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0342_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold161 (.A(\global_SN_gen.Input_2[0] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold162 (.A(\global_SN_gen.Input_1[1] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold163 (.A(\global_input.output_bitcounter_1[7] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0334_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold165 (.A(\global_input.output_bitcounter_2[7] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mul_avg[3] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0408_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold168 (.A(\global_input.output_bitcounter_1[8] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0335_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold170 (.A(\add_up_counter.prob_counter[9] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold171 (.A(\add_up_counter.clk_counter[10] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0001_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold173 (.A(\add_avg[1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold174 (.A(\add_up_counter.prob_counter[11] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0347_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold176 (.A(\smul_output.bitseq[3] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0039_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold178 (.A(\add_up_counter.prob_counter[15] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0287_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold180 (.A(\add_up_counter.clk_counter[7] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0015_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold182 (.A(\global_SN_gen.Input_1[6] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold183 (.A(\add_up_counter.clk_counter[13] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0004_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold185 (.A(\add_up_counter.prob_counter[5] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0341_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mul_output.counter[2] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0403_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold189 (.A(\global_input.output_bitcounter_1[0] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0327_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold191 (.A(\add_output.counter[2] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0416_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold193 (.A(\smul_up_counter.prob_counter[16] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0400_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold195 (.A(\global_input.output_bitcounter_1[4] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold196 (.A(\add_up_counter.prob_counter[14] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0350_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold198 (.A(\add_up_counter.prob_counter[15] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold199 (.A(\add_avg[2] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0282_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold201 (.A(\add_up_counter.prob_counter[13] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0349_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold203 (.A(\add_up_counter.clk_counter[6] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0014_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold205 (.A(\add_avg[3] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold206 (.A(\smul_up_counter.prob_counter[4] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold207 (.A(\add_avg[4] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0284_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold209 (.A(\add_avg[5] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold210 (.A(\mul_output.bitseq[5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0530_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold212 (.A(\global_input.output_bitcounter_1[5] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold213 (.A(\add_up_counter.clk_counter[15] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0583_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0006_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold216 (.A(\add_up_counter.prob_counter[7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold217 (.A(\add_up_counter.prob_counter[12] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold218 (.A(\add_up_counter.clk_counter[16] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0007_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold220 (.A(\add_up_counter.prob_counter[4] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold221 (.A(\smul_up_counter.prob_counter[3] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0387_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold223 (.A(\add_avg[6] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold224 (.A(\add_up_counter.prob_counter[7] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold225 (.A(\smul_up_counter.prob_counter[0] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold226 (.A(\add_output.counter[1] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold227 (.A(\global_input.adjustment[2] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0304_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold229 (.A(\global_input.output_case[2] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0373_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold231 (.A(\smul_output.counter[2] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0291_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold233 (.A(\add_up_counter.prob_counter[10] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0346_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold235 (.A(\add_up_counter.clk_counter[11] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0002_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold237 (.A(\global_SN_gen.Input_1[4] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold238 (.A(\add_up_counter.prob_counter[1] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0337_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold240 (.A(\mul_output.counter[1] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold241 (.A(\smul_up_counter.prob_counter[2] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0386_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold243 (.A(\add_up_counter.clk_counter[8] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0016_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold245 (.A(\add_up_counter.clk_counter[14] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0005_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold247 (.A(\smul_up_counter.prob_counter[1] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold248 (.A(\smul_up_counter.prob_counter[11] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0395_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold250 (.A(\smul_up_counter.prob_counter[15] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0399_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold252 (.A(\smul_up_counter.prob_counter[5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold253 (.A(\add_up_counter.clk_counter[3] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0011_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold255 (.A(\global_SN_gen.Input_1[5] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold256 (.A(\smul_up_counter.prob_counter[8] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0392_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold258 (.A(\smul_up_counter.prob_counter[12] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0396_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0047_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold261 (.A(\add_output.counter[3] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold262 (.A(\smul_up_counter.prob_counter[13] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold263 (.A(\add_up_counter.prob_counter[0] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold264 (.A(\add_up_counter.clk_counter[0] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mul_output.counter[3] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold266 (.A(\smul_up_counter.prob_counter[10] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0394_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold268 (.A(\add_up_counter.clk_counter[1] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold269 (.A(\smul_up_counter.prob_counter[14] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold270 (.A(\add_up_counter.clk_counter[17] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold271 (.A(\smul_up_counter.prob_counter[9] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0393_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold273 (.A(\smul_output.counter[1] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold274 (.A(\mul_up_counter.prob_counter[0] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold275 (.A(\add_up_counter.clk_counter[4] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0012_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold277 (.A(\mul_up_counter.prob_counter[5] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0314_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold279 (.A(\mul_up_counter.prob_counter[6] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0315_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold281 (.A(\mul_up_counter.prob_counter[2] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold282 (.A(\mul_up_counter.prob_counter[15] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0452_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold284 (.A(\add_up_counter.clk_counter[9] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold285 (.A(\mul_up_counter.prob_counter[11] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0462_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold287 (.A(\mul_up_counter.prob_counter[3] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0312_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold289 (.A(\mul_up_counter.prob_counter[8] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold290 (.A(\mul_up_counter.prob_counter[13] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0322_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold292 (.A(\add_up_counter.clk_counter[5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0013_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold294 (.A(\mul_up_counter.prob_counter[7] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold295 (.A(\global_input.output_case[3] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold296 (.A(\mul_up_counter.prob_counter[9] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold297 (.A(\add_up_counter.clk_counter[12] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold298 (.A(\smul_up_counter.prob_counter[7] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold299 (.A(\mul_up_counter.prob_counter[1] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold300 (.A(\mul_up_counter.prob_counter[4] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold301 (.A(\global_SN_gen.Input_1[8] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold302 (.A(SN_Bit_1),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold303 (.A(\add_up_counter.clk_counter[2] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold304 (.A(\mul_up_counter.prob_counter[12] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold305 (.A(\mul_up_counter.prob_counter[14] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold306 (.A(\mul_up_counter.prob_counter[10] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold307 (.A(\global_input.output_case[1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold308 (.A(\global_input.output_case[0] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold309 (.A(\add_up_counter.prob_counter[10] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold310 (.A(\add_up_counter.prob_counter[4] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold311 (.A(\add_up_counter.prob_counter[1] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold312 (.A(\mul_output.counter[3] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0670_),
    .X(net421));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_4 FILLER_20_217 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_285 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_327 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_decap_4 FILLER_21_191 ();
 sg13g2_fill_2 FILLER_21_195 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_4 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_172 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_decap_8 FILLER_23_313 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_8 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_4 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_217 ();
 sg13g2_fill_1 FILLER_25_226 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_decap_8 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_302 ();
 sg13g2_decap_8 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_316 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_4 FILLER_26_168 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_158 ();
 sg13g2_fill_1 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_300 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_decap_8 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_fill_2 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_314 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_211 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_fill_2 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_142 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_334 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_decap_8 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_decap_4 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_decap_8 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_223 ();
 sg13g2_decap_4 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_356 ();
 sg13g2_decap_8 FILLER_33_363 ();
 sg13g2_decap_8 FILLER_33_370 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_decap_4 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_170 ();
 sg13g2_fill_2 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_4 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_116 ();
 sg13g2_fill_2 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_4 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_fill_2 FILLER_38_119 ();
 sg13g2_fill_1 FILLER_38_121 ();
 sg13g2_fill_1 FILLER_38_174 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_fill_2 FILLER_38_214 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_4 FILLER_39_98 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_decap_8 FILLER_39_178 ();
 sg13g2_fill_1 FILLER_39_185 ();
 sg13g2_fill_2 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_226 ();
 sg13g2_decap_8 FILLER_39_233 ();
 sg13g2_decap_8 FILLER_39_326 ();
 sg13g2_decap_8 FILLER_39_333 ();
 sg13g2_decap_8 FILLER_39_340 ();
 sg13g2_decap_8 FILLER_39_347 ();
 sg13g2_fill_1 FILLER_39_354 ();
 sg13g2_decap_8 FILLER_39_358 ();
 sg13g2_decap_8 FILLER_39_365 ();
 sg13g2_decap_8 FILLER_39_372 ();
 sg13g2_decap_8 FILLER_39_379 ();
 sg13g2_decap_8 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_39_400 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_4 FILLER_40_98 ();
 sg13g2_fill_1 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_129 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_fill_1 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_181 ();
 sg13g2_decap_4 FILLER_40_231 ();
 sg13g2_fill_1 FILLER_40_255 ();
 sg13g2_fill_1 FILLER_40_291 ();
 sg13g2_decap_8 FILLER_40_370 ();
 sg13g2_decap_8 FILLER_40_377 ();
 sg13g2_decap_8 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_398 ();
 sg13g2_decap_4 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_fill_2 FILLER_41_98 ();
 sg13g2_fill_1 FILLER_41_100 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_fill_1 FILLER_41_149 ();
 sg13g2_fill_2 FILLER_41_159 ();
 sg13g2_fill_1 FILLER_41_202 ();
 sg13g2_fill_1 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_242 ();
 sg13g2_fill_1 FILLER_41_258 ();
 sg13g2_decap_4 FILLER_41_264 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_272 ();
 sg13g2_fill_1 FILLER_41_278 ();
 sg13g2_fill_2 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_4 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_102 ();
 sg13g2_fill_1 FILLER_42_155 ();
 sg13g2_decap_8 FILLER_42_222 ();
 sg13g2_decap_8 FILLER_42_229 ();
 sg13g2_fill_1 FILLER_42_248 ();
 sg13g2_fill_2 FILLER_42_356 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_4 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_fill_2 FILLER_43_98 ();
 sg13g2_fill_1 FILLER_43_100 ();
 sg13g2_fill_2 FILLER_43_125 ();
 sg13g2_fill_1 FILLER_43_127 ();
 sg13g2_fill_2 FILLER_43_137 ();
 sg13g2_fill_1 FILLER_43_139 ();
 sg13g2_fill_1 FILLER_43_149 ();
 sg13g2_decap_8 FILLER_43_213 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_4 FILLER_43_231 ();
 sg13g2_fill_1 FILLER_43_235 ();
 sg13g2_fill_2 FILLER_43_239 ();
 sg13g2_fill_1 FILLER_43_270 ();
 sg13g2_fill_2 FILLER_43_280 ();
 sg13g2_fill_1 FILLER_43_282 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_390 ();
 sg13g2_fill_2 FILLER_43_397 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_fill_1 FILLER_44_98 ();
 sg13g2_fill_1 FILLER_44_135 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_fill_2 FILLER_44_211 ();
 sg13g2_fill_1 FILLER_44_213 ();
 sg13g2_fill_1 FILLER_44_249 ();
 sg13g2_fill_2 FILLER_44_264 ();
 sg13g2_fill_2 FILLER_44_279 ();
 sg13g2_fill_1 FILLER_44_281 ();
 sg13g2_decap_8 FILLER_44_321 ();
 sg13g2_fill_2 FILLER_44_328 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_4 FILLER_45_91 ();
 sg13g2_fill_1 FILLER_45_95 ();
 sg13g2_fill_1 FILLER_45_156 ();
 sg13g2_fill_1 FILLER_45_183 ();
 sg13g2_decap_8 FILLER_45_225 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_fill_1 FILLER_45_358 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_124 ();
 sg13g2_fill_2 FILLER_46_135 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_fill_1 FILLER_46_234 ();
 sg13g2_decap_8 FILLER_46_283 ();
 sg13g2_decap_8 FILLER_46_290 ();
 sg13g2_fill_2 FILLER_46_302 ();
 sg13g2_fill_2 FILLER_46_330 ();
 sg13g2_fill_2 FILLER_46_361 ();
 sg13g2_fill_1 FILLER_46_363 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_4 FILLER_47_98 ();
 sg13g2_fill_2 FILLER_47_102 ();
 sg13g2_fill_1 FILLER_47_119 ();
 sg13g2_fill_2 FILLER_47_146 ();
 sg13g2_fill_2 FILLER_47_163 ();
 sg13g2_fill_2 FILLER_47_174 ();
 sg13g2_fill_2 FILLER_47_202 ();
 sg13g2_fill_2 FILLER_47_267 ();
 sg13g2_decap_4 FILLER_47_298 ();
 sg13g2_fill_2 FILLER_47_321 ();
 sg13g2_decap_4 FILLER_47_359 ();
 sg13g2_decap_8 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_47_388 ();
 sg13g2_decap_8 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_4 FILLER_48_98 ();
 sg13g2_fill_2 FILLER_48_102 ();
 sg13g2_fill_2 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_fill_2 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_212 ();
 sg13g2_decap_4 FILLER_48_219 ();
 sg13g2_fill_1 FILLER_48_223 ();
 sg13g2_decap_4 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_231 ();
 sg13g2_fill_2 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_316 ();
 sg13g2_fill_2 FILLER_48_357 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_98 ();
 sg13g2_fill_1 FILLER_49_126 ();
 sg13g2_decap_4 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_174 ();
 sg13g2_fill_2 FILLER_49_189 ();
 sg13g2_fill_2 FILLER_49_205 ();
 sg13g2_decap_8 FILLER_49_215 ();
 sg13g2_decap_8 FILLER_49_222 ();
 sg13g2_decap_8 FILLER_49_229 ();
 sg13g2_fill_1 FILLER_49_236 ();
 sg13g2_fill_1 FILLER_49_248 ();
 sg13g2_fill_1 FILLER_49_318 ();
 sg13g2_decap_4 FILLER_49_325 ();
 sg13g2_fill_2 FILLER_49_341 ();
 sg13g2_decap_4 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_fill_2 FILLER_50_98 ();
 sg13g2_fill_2 FILLER_50_148 ();
 sg13g2_decap_4 FILLER_50_159 ();
 sg13g2_fill_1 FILLER_50_163 ();
 sg13g2_decap_8 FILLER_50_229 ();
 sg13g2_decap_8 FILLER_50_236 ();
 sg13g2_decap_8 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_4 FILLER_51_105 ();
 sg13g2_fill_1 FILLER_51_109 ();
 sg13g2_fill_2 FILLER_51_115 ();
 sg13g2_fill_2 FILLER_51_126 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_decap_4 FILLER_51_142 ();
 sg13g2_fill_2 FILLER_51_236 ();
 sg13g2_fill_1 FILLER_51_238 ();
 sg13g2_fill_2 FILLER_51_279 ();
 sg13g2_fill_2 FILLER_51_285 ();
 sg13g2_fill_1 FILLER_51_287 ();
 sg13g2_fill_1 FILLER_51_300 ();
 sg13g2_decap_8 FILLER_51_316 ();
 sg13g2_fill_2 FILLER_51_332 ();
 sg13g2_fill_1 FILLER_51_334 ();
 sg13g2_decap_4 FILLER_51_343 ();
 sg13g2_fill_2 FILLER_51_347 ();
 sg13g2_fill_2 FILLER_51_352 ();
 sg13g2_fill_2 FILLER_51_363 ();
 sg13g2_fill_1 FILLER_51_365 ();
 sg13g2_fill_2 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_4 FILLER_52_112 ();
 sg13g2_fill_1 FILLER_52_116 ();
 sg13g2_decap_8 FILLER_52_129 ();
 sg13g2_fill_2 FILLER_52_136 ();
 sg13g2_fill_1 FILLER_52_138 ();
 sg13g2_fill_2 FILLER_52_180 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_fill_2 FILLER_52_211 ();
 sg13g2_decap_8 FILLER_52_246 ();
 sg13g2_fill_1 FILLER_52_261 ();
 sg13g2_fill_1 FILLER_52_268 ();
 sg13g2_decap_4 FILLER_52_272 ();
 sg13g2_fill_1 FILLER_52_311 ();
 sg13g2_decap_8 FILLER_52_320 ();
 sg13g2_fill_2 FILLER_52_356 ();
 sg13g2_fill_1 FILLER_52_358 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_fill_1 FILLER_53_133 ();
 sg13g2_fill_1 FILLER_53_142 ();
 sg13g2_fill_2 FILLER_53_195 ();
 sg13g2_fill_1 FILLER_53_217 ();
 sg13g2_fill_2 FILLER_53_253 ();
 sg13g2_fill_1 FILLER_53_260 ();
 sg13g2_decap_4 FILLER_53_266 ();
 sg13g2_decap_4 FILLER_53_379 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_fill_2 FILLER_54_119 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_fill_2 FILLER_54_180 ();
 sg13g2_fill_1 FILLER_54_191 ();
 sg13g2_fill_2 FILLER_54_219 ();
 sg13g2_decap_4 FILLER_54_246 ();
 sg13g2_fill_2 FILLER_54_250 ();
 sg13g2_fill_1 FILLER_54_321 ();
 sg13g2_fill_2 FILLER_54_344 ();
 sg13g2_fill_1 FILLER_54_370 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_4 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_123 ();
 sg13g2_decap_8 FILLER_55_268 ();
 sg13g2_fill_2 FILLER_55_292 ();
 sg13g2_fill_1 FILLER_55_303 ();
 sg13g2_decap_4 FILLER_55_343 ();
 sg13g2_fill_2 FILLER_55_355 ();
 sg13g2_fill_1 FILLER_55_357 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_fill_2 FILLER_56_119 ();
 sg13g2_fill_2 FILLER_56_147 ();
 sg13g2_fill_1 FILLER_56_200 ();
 sg13g2_fill_1 FILLER_56_229 ();
 sg13g2_fill_2 FILLER_56_233 ();
 sg13g2_fill_1 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_266 ();
 sg13g2_decap_8 FILLER_56_273 ();
 sg13g2_decap_4 FILLER_56_280 ();
 sg13g2_decap_4 FILLER_56_323 ();
 sg13g2_fill_2 FILLER_56_357 ();
 sg13g2_fill_1 FILLER_56_359 ();
 sg13g2_decap_8 FILLER_56_397 ();
 sg13g2_decap_4 FILLER_56_404 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_fill_1 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_159 ();
 sg13g2_fill_2 FILLER_57_200 ();
 sg13g2_decap_4 FILLER_57_264 ();
 sg13g2_fill_2 FILLER_57_281 ();
 sg13g2_fill_1 FILLER_57_293 ();
 sg13g2_fill_2 FILLER_57_303 ();
 sg13g2_fill_1 FILLER_57_305 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_fill_2 FILLER_57_337 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_4 FILLER_58_112 ();
 sg13g2_fill_2 FILLER_58_116 ();
 sg13g2_fill_2 FILLER_58_300 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_fill_2 FILLER_58_341 ();
 sg13g2_fill_1 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_fill_2 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_145 ();
 sg13g2_fill_2 FILLER_59_182 ();
 sg13g2_fill_2 FILLER_59_193 ();
 sg13g2_fill_1 FILLER_59_207 ();
 sg13g2_fill_2 FILLER_59_222 ();
 sg13g2_fill_2 FILLER_59_236 ();
 sg13g2_fill_1 FILLER_59_238 ();
 sg13g2_fill_1 FILLER_59_267 ();
 sg13g2_fill_1 FILLER_59_285 ();
 sg13g2_fill_2 FILLER_59_324 ();
 sg13g2_decap_8 FILLER_59_340 ();
 sg13g2_fill_1 FILLER_59_376 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_fill_2 FILLER_60_126 ();
 sg13g2_fill_1 FILLER_60_128 ();
 sg13g2_fill_2 FILLER_60_132 ();
 sg13g2_fill_1 FILLER_60_134 ();
 sg13g2_decap_4 FILLER_60_140 ();
 sg13g2_fill_2 FILLER_60_148 ();
 sg13g2_decap_4 FILLER_60_173 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_1 FILLER_60_182 ();
 sg13g2_fill_1 FILLER_60_195 ();
 sg13g2_fill_1 FILLER_60_208 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_fill_1 FILLER_60_238 ();
 sg13g2_fill_2 FILLER_60_250 ();
 sg13g2_fill_2 FILLER_60_283 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_fill_1 FILLER_61_119 ();
 sg13g2_fill_1 FILLER_61_146 ();
 sg13g2_fill_2 FILLER_61_152 ();
 sg13g2_fill_1 FILLER_61_154 ();
 sg13g2_fill_1 FILLER_61_158 ();
 sg13g2_fill_2 FILLER_61_178 ();
 sg13g2_fill_1 FILLER_61_226 ();
 sg13g2_fill_1 FILLER_61_244 ();
 sg13g2_fill_1 FILLER_61_282 ();
 sg13g2_fill_1 FILLER_61_312 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_4 FILLER_62_126 ();
 sg13g2_fill_1 FILLER_62_130 ();
 sg13g2_fill_1 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_299 ();
 sg13g2_fill_1 FILLER_62_392 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_4 FILLER_63_126 ();
 sg13g2_fill_2 FILLER_63_130 ();
 sg13g2_fill_1 FILLER_63_179 ();
 sg13g2_fill_1 FILLER_63_292 ();
 sg13g2_fill_1 FILLER_63_302 ();
 sg13g2_fill_1 FILLER_63_372 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_4 FILLER_64_119 ();
 sg13g2_fill_1 FILLER_64_158 ();
 sg13g2_fill_1 FILLER_64_211 ();
 sg13g2_fill_1 FILLER_64_225 ();
 sg13g2_fill_2 FILLER_64_272 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_fill_1 FILLER_64_323 ();
 sg13g2_fill_1 FILLER_64_340 ();
 sg13g2_fill_1 FILLER_64_353 ();
 sg13g2_fill_1 FILLER_64_369 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_4 FILLER_65_119 ();
 sg13g2_fill_1 FILLER_65_123 ();
 sg13g2_fill_1 FILLER_65_171 ();
 sg13g2_fill_1 FILLER_65_205 ();
 sg13g2_fill_1 FILLER_65_210 ();
 sg13g2_fill_1 FILLER_65_219 ();
 sg13g2_fill_2 FILLER_65_228 ();
 sg13g2_fill_2 FILLER_65_245 ();
 sg13g2_fill_1 FILLER_65_286 ();
 sg13g2_decap_8 FILLER_65_316 ();
 sg13g2_decap_8 FILLER_65_323 ();
 sg13g2_decap_4 FILLER_65_330 ();
 sg13g2_fill_1 FILLER_65_334 ();
 sg13g2_fill_2 FILLER_65_340 ();
 sg13g2_decap_4 FILLER_65_356 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_4 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_166 ();
 sg13g2_fill_1 FILLER_66_233 ();
 sg13g2_fill_2 FILLER_66_254 ();
 sg13g2_fill_1 FILLER_66_296 ();
 sg13g2_decap_4 FILLER_66_323 ();
 sg13g2_fill_1 FILLER_66_327 ();
 sg13g2_fill_2 FILLER_66_338 ();
 sg13g2_fill_1 FILLER_66_340 ();
 sg13g2_decap_4 FILLER_66_344 ();
 sg13g2_fill_2 FILLER_66_348 ();
 sg13g2_fill_2 FILLER_66_365 ();
 sg13g2_fill_2 FILLER_66_396 ();
 sg13g2_fill_1 FILLER_66_398 ();
 sg13g2_decap_8 FILLER_66_402 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_4 FILLER_67_119 ();
 sg13g2_fill_1 FILLER_67_161 ();
 sg13g2_fill_1 FILLER_67_167 ();
 sg13g2_fill_1 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_258 ();
 sg13g2_fill_1 FILLER_67_317 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_fill_2 FILLER_68_197 ();
 sg13g2_fill_2 FILLER_68_227 ();
 sg13g2_fill_1 FILLER_68_297 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_4 FILLER_69_133 ();
 sg13g2_fill_1 FILLER_69_137 ();
 sg13g2_fill_1 FILLER_69_148 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_fill_1 FILLER_69_231 ();
 sg13g2_fill_1 FILLER_69_246 ();
 sg13g2_fill_2 FILLER_69_361 ();
 sg13g2_fill_2 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_fill_1 FILLER_70_258 ();
 sg13g2_fill_1 FILLER_70_305 ();
 sg13g2_fill_1 FILLER_70_351 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_decap_8 FILLER_70_397 ();
 sg13g2_decap_4 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_4 FILLER_71_147 ();
 sg13g2_fill_1 FILLER_71_184 ();
 sg13g2_fill_2 FILLER_71_228 ();
 sg13g2_fill_2 FILLER_71_261 ();
 sg13g2_fill_1 FILLER_71_273 ();
 sg13g2_fill_2 FILLER_71_297 ();
 sg13g2_fill_1 FILLER_71_356 ();
 sg13g2_fill_1 FILLER_71_368 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_fill_2 FILLER_72_161 ();
 sg13g2_fill_1 FILLER_72_284 ();
 sg13g2_fill_1 FILLER_72_337 ();
 sg13g2_fill_1 FILLER_72_369 ();
 sg13g2_decap_4 FILLER_72_385 ();
 sg13g2_fill_1 FILLER_72_389 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_fill_2 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_fill_2 FILLER_73_168 ();
 sg13g2_fill_1 FILLER_73_170 ();
 sg13g2_fill_1 FILLER_73_206 ();
 sg13g2_fill_1 FILLER_73_373 ();
 sg13g2_decap_8 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_fill_2 FILLER_74_175 ();
 sg13g2_fill_1 FILLER_74_177 ();
 sg13g2_fill_2 FILLER_74_195 ();
 sg13g2_fill_2 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_218 ();
 sg13g2_fill_1 FILLER_74_226 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_277 ();
 sg13g2_fill_1 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_298 ();
 sg13g2_fill_2 FILLER_74_316 ();
 sg13g2_fill_1 FILLER_74_318 ();
 sg13g2_fill_1 FILLER_74_352 ();
 sg13g2_decap_4 FILLER_74_405 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_4 FILLER_75_175 ();
 sg13g2_fill_2 FILLER_75_202 ();
 sg13g2_fill_1 FILLER_75_204 ();
 sg13g2_fill_1 FILLER_75_222 ();
 sg13g2_fill_1 FILLER_75_226 ();
 sg13g2_decap_8 FILLER_75_264 ();
 sg13g2_fill_2 FILLER_75_290 ();
 sg13g2_fill_1 FILLER_75_292 ();
 sg13g2_fill_1 FILLER_75_301 ();
 sg13g2_fill_2 FILLER_75_323 ();
 sg13g2_decap_4 FILLER_75_334 ();
 sg13g2_fill_1 FILLER_75_338 ();
 sg13g2_decap_8 FILLER_75_342 ();
 sg13g2_decap_4 FILLER_75_349 ();
 sg13g2_fill_1 FILLER_75_369 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_4 FILLER_76_168 ();
 sg13g2_fill_1 FILLER_76_172 ();
 sg13g2_fill_1 FILLER_76_280 ();
 sg13g2_fill_1 FILLER_76_375 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_4 FILLER_77_161 ();
 sg13g2_fill_2 FILLER_77_165 ();
 sg13g2_fill_2 FILLER_77_214 ();
 sg13g2_fill_1 FILLER_77_242 ();
 sg13g2_fill_1 FILLER_77_258 ();
 sg13g2_fill_1 FILLER_77_300 ();
 sg13g2_fill_2 FILLER_77_323 ();
 sg13g2_fill_1 FILLER_77_371 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_4 FILLER_78_161 ();
 sg13g2_fill_1 FILLER_78_165 ();
 sg13g2_fill_1 FILLER_78_287 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_fill_1 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_390 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_fill_2 FILLER_79_168 ();
 sg13g2_fill_1 FILLER_79_170 ();
 sg13g2_decap_8 FILLER_79_214 ();
 sg13g2_decap_4 FILLER_79_221 ();
 sg13g2_fill_2 FILLER_79_286 ();
 sg13g2_fill_1 FILLER_79_288 ();
 sg13g2_fill_2 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_8 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_fill_2 FILLER_80_172 ();
 sg13g2_fill_1 FILLER_80_174 ();
 sg13g2_decap_8 FILLER_80_214 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_fill_2 FILLER_80_228 ();
 sg13g2_fill_2 FILLER_80_242 ();
 sg13g2_fill_1 FILLER_80_262 ();
 sg13g2_fill_1 FILLER_80_278 ();
 sg13g2_decap_4 FILLER_80_327 ();
 sg13g2_fill_2 FILLER_80_331 ();
 sg13g2_decap_8 FILLER_80_343 ();
 sg13g2_fill_2 FILLER_80_350 ();
 sg13g2_fill_1 FILLER_80_352 ();
 sg13g2_fill_2 FILLER_80_356 ();
 sg13g2_fill_1 FILLER_80_358 ();
 sg13g2_decap_8 FILLER_80_376 ();
 sg13g2_decap_8 FILLER_80_383 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_decap_4 FILLER_80_404 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
 assign uo_out[4] = net19;
 assign uo_out[5] = net20;
 assign uo_out[6] = net21;
 assign uo_out[7] = net22;
endmodule

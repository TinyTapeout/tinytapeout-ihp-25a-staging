module tt_um_histogramming (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire \bin_array[0][0] ;
 wire \bin_array[0][1] ;
 wire \bin_array[0][2] ;
 wire \bin_array[0][3] ;
 wire \bin_array[10][0] ;
 wire \bin_array[10][1] ;
 wire \bin_array[10][2] ;
 wire \bin_array[10][3] ;
 wire \bin_array[11][0] ;
 wire \bin_array[11][1] ;
 wire \bin_array[11][2] ;
 wire \bin_array[11][3] ;
 wire \bin_array[12][0] ;
 wire \bin_array[12][1] ;
 wire \bin_array[12][2] ;
 wire \bin_array[12][3] ;
 wire \bin_array[13][0] ;
 wire \bin_array[13][1] ;
 wire \bin_array[13][2] ;
 wire \bin_array[13][3] ;
 wire \bin_array[14][0] ;
 wire \bin_array[14][1] ;
 wire \bin_array[14][2] ;
 wire \bin_array[14][3] ;
 wire \bin_array[15][0] ;
 wire \bin_array[15][1] ;
 wire \bin_array[15][2] ;
 wire \bin_array[15][3] ;
 wire \bin_array[16][0] ;
 wire \bin_array[16][1] ;
 wire \bin_array[16][2] ;
 wire \bin_array[16][3] ;
 wire \bin_array[17][0] ;
 wire \bin_array[17][1] ;
 wire \bin_array[17][2] ;
 wire \bin_array[17][3] ;
 wire \bin_array[18][0] ;
 wire \bin_array[18][1] ;
 wire \bin_array[18][2] ;
 wire \bin_array[18][3] ;
 wire \bin_array[19][0] ;
 wire \bin_array[19][1] ;
 wire \bin_array[19][2] ;
 wire \bin_array[19][3] ;
 wire \bin_array[1][0] ;
 wire \bin_array[1][1] ;
 wire \bin_array[1][2] ;
 wire \bin_array[1][3] ;
 wire \bin_array[20][0] ;
 wire \bin_array[20][1] ;
 wire \bin_array[20][2] ;
 wire \bin_array[20][3] ;
 wire \bin_array[21][0] ;
 wire \bin_array[21][1] ;
 wire \bin_array[21][2] ;
 wire \bin_array[21][3] ;
 wire \bin_array[22][0] ;
 wire \bin_array[22][1] ;
 wire \bin_array[22][2] ;
 wire \bin_array[22][3] ;
 wire \bin_array[23][0] ;
 wire \bin_array[23][1] ;
 wire \bin_array[23][2] ;
 wire \bin_array[23][3] ;
 wire \bin_array[24][0] ;
 wire \bin_array[24][1] ;
 wire \bin_array[24][2] ;
 wire \bin_array[24][3] ;
 wire \bin_array[25][0] ;
 wire \bin_array[25][1] ;
 wire \bin_array[25][2] ;
 wire \bin_array[25][3] ;
 wire \bin_array[26][0] ;
 wire \bin_array[26][1] ;
 wire \bin_array[26][2] ;
 wire \bin_array[26][3] ;
 wire \bin_array[27][0] ;
 wire \bin_array[27][1] ;
 wire \bin_array[27][2] ;
 wire \bin_array[27][3] ;
 wire \bin_array[28][0] ;
 wire \bin_array[28][1] ;
 wire \bin_array[28][2] ;
 wire \bin_array[28][3] ;
 wire \bin_array[29][0] ;
 wire \bin_array[29][1] ;
 wire \bin_array[29][2] ;
 wire \bin_array[29][3] ;
 wire \bin_array[2][0] ;
 wire \bin_array[2][1] ;
 wire \bin_array[2][2] ;
 wire \bin_array[2][3] ;
 wire \bin_array[30][0] ;
 wire \bin_array[30][1] ;
 wire \bin_array[30][2] ;
 wire \bin_array[30][3] ;
 wire \bin_array[31][0] ;
 wire \bin_array[31][1] ;
 wire \bin_array[31][2] ;
 wire \bin_array[31][3] ;
 wire \bin_array[3][0] ;
 wire \bin_array[3][1] ;
 wire \bin_array[3][2] ;
 wire \bin_array[3][3] ;
 wire \bin_array[4][0] ;
 wire \bin_array[4][1] ;
 wire \bin_array[4][2] ;
 wire \bin_array[4][3] ;
 wire \bin_array[5][0] ;
 wire \bin_array[5][1] ;
 wire \bin_array[5][2] ;
 wire \bin_array[5][3] ;
 wire \bin_array[6][0] ;
 wire \bin_array[6][1] ;
 wire \bin_array[6][2] ;
 wire \bin_array[6][3] ;
 wire \bin_array[7][0] ;
 wire \bin_array[7][1] ;
 wire \bin_array[7][2] ;
 wire \bin_array[7][3] ;
 wire \bin_array[8][0] ;
 wire \bin_array[8][1] ;
 wire \bin_array[8][2] ;
 wire \bin_array[8][3] ;
 wire \bin_array[9][0] ;
 wire \bin_array[9][1] ;
 wire \bin_array[9][2] ;
 wire \bin_array[9][3] ;
 wire last_bin_reg;
 wire ready_reg;
 wire \shift_count[0] ;
 wire \shift_count[1] ;
 wire \shift_count[2] ;
 wire \shift_count[3] ;
 wire \shift_count[4] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire valid_out_reg;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;

 sg13g2_inv_1 _0793_ (.Y(_0150_),
    .A(net535));
 sg13g2_inv_1 _0794_ (.Y(_0151_),
    .A(\state[0] ));
 sg13g2_inv_1 _0795_ (.Y(_0152_),
    .A(net1));
 sg13g2_inv_1 _0796_ (.Y(_0153_),
    .A(\state[2] ));
 sg13g2_inv_1 _0797_ (.Y(_0154_),
    .A(_0005_));
 sg13g2_inv_1 _0798_ (.Y(_0155_),
    .A(net459));
 sg13g2_nor2_1 _0799_ (.A(net539),
    .B(net538),
    .Y(_0156_));
 sg13g2_nor2_2 _0800_ (.A(net536),
    .B(net537),
    .Y(_0157_));
 sg13g2_and3_2 _0801_ (.X(_0158_),
    .A(net518),
    .B(net508),
    .C(net503));
 sg13g2_nand3_1 _0802_ (.B(net505),
    .C(net501),
    .A(net510),
    .Y(_0159_));
 sg13g2_nor2b_1 _0803_ (.A(net537),
    .B_N(net536),
    .Y(_0160_));
 sg13g2_nand2b_1 _0804_ (.Y(_0161_),
    .B(net6),
    .A_N(net5));
 sg13g2_nor4_1 _0805_ (.A(net533),
    .B(net3),
    .C(net4),
    .D(_0161_),
    .Y(_0162_));
 sg13g2_nand4_1 _0806_ (.B(\bin_array[8][2] ),
    .C(net506),
    .A(net514),
    .Y(_0163_),
    .D(net496));
 sg13g2_nor2b_1 _0807_ (.A(net538),
    .B_N(net539),
    .Y(_0164_));
 sg13g2_nand2b_2 _0808_ (.Y(_0165_),
    .B(net3),
    .A_N(net4));
 sg13g2_nor4_1 _0809_ (.A(net533),
    .B(net6),
    .C(net5),
    .D(_0165_),
    .Y(_0166_));
 sg13g2_nand4_1 _0810_ (.B(\bin_array[1][2] ),
    .C(net503),
    .A(net515),
    .Y(_0167_),
    .D(net489));
 sg13g2_and2_1 _0811_ (.A(net539),
    .B(net538),
    .X(_0168_));
 sg13g2_nand2_1 _0812_ (.Y(_0169_),
    .A(net539),
    .B(net538));
 sg13g2_nor2b_2 _0813_ (.A(net536),
    .B_N(net537),
    .Y(_0170_));
 sg13g2_nand2b_2 _0814_ (.Y(_0171_),
    .B(net5),
    .A_N(net536));
 sg13g2_nor3_1 _0815_ (.A(net534),
    .B(_0169_),
    .C(_0171_),
    .Y(_0172_));
 sg13g2_nand4_1 _0816_ (.B(\bin_array[7][2] ),
    .C(net486),
    .A(net514),
    .Y(_0173_),
    .D(net481));
 sg13g2_nor2b_1 _0817_ (.A(net539),
    .B_N(net538),
    .Y(_0174_));
 sg13g2_nand2b_2 _0818_ (.Y(_0175_),
    .B(net4),
    .A_N(net3));
 sg13g2_nor3_1 _0819_ (.A(net533),
    .B(_0171_),
    .C(_0175_),
    .Y(_0176_));
 sg13g2_nand4_1 _0820_ (.B(\bin_array[6][2] ),
    .C(net481),
    .A(net515),
    .Y(_0177_),
    .D(net476));
 sg13g2_nand4_1 _0821_ (.B(_0167_),
    .C(_0173_),
    .A(_0163_),
    .Y(_0178_),
    .D(_0177_));
 sg13g2_nor3_1 _0822_ (.A(net533),
    .B(_0161_),
    .C(_0175_),
    .Y(_0179_));
 sg13g2_nand4_1 _0823_ (.B(\bin_array[10][2] ),
    .C(net496),
    .A(net514),
    .Y(_0180_),
    .D(net476));
 sg13g2_nor4_1 _0824_ (.A(net534),
    .B(net6),
    .C(net537),
    .D(_0169_),
    .Y(_0181_));
 sg13g2_nand4_1 _0825_ (.B(\bin_array[3][2] ),
    .C(net502),
    .A(net516),
    .Y(_0182_),
    .D(net485));
 sg13g2_and2_1 _0826_ (.A(net536),
    .B(net537),
    .X(_0183_));
 sg13g2_nand2_1 _0827_ (.Y(_0184_),
    .A(net536),
    .B(net537));
 sg13g2_nand3_1 _0828_ (.B(net491),
    .C(net468),
    .A(net531),
    .Y(_0185_));
 sg13g2_nand4_1 _0829_ (.B(\bin_array[29][2] ),
    .C(net491),
    .A(net531),
    .Y(_0186_),
    .D(net468));
 sg13g2_nor4_1 _0830_ (.A(net533),
    .B(net536),
    .C(net537),
    .D(_0175_),
    .Y(_0187_));
 sg13g2_nand4_1 _0831_ (.B(\bin_array[2][2] ),
    .C(net503),
    .A(net514),
    .Y(_0188_),
    .D(net476));
 sg13g2_nand4_1 _0832_ (.B(_0182_),
    .C(_0186_),
    .A(_0180_),
    .Y(_0189_),
    .D(_0188_));
 sg13g2_nand3_1 _0833_ (.B(net504),
    .C(net499),
    .A(net521),
    .Y(_0190_));
 sg13g2_nand4_1 _0834_ (.B(\bin_array[16][2] ),
    .C(net507),
    .A(net525),
    .Y(_0191_),
    .D(net502));
 sg13g2_nand3_1 _0835_ (.B(net493),
    .C(net487),
    .A(net522),
    .Y(_0192_));
 sg13g2_nand4_1 _0836_ (.B(\bin_array[25][2] ),
    .C(net497),
    .A(net525),
    .Y(_0193_),
    .D(net489));
 sg13g2_nor3_1 _0837_ (.A(net533),
    .B(_0161_),
    .C(_0169_),
    .Y(_0194_));
 sg13g2_nand4_1 _0838_ (.B(\bin_array[11][2] ),
    .C(net497),
    .A(net517),
    .Y(_0195_),
    .D(net485));
 sg13g2_nand3_1 _0839_ (.B(net499),
    .C(net487),
    .A(net523),
    .Y(_0196_));
 sg13g2_nand4_1 _0840_ (.B(\bin_array[17][2] ),
    .C(net502),
    .A(net525),
    .Y(_0197_),
    .D(net488));
 sg13g2_nand4_1 _0841_ (.B(_0193_),
    .C(_0195_),
    .A(_0191_),
    .Y(_0198_),
    .D(_0197_));
 sg13g2_nor4_1 _0842_ (.A(net534),
    .B(net539),
    .C(net538),
    .D(_0184_),
    .Y(_0199_));
 sg13g2_nand4_1 _0843_ (.B(\bin_array[12][2] ),
    .C(net506),
    .A(net514),
    .Y(_0200_),
    .D(net468));
 sg13g2_nand3_1 _0844_ (.B(net506),
    .C(net468),
    .A(net532),
    .Y(_0201_));
 sg13g2_nand4_1 _0845_ (.B(\bin_array[28][2] ),
    .C(net506),
    .A(net531),
    .Y(_0202_),
    .D(net468));
 sg13g2_nor4_1 _0846_ (.A(net534),
    .B(net539),
    .C(net538),
    .D(_0171_),
    .Y(_0203_));
 sg13g2_nand4_1 _0847_ (.B(\bin_array[4][2] ),
    .C(net506),
    .A(net516),
    .Y(_0204_),
    .D(net481));
 sg13g2_nand3_1 _0848_ (.B(net496),
    .C(net485),
    .A(net532),
    .Y(_0205_));
 sg13g2_nand4_1 _0849_ (.B(\bin_array[27][2] ),
    .C(net496),
    .A(net531),
    .Y(_0206_),
    .D(net485));
 sg13g2_nand4_1 _0850_ (.B(_0202_),
    .C(_0204_),
    .A(_0200_),
    .Y(_0207_),
    .D(_0206_));
 sg13g2_nor4_2 _0851_ (.A(_0178_),
    .B(_0189_),
    .C(_0198_),
    .Y(_0208_),
    .D(_0207_));
 sg13g2_nand3_1 _0852_ (.B(net474),
    .C(net471),
    .A(net529),
    .Y(_0209_));
 sg13g2_nand4_1 _0853_ (.B(\bin_array[30][2] ),
    .C(net474),
    .A(net527),
    .Y(_0210_),
    .D(net471));
 sg13g2_nor3_1 _0854_ (.A(net533),
    .B(_0165_),
    .C(_0171_),
    .Y(_0211_));
 sg13g2_nand4_1 _0855_ (.B(\bin_array[5][2] ),
    .C(net492),
    .A(net511),
    .Y(_0212_),
    .D(net479));
 sg13g2_and4_1 _0856_ (.A(net539),
    .B(net538),
    .C(net536),
    .D(net537),
    .X(_0213_));
 sg13g2_nand3_1 _0857_ (.B(\bin_array[15][2] ),
    .C(net467),
    .A(net511),
    .Y(_0214_));
 sg13g2_nand3_1 _0858_ (.B(net494),
    .C(net472),
    .A(net521),
    .Y(_0215_));
 sg13g2_nand4_1 _0859_ (.B(\bin_array[26][2] ),
    .C(net494),
    .A(net523),
    .Y(_0216_),
    .D(net472));
 sg13g2_nand4_1 _0860_ (.B(_0212_),
    .C(_0214_),
    .A(_0210_),
    .Y(_0217_),
    .D(_0216_));
 sg13g2_nor3_1 _0861_ (.A(net534),
    .B(_0165_),
    .C(_0184_),
    .Y(_0218_));
 sg13g2_nand4_1 _0862_ (.B(\bin_array[13][2] ),
    .C(net490),
    .A(net518),
    .Y(_0219_),
    .D(net470));
 sg13g2_nor3_2 _0863_ (.A(net534),
    .B(_0175_),
    .C(_0184_),
    .Y(_0220_));
 sg13g2_nand4_1 _0864_ (.B(\bin_array[14][2] ),
    .C(net474),
    .A(net511),
    .Y(_0221_),
    .D(net471));
 sg13g2_nand3_1 _0865_ (.B(net502),
    .C(net485),
    .A(net525),
    .Y(_0222_));
 sg13g2_nand4_1 _0866_ (.B(\bin_array[19][2] ),
    .C(net501),
    .A(net529),
    .Y(_0223_),
    .D(net483));
 sg13g2_nand4_1 _0867_ (.B(_0219_),
    .C(_0221_),
    .A(_0159_),
    .Y(_0224_),
    .D(_0223_));
 sg13g2_nand3_1 _0868_ (.B(net499),
    .C(net472),
    .A(net521),
    .Y(_0225_));
 sg13g2_nand4_1 _0869_ (.B(\bin_array[18][2] ),
    .C(net499),
    .A(net522),
    .Y(_0226_),
    .D(net472));
 sg13g2_nand3_1 _0870_ (.B(net504),
    .C(net478),
    .A(net521),
    .Y(_0227_));
 sg13g2_nand4_1 _0871_ (.B(\bin_array[20][2] ),
    .C(net504),
    .A(net522),
    .Y(_0228_),
    .D(net478));
 sg13g2_nor3_1 _0872_ (.A(net533),
    .B(_0161_),
    .C(_0165_),
    .Y(_0229_));
 sg13g2_nand4_1 _0873_ (.B(\bin_array[9][2] ),
    .C(net494),
    .A(net510),
    .Y(_0230_),
    .D(net487));
 sg13g2_nand3_1 _0874_ (.B(net478),
    .C(net472),
    .A(net521),
    .Y(_0231_));
 sg13g2_nand4_1 _0875_ (.B(\bin_array[22][2] ),
    .C(net478),
    .A(net521),
    .Y(_0232_),
    .D(net472));
 sg13g2_nand4_1 _0876_ (.B(_0228_),
    .C(_0230_),
    .A(_0226_),
    .Y(_0233_),
    .D(_0232_));
 sg13g2_nand3_1 _0877_ (.B(net505),
    .C(net495),
    .A(net527),
    .Y(_0234_));
 sg13g2_nand4_1 _0878_ (.B(\bin_array[24][2] ),
    .C(net505),
    .A(net527),
    .Y(_0235_),
    .D(net495));
 sg13g2_nand3_1 _0879_ (.B(net484),
    .C(net479),
    .A(net527),
    .Y(_0236_));
 sg13g2_nand4_1 _0880_ (.B(\bin_array[23][2] ),
    .C(net484),
    .A(net528),
    .Y(_0237_),
    .D(net479));
 sg13g2_nand3_1 _0881_ (.B(\bin_array[31][2] ),
    .C(net467),
    .A(net528),
    .Y(_0238_));
 sg13g2_nand3_1 _0882_ (.B(net492),
    .C(net479),
    .A(net523),
    .Y(_0239_));
 sg13g2_nand4_1 _0883_ (.B(\bin_array[21][2] ),
    .C(net488),
    .A(net527),
    .Y(_0240_),
    .D(net479));
 sg13g2_nand4_1 _0884_ (.B(_0237_),
    .C(_0238_),
    .A(_0235_),
    .Y(_0241_),
    .D(_0240_));
 sg13g2_nor4_2 _0885_ (.A(_0217_),
    .B(_0224_),
    .C(_0233_),
    .Y(_0242_),
    .D(_0241_));
 sg13g2_a22oi_1 _0886_ (.Y(_0243_),
    .B1(_0208_),
    .B2(_0242_),
    .A2(_0158_),
    .A1(_0003_));
 sg13g2_nand4_1 _0887_ (.B(\bin_array[28][3] ),
    .C(net507),
    .A(net531),
    .Y(_0244_),
    .D(net468));
 sg13g2_nand4_1 _0888_ (.B(\bin_array[9][3] ),
    .C(net496),
    .A(net514),
    .Y(_0245_),
    .D(net489));
 sg13g2_nand4_1 _0889_ (.B(\bin_array[5][3] ),
    .C(net489),
    .A(net517),
    .Y(_0246_),
    .D(net481));
 sg13g2_nand4_1 _0890_ (.B(\bin_array[8][3] ),
    .C(net506),
    .A(net515),
    .Y(_0247_),
    .D(net497));
 sg13g2_nand4_1 _0891_ (.B(_0245_),
    .C(_0246_),
    .A(_0244_),
    .Y(_0248_),
    .D(_0247_));
 sg13g2_nand3_1 _0892_ (.B(\bin_array[31][3] ),
    .C(net467),
    .A(net529),
    .Y(_0249_));
 sg13g2_nand4_1 _0893_ (.B(\bin_array[22][3] ),
    .C(net478),
    .A(net521),
    .Y(_0250_),
    .D(net472));
 sg13g2_nand4_1 _0894_ (.B(\bin_array[20][3] ),
    .C(net504),
    .A(net522),
    .Y(_0251_),
    .D(net478));
 sg13g2_nand4_1 _0895_ (.B(\bin_array[16][3] ),
    .C(net504),
    .A(net521),
    .Y(_0252_),
    .D(net499));
 sg13g2_nand4_1 _0896_ (.B(_0250_),
    .C(_0251_),
    .A(_0249_),
    .Y(_0253_),
    .D(_0252_));
 sg13g2_nand4_1 _0897_ (.B(\bin_array[2][3] ),
    .C(net503),
    .A(net515),
    .Y(_0254_),
    .D(net476));
 sg13g2_nand4_1 _0898_ (.B(\bin_array[7][3] ),
    .C(net485),
    .A(net515),
    .Y(_0255_),
    .D(net481));
 sg13g2_nand4_1 _0899_ (.B(\bin_array[21][3] ),
    .C(net489),
    .A(net525),
    .Y(_0256_),
    .D(net481));
 sg13g2_nand4_1 _0900_ (.B(\bin_array[17][3] ),
    .C(net502),
    .A(net531),
    .Y(_0257_),
    .D(net489));
 sg13g2_nand4_1 _0901_ (.B(_0255_),
    .C(_0256_),
    .A(_0254_),
    .Y(_0258_),
    .D(_0257_));
 sg13g2_nand4_1 _0902_ (.B(\bin_array[27][3] ),
    .C(net496),
    .A(net531),
    .Y(_0259_),
    .D(net486));
 sg13g2_nand4_1 _0903_ (.B(\bin_array[6][3] ),
    .C(net481),
    .A(net515),
    .Y(_0260_),
    .D(net476));
 sg13g2_nand4_1 _0904_ (.B(\bin_array[30][3] ),
    .C(net474),
    .A(net527),
    .Y(_0261_),
    .D(net471));
 sg13g2_nand4_1 _0905_ (.B(\bin_array[12][3] ),
    .C(net506),
    .A(net517),
    .Y(_0262_),
    .D(net468));
 sg13g2_nand4_1 _0906_ (.B(_0260_),
    .C(_0261_),
    .A(_0259_),
    .Y(_0263_),
    .D(_0262_));
 sg13g2_nor4_2 _0907_ (.A(_0248_),
    .B(_0253_),
    .C(_0258_),
    .Y(_0264_),
    .D(_0263_));
 sg13g2_nand4_1 _0908_ (.B(\bin_array[23][3] ),
    .C(net483),
    .A(net528),
    .Y(_0265_),
    .D(net479));
 sg13g2_nand4_1 _0909_ (.B(\bin_array[18][3] ),
    .C(net501),
    .A(net523),
    .Y(_0266_),
    .D(net474));
 sg13g2_nand4_1 _0910_ (.B(\bin_array[24][3] ),
    .C(net505),
    .A(net527),
    .Y(_0267_),
    .D(net495));
 sg13g2_nand3_1 _0911_ (.B(\bin_array[15][3] ),
    .C(net467),
    .A(net511),
    .Y(_0268_));
 sg13g2_nand4_1 _0912_ (.B(_0266_),
    .C(_0267_),
    .A(_0265_),
    .Y(_0269_),
    .D(_0268_));
 sg13g2_nand4_1 _0913_ (.B(\bin_array[26][3] ),
    .C(net493),
    .A(net524),
    .Y(_0270_),
    .D(net473));
 sg13g2_nand4_1 _0914_ (.B(\bin_array[29][3] ),
    .C(net489),
    .A(net525),
    .Y(_0271_),
    .D(net469));
 sg13g2_nand4_1 _0915_ (.B(\bin_array[19][3] ),
    .C(net502),
    .A(net525),
    .Y(_0272_),
    .D(net483));
 sg13g2_nand4_1 _0916_ (.B(_0270_),
    .C(_0271_),
    .A(_0159_),
    .Y(_0273_),
    .D(_0272_));
 sg13g2_nand4_1 _0917_ (.B(\bin_array[13][3] ),
    .C(net490),
    .A(net519),
    .Y(_0274_),
    .D(net470));
 sg13g2_nand4_1 _0918_ (.B(\bin_array[10][3] ),
    .C(net498),
    .A(net520),
    .Y(_0275_),
    .D(net477));
 sg13g2_nand4_1 _0919_ (.B(\bin_array[25][3] ),
    .C(net498),
    .A(net532),
    .Y(_0276_),
    .D(net491));
 sg13g2_nand4_1 _0920_ (.B(\bin_array[11][3] ),
    .C(net498),
    .A(net519),
    .Y(_0277_),
    .D(net486));
 sg13g2_nand4_1 _0921_ (.B(_0275_),
    .C(_0276_),
    .A(_0274_),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_nand4_1 _0922_ (.B(\bin_array[3][3] ),
    .C(net503),
    .A(net518),
    .Y(_0279_),
    .D(net486));
 sg13g2_nand4_1 _0923_ (.B(\bin_array[4][3] ),
    .C(net508),
    .A(net518),
    .Y(_0280_),
    .D(net482));
 sg13g2_nand4_1 _0924_ (.B(\bin_array[14][3] ),
    .C(net475),
    .A(net512),
    .Y(_0281_),
    .D(net471));
 sg13g2_nand4_1 _0925_ (.B(\bin_array[1][3] ),
    .C(net501),
    .A(net512),
    .Y(_0282_),
    .D(net488));
 sg13g2_nand4_1 _0926_ (.B(_0280_),
    .C(_0281_),
    .A(_0279_),
    .Y(_0283_),
    .D(_0282_));
 sg13g2_nor4_2 _0927_ (.A(_0269_),
    .B(_0273_),
    .C(_0278_),
    .Y(_0284_),
    .D(_0283_));
 sg13g2_a22oi_1 _0928_ (.Y(_0285_),
    .B1(_0264_),
    .B2(_0284_),
    .A2(_0158_),
    .A1(_0004_));
 sg13g2_inv_1 _0929_ (.Y(_0286_),
    .A(_0285_));
 sg13g2_and2_1 _0930_ (.A(_0243_),
    .B(_0285_),
    .X(_0287_));
 sg13g2_nand4_1 _0931_ (.B(\bin_array[18][0] ),
    .C(net501),
    .A(net523),
    .Y(_0288_),
    .D(net473));
 sg13g2_nand4_1 _0932_ (.B(\bin_array[3][0] ),
    .C(net501),
    .A(net511),
    .Y(_0289_),
    .D(net484));
 sg13g2_nand4_1 _0933_ (.B(\bin_array[7][0] ),
    .C(net483),
    .A(net510),
    .Y(_0290_),
    .D(net478));
 sg13g2_nand4_1 _0934_ (.B(\bin_array[8][0] ),
    .C(net504),
    .A(net510),
    .Y(_0291_),
    .D(net493));
 sg13g2_nand4_1 _0935_ (.B(\bin_array[21][0] ),
    .C(net488),
    .A(net523),
    .Y(_0292_),
    .D(net480));
 sg13g2_nand4_1 _0936_ (.B(\bin_array[27][0] ),
    .C(net494),
    .A(net526),
    .Y(_0293_),
    .D(net483));
 sg13g2_nand4_1 _0937_ (.B(\bin_array[26][0] ),
    .C(net493),
    .A(net524),
    .Y(_0294_),
    .D(net473));
 sg13g2_nand4_1 _0938_ (.B(\bin_array[6][0] ),
    .C(net479),
    .A(net512),
    .Y(_0295_),
    .D(net474));
 sg13g2_nand4_1 _0939_ (.B(\bin_array[20][0] ),
    .C(net504),
    .A(net522),
    .Y(_0296_),
    .D(net478));
 sg13g2_nand4_1 _0940_ (.B(\bin_array[17][0] ),
    .C(net499),
    .A(net522),
    .Y(_0297_),
    .D(net487));
 sg13g2_nand4_1 _0941_ (.B(\bin_array[23][0] ),
    .C(net483),
    .A(net528),
    .Y(_0298_),
    .D(net479));
 sg13g2_nand4_1 _0942_ (.B(\bin_array[16][0] ),
    .C(net505),
    .A(net530),
    .Y(_0299_),
    .D(_0157_));
 sg13g2_nand4_1 _0943_ (.B(\bin_array[24][0] ),
    .C(net508),
    .A(net526),
    .Y(_0300_),
    .D(net498));
 sg13g2_nand4_1 _0944_ (.B(\bin_array[12][0] ),
    .C(net508),
    .A(net516),
    .Y(_0301_),
    .D(net470));
 sg13g2_nand4_1 _0945_ (.B(\bin_array[28][0] ),
    .C(net509),
    .A(net532),
    .Y(_0302_),
    .D(net470));
 sg13g2_nand4_1 _0946_ (.B(\bin_array[4][0] ),
    .C(net508),
    .A(net519),
    .Y(_0303_),
    .D(net482));
 sg13g2_nand4_1 _0947_ (.B(\bin_array[22][0] ),
    .C(net480),
    .A(net523),
    .Y(_0304_),
    .D(net473));
 sg13g2_nand4_1 _0948_ (.B(\bin_array[25][0] ),
    .C(net493),
    .A(net526),
    .Y(_0305_),
    .D(net487));
 sg13g2_nand3_1 _0949_ (.B(\bin_array[31][0] ),
    .C(net467),
    .A(net528),
    .Y(_0306_));
 sg13g2_nand4_1 _0950_ (.B(\bin_array[5][0] ),
    .C(net488),
    .A(net510),
    .Y(_0307_),
    .D(net480));
 sg13g2_nand4_1 _0951_ (.B(\bin_array[1][0] ),
    .C(net499),
    .A(net510),
    .Y(_0308_),
    .D(net487));
 sg13g2_nand3_1 _0952_ (.B(\bin_array[15][0] ),
    .C(net467),
    .A(net512),
    .Y(_0309_));
 sg13g2_nand4_1 _0953_ (.B(\bin_array[10][0] ),
    .C(net495),
    .A(net510),
    .Y(_0310_),
    .D(net472));
 sg13g2_nand4_1 _0954_ (.B(\bin_array[9][0] ),
    .C(net493),
    .A(net513),
    .Y(_0311_),
    .D(net487));
 sg13g2_nand4_1 _0955_ (.B(\bin_array[30][0] ),
    .C(net474),
    .A(net527),
    .Y(_0312_),
    .D(net471));
 sg13g2_nand4_1 _0956_ (.B(\bin_array[19][0] ),
    .C(net499),
    .A(net522),
    .Y(_0313_),
    .D(net483));
 sg13g2_nand4_1 _0957_ (.B(\bin_array[14][0] ),
    .C(net477),
    .A(net518),
    .Y(_0314_),
    .D(net470));
 sg13g2_nand4_1 _0958_ (.B(\bin_array[2][0] ),
    .C(net502),
    .A(net516),
    .Y(_0315_),
    .D(net476));
 sg13g2_nand4_1 _0959_ (.B(\bin_array[13][0] ),
    .C(net490),
    .A(net520),
    .Y(_0316_),
    .D(net470));
 sg13g2_nand4_1 _0960_ (.B(\bin_array[29][0] ),
    .C(net490),
    .A(net532),
    .Y(_0317_),
    .D(net469));
 sg13g2_nand4_1 _0961_ (.B(\bin_array[11][0] ),
    .C(net495),
    .A(net511),
    .Y(_0318_),
    .D(net484));
 sg13g2_nand4_1 _0962_ (.B(_0293_),
    .C(_0308_),
    .A(_0292_),
    .Y(_0319_),
    .D(_0310_));
 sg13g2_nand4_1 _0963_ (.B(_0289_),
    .C(_0307_),
    .A(_0288_),
    .Y(_0320_),
    .D(_0318_));
 sg13g2_nand4_1 _0964_ (.B(_0290_),
    .C(_0304_),
    .A(_0159_),
    .Y(_0321_),
    .D(_0306_));
 sg13g2_nand4_1 _0965_ (.B(_0296_),
    .C(_0297_),
    .A(_0291_),
    .Y(_0322_),
    .D(_0313_));
 sg13g2_nor4_2 _0966_ (.A(_0319_),
    .B(_0320_),
    .C(_0321_),
    .Y(_0323_),
    .D(_0322_));
 sg13g2_nand4_1 _0967_ (.B(_0305_),
    .C(_0309_),
    .A(_0294_),
    .Y(_0324_),
    .D(_0311_));
 sg13g2_nand4_1 _0968_ (.B(_0298_),
    .C(_0299_),
    .A(_0295_),
    .Y(_0325_),
    .D(_0312_));
 sg13g2_nand4_1 _0969_ (.B(_0315_),
    .C(_0316_),
    .A(_0300_),
    .Y(_0326_),
    .D(_0317_));
 sg13g2_nand4_1 _0970_ (.B(_0302_),
    .C(_0303_),
    .A(_0301_),
    .Y(_0327_),
    .D(_0314_));
 sg13g2_nor4_2 _0971_ (.A(_0324_),
    .B(_0325_),
    .C(_0326_),
    .Y(_0328_),
    .D(_0327_));
 sg13g2_nor2_1 _0972_ (.A(\bin_array[0][0] ),
    .B(_0159_),
    .Y(_0329_));
 sg13g2_a21oi_2 _0973_ (.B1(_0329_),
    .Y(_0330_),
    .A2(_0328_),
    .A1(_0323_));
 sg13g2_a21o_1 _0974_ (.A2(_0328_),
    .A1(_0323_),
    .B1(_0329_),
    .X(_0331_));
 sg13g2_nand4_1 _0975_ (.B(\bin_array[30][1] ),
    .C(net475),
    .A(net529),
    .Y(_0332_),
    .D(net471));
 sg13g2_nand4_1 _0976_ (.B(\bin_array[20][1] ),
    .C(net505),
    .A(net530),
    .Y(_0333_),
    .D(net480));
 sg13g2_nand4_1 _0977_ (.B(\bin_array[7][1] ),
    .C(net486),
    .A(net518),
    .Y(_0334_),
    .D(net482));
 sg13g2_nand4_1 _0978_ (.B(\bin_array[4][1] ),
    .C(net508),
    .A(net518),
    .Y(_0335_),
    .D(net482));
 sg13g2_nand4_1 _0979_ (.B(_0333_),
    .C(_0334_),
    .A(_0332_),
    .Y(_0336_),
    .D(_0335_));
 sg13g2_nand4_1 _0980_ (.B(\bin_array[29][1] ),
    .C(net490),
    .A(net529),
    .Y(_0337_),
    .D(_0183_));
 sg13g2_nand4_1 _0981_ (.B(\bin_array[19][1] ),
    .C(net503),
    .A(net529),
    .Y(_0338_),
    .D(net486));
 sg13g2_nand4_1 _0982_ (.B(\bin_array[14][1] ),
    .C(net474),
    .A(net512),
    .Y(_0339_),
    .D(net471));
 sg13g2_nand4_1 _0983_ (.B(\bin_array[6][1] ),
    .C(net482),
    .A(net519),
    .Y(_0340_),
    .D(net477));
 sg13g2_nand4_1 _0984_ (.B(_0338_),
    .C(_0339_),
    .A(_0337_),
    .Y(_0341_),
    .D(_0340_));
 sg13g2_nand3_1 _0985_ (.B(\bin_array[15][1] ),
    .C(_0213_),
    .A(net511),
    .Y(_0342_));
 sg13g2_nand4_1 _0986_ (.B(\bin_array[10][1] ),
    .C(net498),
    .A(net518),
    .Y(_0343_),
    .D(net476));
 sg13g2_nand4_1 _0987_ (.B(\bin_array[23][1] ),
    .C(net483),
    .A(net529),
    .Y(_0344_),
    .D(net480));
 sg13g2_nand3_1 _0988_ (.B(\bin_array[31][1] ),
    .C(_0213_),
    .A(net528),
    .Y(_0345_));
 sg13g2_nand4_1 _0989_ (.B(_0343_),
    .C(_0344_),
    .A(_0342_),
    .Y(_0346_),
    .D(_0345_));
 sg13g2_nand4_1 _0990_ (.B(\bin_array[24][1] ),
    .C(net508),
    .A(net535),
    .Y(_0347_),
    .D(net498));
 sg13g2_nand4_1 _0991_ (.B(\bin_array[5][1] ),
    .C(net490),
    .A(net519),
    .Y(_0348_),
    .D(net482));
 sg13g2_nand4_1 _0992_ (.B(\bin_array[3][1] ),
    .C(net503),
    .A(net519),
    .Y(_0349_),
    .D(net486));
 sg13g2_nand4_1 _0993_ (.B(\bin_array[12][1] ),
    .C(net508),
    .A(net519),
    .Y(_0350_),
    .D(net470));
 sg13g2_nand4_1 _0994_ (.B(_0348_),
    .C(_0349_),
    .A(_0347_),
    .Y(_0351_),
    .D(_0350_));
 sg13g2_nor4_2 _0995_ (.A(_0336_),
    .B(_0341_),
    .C(_0346_),
    .Y(_0352_),
    .D(_0351_));
 sg13g2_nand4_1 _0996_ (.B(\bin_array[13][1] ),
    .C(net490),
    .A(net517),
    .Y(_0353_),
    .D(net469));
 sg13g2_nand4_1 _0997_ (.B(\bin_array[8][1] ),
    .C(net507),
    .A(net517),
    .Y(_0354_),
    .D(net497));
 sg13g2_nand4_1 _0998_ (.B(\bin_array[26][1] ),
    .C(net493),
    .A(net524),
    .Y(_0355_),
    .D(net473));
 sg13g2_nand4_1 _0999_ (.B(\bin_array[21][1] ),
    .C(net490),
    .A(net526),
    .Y(_0356_),
    .D(net481));
 sg13g2_nand4_1 _1000_ (.B(_0354_),
    .C(_0355_),
    .A(_0353_),
    .Y(_0357_),
    .D(_0356_));
 sg13g2_nand4_1 _1001_ (.B(\bin_array[17][1] ),
    .C(net500),
    .A(net524),
    .Y(_0358_),
    .D(net488));
 sg13g2_nand4_1 _1002_ (.B(\bin_array[27][1] ),
    .C(net497),
    .A(net525),
    .Y(_0359_),
    .D(net485));
 sg13g2_nand4_1 _1003_ (.B(\bin_array[1][1] ),
    .C(net500),
    .A(net510),
    .Y(_0360_),
    .D(net487));
 sg13g2_nand4_1 _1004_ (.B(_0358_),
    .C(_0359_),
    .A(_0159_),
    .Y(_0361_),
    .D(_0360_));
 sg13g2_nand4_1 _1005_ (.B(\bin_array[22][1] ),
    .C(net480),
    .A(net524),
    .Y(_0362_),
    .D(net473));
 sg13g2_nand4_1 _1006_ (.B(\bin_array[16][1] ),
    .C(net504),
    .A(net524),
    .Y(_0363_),
    .D(net500));
 sg13g2_nand4_1 _1007_ (.B(\bin_array[18][1] ),
    .C(net500),
    .A(net524),
    .Y(_0364_),
    .D(net473));
 sg13g2_nand4_1 _1008_ (.B(\bin_array[25][1] ),
    .C(net493),
    .A(net524),
    .Y(_0365_),
    .D(net488));
 sg13g2_nand4_1 _1009_ (.B(_0363_),
    .C(_0364_),
    .A(_0362_),
    .Y(_0366_),
    .D(_0365_));
 sg13g2_nand4_1 _1010_ (.B(\bin_array[28][1] ),
    .C(net506),
    .A(net531),
    .Y(_0367_),
    .D(net468));
 sg13g2_nand4_1 _1011_ (.B(\bin_array[11][1] ),
    .C(net496),
    .A(net515),
    .Y(_0368_),
    .D(net485));
 sg13g2_nand4_1 _1012_ (.B(\bin_array[2][1] ),
    .C(net502),
    .A(net514),
    .Y(_0369_),
    .D(net476));
 sg13g2_nand4_1 _1013_ (.B(\bin_array[9][1] ),
    .C(net496),
    .A(net514),
    .Y(_0370_),
    .D(net489));
 sg13g2_nand4_1 _1014_ (.B(_0368_),
    .C(_0369_),
    .A(_0367_),
    .Y(_0371_),
    .D(_0370_));
 sg13g2_nor4_2 _1015_ (.A(_0357_),
    .B(_0361_),
    .C(_0366_),
    .Y(_0372_),
    .D(_0371_));
 sg13g2_a22oi_1 _1016_ (.Y(_0373_),
    .B1(_0352_),
    .B2(_0372_),
    .A2(_0158_),
    .A1(_0002_));
 sg13g2_a221oi_1 _1017_ (.B2(_0372_),
    .C1(_0152_),
    .B1(_0352_),
    .A1(_0002_),
    .Y(_0374_),
    .A2(_0158_));
 sg13g2_nand4_1 _1018_ (.B(_0285_),
    .C(_0331_),
    .A(_0243_),
    .Y(_0375_),
    .D(_0374_));
 sg13g2_nand3_1 _1019_ (.B(net7),
    .C(net2),
    .A(ready_reg),
    .Y(_0376_));
 sg13g2_and2_1 _1020_ (.A(net31),
    .B(_0376_),
    .X(_0377_));
 sg13g2_nand2_1 _1021_ (.Y(_0378_),
    .A(\state[0] ),
    .B(_0376_));
 sg13g2_a221oi_1 _1022_ (.B2(net31),
    .C1(_0377_),
    .B1(_0375_),
    .A1(net29),
    .Y(_0009_),
    .A2(net1));
 sg13g2_nor2_1 _1023_ (.A(_0151_),
    .B(_0376_),
    .Y(_0379_));
 sg13g2_or2_1 _1024_ (.X(_0380_),
    .B(_0376_),
    .A(_0151_));
 sg13g2_nand2_2 _1025_ (.Y(_0381_),
    .A(\shift_count[1] ),
    .B(\shift_count[0] ));
 sg13g2_nand2_2 _1026_ (.Y(_0382_),
    .A(net464),
    .B(net466));
 sg13g2_nand3_1 _1027_ (.B(\shift_count[0] ),
    .C(net466),
    .A(\shift_count[1] ),
    .Y(_0383_));
 sg13g2_nor2_2 _1028_ (.A(_0381_),
    .B(_0382_),
    .Y(_0384_));
 sg13g2_and2_2 _1029_ (.A(net462),
    .B(_0384_),
    .X(_0385_));
 sg13g2_nand2_2 _1030_ (.Y(_0386_),
    .A(net462),
    .B(_0384_));
 sg13g2_o21ai_1 _1031_ (.B1(net177),
    .Y(_0387_),
    .A1(_0152_),
    .A2(_0386_));
 sg13g2_o21ai_1 _1032_ (.B1(_0387_),
    .Y(_0001_),
    .A1(_0375_),
    .A2(net453));
 sg13g2_nor2_1 _1033_ (.A(_0152_),
    .B(_0153_),
    .Y(_0388_));
 sg13g2_nand2_2 _1034_ (.Y(_0389_),
    .A(net1),
    .B(\state[2] ));
 sg13g2_nand2_1 _1035_ (.Y(_0390_),
    .A(net29),
    .B(_0152_));
 sg13g2_o21ai_1 _1036_ (.B1(_0390_),
    .Y(_0000_),
    .A1(_0386_),
    .A2(_0389_));
 sg13g2_o21ai_1 _1037_ (.B1(net1),
    .Y(_0391_),
    .A1(\state[0] ),
    .A2(\state[2] ));
 sg13g2_nand2_1 _1038_ (.Y(_0392_),
    .A(net42),
    .B(_0391_));
 sg13g2_nand2b_2 _1039_ (.Y(_0393_),
    .B(\shift_count[1] ),
    .A_N(\shift_count[0] ));
 sg13g2_nand2b_2 _1040_ (.Y(_0394_),
    .B(net465),
    .A_N(net463));
 sg13g2_nor3_2 _1041_ (.A(net457),
    .B(_0393_),
    .C(_0394_),
    .Y(_0395_));
 sg13g2_or2_1 _1042_ (.X(_0396_),
    .B(\shift_count[0] ),
    .A(\shift_count[1] ));
 sg13g2_nor3_2 _1043_ (.A(net457),
    .B(_0382_),
    .C(net456),
    .Y(_0397_));
 sg13g2_nand2b_2 _1044_ (.Y(_0398_),
    .B(net463),
    .A_N(net465));
 sg13g2_nor3_2 _1045_ (.A(net457),
    .B(_0381_),
    .C(_0398_),
    .Y(_0399_));
 sg13g2_nand2b_2 _1046_ (.Y(_0400_),
    .B(\shift_count[0] ),
    .A_N(\shift_count[1] ));
 sg13g2_nor3_2 _1047_ (.A(net460),
    .B(_0398_),
    .C(_0400_),
    .Y(_0401_));
 sg13g2_nor3_2 _1048_ (.A(net461),
    .B(_0394_),
    .C(net456),
    .Y(_0402_));
 sg13g2_nor3_2 _1049_ (.A(_0155_),
    .B(_0381_),
    .C(_0382_),
    .Y(_0403_));
 sg13g2_or3_2 _1050_ (.A(net463),
    .B(net465),
    .C(net458),
    .X(_0404_));
 sg13g2_nor2_2 _1051_ (.A(_0381_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_nor3_2 _1052_ (.A(net461),
    .B(_0393_),
    .C(_0398_),
    .Y(_0406_));
 sg13g2_nor3_2 _1053_ (.A(net460),
    .B(_0394_),
    .C(_0400_),
    .Y(_0407_));
 sg13g2_nor4_2 _1054_ (.A(net463),
    .B(net465),
    .C(net461),
    .Y(_0408_),
    .D(_0393_));
 sg13g2_nor3_2 _1055_ (.A(net457),
    .B(_0393_),
    .C(_0398_),
    .Y(_0409_));
 sg13g2_nor4_2 _1056_ (.A(net463),
    .B(net465),
    .C(net461),
    .Y(_0410_),
    .D(_0400_));
 sg13g2_nor3_1 _1057_ (.A(net464),
    .B(net466),
    .C(_0396_),
    .Y(_0411_));
 sg13g2_nor2_2 _1058_ (.A(net456),
    .B(_0404_),
    .Y(_0412_));
 sg13g2_nor3_2 _1059_ (.A(net460),
    .B(_0393_),
    .C(_0394_),
    .Y(_0413_));
 sg13g2_nor3_2 _1060_ (.A(net463),
    .B(net460),
    .C(_0383_),
    .Y(_0414_));
 sg13g2_nand3_1 _1061_ (.B(net464),
    .C(net466),
    .A(\shift_count[1] ),
    .Y(_0415_));
 sg13g2_a21o_1 _1062_ (.A2(_0415_),
    .A1(net462),
    .B1(_0411_),
    .X(_0416_));
 sg13g2_nor2_1 _1063_ (.A(net462),
    .B(net459),
    .Y(_0417_));
 sg13g2_a22oi_1 _1064_ (.Y(_0418_),
    .B1(_0417_),
    .B2(_0384_),
    .A2(_0416_),
    .A1(net459));
 sg13g2_inv_1 _1065_ (.Y(_0419_),
    .A(_0418_));
 sg13g2_nor3_2 _1066_ (.A(net463),
    .B(net458),
    .C(_0383_),
    .Y(_0420_));
 sg13g2_nor3_2 _1067_ (.A(net457),
    .B(_0394_),
    .C(_0400_),
    .Y(_0421_));
 sg13g2_nor2_2 _1068_ (.A(_0393_),
    .B(_0404_),
    .Y(_0422_));
 sg13g2_nand2_1 _1069_ (.Y(_0423_),
    .A(\bin_array[18][0] ),
    .B(_0422_));
 sg13g2_nor4_2 _1070_ (.A(net463),
    .B(net465),
    .C(net460),
    .Y(_0424_),
    .D(_0381_));
 sg13g2_nor3_2 _1071_ (.A(net458),
    .B(net456),
    .C(_0398_),
    .Y(_0425_));
 sg13g2_nor3_2 _1072_ (.A(_0155_),
    .B(_0382_),
    .C(_0393_),
    .Y(_0426_));
 sg13g2_nor3_2 _1073_ (.A(net459),
    .B(_0382_),
    .C(_0393_),
    .Y(_0427_));
 sg13g2_nor3_2 _1074_ (.A(net460),
    .B(_0382_),
    .C(net456),
    .Y(_0428_));
 sg13g2_nor3_2 _1075_ (.A(net457),
    .B(_0382_),
    .C(_0400_),
    .Y(_0429_));
 sg13g2_a22oi_1 _1076_ (.Y(_0430_),
    .B1(_0429_),
    .B2(\bin_array[29][0] ),
    .A2(_0428_),
    .A1(\bin_array[12][0] ));
 sg13g2_nor2_2 _1077_ (.A(_0400_),
    .B(_0404_),
    .Y(_0431_));
 sg13g2_nor3_2 _1078_ (.A(net460),
    .B(_0381_),
    .C(_0398_),
    .Y(_0432_));
 sg13g2_nor3_2 _1079_ (.A(net461),
    .B(_0382_),
    .C(_0400_),
    .Y(_0433_));
 sg13g2_nor3_2 _1080_ (.A(net457),
    .B(_0394_),
    .C(net456),
    .Y(_0434_));
 sg13g2_nor3_2 _1081_ (.A(net460),
    .B(net456),
    .C(_0398_),
    .Y(_0435_));
 sg13g2_nor3_2 _1082_ (.A(net457),
    .B(_0398_),
    .C(_0400_),
    .Y(_0436_));
 sg13g2_a22oi_1 _1083_ (.Y(_0437_),
    .B1(_0433_),
    .B2(\bin_array[13][0] ),
    .A2(_0402_),
    .A1(\bin_array[4][0] ));
 sg13g2_a22oi_1 _1084_ (.Y(_0438_),
    .B1(_0424_),
    .B2(\bin_array[3][0] ),
    .A2(_0421_),
    .A1(\bin_array[21][0] ));
 sg13g2_a22oi_1 _1085_ (.Y(_0439_),
    .B1(_0431_),
    .B2(\bin_array[17][0] ),
    .A2(_0395_),
    .A1(\bin_array[22][0] ));
 sg13g2_a22oi_1 _1086_ (.Y(_0440_),
    .B1(_0434_),
    .B2(\bin_array[20][0] ),
    .A2(_0405_),
    .A1(\bin_array[19][0] ));
 sg13g2_nand4_1 _1087_ (.B(_0438_),
    .C(_0439_),
    .A(_0437_),
    .Y(_0441_),
    .D(_0440_));
 sg13g2_a22oi_1 _1088_ (.Y(_0442_),
    .B1(_0425_),
    .B2(\bin_array[24][0] ),
    .A2(_0407_),
    .A1(\bin_array[5][0] ));
 sg13g2_nand3_1 _1089_ (.B(_0423_),
    .C(_0442_),
    .A(_0418_),
    .Y(_0443_));
 sg13g2_a22oi_1 _1090_ (.Y(_0444_),
    .B1(_0435_),
    .B2(\bin_array[8][0] ),
    .A2(_0409_),
    .A1(\bin_array[26][0] ));
 sg13g2_a22oi_1 _1091_ (.Y(_0445_),
    .B1(_0412_),
    .B2(\bin_array[16][0] ),
    .A2(_0410_),
    .A1(\bin_array[1][0] ));
 sg13g2_a22oi_1 _1092_ (.Y(_0446_),
    .B1(_0420_),
    .B2(\bin_array[23][0] ),
    .A2(_0399_),
    .A1(\bin_array[27][0] ));
 sg13g2_nand3_1 _1093_ (.B(_0445_),
    .C(_0446_),
    .A(_0444_),
    .Y(_0447_));
 sg13g2_a221oi_1 _1094_ (.B2(\bin_array[10][0] ),
    .C1(_0447_),
    .B1(_0406_),
    .A1(\bin_array[28][0] ),
    .Y(_0448_),
    .A2(_0397_));
 sg13g2_a22oi_1 _1095_ (.Y(_0449_),
    .B1(_0408_),
    .B2(\bin_array[2][0] ),
    .A2(_0401_),
    .A1(\bin_array[9][0] ));
 sg13g2_a22oi_1 _1096_ (.Y(_0450_),
    .B1(_0436_),
    .B2(\bin_array[25][0] ),
    .A2(_0414_),
    .A1(\bin_array[7][0] ));
 sg13g2_nand3_1 _1097_ (.B(_0449_),
    .C(_0450_),
    .A(_0430_),
    .Y(_0451_));
 sg13g2_a221oi_1 _1098_ (.B2(\bin_array[11][0] ),
    .C1(_0451_),
    .B1(_0432_),
    .A1(\bin_array[6][0] ),
    .Y(_0452_),
    .A2(_0413_));
 sg13g2_a22oi_1 _1099_ (.Y(_0453_),
    .B1(_0426_),
    .B2(\bin_array[14][0] ),
    .A2(_0403_),
    .A1(\bin_array[15][0] ));
 sg13g2_a22oi_1 _1100_ (.Y(_0454_),
    .B1(_0427_),
    .B2(\bin_array[30][0] ),
    .A2(_0385_),
    .A1(\bin_array[31][0] ));
 sg13g2_nand4_1 _1101_ (.B(_0452_),
    .C(_0453_),
    .A(_0448_),
    .Y(_0455_),
    .D(_0454_));
 sg13g2_nor3_2 _1102_ (.A(_0441_),
    .B(_0443_),
    .C(_0455_),
    .Y(_0456_));
 sg13g2_o21ai_1 _1103_ (.B1(_0388_),
    .Y(_0457_),
    .A1(\bin_array[0][0] ),
    .A2(_0418_));
 sg13g2_o21ai_1 _1104_ (.B1(net43),
    .Y(_0010_),
    .A1(_0456_),
    .A2(_0457_));
 sg13g2_nand2_1 _1105_ (.Y(_0458_),
    .A(\bin_array[23][1] ),
    .B(_0420_));
 sg13g2_a22oi_1 _1106_ (.Y(_0459_),
    .B1(_0433_),
    .B2(\bin_array[13][1] ),
    .A2(_0407_),
    .A1(\bin_array[5][1] ));
 sg13g2_a22oi_1 _1107_ (.Y(_0460_),
    .B1(_0414_),
    .B2(\bin_array[7][1] ),
    .A2(_0395_),
    .A1(\bin_array[22][1] ));
 sg13g2_a22oi_1 _1108_ (.Y(_0461_),
    .B1(_0412_),
    .B2(\bin_array[16][1] ),
    .A2(_0409_),
    .A1(\bin_array[26][1] ));
 sg13g2_a22oi_1 _1109_ (.Y(_0462_),
    .B1(_0408_),
    .B2(\bin_array[2][1] ),
    .A2(_0399_),
    .A1(\bin_array[27][1] ));
 sg13g2_a22oi_1 _1110_ (.Y(_0463_),
    .B1(_0434_),
    .B2(\bin_array[20][1] ),
    .A2(_0422_),
    .A1(\bin_array[18][1] ));
 sg13g2_nand4_1 _1111_ (.B(_0460_),
    .C(_0462_),
    .A(_0459_),
    .Y(_0464_),
    .D(_0463_));
 sg13g2_nand3_1 _1112_ (.B(_0458_),
    .C(_0461_),
    .A(_0418_),
    .Y(_0465_));
 sg13g2_nor2_1 _1113_ (.A(_0464_),
    .B(_0465_),
    .Y(_0466_));
 sg13g2_a22oi_1 _1114_ (.Y(_0467_),
    .B1(_0431_),
    .B2(\bin_array[17][1] ),
    .A2(_0410_),
    .A1(\bin_array[1][1] ));
 sg13g2_a22oi_1 _1115_ (.Y(_0468_),
    .B1(_0401_),
    .B2(\bin_array[9][1] ),
    .A2(_0397_),
    .A1(\bin_array[28][1] ));
 sg13g2_a22oi_1 _1116_ (.Y(_0469_),
    .B1(_0436_),
    .B2(\bin_array[25][1] ),
    .A2(_0429_),
    .A1(\bin_array[29][1] ));
 sg13g2_a22oi_1 _1117_ (.Y(_0470_),
    .B1(_0424_),
    .B2(\bin_array[3][1] ),
    .A2(_0406_),
    .A1(\bin_array[10][1] ));
 sg13g2_nand4_1 _1118_ (.B(_0468_),
    .C(_0469_),
    .A(_0467_),
    .Y(_0471_),
    .D(_0470_));
 sg13g2_a22oi_1 _1119_ (.Y(_0472_),
    .B1(_0428_),
    .B2(\bin_array[12][1] ),
    .A2(_0405_),
    .A1(\bin_array[19][1] ));
 sg13g2_a22oi_1 _1120_ (.Y(_0473_),
    .B1(_0425_),
    .B2(\bin_array[24][1] ),
    .A2(_0402_),
    .A1(\bin_array[4][1] ));
 sg13g2_a22oi_1 _1121_ (.Y(_0474_),
    .B1(_0421_),
    .B2(\bin_array[21][1] ),
    .A2(_0413_),
    .A1(\bin_array[6][1] ));
 sg13g2_a22oi_1 _1122_ (.Y(_0475_),
    .B1(_0435_),
    .B2(\bin_array[8][1] ),
    .A2(_0432_),
    .A1(\bin_array[11][1] ));
 sg13g2_nand4_1 _1123_ (.B(_0473_),
    .C(_0474_),
    .A(_0472_),
    .Y(_0476_),
    .D(_0475_));
 sg13g2_a22oi_1 _1124_ (.Y(_0477_),
    .B1(_0426_),
    .B2(\bin_array[14][1] ),
    .A2(_0385_),
    .A1(\bin_array[31][1] ));
 sg13g2_a22oi_1 _1125_ (.Y(_0478_),
    .B1(_0427_),
    .B2(\bin_array[30][1] ),
    .A2(_0403_),
    .A1(\bin_array[15][1] ));
 sg13g2_nand2_1 _1126_ (.Y(_0479_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_nor3_1 _1127_ (.A(_0471_),
    .B(_0476_),
    .C(_0479_),
    .Y(_0480_));
 sg13g2_a221oi_1 _1128_ (.B2(_0480_),
    .C1(_0389_),
    .B1(_0466_),
    .A1(_0002_),
    .Y(_0481_),
    .A2(_0419_));
 sg13g2_a21o_1 _1129_ (.A2(_0391_),
    .A1(net93),
    .B1(_0481_),
    .X(_0011_));
 sg13g2_a22oi_1 _1130_ (.Y(_0482_),
    .B1(_0421_),
    .B2(\bin_array[21][2] ),
    .A2(_0397_),
    .A1(\bin_array[28][2] ));
 sg13g2_nand2_1 _1131_ (.Y(_0483_),
    .A(\bin_array[23][2] ),
    .B(_0420_));
 sg13g2_a22oi_1 _1132_ (.Y(_0484_),
    .B1(_0428_),
    .B2(\bin_array[12][2] ),
    .A2(_0399_),
    .A1(\bin_array[27][2] ));
 sg13g2_a22oi_1 _1133_ (.Y(_0485_),
    .B1(_0432_),
    .B2(\bin_array[11][2] ),
    .A2(_0425_),
    .A1(\bin_array[24][2] ));
 sg13g2_a22oi_1 _1134_ (.Y(_0486_),
    .B1(_0434_),
    .B2(\bin_array[20][2] ),
    .A2(_0410_),
    .A1(\bin_array[1][2] ));
 sg13g2_a22oi_1 _1135_ (.Y(_0487_),
    .B1(_0433_),
    .B2(\bin_array[13][2] ),
    .A2(_0413_),
    .A1(\bin_array[6][2] ));
 sg13g2_a22oi_1 _1136_ (.Y(_0488_),
    .B1(_0414_),
    .B2(\bin_array[7][2] ),
    .A2(_0408_),
    .A1(\bin_array[2][2] ));
 sg13g2_nand4_1 _1137_ (.B(_0486_),
    .C(_0487_),
    .A(_0484_),
    .Y(_0489_),
    .D(_0488_));
 sg13g2_nand3_1 _1138_ (.B(_0483_),
    .C(_0485_),
    .A(_0418_),
    .Y(_0490_));
 sg13g2_nor2_1 _1139_ (.A(_0489_),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_a22oi_1 _1140_ (.Y(_0492_),
    .B1(_0424_),
    .B2(\bin_array[3][2] ),
    .A2(_0406_),
    .A1(\bin_array[10][2] ));
 sg13g2_a22oi_1 _1141_ (.Y(_0493_),
    .B1(_0422_),
    .B2(\bin_array[18][2] ),
    .A2(_0407_),
    .A1(\bin_array[5][2] ));
 sg13g2_a22oi_1 _1142_ (.Y(_0494_),
    .B1(_0405_),
    .B2(\bin_array[19][2] ),
    .A2(_0402_),
    .A1(\bin_array[4][2] ));
 sg13g2_nand4_1 _1143_ (.B(_0492_),
    .C(_0493_),
    .A(_0482_),
    .Y(_0495_),
    .D(_0494_));
 sg13g2_a22oi_1 _1144_ (.Y(_0496_),
    .B1(_0436_),
    .B2(\bin_array[25][2] ),
    .A2(_0435_),
    .A1(\bin_array[8][2] ));
 sg13g2_a22oi_1 _1145_ (.Y(_0497_),
    .B1(_0431_),
    .B2(\bin_array[17][2] ),
    .A2(_0412_),
    .A1(\bin_array[16][2] ));
 sg13g2_a22oi_1 _1146_ (.Y(_0498_),
    .B1(_0409_),
    .B2(\bin_array[26][2] ),
    .A2(_0401_),
    .A1(\bin_array[9][2] ));
 sg13g2_a22oi_1 _1147_ (.Y(_0499_),
    .B1(_0429_),
    .B2(\bin_array[29][2] ),
    .A2(_0395_),
    .A1(\bin_array[22][2] ));
 sg13g2_nand4_1 _1148_ (.B(_0497_),
    .C(_0498_),
    .A(_0496_),
    .Y(_0500_),
    .D(_0499_));
 sg13g2_a22oi_1 _1149_ (.Y(_0501_),
    .B1(_0427_),
    .B2(\bin_array[30][2] ),
    .A2(_0385_),
    .A1(\bin_array[31][2] ));
 sg13g2_a22oi_1 _1150_ (.Y(_0502_),
    .B1(_0426_),
    .B2(\bin_array[14][2] ),
    .A2(_0403_),
    .A1(\bin_array[15][2] ));
 sg13g2_nand2_1 _1151_ (.Y(_0503_),
    .A(_0501_),
    .B(_0502_));
 sg13g2_nor3_1 _1152_ (.A(_0495_),
    .B(_0500_),
    .C(_0503_),
    .Y(_0504_));
 sg13g2_a221oi_1 _1153_ (.B2(_0504_),
    .C1(_0389_),
    .B1(_0491_),
    .A1(_0003_),
    .Y(_0505_),
    .A2(_0419_));
 sg13g2_a21o_1 _1154_ (.A2(_0391_),
    .A1(net60),
    .B1(_0505_),
    .X(_0012_));
 sg13g2_nand2_1 _1155_ (.Y(_0506_),
    .A(\bin_array[11][3] ),
    .B(_0432_));
 sg13g2_a22oi_1 _1156_ (.Y(_0507_),
    .B1(_0434_),
    .B2(\bin_array[20][3] ),
    .A2(_0428_),
    .A1(\bin_array[12][3] ));
 sg13g2_a22oi_1 _1157_ (.Y(_0508_),
    .B1(_0429_),
    .B2(\bin_array[29][3] ),
    .A2(_0412_),
    .A1(\bin_array[16][3] ));
 sg13g2_a22oi_1 _1158_ (.Y(_0509_),
    .B1(_0424_),
    .B2(\bin_array[3][3] ),
    .A2(_0414_),
    .A1(\bin_array[7][3] ));
 sg13g2_a22oi_1 _1159_ (.Y(_0510_),
    .B1(_0406_),
    .B2(\bin_array[10][3] ),
    .A2(_0397_),
    .A1(\bin_array[28][3] ));
 sg13g2_nand4_1 _1160_ (.B(_0508_),
    .C(_0509_),
    .A(_0507_),
    .Y(_0511_),
    .D(_0510_));
 sg13g2_a22oi_1 _1161_ (.Y(_0512_),
    .B1(_0409_),
    .B2(\bin_array[26][3] ),
    .A2(_0395_),
    .A1(\bin_array[22][3] ));
 sg13g2_nand3_1 _1162_ (.B(_0506_),
    .C(_0512_),
    .A(_0418_),
    .Y(_0513_));
 sg13g2_nor2_1 _1163_ (.A(_0511_),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_a22oi_1 _1164_ (.Y(_0515_),
    .B1(_0420_),
    .B2(\bin_array[23][3] ),
    .A2(_0410_),
    .A1(\bin_array[1][3] ));
 sg13g2_a22oi_1 _1165_ (.Y(_0516_),
    .B1(_0421_),
    .B2(\bin_array[21][3] ),
    .A2(_0407_),
    .A1(\bin_array[5][3] ));
 sg13g2_a22oi_1 _1166_ (.Y(_0517_),
    .B1(_0433_),
    .B2(\bin_array[13][3] ),
    .A2(_0402_),
    .A1(\bin_array[4][3] ));
 sg13g2_a22oi_1 _1167_ (.Y(_0518_),
    .B1(_0435_),
    .B2(\bin_array[8][3] ),
    .A2(_0425_),
    .A1(\bin_array[24][3] ));
 sg13g2_nand4_1 _1168_ (.B(_0516_),
    .C(_0517_),
    .A(_0515_),
    .Y(_0519_),
    .D(_0518_));
 sg13g2_a22oi_1 _1169_ (.Y(_0520_),
    .B1(_0431_),
    .B2(\bin_array[17][3] ),
    .A2(_0413_),
    .A1(\bin_array[6][3] ));
 sg13g2_a22oi_1 _1170_ (.Y(_0521_),
    .B1(_0401_),
    .B2(\bin_array[9][3] ),
    .A2(_0399_),
    .A1(\bin_array[27][3] ));
 sg13g2_a22oi_1 _1171_ (.Y(_0522_),
    .B1(_0408_),
    .B2(\bin_array[2][3] ),
    .A2(_0405_),
    .A1(\bin_array[19][3] ));
 sg13g2_a22oi_1 _1172_ (.Y(_0523_),
    .B1(_0436_),
    .B2(\bin_array[25][3] ),
    .A2(_0422_),
    .A1(\bin_array[18][3] ));
 sg13g2_nand4_1 _1173_ (.B(_0521_),
    .C(_0522_),
    .A(_0520_),
    .Y(_0524_),
    .D(_0523_));
 sg13g2_a22oi_1 _1174_ (.Y(_0525_),
    .B1(_0427_),
    .B2(\bin_array[30][3] ),
    .A2(_0385_),
    .A1(\bin_array[31][3] ));
 sg13g2_a22oi_1 _1175_ (.Y(_0526_),
    .B1(_0426_),
    .B2(\bin_array[14][3] ),
    .A2(_0403_),
    .A1(\bin_array[15][3] ));
 sg13g2_nand2_1 _1176_ (.Y(_0527_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_nor3_1 _1177_ (.A(_0519_),
    .B(_0524_),
    .C(_0527_),
    .Y(_0528_));
 sg13g2_a221oi_1 _1178_ (.B2(_0528_),
    .C1(_0389_),
    .B1(_0514_),
    .A1(_0004_),
    .Y(_0529_),
    .A2(_0419_));
 sg13g2_a21o_1 _1179_ (.A2(_0391_),
    .A1(net86),
    .B1(_0529_),
    .X(_0013_));
 sg13g2_or2_1 _1180_ (.X(_0530_),
    .B(net31),
    .A(net29));
 sg13g2_nand2_1 _1181_ (.Y(_0531_),
    .A(_0378_),
    .B(_0530_));
 sg13g2_nand2_2 _1182_ (.Y(_0532_),
    .A(net1),
    .B(_0530_));
 sg13g2_nor2_1 _1183_ (.A(_0377_),
    .B(_0532_),
    .Y(_0533_));
 sg13g2_nand2b_1 _1184_ (.Y(_0534_),
    .B(_0378_),
    .A_N(_0532_));
 sg13g2_a21oi_1 _1185_ (.A1(net528),
    .A2(net467),
    .Y(_0535_),
    .B1(net453));
 sg13g2_nor2_2 _1186_ (.A(net446),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_nor2_1 _1187_ (.A(net64),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_nand2_1 _1188_ (.Y(_0538_),
    .A(_0005_),
    .B(_0331_));
 sg13g2_a21oi_1 _1189_ (.A1(_0536_),
    .A2(net444),
    .Y(_0014_),
    .B1(_0537_));
 sg13g2_and2_1 _1190_ (.A(_0330_),
    .B(_0373_),
    .X(_0539_));
 sg13g2_o21ai_1 _1191_ (.B1(_0005_),
    .Y(_0540_),
    .A1(_0330_),
    .A2(_0373_));
 sg13g2_nor2_1 _1192_ (.A(_0539_),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_mux2_1 _1193_ (.A0(net85),
    .A1(net436),
    .S(_0536_),
    .X(_0015_));
 sg13g2_a21o_1 _1194_ (.A2(_0373_),
    .A1(_0330_),
    .B1(_0243_),
    .X(_0542_));
 sg13g2_nand3_1 _1195_ (.B(_0330_),
    .C(_0373_),
    .A(_0243_),
    .Y(_0543_));
 sg13g2_nand3_1 _1196_ (.B(_0542_),
    .C(_0543_),
    .A(_0005_),
    .Y(_0544_));
 sg13g2_nor2_1 _1197_ (.A(net75),
    .B(_0536_),
    .Y(_0545_));
 sg13g2_a21oi_1 _1198_ (.A1(_0536_),
    .A2(net430),
    .Y(_0016_),
    .B1(_0545_));
 sg13g2_a221oi_1 _1199_ (.B2(_0286_),
    .C1(_0154_),
    .B1(_0543_),
    .A1(_0287_),
    .Y(_0546_),
    .A2(_0539_));
 sg13g2_mux2_1 _1200_ (.A0(net59),
    .A1(net426),
    .S(_0536_),
    .X(_0017_));
 sg13g2_nand2_1 _1201_ (.Y(_0547_),
    .A(net1),
    .B(net453));
 sg13g2_nand2_1 _1202_ (.Y(_0548_),
    .A(\state[2] ),
    .B(_0378_));
 sg13g2_a22oi_1 _1203_ (.Y(_0549_),
    .B1(_0548_),
    .B2(_0531_),
    .A2(_0547_),
    .A1(_0375_));
 sg13g2_nor2_1 _1204_ (.A(_0153_),
    .B(net179),
    .Y(_0550_));
 sg13g2_mux2_1 _1205_ (.A0(net179),
    .A1(_0550_),
    .S(_0549_),
    .X(_0018_));
 sg13g2_and3_1 _1206_ (.X(_0551_),
    .A(\state[2] ),
    .B(_0381_),
    .C(net456));
 sg13g2_mux2_1 _1207_ (.A0(net175),
    .A1(_0551_),
    .S(_0549_),
    .X(_0019_));
 sg13g2_nand2b_1 _1208_ (.Y(_0552_),
    .B(_0381_),
    .A_N(net465));
 sg13g2_and3_1 _1209_ (.X(_0553_),
    .A(net177),
    .B(_0383_),
    .C(_0552_));
 sg13g2_mux2_1 _1210_ (.A0(net465),
    .A1(_0553_),
    .S(_0549_),
    .X(_0020_));
 sg13g2_nor2b_1 _1211_ (.A(net464),
    .B_N(_0383_),
    .Y(_0554_));
 sg13g2_nor3_1 _1212_ (.A(_0153_),
    .B(_0384_),
    .C(_0554_),
    .Y(_0555_));
 sg13g2_mux2_1 _1213_ (.A0(net464),
    .A1(_0555_),
    .S(_0549_),
    .X(_0021_));
 sg13g2_nor2_1 _1214_ (.A(net462),
    .B(_0384_),
    .Y(_0556_));
 sg13g2_nor3_1 _1215_ (.A(_0153_),
    .B(_0385_),
    .C(_0556_),
    .Y(_0557_));
 sg13g2_mux2_1 _1216_ (.A0(net462),
    .A1(_0557_),
    .S(_0549_),
    .X(_0022_));
 sg13g2_o21ai_1 _1217_ (.B1(_0532_),
    .Y(_0558_),
    .A1(net89),
    .A2(_0388_));
 sg13g2_inv_1 _1218_ (.Y(_0023_),
    .A(_0558_));
 sg13g2_nor3_1 _1219_ (.A(_0386_),
    .B(_0389_),
    .C(_0530_),
    .Y(_0559_));
 sg13g2_a22oi_1 _1220_ (.Y(_0560_),
    .B1(_0389_),
    .B2(_0532_),
    .A2(_0386_),
    .A1(\state[2] ));
 sg13g2_nand2b_1 _1221_ (.Y(_0561_),
    .B(net34),
    .A_N(_0560_));
 sg13g2_nand2b_1 _1222_ (.Y(_0024_),
    .B(net35),
    .A_N(_0559_));
 sg13g2_a21oi_1 _1223_ (.A1(_0375_),
    .A2(_0547_),
    .Y(_0562_),
    .B1(_0531_));
 sg13g2_mux2_1 _1224_ (.A0(net27),
    .A1(_0005_),
    .S(_0562_),
    .X(_0025_));
 sg13g2_o21ai_1 _1225_ (.B1(net450),
    .Y(_0563_),
    .A1(_0158_),
    .A2(net453));
 sg13g2_nand2_1 _1226_ (.Y(_0564_),
    .A(net50),
    .B(_0563_));
 sg13g2_o21ai_1 _1227_ (.B1(_0564_),
    .Y(_0026_),
    .A1(net441),
    .A2(_0563_));
 sg13g2_mux2_1 _1228_ (.A0(net439),
    .A1(net45),
    .S(_0563_),
    .X(_0027_));
 sg13g2_nand2_1 _1229_ (.Y(_0565_),
    .A(net25),
    .B(_0563_));
 sg13g2_o21ai_1 _1230_ (.B1(_0565_),
    .Y(_0028_),
    .A1(net434),
    .A2(_0563_));
 sg13g2_mux2_1 _1231_ (.A0(net425),
    .A1(net37),
    .S(_0563_),
    .X(_0029_));
 sg13g2_o21ai_1 _1232_ (.B1(net448),
    .Y(_0566_),
    .A1(_0166_),
    .A2(net451));
 sg13g2_nand2_1 _1233_ (.Y(_0567_),
    .A(net33),
    .B(_0566_));
 sg13g2_o21ai_1 _1234_ (.B1(_0567_),
    .Y(_0030_),
    .A1(net441),
    .A2(_0566_));
 sg13g2_mux2_1 _1235_ (.A0(net435),
    .A1(net134),
    .S(_0566_),
    .X(_0031_));
 sg13g2_nand2_1 _1236_ (.Y(_0568_),
    .A(net68),
    .B(_0566_));
 sg13g2_o21ai_1 _1237_ (.B1(_0568_),
    .Y(_0032_),
    .A1(net431),
    .A2(_0566_));
 sg13g2_mux2_1 _1238_ (.A0(net426),
    .A1(net107),
    .S(_0566_),
    .X(_0033_));
 sg13g2_o21ai_1 _1239_ (.B1(net449),
    .Y(_0569_),
    .A1(_0187_),
    .A2(net452));
 sg13g2_nand2_1 _1240_ (.Y(_0570_),
    .A(net80),
    .B(_0569_));
 sg13g2_o21ai_1 _1241_ (.B1(_0570_),
    .Y(_0034_),
    .A1(net442),
    .A2(_0569_));
 sg13g2_mux2_1 _1242_ (.A0(net438),
    .A1(net172),
    .S(_0569_),
    .X(_0035_));
 sg13g2_nand2_1 _1243_ (.Y(_0571_),
    .A(net53),
    .B(_0569_));
 sg13g2_o21ai_1 _1244_ (.B1(_0571_),
    .Y(_0036_),
    .A1(net433),
    .A2(_0569_));
 sg13g2_mux2_1 _1245_ (.A0(net427),
    .A1(net163),
    .S(_0569_),
    .X(_0037_));
 sg13g2_o21ai_1 _1246_ (.B1(net449),
    .Y(_0572_),
    .A1(_0181_),
    .A2(net452));
 sg13g2_nand2_1 _1247_ (.Y(_0573_),
    .A(net168),
    .B(_0572_));
 sg13g2_o21ai_1 _1248_ (.B1(_0573_),
    .Y(_0038_),
    .A1(net443),
    .A2(_0572_));
 sg13g2_mux2_1 _1249_ (.A0(net438),
    .A1(net156),
    .S(_0572_),
    .X(_0039_));
 sg13g2_nand2_1 _1250_ (.Y(_0574_),
    .A(net136),
    .B(_0572_));
 sg13g2_o21ai_1 _1251_ (.B1(_0574_),
    .Y(_0040_),
    .A1(net433),
    .A2(_0572_));
 sg13g2_mux2_1 _1252_ (.A0(net428),
    .A1(net180),
    .S(_0572_),
    .X(_0041_));
 sg13g2_o21ai_1 _1253_ (.B1(net449),
    .Y(_0575_),
    .A1(_0203_),
    .A2(net452));
 sg13g2_nand2_1 _1254_ (.Y(_0576_),
    .A(net116),
    .B(_0575_));
 sg13g2_o21ai_1 _1255_ (.B1(_0576_),
    .Y(_0042_),
    .A1(net443),
    .A2(_0575_));
 sg13g2_mux2_1 _1256_ (.A0(net437),
    .A1(net169),
    .S(_0575_),
    .X(_0043_));
 sg13g2_nand2_1 _1257_ (.Y(_0577_),
    .A(net142),
    .B(_0575_));
 sg13g2_o21ai_1 _1258_ (.B1(_0577_),
    .Y(_0044_),
    .A1(net433),
    .A2(_0575_));
 sg13g2_mux2_1 _1259_ (.A0(net428),
    .A1(net166),
    .S(_0575_),
    .X(_0045_));
 sg13g2_o21ai_1 _1260_ (.B1(net448),
    .Y(_0578_),
    .A1(_0211_),
    .A2(net451));
 sg13g2_nand2_1 _1261_ (.Y(_0579_),
    .A(net46),
    .B(_0578_));
 sg13g2_o21ai_1 _1262_ (.B1(_0579_),
    .Y(_0046_),
    .A1(net441),
    .A2(_0578_));
 sg13g2_mux2_1 _1263_ (.A0(net437),
    .A1(net129),
    .S(_0578_),
    .X(_0047_));
 sg13g2_nand2_1 _1264_ (.Y(_0580_),
    .A(net40),
    .B(_0578_));
 sg13g2_o21ai_1 _1265_ (.B1(_0580_),
    .Y(_0048_),
    .A1(net430),
    .A2(_0578_));
 sg13g2_mux2_1 _1266_ (.A0(net424),
    .A1(net162),
    .S(_0578_),
    .X(_0049_));
 sg13g2_o21ai_1 _1267_ (.B1(net449),
    .Y(_0581_),
    .A1(_0176_),
    .A2(net451));
 sg13g2_nand2_1 _1268_ (.Y(_0582_),
    .A(net110),
    .B(_0581_));
 sg13g2_o21ai_1 _1269_ (.B1(_0582_),
    .Y(_0050_),
    .A1(net443),
    .A2(_0581_));
 sg13g2_mux2_1 _1270_ (.A0(net437),
    .A1(net167),
    .S(_0581_),
    .X(_0051_));
 sg13g2_nand2_1 _1271_ (.Y(_0583_),
    .A(net49),
    .B(_0581_));
 sg13g2_o21ai_1 _1272_ (.B1(_0583_),
    .Y(_0052_),
    .A1(net432),
    .A2(_0581_));
 sg13g2_mux2_1 _1273_ (.A0(net427),
    .A1(net152),
    .S(_0581_),
    .X(_0053_));
 sg13g2_o21ai_1 _1274_ (.B1(net448),
    .Y(_0584_),
    .A1(_0172_),
    .A2(net451));
 sg13g2_nand2_1 _1275_ (.Y(_0585_),
    .A(net79),
    .B(_0584_));
 sg13g2_o21ai_1 _1276_ (.B1(_0585_),
    .Y(_0054_),
    .A1(net442),
    .A2(_0584_));
 sg13g2_mux2_1 _1277_ (.A0(net437),
    .A1(net173),
    .S(_0584_),
    .X(_0055_));
 sg13g2_nand2_1 _1278_ (.Y(_0586_),
    .A(net47),
    .B(_0584_));
 sg13g2_o21ai_1 _1279_ (.B1(_0586_),
    .Y(_0056_),
    .A1(net433),
    .A2(_0584_));
 sg13g2_mux2_1 _1280_ (.A0(net427),
    .A1(net155),
    .S(_0584_),
    .X(_0057_));
 sg13g2_o21ai_1 _1281_ (.B1(net448),
    .Y(_0587_),
    .A1(_0162_),
    .A2(net451));
 sg13g2_nand2_1 _1282_ (.Y(_0588_),
    .A(net66),
    .B(_0587_));
 sg13g2_o21ai_1 _1283_ (.B1(_0588_),
    .Y(_0058_),
    .A1(net442),
    .A2(_0587_));
 sg13g2_mux2_1 _1284_ (.A0(net438),
    .A1(net139),
    .S(_0587_),
    .X(_0059_));
 sg13g2_nand2_1 _1285_ (.Y(_0589_),
    .A(net54),
    .B(_0587_));
 sg13g2_o21ai_1 _1286_ (.B1(_0589_),
    .Y(_0060_),
    .A1(net432),
    .A2(_0587_));
 sg13g2_mux2_1 _1287_ (.A0(net427),
    .A1(net170),
    .S(_0587_),
    .X(_0061_));
 sg13g2_o21ai_1 _1288_ (.B1(net448),
    .Y(_0590_),
    .A1(_0229_),
    .A2(net451));
 sg13g2_nand2_1 _1289_ (.Y(_0591_),
    .A(net58),
    .B(_0590_));
 sg13g2_o21ai_1 _1290_ (.B1(_0591_),
    .Y(_0062_),
    .A1(net442),
    .A2(_0590_));
 sg13g2_mux2_1 _1291_ (.A0(net438),
    .A1(net126),
    .S(_0590_),
    .X(_0063_));
 sg13g2_nand2_1 _1292_ (.Y(_0592_),
    .A(net76),
    .B(_0590_));
 sg13g2_o21ai_1 _1293_ (.B1(_0592_),
    .Y(_0064_),
    .A1(net432),
    .A2(_0590_));
 sg13g2_mux2_1 _1294_ (.A0(net427),
    .A1(net114),
    .S(_0590_),
    .X(_0065_));
 sg13g2_o21ai_1 _1295_ (.B1(net448),
    .Y(_0593_),
    .A1(_0179_),
    .A2(net452));
 sg13g2_nand2_1 _1296_ (.Y(_0594_),
    .A(net115),
    .B(_0593_));
 sg13g2_o21ai_1 _1297_ (.B1(_0594_),
    .Y(_0066_),
    .A1(net443),
    .A2(_0593_));
 sg13g2_mux2_1 _1298_ (.A0(net437),
    .A1(net141),
    .S(_0593_),
    .X(_0067_));
 sg13g2_nand2_1 _1299_ (.Y(_0595_),
    .A(net51),
    .B(_0593_));
 sg13g2_o21ai_1 _1300_ (.B1(_0595_),
    .Y(_0068_),
    .A1(net432),
    .A2(_0593_));
 sg13g2_mux2_1 _1301_ (.A0(net428),
    .A1(net160),
    .S(_0593_),
    .X(_0069_));
 sg13g2_o21ai_1 _1302_ (.B1(net448),
    .Y(_0596_),
    .A1(_0194_),
    .A2(net451));
 sg13g2_nand2_1 _1303_ (.Y(_0597_),
    .A(net90),
    .B(_0596_));
 sg13g2_o21ai_1 _1304_ (.B1(_0597_),
    .Y(_0070_),
    .A1(net443),
    .A2(_0596_));
 sg13g2_mux2_1 _1305_ (.A0(net437),
    .A1(net174),
    .S(_0596_),
    .X(_0071_));
 sg13g2_nand2_1 _1306_ (.Y(_0598_),
    .A(net132),
    .B(_0596_));
 sg13g2_o21ai_1 _1307_ (.B1(_0598_),
    .Y(_0072_),
    .A1(net433),
    .A2(_0596_));
 sg13g2_mux2_1 _1308_ (.A0(net428),
    .A1(net153),
    .S(_0596_),
    .X(_0073_));
 sg13g2_o21ai_1 _1309_ (.B1(net448),
    .Y(_0599_),
    .A1(_0199_),
    .A2(net451));
 sg13g2_nand2_1 _1310_ (.Y(_0600_),
    .A(net55),
    .B(_0599_));
 sg13g2_o21ai_1 _1311_ (.B1(_0600_),
    .Y(_0074_),
    .A1(net442),
    .A2(_0599_));
 sg13g2_mux2_1 _1312_ (.A0(net437),
    .A1(net164),
    .S(_0599_),
    .X(_0075_));
 sg13g2_nand2_1 _1313_ (.Y(_0601_),
    .A(net52),
    .B(_0599_));
 sg13g2_o21ai_1 _1314_ (.B1(_0601_),
    .Y(_0076_),
    .A1(net433),
    .A2(_0599_));
 sg13g2_mux2_1 _1315_ (.A0(net427),
    .A1(net151),
    .S(_0599_),
    .X(_0077_));
 sg13g2_o21ai_1 _1316_ (.B1(net449),
    .Y(_0602_),
    .A1(_0218_),
    .A2(net452));
 sg13g2_nand2_1 _1317_ (.Y(_0603_),
    .A(net125),
    .B(_0602_));
 sg13g2_o21ai_1 _1318_ (.B1(_0603_),
    .Y(_0078_),
    .A1(net443),
    .A2(_0602_));
 sg13g2_mux2_1 _1319_ (.A0(net437),
    .A1(net171),
    .S(_0602_),
    .X(_0079_));
 sg13g2_nand2_1 _1320_ (.Y(_0604_),
    .A(net117),
    .B(_0602_));
 sg13g2_o21ai_1 _1321_ (.B1(_0604_),
    .Y(_0080_),
    .A1(net433),
    .A2(_0602_));
 sg13g2_mux2_1 _1322_ (.A0(net428),
    .A1(net161),
    .S(_0602_),
    .X(_0081_));
 sg13g2_o21ai_1 _1323_ (.B1(net450),
    .Y(_0605_),
    .A1(_0220_),
    .A2(net453));
 sg13g2_nand2_1 _1324_ (.Y(_0606_),
    .A(net98),
    .B(_0605_));
 sg13g2_o21ai_1 _1325_ (.B1(_0606_),
    .Y(_0082_),
    .A1(net441),
    .A2(_0605_));
 sg13g2_mux2_1 _1326_ (.A0(net436),
    .A1(net138),
    .S(_0605_),
    .X(_0083_));
 sg13g2_nand2_1 _1327_ (.Y(_0607_),
    .A(net41),
    .B(_0605_));
 sg13g2_o21ai_1 _1328_ (.B1(_0607_),
    .Y(_0084_),
    .A1(net430),
    .A2(_0605_));
 sg13g2_mux2_1 _1329_ (.A0(net425),
    .A1(net120),
    .S(_0605_),
    .X(_0085_));
 sg13g2_a21oi_1 _1330_ (.A1(net511),
    .A2(net467),
    .Y(_0608_),
    .B1(net453));
 sg13g2_nand2b_2 _1331_ (.Y(_0609_),
    .B(net450),
    .A_N(_0608_));
 sg13g2_nand2_1 _1332_ (.Y(_0610_),
    .A(net39),
    .B(_0609_));
 sg13g2_o21ai_1 _1333_ (.B1(_0610_),
    .Y(_0086_),
    .A1(net441),
    .A2(_0609_));
 sg13g2_mux2_1 _1334_ (.A0(net436),
    .A1(net131),
    .S(_0609_),
    .X(_0087_));
 sg13g2_nand2_1 _1335_ (.Y(_0611_),
    .A(net38),
    .B(_0609_));
 sg13g2_o21ai_1 _1336_ (.B1(_0611_),
    .Y(_0088_),
    .A1(net430),
    .A2(_0609_));
 sg13g2_mux2_1 _1337_ (.A0(net426),
    .A1(net82),
    .S(_0609_),
    .X(_0089_));
 sg13g2_a21oi_2 _1338_ (.B1(net445),
    .Y(_0612_),
    .A2(net454),
    .A1(_0190_));
 sg13g2_nor2_1 _1339_ (.A(net130),
    .B(_0612_),
    .Y(_0613_));
 sg13g2_a21oi_1 _1340_ (.A1(net441),
    .A2(_0612_),
    .Y(_0090_),
    .B1(_0613_));
 sg13g2_mux2_1 _1341_ (.A0(net102),
    .A1(net435),
    .S(_0612_),
    .X(_0091_));
 sg13g2_nor2_1 _1342_ (.A(net144),
    .B(_0612_),
    .Y(_0614_));
 sg13g2_a21oi_1 _1343_ (.A1(net431),
    .A2(_0612_),
    .Y(_0092_),
    .B1(_0614_));
 sg13g2_mux2_1 _1344_ (.A0(net99),
    .A1(net424),
    .S(_0612_),
    .X(_0093_));
 sg13g2_a21oi_2 _1345_ (.B1(net445),
    .Y(_0615_),
    .A2(net454),
    .A1(_0196_));
 sg13g2_nor2_1 _1346_ (.A(net74),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_a21oi_1 _1347_ (.A1(net440),
    .A2(_0615_),
    .Y(_0094_),
    .B1(_0616_));
 sg13g2_mux2_1 _1348_ (.A0(net84),
    .A1(net435),
    .S(_0615_),
    .X(_0095_));
 sg13g2_nor2_1 _1349_ (.A(net73),
    .B(_0615_),
    .Y(_0617_));
 sg13g2_a21oi_1 _1350_ (.A1(net431),
    .A2(_0615_),
    .Y(_0096_),
    .B1(_0617_));
 sg13g2_mux2_1 _1351_ (.A0(net106),
    .A1(net425),
    .S(_0615_),
    .X(_0097_));
 sg13g2_a21oi_2 _1352_ (.B1(net445),
    .Y(_0618_),
    .A2(net454),
    .A1(_0225_));
 sg13g2_nor2_1 _1353_ (.A(net105),
    .B(_0618_),
    .Y(_0619_));
 sg13g2_a21oi_1 _1354_ (.A1(net440),
    .A2(_0618_),
    .Y(_0098_),
    .B1(_0619_));
 sg13g2_mux2_1 _1355_ (.A0(net112),
    .A1(net435),
    .S(_0618_),
    .X(_0099_));
 sg13g2_nor2_1 _1356_ (.A(net92),
    .B(_0618_),
    .Y(_0620_));
 sg13g2_a21oi_1 _1357_ (.A1(net431),
    .A2(_0618_),
    .Y(_0100_),
    .B1(_0620_));
 sg13g2_mux2_1 _1358_ (.A0(net143),
    .A1(net424),
    .S(_0618_),
    .X(_0101_));
 sg13g2_a21oi_2 _1359_ (.B1(net447),
    .Y(_0621_),
    .A2(net455),
    .A1(_0222_));
 sg13g2_nor2_1 _1360_ (.A(net78),
    .B(_0621_),
    .Y(_0622_));
 sg13g2_a21oi_1 _1361_ (.A1(net440),
    .A2(_0621_),
    .Y(_0102_),
    .B1(_0622_));
 sg13g2_mux2_1 _1362_ (.A0(net145),
    .A1(net438),
    .S(_0621_),
    .X(_0103_));
 sg13g2_nor2_1 _1363_ (.A(net159),
    .B(_0621_),
    .Y(_0623_));
 sg13g2_a21oi_1 _1364_ (.A1(net431),
    .A2(_0621_),
    .Y(_0104_),
    .B1(_0623_));
 sg13g2_mux2_1 _1365_ (.A0(net81),
    .A1(net424),
    .S(_0621_),
    .X(_0105_));
 sg13g2_a21oi_2 _1366_ (.B1(net445),
    .Y(_0624_),
    .A2(net454),
    .A1(_0227_));
 sg13g2_nor2_1 _1367_ (.A(net113),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_a21oi_1 _1368_ (.A1(net440),
    .A2(_0624_),
    .Y(_0106_),
    .B1(_0625_));
 sg13g2_mux2_1 _1369_ (.A0(net148),
    .A1(net435),
    .S(_0624_),
    .X(_0107_));
 sg13g2_nor2_1 _1370_ (.A(net77),
    .B(_0624_),
    .Y(_0626_));
 sg13g2_a21oi_1 _1371_ (.A1(net431),
    .A2(_0624_),
    .Y(_0108_),
    .B1(_0626_));
 sg13g2_mux2_1 _1372_ (.A0(net122),
    .A1(net424),
    .S(_0624_),
    .X(_0109_));
 sg13g2_a21oi_2 _1373_ (.B1(net445),
    .Y(_0627_),
    .A2(net455),
    .A1(_0239_));
 sg13g2_nor2_1 _1374_ (.A(net109),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_a21oi_1 _1375_ (.A1(net440),
    .A2(_0627_),
    .Y(_0110_),
    .B1(_0628_));
 sg13g2_mux2_1 _1376_ (.A0(net158),
    .A1(net436),
    .S(_0627_),
    .X(_0111_));
 sg13g2_nor2_1 _1377_ (.A(net128),
    .B(_0627_),
    .Y(_0629_));
 sg13g2_a21oi_1 _1378_ (.A1(net430),
    .A2(_0627_),
    .Y(_0112_),
    .B1(_0629_));
 sg13g2_mux2_1 _1379_ (.A0(net149),
    .A1(net424),
    .S(_0627_),
    .X(_0113_));
 sg13g2_a21oi_2 _1380_ (.B1(net445),
    .Y(_0630_),
    .A2(net454),
    .A1(_0231_));
 sg13g2_nor2_1 _1381_ (.A(net127),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_a21oi_1 _1382_ (.A1(net440),
    .A2(_0630_),
    .Y(_0114_),
    .B1(_0631_));
 sg13g2_mux2_1 _1383_ (.A0(net150),
    .A1(net435),
    .S(_0630_),
    .X(_0115_));
 sg13g2_nor2_1 _1384_ (.A(net154),
    .B(_0630_),
    .Y(_0632_));
 sg13g2_a21oi_1 _1385_ (.A1(net431),
    .A2(_0630_),
    .Y(_0116_),
    .B1(_0632_));
 sg13g2_mux2_1 _1386_ (.A0(net101),
    .A1(net424),
    .S(_0630_),
    .X(_0117_));
 sg13g2_a21oi_2 _1387_ (.B1(net446),
    .Y(_0633_),
    .A2(net455),
    .A1(_0236_));
 sg13g2_nor2_1 _1388_ (.A(net118),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_a21oi_1 _1389_ (.A1(net444),
    .A2(_0633_),
    .Y(_0118_),
    .B1(_0634_));
 sg13g2_mux2_1 _1390_ (.A0(net121),
    .A1(net436),
    .S(_0633_),
    .X(_0119_));
 sg13g2_nor2_1 _1391_ (.A(net91),
    .B(_0633_),
    .Y(_0635_));
 sg13g2_a21oi_1 _1392_ (.A1(net430),
    .A2(_0633_),
    .Y(_0120_),
    .B1(_0635_));
 sg13g2_mux2_1 _1393_ (.A0(net88),
    .A1(net426),
    .S(_0633_),
    .X(_0121_));
 sg13g2_a21oi_2 _1394_ (.B1(net446),
    .Y(_0636_),
    .A2(net455),
    .A1(_0234_));
 sg13g2_nor2_1 _1395_ (.A(net103),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_a21oi_1 _1396_ (.A1(net444),
    .A2(_0636_),
    .Y(_0122_),
    .B1(_0637_));
 sg13g2_mux2_1 _1397_ (.A0(net146),
    .A1(net436),
    .S(_0636_),
    .X(_0123_));
 sg13g2_nor2_1 _1398_ (.A(net96),
    .B(_0636_),
    .Y(_0638_));
 sg13g2_a21oi_1 _1399_ (.A1(net430),
    .A2(_0636_),
    .Y(_0124_),
    .B1(_0638_));
 sg13g2_mux2_1 _1400_ (.A0(net95),
    .A1(net425),
    .S(_0636_),
    .X(_0125_));
 sg13g2_a21oi_2 _1401_ (.B1(net445),
    .Y(_0639_),
    .A2(net454),
    .A1(_0192_));
 sg13g2_nor2_1 _1402_ (.A(net133),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_a21oi_1 _1403_ (.A1(net440),
    .A2(_0639_),
    .Y(_0126_),
    .B1(_0640_));
 sg13g2_mux2_1 _1404_ (.A0(net157),
    .A1(net435),
    .S(_0639_),
    .X(_0127_));
 sg13g2_nor2_1 _1405_ (.A(net63),
    .B(_0639_),
    .Y(_0641_));
 sg13g2_a21oi_1 _1406_ (.A1(net432),
    .A2(_0639_),
    .Y(_0128_),
    .B1(_0641_));
 sg13g2_mux2_1 _1407_ (.A0(net147),
    .A1(net425),
    .S(_0639_),
    .X(_0129_));
 sg13g2_a21oi_2 _1408_ (.B1(net445),
    .Y(_0642_),
    .A2(net454),
    .A1(_0215_));
 sg13g2_nor2_1 _1409_ (.A(net100),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_a21oi_1 _1410_ (.A1(net440),
    .A2(_0642_),
    .Y(_0130_),
    .B1(_0643_));
 sg13g2_mux2_1 _1411_ (.A0(net62),
    .A1(net435),
    .S(_0642_),
    .X(_0131_));
 sg13g2_nor2_1 _1412_ (.A(net111),
    .B(_0642_),
    .Y(_0644_));
 sg13g2_a21oi_1 _1413_ (.A1(net431),
    .A2(_0642_),
    .Y(_0132_),
    .B1(_0644_));
 sg13g2_mux2_1 _1414_ (.A0(net67),
    .A1(net424),
    .S(_0642_),
    .X(_0133_));
 sg13g2_a21oi_2 _1415_ (.B1(net447),
    .Y(_0645_),
    .A2(net455),
    .A1(_0205_));
 sg13g2_nor2_1 _1416_ (.A(net108),
    .B(_0645_),
    .Y(_0646_));
 sg13g2_a21oi_1 _1417_ (.A1(net442),
    .A2(_0645_),
    .Y(_0134_),
    .B1(_0646_));
 sg13g2_mux2_1 _1418_ (.A0(net71),
    .A1(net438),
    .S(_0645_),
    .X(_0135_));
 sg13g2_nor2_1 _1419_ (.A(net56),
    .B(_0645_),
    .Y(_0647_));
 sg13g2_a21oi_1 _1420_ (.A1(net432),
    .A2(_0645_),
    .Y(_0136_),
    .B1(_0647_));
 sg13g2_mux2_1 _1421_ (.A0(net57),
    .A1(net427),
    .S(_0645_),
    .X(_0137_));
 sg13g2_a21oi_2 _1422_ (.B1(net447),
    .Y(_0648_),
    .A2(net455),
    .A1(_0201_));
 sg13g2_nor2_1 _1423_ (.A(net140),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_a21oi_1 _1424_ (.A1(net442),
    .A2(_0648_),
    .Y(_0138_),
    .B1(_0649_));
 sg13g2_mux2_1 _1425_ (.A0(net83),
    .A1(net438),
    .S(_0648_),
    .X(_0139_));
 sg13g2_nor2_1 _1426_ (.A(net137),
    .B(_0648_),
    .Y(_0650_));
 sg13g2_a21oi_1 _1427_ (.A1(net432),
    .A2(_0648_),
    .Y(_0140_),
    .B1(_0650_));
 sg13g2_mux2_1 _1428_ (.A0(net135),
    .A1(net427),
    .S(_0648_),
    .X(_0141_));
 sg13g2_a21oi_2 _1429_ (.B1(net447),
    .Y(_0651_),
    .A2(net455),
    .A1(_0185_));
 sg13g2_nor2_1 _1430_ (.A(net97),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_a21oi_1 _1431_ (.A1(net442),
    .A2(_0651_),
    .Y(_0142_),
    .B1(_0652_));
 sg13g2_mux2_1 _1432_ (.A0(net165),
    .A1(net438),
    .S(_0651_),
    .X(_0143_));
 sg13g2_nor2_1 _1433_ (.A(net124),
    .B(_0651_),
    .Y(_0653_));
 sg13g2_a21oi_1 _1434_ (.A1(net432),
    .A2(_0651_),
    .Y(_0144_),
    .B1(_0653_));
 sg13g2_mux2_1 _1435_ (.A0(net69),
    .A1(net425),
    .S(_0651_),
    .X(_0145_));
 sg13g2_a21oi_2 _1436_ (.B1(net446),
    .Y(_0654_),
    .A2(net454),
    .A1(_0209_));
 sg13g2_nor2_1 _1437_ (.A(net48),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_a21oi_1 _1438_ (.A1(net441),
    .A2(_0654_),
    .Y(_0146_),
    .B1(_0655_));
 sg13g2_mux2_1 _1439_ (.A0(net123),
    .A1(net436),
    .S(_0654_),
    .X(_0147_));
 sg13g2_nor2_1 _1440_ (.A(net72),
    .B(_0654_),
    .Y(_0656_));
 sg13g2_a21oi_1 _1441_ (.A1(net430),
    .A2(_0654_),
    .Y(_0148_),
    .B1(_0656_));
 sg13g2_mux2_1 _1442_ (.A0(net70),
    .A1(net425),
    .S(_0654_),
    .X(_0149_));
 sg13g2_dfrbp_1 _1443_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net559),
    .D(net32),
    .Q_N(\state[0] ),
    .Q(_0007_));
 sg13g2_dfrbp_1 _1444_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net558),
    .D(net30),
    .Q_N(_0005_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _1445_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net559),
    .D(net178),
    .Q_N(_0792_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _1446_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net558),
    .D(net44),
    .Q_N(_0791_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1447_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net558),
    .D(net94),
    .Q_N(_0790_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1448_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net558),
    .D(net61),
    .Q_N(_0789_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1449_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net550),
    .D(net87),
    .Q_N(_0788_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1450_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net548),
    .D(net65),
    .Q_N(_0787_),
    .Q(\bin_array[31][0] ));
 sg13g2_dfrbp_1 _1451_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net548),
    .D(_0015_),
    .Q_N(_0786_),
    .Q(\bin_array[31][1] ));
 sg13g2_dfrbp_1 _1452_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net548),
    .D(_0016_),
    .Q_N(_0785_),
    .Q(\bin_array[31][2] ));
 sg13g2_dfrbp_1 _1453_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net548),
    .D(_0017_),
    .Q_N(_0784_),
    .Q(\bin_array[31][3] ));
 sg13g2_dfrbp_1 _1454_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net559),
    .D(_0018_),
    .Q_N(_0783_),
    .Q(\shift_count[0] ));
 sg13g2_dfrbp_1 _1455_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net559),
    .D(net176),
    .Q_N(_0782_),
    .Q(\shift_count[1] ));
 sg13g2_dfrbp_1 _1456_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net558),
    .D(_0020_),
    .Q_N(_0781_),
    .Q(\shift_count[2] ));
 sg13g2_dfrbp_1 _1457_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net558),
    .D(_0021_),
    .Q_N(_0780_),
    .Q(\shift_count[3] ));
 sg13g2_dfrbp_1 _1458_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net558),
    .D(_0022_),
    .Q_N(_0006_),
    .Q(\shift_count[4] ));
 sg13g2_dfrbp_1 _1459_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net549),
    .D(_0023_),
    .Q_N(_0779_),
    .Q(valid_out_reg));
 sg13g2_dfrbp_1 _1460_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net549),
    .D(net36),
    .Q_N(_0778_),
    .Q(last_bin_reg));
 sg13g2_dfrbp_1 _1461_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net559),
    .D(net28),
    .Q_N(ready_reg),
    .Q(_0008_));
 sg13g2_dfrbp_1 _1462_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net549),
    .D(_0026_),
    .Q_N(_0777_),
    .Q(\bin_array[0][0] ));
 sg13g2_dfrbp_1 _1463_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net558),
    .D(_0027_),
    .Q_N(_0002_),
    .Q(\bin_array[0][1] ));
 sg13g2_dfrbp_1 _1464_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net550),
    .D(net26),
    .Q_N(_0003_),
    .Q(\bin_array[0][2] ));
 sg13g2_dfrbp_1 _1465_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net550),
    .D(_0029_),
    .Q_N(_0004_),
    .Q(\bin_array[0][3] ));
 sg13g2_dfrbp_1 _1466_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net545),
    .D(_0030_),
    .Q_N(_0776_),
    .Q(\bin_array[1][0] ));
 sg13g2_dfrbp_1 _1467_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net541),
    .D(_0031_),
    .Q_N(_0775_),
    .Q(\bin_array[1][1] ));
 sg13g2_dfrbp_1 _1468_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net541),
    .D(_0032_),
    .Q_N(_0774_),
    .Q(\bin_array[1][2] ));
 sg13g2_dfrbp_1 _1469_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net547),
    .D(_0033_),
    .Q_N(_0773_),
    .Q(\bin_array[1][3] ));
 sg13g2_dfrbp_1 _1470_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net554),
    .D(_0034_),
    .Q_N(_0772_),
    .Q(\bin_array[2][0] ));
 sg13g2_dfrbp_1 _1471_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net554),
    .D(_0035_),
    .Q_N(_0771_),
    .Q(\bin_array[2][1] ));
 sg13g2_dfrbp_1 _1472_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net554),
    .D(_0036_),
    .Q_N(_0770_),
    .Q(\bin_array[2][2] ));
 sg13g2_dfrbp_1 _1473_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net554),
    .D(_0037_),
    .Q_N(_0769_),
    .Q(\bin_array[2][3] ));
 sg13g2_dfrbp_1 _1474_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net561),
    .D(_0038_),
    .Q_N(_0768_),
    .Q(\bin_array[3][0] ));
 sg13g2_dfrbp_1 _1475_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net561),
    .D(_0039_),
    .Q_N(_0767_),
    .Q(\bin_array[3][1] ));
 sg13g2_dfrbp_1 _1476_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net561),
    .D(_0040_),
    .Q_N(_0766_),
    .Q(\bin_array[3][2] ));
 sg13g2_dfrbp_1 _1477_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net561),
    .D(_0041_),
    .Q_N(_0765_),
    .Q(\bin_array[3][3] ));
 sg13g2_dfrbp_1 _1478_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net561),
    .D(_0042_),
    .Q_N(_0764_),
    .Q(\bin_array[4][0] ));
 sg13g2_dfrbp_1 _1479_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net562),
    .D(_0043_),
    .Q_N(_0763_),
    .Q(\bin_array[4][1] ));
 sg13g2_dfrbp_1 _1480_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net562),
    .D(_0044_),
    .Q_N(_0762_),
    .Q(\bin_array[4][2] ));
 sg13g2_dfrbp_1 _1481_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net562),
    .D(_0045_),
    .Q_N(_0761_),
    .Q(\bin_array[4][3] ));
 sg13g2_dfrbp_1 _1482_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net547),
    .D(_0046_),
    .Q_N(_0760_),
    .Q(\bin_array[5][0] ));
 sg13g2_dfrbp_1 _1483_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net560),
    .D(_0047_),
    .Q_N(_0759_),
    .Q(\bin_array[5][1] ));
 sg13g2_dfrbp_1 _1484_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net551),
    .D(_0048_),
    .Q_N(_0758_),
    .Q(\bin_array[5][2] ));
 sg13g2_dfrbp_1 _1485_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net541),
    .D(_0049_),
    .Q_N(_0757_),
    .Q(\bin_array[5][3] ));
 sg13g2_dfrbp_1 _1486_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net563),
    .D(_0050_),
    .Q_N(_0756_),
    .Q(\bin_array[6][0] ));
 sg13g2_dfrbp_1 _1487_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net563),
    .D(_0051_),
    .Q_N(_0755_),
    .Q(\bin_array[6][1] ));
 sg13g2_dfrbp_1 _1488_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net555),
    .D(_0052_),
    .Q_N(_0754_),
    .Q(\bin_array[6][2] ));
 sg13g2_dfrbp_1 _1489_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net555),
    .D(_0053_),
    .Q_N(_0753_),
    .Q(\bin_array[6][3] ));
 sg13g2_dfrbp_1 _1490_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net555),
    .D(_0054_),
    .Q_N(_0752_),
    .Q(\bin_array[7][0] ));
 sg13g2_dfrbp_1 _1491_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net560),
    .D(_0055_),
    .Q_N(_0751_),
    .Q(\bin_array[7][1] ));
 sg13g2_dfrbp_1 _1492_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net555),
    .D(_0056_),
    .Q_N(_0750_),
    .Q(\bin_array[7][2] ));
 sg13g2_dfrbp_1 _1493_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net555),
    .D(_0057_),
    .Q_N(_0749_),
    .Q(\bin_array[7][3] ));
 sg13g2_dfrbp_1 _1494_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net556),
    .D(_0058_),
    .Q_N(_0748_),
    .Q(\bin_array[8][0] ));
 sg13g2_dfrbp_1 _1495_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net556),
    .D(_0059_),
    .Q_N(_0747_),
    .Q(\bin_array[8][1] ));
 sg13g2_dfrbp_1 _1496_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net556),
    .D(_0060_),
    .Q_N(_0746_),
    .Q(\bin_array[8][2] ));
 sg13g2_dfrbp_1 _1497_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net556),
    .D(_0061_),
    .Q_N(_0745_),
    .Q(\bin_array[8][3] ));
 sg13g2_dfrbp_1 _1498_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net556),
    .D(_0062_),
    .Q_N(_0744_),
    .Q(\bin_array[9][0] ));
 sg13g2_dfrbp_1 _1499_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net554),
    .D(_0063_),
    .Q_N(_0743_),
    .Q(\bin_array[9][1] ));
 sg13g2_dfrbp_1 _1500_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net557),
    .D(_0064_),
    .Q_N(_0742_),
    .Q(\bin_array[9][2] ));
 sg13g2_dfrbp_1 _1501_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net554),
    .D(_0065_),
    .Q_N(_0741_),
    .Q(\bin_array[9][3] ));
 sg13g2_dfrbp_1 _1502_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net560),
    .D(_0066_),
    .Q_N(_0740_),
    .Q(\bin_array[10][0] ));
 sg13g2_dfrbp_1 _1503_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net560),
    .D(_0067_),
    .Q_N(_0739_),
    .Q(\bin_array[10][1] ));
 sg13g2_dfrbp_1 _1504_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net556),
    .D(_0068_),
    .Q_N(_0738_),
    .Q(\bin_array[10][2] ));
 sg13g2_dfrbp_1 _1505_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net560),
    .D(_0069_),
    .Q_N(_0737_),
    .Q(\bin_array[10][3] ));
 sg13g2_dfrbp_1 _1506_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net560),
    .D(_0070_),
    .Q_N(_0736_),
    .Q(\bin_array[11][0] ));
 sg13g2_dfrbp_1 _1507_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net557),
    .D(_0071_),
    .Q_N(_0735_),
    .Q(\bin_array[11][1] ));
 sg13g2_dfrbp_1 _1508_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net555),
    .D(_0072_),
    .Q_N(_0734_),
    .Q(\bin_array[11][2] ));
 sg13g2_dfrbp_1 _1509_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net563),
    .D(_0073_),
    .Q_N(_0733_),
    .Q(\bin_array[11][3] ));
 sg13g2_dfrbp_1 _1510_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net556),
    .D(_0074_),
    .Q_N(_0732_),
    .Q(\bin_array[12][0] ));
 sg13g2_dfrbp_1 _1511_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net560),
    .D(_0075_),
    .Q_N(_0731_),
    .Q(\bin_array[12][1] ));
 sg13g2_dfrbp_1 _1512_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net555),
    .D(_0076_),
    .Q_N(_0730_),
    .Q(\bin_array[12][2] ));
 sg13g2_dfrbp_1 _1513_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net555),
    .D(_0077_),
    .Q_N(_0729_),
    .Q(\bin_array[12][3] ));
 sg13g2_dfrbp_1 _1514_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net561),
    .D(_0078_),
    .Q_N(_0728_),
    .Q(\bin_array[13][0] ));
 sg13g2_dfrbp_1 _1515_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net561),
    .D(_0079_),
    .Q_N(_0727_),
    .Q(\bin_array[13][1] ));
 sg13g2_dfrbp_1 _1516_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net561),
    .D(_0080_),
    .Q_N(_0726_),
    .Q(\bin_array[13][2] ));
 sg13g2_dfrbp_1 _1517_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net560),
    .D(_0081_),
    .Q_N(_0725_),
    .Q(\bin_array[13][3] ));
 sg13g2_dfrbp_1 _1518_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net549),
    .D(_0082_),
    .Q_N(_0724_),
    .Q(\bin_array[14][0] ));
 sg13g2_dfrbp_1 _1519_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net549),
    .D(_0083_),
    .Q_N(_0723_),
    .Q(\bin_array[14][1] ));
 sg13g2_dfrbp_1 _1520_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net549),
    .D(_0084_),
    .Q_N(_0722_),
    .Q(\bin_array[14][2] ));
 sg13g2_dfrbp_1 _1521_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net550),
    .D(_0085_),
    .Q_N(_0721_),
    .Q(\bin_array[14][3] ));
 sg13g2_dfrbp_1 _1522_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net551),
    .D(_0086_),
    .Q_N(_0720_),
    .Q(\bin_array[15][0] ));
 sg13g2_dfrbp_1 _1523_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net549),
    .D(_0087_),
    .Q_N(_0719_),
    .Q(\bin_array[15][1] ));
 sg13g2_dfrbp_1 _1524_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net549),
    .D(_0088_),
    .Q_N(_0718_),
    .Q(\bin_array[15][2] ));
 sg13g2_dfrbp_1 _1525_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net551),
    .D(_0089_),
    .Q_N(_0717_),
    .Q(\bin_array[15][3] ));
 sg13g2_dfrbp_1 _1526_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net543),
    .D(_0090_),
    .Q_N(_0716_),
    .Q(\bin_array[16][0] ));
 sg13g2_dfrbp_1 _1527_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net543),
    .D(_0091_),
    .Q_N(_0715_),
    .Q(\bin_array[16][1] ));
 sg13g2_dfrbp_1 _1528_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net542),
    .D(_0092_),
    .Q_N(_0714_),
    .Q(\bin_array[16][2] ));
 sg13g2_dfrbp_1 _1529_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net542),
    .D(_0093_),
    .Q_N(_0713_),
    .Q(\bin_array[16][3] ));
 sg13g2_dfrbp_1 _1530_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net543),
    .D(_0094_),
    .Q_N(_0712_),
    .Q(\bin_array[17][0] ));
 sg13g2_dfrbp_1 _1531_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net544),
    .D(_0095_),
    .Q_N(_0711_),
    .Q(\bin_array[17][1] ));
 sg13g2_dfrbp_1 _1532_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net543),
    .D(_0096_),
    .Q_N(_0710_),
    .Q(\bin_array[17][2] ));
 sg13g2_dfrbp_1 _1533_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net544),
    .D(_0097_),
    .Q_N(_0709_),
    .Q(\bin_array[17][3] ));
 sg13g2_dfrbp_1 _1534_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net540),
    .D(_0098_),
    .Q_N(_0708_),
    .Q(\bin_array[18][0] ));
 sg13g2_dfrbp_1 _1535_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net540),
    .D(_0099_),
    .Q_N(_0707_),
    .Q(\bin_array[18][1] ));
 sg13g2_dfrbp_1 _1536_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net541),
    .D(_0100_),
    .Q_N(_0706_),
    .Q(\bin_array[18][2] ));
 sg13g2_dfrbp_1 _1537_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net541),
    .D(_0101_),
    .Q_N(_0705_),
    .Q(\bin_array[18][3] ));
 sg13g2_dfrbp_1 _1538_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net543),
    .D(_0102_),
    .Q_N(_0704_),
    .Q(\bin_array[19][0] ));
 sg13g2_dfrbp_1 _1539_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net552),
    .D(_0103_),
    .Q_N(_0703_),
    .Q(\bin_array[19][1] ));
 sg13g2_dfrbp_1 _1540_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net543),
    .D(_0104_),
    .Q_N(_0702_),
    .Q(\bin_array[19][2] ));
 sg13g2_dfrbp_1 _1541_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net552),
    .D(_0105_),
    .Q_N(_0701_),
    .Q(\bin_array[19][3] ));
 sg13g2_dfrbp_1 _1542_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net540),
    .D(_0106_),
    .Q_N(_0700_),
    .Q(\bin_array[20][0] ));
 sg13g2_dfrbp_1 _1543_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net540),
    .D(_0107_),
    .Q_N(_0699_),
    .Q(\bin_array[20][1] ));
 sg13g2_dfrbp_1 _1544_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net540),
    .D(_0108_),
    .Q_N(_0698_),
    .Q(\bin_array[20][2] ));
 sg13g2_dfrbp_1 _1545_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net541),
    .D(_0109_),
    .Q_N(_0697_),
    .Q(\bin_array[20][3] ));
 sg13g2_dfrbp_1 _1546_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net540),
    .D(_0110_),
    .Q_N(_0696_),
    .Q(\bin_array[21][0] ));
 sg13g2_dfrbp_1 _1547_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net540),
    .D(_0111_),
    .Q_N(_0695_),
    .Q(\bin_array[21][1] ));
 sg13g2_dfrbp_1 _1548_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net546),
    .D(_0112_),
    .Q_N(_0694_),
    .Q(\bin_array[21][2] ));
 sg13g2_dfrbp_1 _1549_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net541),
    .D(_0113_),
    .Q_N(_0693_),
    .Q(\bin_array[21][3] ));
 sg13g2_dfrbp_1 _1550_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net542),
    .D(_0114_),
    .Q_N(_0692_),
    .Q(\bin_array[22][0] ));
 sg13g2_dfrbp_1 _1551_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net540),
    .D(_0115_),
    .Q_N(_0691_),
    .Q(\bin_array[22][1] ));
 sg13g2_dfrbp_1 _1552_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net542),
    .D(_0116_),
    .Q_N(_0690_),
    .Q(\bin_array[22][2] ));
 sg13g2_dfrbp_1 _1553_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net542),
    .D(_0117_),
    .Q_N(_0689_),
    .Q(\bin_array[22][3] ));
 sg13g2_dfrbp_1 _1554_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net546),
    .D(net119),
    .Q_N(_0688_),
    .Q(\bin_array[23][0] ));
 sg13g2_dfrbp_1 _1555_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net546),
    .D(_0119_),
    .Q_N(_0687_),
    .Q(\bin_array[23][1] ));
 sg13g2_dfrbp_1 _1556_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net546),
    .D(_0120_),
    .Q_N(_0686_),
    .Q(\bin_array[23][2] ));
 sg13g2_dfrbp_1 _1557_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net547),
    .D(_0121_),
    .Q_N(_0685_),
    .Q(\bin_array[23][3] ));
 sg13g2_dfrbp_1 _1558_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net546),
    .D(net104),
    .Q_N(_0684_),
    .Q(\bin_array[24][0] ));
 sg13g2_dfrbp_1 _1559_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net546),
    .D(_0123_),
    .Q_N(_0683_),
    .Q(\bin_array[24][1] ));
 sg13g2_dfrbp_1 _1560_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net546),
    .D(_0124_),
    .Q_N(_0682_),
    .Q(\bin_array[24][2] ));
 sg13g2_dfrbp_1 _1561_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net547),
    .D(_0125_),
    .Q_N(_0681_),
    .Q(\bin_array[24][3] ));
 sg13g2_dfrbp_1 _1562_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net544),
    .D(_0126_),
    .Q_N(_0680_),
    .Q(\bin_array[25][0] ));
 sg13g2_dfrbp_1 _1563_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net544),
    .D(_0127_),
    .Q_N(_0679_),
    .Q(\bin_array[25][1] ));
 sg13g2_dfrbp_1 _1564_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net552),
    .D(_0128_),
    .Q_N(_0678_),
    .Q(\bin_array[25][2] ));
 sg13g2_dfrbp_1 _1565_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net552),
    .D(_0129_),
    .Q_N(_0677_),
    .Q(\bin_array[25][3] ));
 sg13g2_dfrbp_1 _1566_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net542),
    .D(_0130_),
    .Q_N(_0676_),
    .Q(\bin_array[26][0] ));
 sg13g2_dfrbp_1 _1567_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net543),
    .D(_0131_),
    .Q_N(_0675_),
    .Q(\bin_array[26][1] ));
 sg13g2_dfrbp_1 _1568_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net542),
    .D(_0132_),
    .Q_N(_0674_),
    .Q(\bin_array[26][2] ));
 sg13g2_dfrbp_1 _1569_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net543),
    .D(_0133_),
    .Q_N(_0673_),
    .Q(\bin_array[26][3] ));
 sg13g2_dfrbp_1 _1570_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net552),
    .D(_0134_),
    .Q_N(_0672_),
    .Q(\bin_array[27][0] ));
 sg13g2_dfrbp_1 _1571_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net553),
    .D(_0135_),
    .Q_N(_0671_),
    .Q(\bin_array[27][1] ));
 sg13g2_dfrbp_1 _1572_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net553),
    .D(_0136_),
    .Q_N(_0670_),
    .Q(\bin_array[27][2] ));
 sg13g2_dfrbp_1 _1573_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net553),
    .D(_0137_),
    .Q_N(_0669_),
    .Q(\bin_array[27][3] ));
 sg13g2_dfrbp_1 _1574_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net554),
    .D(_0138_),
    .Q_N(_0668_),
    .Q(\bin_array[28][0] ));
 sg13g2_dfrbp_1 _1575_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net553),
    .D(_0139_),
    .Q_N(_0667_),
    .Q(\bin_array[28][1] ));
 sg13g2_dfrbp_1 _1576_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net553),
    .D(_0140_),
    .Q_N(_0666_),
    .Q(\bin_array[28][2] ));
 sg13g2_dfrbp_1 _1577_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net554),
    .D(_0141_),
    .Q_N(_0665_),
    .Q(\bin_array[28][3] ));
 sg13g2_dfrbp_1 _1578_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net552),
    .D(_0142_),
    .Q_N(_0664_),
    .Q(\bin_array[29][0] ));
 sg13g2_dfrbp_1 _1579_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net552),
    .D(_0143_),
    .Q_N(_0663_),
    .Q(\bin_array[29][1] ));
 sg13g2_dfrbp_1 _1580_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net553),
    .D(_0144_),
    .Q_N(_0662_),
    .Q(\bin_array[29][2] ));
 sg13g2_dfrbp_1 _1581_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net552),
    .D(_0145_),
    .Q_N(_0661_),
    .Q(\bin_array[29][3] ));
 sg13g2_dfrbp_1 _1582_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net547),
    .D(_0146_),
    .Q_N(_0660_),
    .Q(\bin_array[30][0] ));
 sg13g2_dfrbp_1 _1583_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net546),
    .D(_0147_),
    .Q_N(_0659_),
    .Q(\bin_array[30][1] ));
 sg13g2_dfrbp_1 _1584_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net547),
    .D(_0148_),
    .Q_N(_0658_),
    .Q(\bin_array[30][2] ));
 sg13g2_dfrbp_1 _1585_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net547),
    .D(_0149_),
    .Q_N(_0657_),
    .Q(\bin_array[30][3] ));
 sg13g2_tiehi tt_um_histogramming_18 (.L_HI(net18));
 sg13g2_tiehi tt_um_histogramming_19 (.L_HI(net19));
 sg13g2_tiehi tt_um_histogramming_20 (.L_HI(net20));
 sg13g2_tiehi tt_um_histogramming_21 (.L_HI(net21));
 sg13g2_tiehi tt_um_histogramming_22 (.L_HI(net22));
 sg13g2_tiehi tt_um_histogramming_23 (.L_HI(net23));
 sg13g2_tiehi tt_um_histogramming_24 (.L_HI(net24));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_histogramming_9 (.L_LO(net9));
 sg13g2_tielo tt_um_histogramming_10 (.L_LO(net10));
 sg13g2_tielo tt_um_histogramming_11 (.L_LO(net11));
 sg13g2_tielo tt_um_histogramming_12 (.L_LO(net12));
 sg13g2_tielo tt_um_histogramming_13 (.L_LO(net13));
 sg13g2_tielo tt_um_histogramming_14 (.L_LO(net14));
 sg13g2_tielo tt_um_histogramming_15 (.L_LO(net15));
 sg13g2_tielo tt_um_histogramming_16 (.L_LO(net16));
 sg13g2_tiehi tt_um_histogramming_17 (.L_HI(net17));
 sg13g2_buf_1 _1603_ (.A(ready_reg),
    .X(uio_out[2]));
 sg13g2_buf_1 _1604_ (.A(last_bin_reg),
    .X(uio_out[3]));
 sg13g2_buf_1 _1605_ (.A(valid_out_reg),
    .X(uio_out[4]));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(net425));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(net429));
 sg13g2_buf_1 fanout426 (.A(net429),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(net429),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(net429),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_0546_),
    .X(net429));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(net434));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(net434));
 sg13g2_buf_4 fanout432 (.X(net432),
    .A(net433));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(net434));
 sg13g2_buf_2 fanout434 (.A(_0544_),
    .X(net434));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(net439));
 sg13g2_buf_2 fanout436 (.A(net439),
    .X(net436));
 sg13g2_buf_4 fanout437 (.X(net437),
    .A(net439));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(net439));
 sg13g2_buf_2 fanout439 (.A(_0541_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(net441),
    .X(net440));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(net444));
 sg13g2_buf_4 fanout442 (.X(net442),
    .A(net444));
 sg13g2_buf_2 fanout443 (.A(net444),
    .X(net443));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(_0538_));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(net447));
 sg13g2_buf_2 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_4 fanout447 (.X(net447),
    .A(_0534_));
 sg13g2_buf_2 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_0533_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(net453),
    .X(net452));
 sg13g2_buf_4 fanout453 (.X(net453),
    .A(_0380_));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(net455));
 sg13g2_buf_8 fanout455 (.A(_0379_),
    .X(net455));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(_0396_));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(net458));
 sg13g2_buf_2 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_0006_),
    .X(net459));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(net461));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(net462));
 sg13g2_buf_2 fanout462 (.A(net181),
    .X(net462));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(\shift_count[3] ));
 sg13g2_buf_2 fanout464 (.A(net182),
    .X(net464));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(net183));
 sg13g2_buf_1 fanout466 (.A(\shift_count[2] ),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_0213_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(net469),
    .X(net468));
 sg13g2_buf_1 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_0183_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_0183_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(net475),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net475),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net477),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(net477),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_0174_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(net480),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_0170_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_0170_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_0170_),
    .X(net482));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(_0168_));
 sg13g2_buf_1 fanout484 (.A(_0168_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_0168_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net492),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(net491),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(net492),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_0164_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(net495),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_0160_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_0160_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(net501),
    .X(net499));
 sg13g2_buf_1 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_0157_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(net503),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_0157_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(net509),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net509),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_1 fanout507 (.A(net509),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_0156_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(net513),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net513),
    .X(net511));
 sg13g2_buf_1 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_1 fanout513 (.A(_0150_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_1 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(net520),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(net519),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_1 fanout520 (.A(_0150_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net523),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net530),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(net526),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net530),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_1 fanout530 (.A(ui_in[5]),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(net535),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_1 fanout535 (.A(ui_in[5]),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net6),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(net5),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(net4),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net3),
    .X(net539));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net541));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(net542));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(net545));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(net545));
 sg13g2_buf_2 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net565),
    .X(net545));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(net547));
 sg13g2_buf_4 fanout547 (.X(net547),
    .A(net548));
 sg13g2_buf_2 fanout548 (.A(net565),
    .X(net548));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(net551));
 sg13g2_buf_2 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net565),
    .X(net551));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(net564));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(net564));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(net557));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(net556));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(net557));
 sg13g2_buf_2 fanout557 (.A(net564),
    .X(net557));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(net564));
 sg13g2_buf_2 fanout559 (.A(net564),
    .X(net559));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(net563));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(net562));
 sg13g2_buf_2 fanout562 (.A(net563),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(net565));
 sg13g2_buf_2 fanout565 (.A(rst_n),
    .X(net565));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_tielo tt_um_histogramming_8 (.L_LO(net8));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\bin_array[0][2] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0028_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0008_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0025_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold5 (.A(\state[1] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0000_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold7 (.A(\state[0] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0009_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold9 (.A(\bin_array[1][0] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold10 (.A(last_bin_reg),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0561_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0024_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold13 (.A(\bin_array[0][3] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold14 (.A(\bin_array[15][2] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold15 (.A(\bin_array[15][0] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold16 (.A(\bin_array[5][2] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold17 (.A(\bin_array[14][2] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold18 (.A(uo_out[0]),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0392_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0010_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold21 (.A(\bin_array[0][1] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold22 (.A(\bin_array[5][0] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold23 (.A(\bin_array[7][2] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold24 (.A(\bin_array[30][0] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold25 (.A(\bin_array[6][2] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold26 (.A(\bin_array[0][0] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold27 (.A(\bin_array[10][2] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold28 (.A(\bin_array[12][2] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold29 (.A(\bin_array[2][2] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold30 (.A(\bin_array[8][2] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold31 (.A(\bin_array[12][0] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold32 (.A(\bin_array[27][2] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold33 (.A(\bin_array[27][3] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold34 (.A(\bin_array[9][0] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold35 (.A(\bin_array[31][3] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold36 (.A(uo_out[2]),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0012_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold38 (.A(\bin_array[26][1] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold39 (.A(\bin_array[25][2] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold40 (.A(\bin_array[31][0] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0014_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold42 (.A(\bin_array[8][0] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold43 (.A(\bin_array[26][3] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold44 (.A(\bin_array[1][2] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold45 (.A(\bin_array[29][3] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold46 (.A(\bin_array[30][3] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold47 (.A(\bin_array[27][1] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold48 (.A(\bin_array[30][2] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold49 (.A(\bin_array[17][2] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold50 (.A(\bin_array[17][0] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold51 (.A(\bin_array[31][2] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold52 (.A(\bin_array[9][2] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold53 (.A(\bin_array[20][2] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold54 (.A(\bin_array[19][0] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold55 (.A(\bin_array[7][0] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold56 (.A(\bin_array[2][0] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold57 (.A(\bin_array[19][3] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold58 (.A(\bin_array[15][3] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold59 (.A(\bin_array[28][1] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold60 (.A(\bin_array[17][1] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold61 (.A(\bin_array[31][1] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold62 (.A(uo_out[3]),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0013_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold64 (.A(\bin_array[23][3] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold65 (.A(valid_out_reg),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold66 (.A(\bin_array[11][0] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold67 (.A(\bin_array[23][2] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold68 (.A(\bin_array[18][2] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold69 (.A(uo_out[1]),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0011_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold71 (.A(\bin_array[24][3] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold72 (.A(\bin_array[24][2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold73 (.A(\bin_array[29][0] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold74 (.A(\bin_array[14][0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold75 (.A(\bin_array[16][3] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold76 (.A(\bin_array[26][0] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold77 (.A(\bin_array[22][3] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold78 (.A(\bin_array[16][1] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold79 (.A(\bin_array[24][0] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0122_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold81 (.A(\bin_array[18][0] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold82 (.A(\bin_array[17][3] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold83 (.A(\bin_array[1][3] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold84 (.A(\bin_array[27][0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold85 (.A(\bin_array[21][0] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold86 (.A(\bin_array[6][0] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold87 (.A(\bin_array[26][2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold88 (.A(\bin_array[18][1] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold89 (.A(\bin_array[20][0] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold90 (.A(\bin_array[9][3] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold91 (.A(\bin_array[10][0] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold92 (.A(\bin_array[4][0] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold93 (.A(\bin_array[13][2] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold94 (.A(\bin_array[23][0] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0118_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold96 (.A(\bin_array[14][3] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold97 (.A(\bin_array[23][1] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold98 (.A(\bin_array[20][3] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold99 (.A(\bin_array[30][1] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold100 (.A(\bin_array[29][2] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold101 (.A(\bin_array[13][0] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold102 (.A(\bin_array[9][1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold103 (.A(\bin_array[22][0] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold104 (.A(\bin_array[21][2] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold105 (.A(\bin_array[5][1] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold106 (.A(\bin_array[16][0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold107 (.A(\bin_array[15][1] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold108 (.A(\bin_array[11][2] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold109 (.A(\bin_array[25][0] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold110 (.A(\bin_array[1][1] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold111 (.A(\bin_array[28][3] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold112 (.A(\bin_array[3][2] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold113 (.A(\bin_array[28][2] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold114 (.A(\bin_array[14][1] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold115 (.A(\bin_array[8][1] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold116 (.A(\bin_array[28][0] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold117 (.A(\bin_array[10][1] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold118 (.A(\bin_array[4][2] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold119 (.A(\bin_array[18][3] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold120 (.A(\bin_array[16][2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold121 (.A(\bin_array[19][1] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold122 (.A(\bin_array[24][1] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold123 (.A(\bin_array[25][3] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold124 (.A(\bin_array[20][1] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold125 (.A(\bin_array[21][3] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold126 (.A(\bin_array[22][1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold127 (.A(\bin_array[12][3] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold128 (.A(\bin_array[6][3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold129 (.A(\bin_array[11][3] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold130 (.A(\bin_array[22][2] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold131 (.A(\bin_array[7][3] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold132 (.A(\bin_array[3][1] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold133 (.A(\bin_array[25][1] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold134 (.A(\bin_array[21][1] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold135 (.A(\bin_array[19][2] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold136 (.A(\bin_array[10][3] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold137 (.A(\bin_array[13][3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold138 (.A(\bin_array[5][3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold139 (.A(\bin_array[2][3] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold140 (.A(\bin_array[12][1] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold141 (.A(\bin_array[29][1] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold142 (.A(\bin_array[4][3] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold143 (.A(\bin_array[6][1] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold144 (.A(\bin_array[3][0] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold145 (.A(\bin_array[4][1] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold146 (.A(\bin_array[8][3] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold147 (.A(\bin_array[13][1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold148 (.A(\bin_array[2][1] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold149 (.A(\bin_array[7][1] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold150 (.A(\bin_array[11][1] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold151 (.A(\shift_count[1] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0019_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold153 (.A(\state[2] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0001_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold155 (.A(\shift_count[0] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold156 (.A(\bin_array[3][3] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold157 (.A(\shift_count[4] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold158 (.A(\shift_count[3] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold159 (.A(\shift_count[2] ),
    .X(net183));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_4 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_199 ();
 sg13g2_decap_8 FILLER_6_206 ();
 sg13g2_decap_8 FILLER_6_213 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_decap_8 FILLER_6_227 ();
 sg13g2_decap_8 FILLER_6_234 ();
 sg13g2_decap_8 FILLER_6_241 ();
 sg13g2_decap_8 FILLER_6_248 ();
 sg13g2_decap_8 FILLER_6_255 ();
 sg13g2_decap_8 FILLER_6_262 ();
 sg13g2_decap_8 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_276 ();
 sg13g2_decap_8 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_290 ();
 sg13g2_decap_8 FILLER_6_297 ();
 sg13g2_decap_8 FILLER_6_304 ();
 sg13g2_decap_8 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_4 FILLER_7_141 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_229 ();
 sg13g2_decap_4 FILLER_7_236 ();
 sg13g2_fill_2 FILLER_7_240 ();
 sg13g2_fill_2 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_275 ();
 sg13g2_decap_8 FILLER_7_282 ();
 sg13g2_decap_4 FILLER_7_289 ();
 sg13g2_fill_2 FILLER_7_293 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_fill_2 FILLER_8_105 ();
 sg13g2_decap_4 FILLER_8_120 ();
 sg13g2_fill_2 FILLER_8_124 ();
 sg13g2_fill_2 FILLER_8_312 ();
 sg13g2_fill_1 FILLER_8_314 ();
 sg13g2_decap_4 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_327 ();
 sg13g2_fill_1 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_4 FILLER_9_91 ();
 sg13g2_fill_2 FILLER_9_95 ();
 sg13g2_fill_1 FILLER_9_132 ();
 sg13g2_fill_1 FILLER_9_190 ();
 sg13g2_decap_8 FILLER_9_219 ();
 sg13g2_decap_4 FILLER_9_226 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_236 ();
 sg13g2_fill_1 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_348 ();
 sg13g2_decap_4 FILLER_9_355 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_fill_1 FILLER_10_63 ();
 sg13g2_fill_2 FILLER_10_69 ();
 sg13g2_fill_1 FILLER_10_80 ();
 sg13g2_fill_1 FILLER_10_89 ();
 sg13g2_fill_2 FILLER_10_112 ();
 sg13g2_fill_2 FILLER_10_127 ();
 sg13g2_fill_2 FILLER_10_164 ();
 sg13g2_fill_2 FILLER_10_292 ();
 sg13g2_fill_1 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_324 ();
 sg13g2_fill_1 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_25 ();
 sg13g2_decap_4 FILLER_11_53 ();
 sg13g2_fill_2 FILLER_11_101 ();
 sg13g2_fill_1 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_2 FILLER_11_209 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_fill_1 FILLER_11_235 ();
 sg13g2_fill_2 FILLER_11_343 ();
 sg13g2_decap_4 FILLER_11_349 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_105 ();
 sg13g2_fill_2 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_158 ();
 sg13g2_fill_2 FILLER_12_195 ();
 sg13g2_fill_2 FILLER_12_254 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_decap_4 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_decap_4 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_decap_4 FILLER_13_233 ();
 sg13g2_fill_1 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_fill_2 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_18 ();
 sg13g2_fill_1 FILLER_14_50 ();
 sg13g2_decap_8 FILLER_14_61 ();
 sg13g2_fill_2 FILLER_14_94 ();
 sg13g2_fill_2 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_2 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_197 ();
 sg13g2_fill_2 FILLER_14_204 ();
 sg13g2_fill_1 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_fill_2 FILLER_14_232 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_265 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_fill_1 FILLER_14_310 ();
 sg13g2_fill_2 FILLER_14_324 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_2 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_fill_2 FILLER_15_115 ();
 sg13g2_fill_1 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_170 ();
 sg13g2_fill_2 FILLER_15_177 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_decap_4 FILLER_15_228 ();
 sg13g2_fill_1 FILLER_15_232 ();
 sg13g2_fill_1 FILLER_15_239 ();
 sg13g2_decap_4 FILLER_15_269 ();
 sg13g2_fill_2 FILLER_15_273 ();
 sg13g2_decap_4 FILLER_15_299 ();
 sg13g2_fill_2 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_340 ();
 sg13g2_fill_1 FILLER_15_367 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_144 ();
 sg13g2_decap_4 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_185 ();
 sg13g2_fill_1 FILLER_16_187 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_fill_1 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_decap_4 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_233 ();
 sg13g2_fill_1 FILLER_17_235 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_fill_2 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_305 ();
 sg13g2_fill_2 FILLER_17_369 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_111 ();
 sg13g2_decap_8 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_decap_4 FILLER_18_141 ();
 sg13g2_fill_1 FILLER_18_145 ();
 sg13g2_decap_4 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_211 ();
 sg13g2_decap_4 FILLER_18_218 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_fill_2 FILLER_18_239 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_decap_4 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_372 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_decap_4 FILLER_19_116 ();
 sg13g2_decap_4 FILLER_19_148 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_decap_8 FILLER_19_171 ();
 sg13g2_fill_2 FILLER_19_178 ();
 sg13g2_fill_1 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_decap_4 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_298 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_47 ();
 sg13g2_fill_1 FILLER_20_68 ();
 sg13g2_fill_2 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_139 ();
 sg13g2_decap_4 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_171 ();
 sg13g2_decap_4 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_259 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_decap_4 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_314 ();
 sg13g2_fill_1 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_110 ();
 sg13g2_decap_4 FILLER_21_121 ();
 sg13g2_decap_8 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_167 ();
 sg13g2_decap_4 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_184 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_decap_4 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_38 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_fill_1 FILLER_22_115 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_decap_8 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_155 ();
 sg13g2_fill_2 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_199 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_219 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_277 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_29 ();
 sg13g2_fill_1 FILLER_23_31 ();
 sg13g2_fill_2 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_124 ();
 sg13g2_fill_1 FILLER_23_131 ();
 sg13g2_decap_8 FILLER_23_155 ();
 sg13g2_decap_4 FILLER_23_173 ();
 sg13g2_decap_4 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_decap_4 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_215 ();
 sg13g2_decap_4 FILLER_23_224 ();
 sg13g2_decap_4 FILLER_23_252 ();
 sg13g2_decap_4 FILLER_23_279 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_2 FILLER_23_300 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_fill_1 FILLER_24_54 ();
 sg13g2_fill_2 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_76 ();
 sg13g2_fill_2 FILLER_24_109 ();
 sg13g2_decap_4 FILLER_24_131 ();
 sg13g2_fill_2 FILLER_24_146 ();
 sg13g2_fill_1 FILLER_24_148 ();
 sg13g2_decap_4 FILLER_24_169 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_fill_1 FILLER_24_229 ();
 sg13g2_fill_2 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_fill_1 FILLER_24_252 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_356 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_113 ();
 sg13g2_fill_2 FILLER_25_131 ();
 sg13g2_decap_4 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_decap_4 FILLER_25_176 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_4 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_decap_4 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_168 ();
 sg13g2_decap_4 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_decap_4 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_1 FILLER_26_261 ();
 sg13g2_fill_1 FILLER_26_274 ();
 sg13g2_fill_2 FILLER_26_280 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_346 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_fill_1 FILLER_27_69 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_decap_4 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_160 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_fill_2 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_100 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_decap_4 FILLER_28_184 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_4 FILLER_28_224 ();
 sg13g2_decap_4 FILLER_28_240 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_52 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_2 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_180 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_fill_1 FILLER_29_192 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_25 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_69 ();
 sg13g2_fill_2 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_fill_1 FILLER_30_153 ();
 sg13g2_fill_2 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_fill_1 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_fill_1 FILLER_31_50 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_decap_4 FILLER_31_152 ();
 sg13g2_decap_4 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_1 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_85 ();
 sg13g2_decap_4 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_283 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_381 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_fill_1 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_2 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_60 ();
 sg13g2_decap_8 FILLER_34_82 ();
 sg13g2_decap_4 FILLER_34_89 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_2 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_fill_2 FILLER_34_331 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_105 ();
 sg13g2_fill_1 FILLER_35_107 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_151 ();
 sg13g2_fill_2 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_190 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_381 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_162 ();
 sg13g2_fill_1 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_fill_2 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_362 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[5] = net10;
 assign uio_out[6] = net11;
 assign uio_out[7] = net12;
 assign uo_out[4] = net13;
 assign uo_out[5] = net14;
 assign uo_out[6] = net15;
 assign uo_out[7] = net16;
endmodule

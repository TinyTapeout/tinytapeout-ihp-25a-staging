module tt_um_MichaelBell_mandelbrot (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire clk_regs;
 wire \i_coord.demo_update ;
 wire \i_coord.demo_update_delay ;
 wire \i_coord.l_xip.gated_clk ;
 wire \i_coord.l_xip.genblk2[0].state.D ;
 wire \i_coord.l_xip.genblk2[0].state.Q ;
 wire \i_coord.l_xip.genblk2[1].state.D ;
 wire \i_coord.l_xip.genblk2[1].state.Q ;
 wire \i_coord.l_xip.genblk2[2].state.D ;
 wire \i_coord.l_xip.genblk2[2].state.Q ;
 wire \i_coord.l_xip.genblk2[3].state.D ;
 wire \i_coord.l_xip.genblk2[3].state.Q ;
 wire \i_coord.l_xip.genblk2[4].state.D ;
 wire \i_coord.l_xip.genblk2[4].state.Q ;
 wire \i_coord.l_xip.genblk2[5].state.D ;
 wire \i_coord.l_xip.genblk2[5].state.Q ;
 wire \i_coord.l_xip.genblk2[6].state.D ;
 wire \i_coord.l_xip.genblk2[6].state.Q ;
 wire \i_coord.l_xip.genblk2[7].state.D ;
 wire \i_coord.l_xip.genblk2[7].state.Q ;
 wire \i_coord.l_xip.genblk2[8].state.D ;
 wire \i_coord.l_xip.genblk2[8].state.Q ;
 wire \i_coord.l_xip.genblk2[9].state.D ;
 wire \i_coord.l_xip.genblk2[9].state.Q ;
 wire \i_coord.l_xir.gated_clk ;
 wire \i_coord.l_xir.genblk2[0].state.D ;
 wire \i_coord.l_xir.genblk2[0].state.Q ;
 wire \i_coord.l_xir.genblk2[1].state.D ;
 wire \i_coord.l_xir.genblk2[1].state.Q ;
 wire \i_coord.l_xir.genblk2[2].state.D ;
 wire \i_coord.l_xir.genblk2[2].state.Q ;
 wire \i_coord.l_xir.genblk2[3].state.D ;
 wire \i_coord.l_xir.genblk2[3].state.Q ;
 wire \i_coord.l_xir.genblk2[4].state.D ;
 wire \i_coord.l_xir.genblk2[4].state.Q ;
 wire \i_coord.l_xir.genblk2[5].state.D ;
 wire \i_coord.l_xir.genblk2[5].state.Q ;
 wire \i_coord.l_xir.genblk2[6].state.D ;
 wire \i_coord.l_xir.genblk2[6].state.Q ;
 wire \i_coord.l_xir.genblk2[7].state.D ;
 wire \i_coord.l_xir.genblk2[7].state.Q ;
 wire \i_coord.l_xl.gated_clk ;
 wire \i_coord.l_xl.genblk2[10].state.Q ;
 wire \i_coord.l_xl.genblk2[11].state.D ;
 wire \i_coord.l_xl.genblk2[11].state.Q ;
 wire \i_coord.l_xl.genblk2[12].state.D ;
 wire \i_coord.l_xl.genblk2[12].state.Q ;
 wire \i_coord.l_xl.genblk2[13].state.D ;
 wire \i_coord.l_xl.genblk2[13].state.Q ;
 wire \i_coord.l_xl.genblk2[14].state.D ;
 wire \i_coord.l_xl.genblk2[14].state.Q ;
 wire \i_coord.l_xl.genblk2[15].state.D ;
 wire \i_coord.l_xl.genblk2[15].state.Q ;
 wire \i_coord.l_xl.genblk2[3].state.Q ;
 wire \i_coord.l_xl.genblk2[4].state.Q ;
 wire \i_coord.l_xl.genblk2[5].state.Q ;
 wire \i_coord.l_xl.genblk2[6].state.Q ;
 wire \i_coord.l_xl.genblk2[7].state.Q ;
 wire \i_coord.l_xl.genblk2[8].state.Q ;
 wire \i_coord.l_xl.genblk2[9].state.Q ;
 wire \i_coord.l_yip.gated_clk ;
 wire \i_coord.l_yip.genblk2[0].state.Q ;
 wire \i_coord.l_yip.genblk2[1].state.Q ;
 wire \i_coord.l_yip.genblk2[2].state.Q ;
 wire \i_coord.l_yip.genblk2[3].state.Q ;
 wire \i_coord.l_yip.genblk2[4].state.Q ;
 wire \i_coord.l_yip.genblk2[5].state.Q ;
 wire \i_coord.l_yip.genblk2[6].state.Q ;
 wire \i_coord.l_yip.genblk2[7].state.Q ;
 wire \i_coord.l_yip.genblk2[8].state.Q ;
 wire \i_coord.l_yip.genblk2[9].state.Q ;
 wire \i_coord.l_yt.gated_clk ;
 wire \i_coord.l_yt.genblk2[0].state.D ;
 wire \i_coord.l_yt.genblk2[0].state.Q ;
 wire \i_coord.l_yt.genblk2[10].state.D ;
 wire \i_coord.l_yt.genblk2[10].state.Q ;
 wire \i_coord.l_yt.genblk2[11].state.D ;
 wire \i_coord.l_yt.genblk2[11].state.Q ;
 wire \i_coord.l_yt.genblk2[12].state.D ;
 wire \i_coord.l_yt.genblk2[12].state.Q ;
 wire \i_coord.l_yt.genblk2[13].state.D ;
 wire \i_coord.l_yt.genblk2[13].state.Q ;
 wire \i_coord.l_yt.genblk2[14].state.D ;
 wire \i_coord.l_yt.genblk2[14].state.Q ;
 wire \i_coord.l_yt.genblk2[1].state.D ;
 wire \i_coord.l_yt.genblk2[1].state.Q ;
 wire \i_coord.l_yt.genblk2[2].state.D ;
 wire \i_coord.l_yt.genblk2[2].state.Q ;
 wire \i_coord.l_yt.genblk2[3].state.D ;
 wire \i_coord.l_yt.genblk2[3].state.Q ;
 wire \i_coord.l_yt.genblk2[4].state.D ;
 wire \i_coord.l_yt.genblk2[4].state.Q ;
 wire \i_coord.l_yt.genblk2[5].state.D ;
 wire \i_coord.l_yt.genblk2[5].state.Q ;
 wire \i_coord.l_yt.genblk2[6].state.D ;
 wire \i_coord.l_yt.genblk2[6].state.Q ;
 wire \i_coord.l_yt.genblk2[7].state.D ;
 wire \i_coord.l_yt.genblk2[7].state.Q ;
 wire \i_coord.l_yt.genblk2[8].state.D ;
 wire \i_coord.l_yt.genblk2[8].state.Q ;
 wire \i_coord.l_yt.genblk2[9].state.D ;
 wire \i_coord.l_yt.genblk2[9].state.Q ;
 wire \i_coord.x0[-10] ;
 wire \i_coord.x0[-11] ;
 wire \i_coord.x0[-12] ;
 wire \i_coord.x0[-13] ;
 wire \i_coord.x0[-1] ;
 wire \i_coord.x0[-2] ;
 wire \i_coord.x0[-3] ;
 wire \i_coord.x0[-4] ;
 wire \i_coord.x0[-5] ;
 wire \i_coord.x0[-6] ;
 wire \i_coord.x0[-7] ;
 wire \i_coord.x0[-8] ;
 wire \i_coord.x0[-9] ;
 wire \i_coord.x0[0] ;
 wire \i_coord.x0[1] ;
 wire \i_coord.x0[2] ;
 wire \i_coord.x_row_start[-10] ;
 wire \i_coord.x_row_start[-11] ;
 wire \i_coord.x_row_start[-12] ;
 wire \i_coord.x_row_start[-13] ;
 wire \i_coord.x_row_start[-1] ;
 wire \i_coord.x_row_start[-2] ;
 wire \i_coord.x_row_start[-3] ;
 wire \i_coord.x_row_start[-4] ;
 wire \i_coord.x_row_start[-5] ;
 wire \i_coord.x_row_start[-6] ;
 wire \i_coord.x_row_start[-7] ;
 wire \i_coord.x_row_start[-8] ;
 wire \i_coord.x_row_start[-9] ;
 wire \i_coord.x_row_start[0] ;
 wire \i_coord.x_row_start[1] ;
 wire \i_coord.x_row_start[2] ;
 wire \i_coord.y0[-10] ;
 wire \i_coord.y0[-11] ;
 wire \i_coord.y0[-12] ;
 wire \i_coord.y0[-13] ;
 wire \i_coord.y0[-1] ;
 wire \i_coord.y0[-2] ;
 wire \i_coord.y0[-3] ;
 wire \i_coord.y0[-4] ;
 wire \i_coord.y0[-5] ;
 wire \i_coord.y0[-6] ;
 wire \i_coord.y0[-7] ;
 wire \i_coord.y0[-8] ;
 wire \i_coord.y0[-9] ;
 wire \i_coord.y0[0] ;
 wire \i_coord.y0[1] ;
 wire \i_coord.y_inc_row[-10] ;
 wire \i_coord.y_inc_row[-11] ;
 wire \i_coord.y_inc_row[-12] ;
 wire \i_coord.y_inc_row[-13] ;
 wire \i_coord.y_inc_row[-6] ;
 wire \i_coord.y_inc_row[-7] ;
 wire \i_coord.y_inc_row[-8] ;
 wire \i_coord.y_inc_row[-9] ;
 wire \i_coord.y_row_start[-10] ;
 wire \i_coord.y_row_start[-11] ;
 wire \i_coord.y_row_start[-12] ;
 wire \i_coord.y_row_start[-13] ;
 wire \i_coord.y_row_start[-1] ;
 wire \i_coord.y_row_start[-2] ;
 wire \i_coord.y_row_start[-3] ;
 wire \i_coord.y_row_start[-4] ;
 wire \i_coord.y_row_start[-5] ;
 wire \i_coord.y_row_start[-6] ;
 wire \i_coord.y_row_start[-7] ;
 wire \i_coord.y_row_start[-8] ;
 wire \i_coord.y_row_start[-9] ;
 wire \i_coord.y_row_start[0] ;
 wire \i_coord.y_row_start[1] ;
 wire \i_mandel.i_xy.hc.gated_clk ;
 wire \i_mandel.i_xy.hc.genblk1.genblk1.CG.GATE ;
 wire \i_mandel.i_xy.hc.genblk2[0].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[0].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[10].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[10].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[11].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[11].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[1].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[1].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[2].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[2].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[3].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[3].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[4].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[4].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[5].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[5].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[6].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[6].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[7].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[7].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[8].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[8].state.Q ;
 wire \i_mandel.i_xy.hc.genblk2[9].state.D ;
 wire \i_mandel.i_xy.hc.genblk2[9].state.Q ;
 wire \i_mandel.i_xy.phase ;
 wire \i_mandel.i_xy.x[-10] ;
 wire \i_mandel.i_xy.x[-11] ;
 wire \i_mandel.i_xy.x[-12] ;
 wire \i_mandel.i_xy.x[-13] ;
 wire \i_mandel.i_xy.x[-1] ;
 wire \i_mandel.i_xy.x[-2] ;
 wire \i_mandel.i_xy.x[-3] ;
 wire \i_mandel.i_xy.x[-4] ;
 wire \i_mandel.i_xy.x[-5] ;
 wire \i_mandel.i_xy.x[-6] ;
 wire \i_mandel.i_xy.x[-7] ;
 wire \i_mandel.i_xy.x[-8] ;
 wire \i_mandel.i_xy.x[-9] ;
 wire \i_mandel.i_xy.x[0] ;
 wire \i_mandel.i_xy.x[1] ;
 wire \i_mandel.i_xy.x[2] ;
 wire \i_mandel.i_xy.y[-10] ;
 wire \i_mandel.i_xy.y[-11] ;
 wire \i_mandel.i_xy.y[-12] ;
 wire \i_mandel.i_xy.y[-13] ;
 wire \i_mandel.i_xy.y[-1] ;
 wire \i_mandel.i_xy.y[-2] ;
 wire \i_mandel.i_xy.y[-3] ;
 wire \i_mandel.i_xy.y[-4] ;
 wire \i_mandel.i_xy.y[-5] ;
 wire \i_mandel.i_xy.y[-6] ;
 wire \i_mandel.i_xy.y[-7] ;
 wire \i_mandel.i_xy.y[-8] ;
 wire \i_mandel.i_xy.y[-9] ;
 wire \i_mandel.i_xy.y[0] ;
 wire \i_mandel.i_xy.y[1] ;
 wire \i_mandel.i_xy.y[2] ;
 wire \i_mandel.l_sq.genblk2[0].state.D ;
 wire \i_mandel.l_sq.genblk2[0].state.Q ;
 wire \i_mandel.l_sq.genblk2[10].state.D ;
 wire \i_mandel.l_sq.genblk2[10].state.Q ;
 wire \i_mandel.l_sq.genblk2[11].state.D ;
 wire \i_mandel.l_sq.genblk2[11].state.Q ;
 wire \i_mandel.l_sq.genblk2[12].state.D ;
 wire \i_mandel.l_sq.genblk2[12].state.Q ;
 wire \i_mandel.l_sq.genblk2[13].state.D ;
 wire \i_mandel.l_sq.genblk2[13].state.Q ;
 wire \i_mandel.l_sq.genblk2[14].state.D ;
 wire \i_mandel.l_sq.genblk2[14].state.Q ;
 wire \i_mandel.l_sq.genblk2[15].state.D ;
 wire \i_mandel.l_sq.genblk2[15].state.Q ;
 wire \i_mandel.l_sq.genblk2[16].state.D ;
 wire \i_mandel.l_sq.genblk2[16].state.Q ;
 wire \i_mandel.l_sq.genblk2[17].state.D ;
 wire \i_mandel.l_sq.genblk2[17].state.Q ;
 wire \i_mandel.l_sq.genblk2[18].state.D ;
 wire \i_mandel.l_sq.genblk2[18].state.Q ;
 wire \i_mandel.l_sq.genblk2[1].state.D ;
 wire \i_mandel.l_sq.genblk2[1].state.Q ;
 wire \i_mandel.l_sq.genblk2[2].state.D ;
 wire \i_mandel.l_sq.genblk2[2].state.Q ;
 wire \i_mandel.l_sq.genblk2[3].state.D ;
 wire \i_mandel.l_sq.genblk2[3].state.Q ;
 wire \i_mandel.l_sq.genblk2[4].state.D ;
 wire \i_mandel.l_sq.genblk2[4].state.Q ;
 wire \i_mandel.l_sq.genblk2[5].state.D ;
 wire \i_mandel.l_sq.genblk2[5].state.Q ;
 wire \i_mandel.l_sq.genblk2[6].state.D ;
 wire \i_mandel.l_sq.genblk2[6].state.Q ;
 wire \i_mandel.l_sq.genblk2[7].state.D ;
 wire \i_mandel.l_sq.genblk2[7].state.Q ;
 wire \i_mandel.l_sq.genblk2[8].state.D ;
 wire \i_mandel.l_sq.genblk2[8].state.Q ;
 wire \i_mandel.l_sq.genblk2[9].state.D ;
 wire \i_mandel.l_sq.genblk2[9].state.Q ;
 wire \i_vga.hsync ;
 wire \i_vga.timing_hor.counter[0] ;
 wire \i_vga.timing_hor.counter[10] ;
 wire \i_vga.timing_hor.counter[1] ;
 wire \i_vga.timing_hor.counter[2] ;
 wire \i_vga.timing_hor.counter[3] ;
 wire \i_vga.timing_hor.counter[4] ;
 wire \i_vga.timing_hor.counter[5] ;
 wire \i_vga.timing_hor.counter[6] ;
 wire \i_vga.timing_hor.counter[7] ;
 wire \i_vga.timing_hor.counter[8] ;
 wire \i_vga.timing_hor.counter[9] ;
 wire \i_vga.timing_ver.blank ;
 wire \i_vga.timing_ver.counter[0] ;
 wire \i_vga.timing_ver.counter[1] ;
 wire \i_vga.timing_ver.counter[2] ;
 wire \i_vga.timing_ver.counter[3] ;
 wire \i_vga.timing_ver.counter[4] ;
 wire \i_vga.timing_ver.counter[5] ;
 wire \i_vga.timing_ver.counter[6] ;
 wire \i_vga.timing_ver.counter[7] ;
 wire \i_vga.timing_ver.counter[8] ;
 wire \i_vga.timing_ver.counter[9] ;
 wire \i_vga.timing_ver.sync ;
 wire \i_vga.timing_ver.sync_tmp ;
 wire \i_vga.vblank ;
 wire \iter[0] ;
 wire \iter[1] ;
 wire \iter[2] ;
 wire \iter[3] ;
 wire \last_iter[0] ;
 wire \last_iter[1] ;
 wire \last_iter[2] ;
 wire \last_iter[3] ;
 wire \step[1] ;
 wire \step[2] ;
 wire \step[3] ;
 wire \step[4] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire \video_colour[0] ;
 wire \video_colour[1] ;
 wire \video_colour[2] ;
 wire \video_colour[3] ;
 wire \video_colour[4] ;
 wire \video_colour[5] ;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire \clknet_0_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_3_0__leaf_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_3_1__leaf_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_3_2__leaf_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_3_3__leaf_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_3_4__leaf_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_3_5__leaf_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_3_6__leaf_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_3_7__leaf_i_mandel.i_xy.hc.gated_clk ;
 wire \clknet_0_i_coord.l_xl.gated_clk ;
 wire \clknet_1_0__leaf_i_coord.l_xl.gated_clk ;
 wire \clknet_1_1__leaf_i_coord.l_xl.gated_clk ;
 wire \clknet_0_i_coord.l_yt.gated_clk ;
 wire \clknet_2_0__leaf_i_coord.l_yt.gated_clk ;
 wire \clknet_2_1__leaf_i_coord.l_yt.gated_clk ;
 wire \clknet_2_2__leaf_i_coord.l_yt.gated_clk ;
 wire \clknet_2_3__leaf_i_coord.l_yt.gated_clk ;
 wire \clknet_0_i_coord.l_xip.gated_clk ;
 wire \clknet_1_0__leaf_i_coord.l_xip.gated_clk ;
 wire \clknet_1_1__leaf_i_coord.l_xip.gated_clk ;
 wire \clknet_0_i_coord.l_yip.gated_clk ;
 wire \clknet_1_0__leaf_i_coord.l_yip.gated_clk ;
 wire \clknet_1_1__leaf_i_coord.l_yip.gated_clk ;
 wire \clknet_0_i_coord.l_xir.gated_clk ;
 wire \clknet_1_0__leaf_i_coord.l_xir.gated_clk ;
 wire \clknet_1_1__leaf_i_coord.l_xir.gated_clk ;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net319;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;

 sg13g2_inv_1 _3796_ (.Y(_3084_),
    .A(\i_vga.timing_hor.counter[10] ));
 sg13g2_inv_1 _3797_ (.Y(_3085_),
    .A(net235));
 sg13g2_inv_1 _3798_ (.Y(_3086_),
    .A(net280));
 sg13g2_inv_1 _3799_ (.Y(_3087_),
    .A(net322));
 sg13g2_inv_1 _3800_ (.Y(_3088_),
    .A(net182));
 sg13g2_inv_1 _3801_ (.Y(_3089_),
    .A(\i_mandel.l_sq.genblk2[14].state.Q ));
 sg13g2_inv_1 _3802_ (.Y(_3090_),
    .A(\i_mandel.l_sq.genblk2[13].state.Q ));
 sg13g2_inv_1 _3803_ (.Y(_3091_),
    .A(\i_mandel.l_sq.genblk2[9].state.Q ));
 sg13g2_inv_1 _3804_ (.Y(_3092_),
    .A(\i_mandel.l_sq.genblk2[7].state.Q ));
 sg13g2_inv_1 _3805_ (.Y(_3093_),
    .A(net3));
 sg13g2_inv_1 _3806_ (.Y(_3094_),
    .A(net367));
 sg13g2_inv_1 _3807_ (.Y(_3095_),
    .A(net940));
 sg13g2_inv_1 _3808_ (.Y(_3096_),
    .A(net6));
 sg13g2_inv_1 _3809_ (.Y(_3097_),
    .A(net7));
 sg13g2_inv_1 _3810_ (.Y(_3098_),
    .A(net258));
 sg13g2_inv_1 _3811_ (.Y(_3099_),
    .A(net237));
 sg13g2_inv_1 _3812_ (.Y(_3100_),
    .A(net265));
 sg13g2_inv_1 _3813_ (.Y(_3101_),
    .A(net239));
 sg13g2_inv_1 _3814_ (.Y(_3102_),
    .A(net806));
 sg13g2_inv_1 _3815_ (.Y(_3103_),
    .A(net218));
 sg13g2_inv_1 _3816_ (.Y(_3104_),
    .A(net268));
 sg13g2_inv_1 _3817_ (.Y(_3105_),
    .A(net259));
 sg13g2_inv_1 _3818_ (.Y(_3106_),
    .A(net257));
 sg13g2_inv_1 _3819_ (.Y(_3107_),
    .A(net238));
 sg13g2_inv_1 _3820_ (.Y(_3108_),
    .A(net281));
 sg13g2_inv_1 _3821_ (.Y(_3109_),
    .A(net269));
 sg13g2_inv_1 _3822_ (.Y(_3110_),
    .A(net251));
 sg13g2_inv_1 _3823_ (.Y(_3111_),
    .A(net225));
 sg13g2_inv_1 _3824_ (.Y(_3112_),
    .A(net270));
 sg13g2_inv_1 _3825_ (.Y(_3113_),
    .A(net232));
 sg13g2_inv_1 _3826_ (.Y(_3114_),
    .A(\i_coord.l_yt.genblk2[14].state.Q ));
 sg13g2_inv_1 _3827_ (.Y(_3115_),
    .A(net961));
 sg13g2_inv_1 _3828_ (.Y(_3116_),
    .A(net246));
 sg13g2_inv_1 _3829_ (.Y(_3117_),
    .A(net250));
 sg13g2_inv_1 _3830_ (.Y(_3118_),
    .A(net304));
 sg13g2_inv_1 _3831_ (.Y(_3119_),
    .A(net361));
 sg13g2_inv_1 _3832_ (.Y(_3120_),
    .A(net207));
 sg13g2_inv_1 _3833_ (.Y(_3121_),
    .A(\i_coord.y0[-7] ));
 sg13g2_inv_1 _3834_ (.Y(_3122_),
    .A(net341));
 sg13g2_inv_2 _3835_ (.Y(_3123_),
    .A(net314));
 sg13g2_inv_1 _3836_ (.Y(_3124_),
    .A(net349));
 sg13g2_inv_1 _3837_ (.Y(_3125_),
    .A(net307));
 sg13g2_inv_2 _3838_ (.Y(_3126_),
    .A(net14));
 sg13g2_inv_2 _3839_ (.Y(_3127_),
    .A(net309));
 sg13g2_inv_2 _3840_ (.Y(_3128_),
    .A(net15));
 sg13g2_inv_1 _3841_ (.Y(_3129_),
    .A(net288));
 sg13g2_inv_1 _3842_ (.Y(_3130_),
    .A(_0020_));
 sg13g2_inv_1 _3843_ (.Y(_3131_),
    .A(net894));
 sg13g2_inv_1 _3844_ (.Y(_3132_),
    .A(net884));
 sg13g2_inv_2 _3845_ (.Y(_3133_),
    .A(net911));
 sg13g2_inv_1 _3846_ (.Y(_3134_),
    .A(\i_coord.l_yip.genblk2[7].state.Q ));
 sg13g2_inv_1 _3847_ (.Y(_3135_),
    .A(\i_mandel.i_xy.y[2] ));
 sg13g2_inv_1 _3848_ (.Y(_3136_),
    .A(net803));
 sg13g2_inv_1 _3849_ (.Y(_3137_),
    .A(net189));
 sg13g2_inv_1 _3850_ (.Y(_3138_),
    .A(net350));
 sg13g2_inv_1 _3851_ (.Y(_3139_),
    .A(net294));
 sg13g2_inv_1 _3852_ (.Y(_3140_),
    .A(\i_mandel.l_sq.genblk2[0].state.Q ));
 sg13g2_inv_1 _3853_ (.Y(_3141_),
    .A(net277));
 sg13g2_inv_1 _3854_ (.Y(_3142_),
    .A(net300));
 sg13g2_inv_1 _3855_ (.Y(_3143_),
    .A(net289));
 sg13g2_inv_1 _3856_ (.Y(_3144_),
    .A(\i_coord.x0[-6] ));
 sg13g2_inv_1 _3857_ (.Y(_3145_),
    .A(\i_coord.x0[1] ));
 sg13g2_inv_1 _3858_ (.Y(_3146_),
    .A(net348));
 sg13g2_and3_1 _3859_ (.X(_3147_),
    .A(\i_vga.timing_ver.counter[8] ),
    .B(\i_vga.timing_ver.counter[7] ),
    .C(\i_vga.timing_ver.counter[6] ));
 sg13g2_nand4_1 _3860_ (.B(\i_vga.timing_ver.counter[5] ),
    .C(\i_vga.timing_ver.counter[4] ),
    .A(\i_vga.timing_ver.counter[9] ),
    .Y(_3148_),
    .D(_3147_));
 sg13g2_o21ai_1 _3861_ (.B1(\i_vga.timing_ver.counter[3] ),
    .Y(_3149_),
    .A1(\i_vga.timing_ver.counter[2] ),
    .A2(\i_vga.timing_ver.counter[1] ));
 sg13g2_inv_1 _3862_ (.Y(_3150_),
    .A(_3149_));
 sg13g2_nor3_1 _3863_ (.A(net180),
    .B(_3148_),
    .C(_3150_),
    .Y(\i_vga.timing_ver.sync_tmp ));
 sg13g2_nor2_1 _3864_ (.A(\i_vga.timing_hor.counter[10] ),
    .B(\i_vga.vblank ),
    .Y(_3151_));
 sg13g2_or2_1 _3865_ (.X(_3152_),
    .B(\i_vga.vblank ),
    .A(\i_vga.timing_hor.counter[10] ));
 sg13g2_and2_1 _3866_ (.A(\video_colour[5] ),
    .B(net873),
    .X(uo_out[0]));
 sg13g2_and2_1 _3867_ (.A(\video_colour[3] ),
    .B(net873),
    .X(uo_out[1]));
 sg13g2_and2_1 _3868_ (.A(\video_colour[1] ),
    .B(net873),
    .X(uo_out[2]));
 sg13g2_and2_1 _3869_ (.A(\video_colour[4] ),
    .B(net872),
    .X(uo_out[4]));
 sg13g2_and2_1 _3870_ (.A(\video_colour[2] ),
    .B(net872),
    .X(uo_out[5]));
 sg13g2_and2_1 _3871_ (.A(\video_colour[0] ),
    .B(net872),
    .X(uo_out[6]));
 sg13g2_nor2_2 _3872_ (.A(net940),
    .B(net959),
    .Y(_3153_));
 sg13g2_and2_1 _3873_ (.A(net4),
    .B(net965),
    .X(\i_coord.l_xir.genblk2[0].state.D ));
 sg13g2_and2_1 _3874_ (.A(net881),
    .B(\i_coord.l_xir.genblk2[0].state.D ),
    .X(\i_coord.l_xip.genblk2[0].state.D ));
 sg13g2_and2_1 _3875_ (.A(net5),
    .B(net964),
    .X(\i_coord.l_xir.genblk2[1].state.D ));
 sg13g2_and2_1 _3876_ (.A(net881),
    .B(\i_coord.l_xir.genblk2[1].state.D ),
    .X(\i_coord.l_xip.genblk2[1].state.D ));
 sg13g2_nor2_2 _3877_ (.A(_3096_),
    .B(net959),
    .Y(\i_coord.l_xir.genblk2[2].state.D ));
 sg13g2_o21ai_1 _3878_ (.B1(net965),
    .Y(_3154_),
    .A1(net938),
    .A2(net6));
 sg13g2_nand2_1 _3879_ (.Y(_3155_),
    .A(\i_coord.y_inc_row[-8] ),
    .B(\i_coord.y_inc_row[-9] ));
 sg13g2_nor3_1 _3880_ (.A(\i_coord.y_inc_row[-10] ),
    .B(\i_coord.y_inc_row[-11] ),
    .C(_3155_),
    .Y(_3156_));
 sg13g2_nand2_1 _3881_ (.Y(_3157_),
    .A(net946),
    .B(net947));
 sg13g2_nor2_1 _3882_ (.A(net945),
    .B(\i_coord.y_inc_row[-7] ),
    .Y(_3158_));
 sg13g2_and4_2 _3883_ (.A(net946),
    .B(net947),
    .C(_3156_),
    .D(_3158_),
    .X(_3159_));
 sg13g2_nand4_1 _3884_ (.B(net947),
    .C(_3156_),
    .A(net946),
    .Y(_3160_),
    .D(_3158_));
 sg13g2_nand3_1 _3885_ (.B(net946),
    .C(net947),
    .A(\i_coord.y_inc_row[-11] ),
    .Y(_3161_));
 sg13g2_nand4_1 _3886_ (.B(\i_coord.y_inc_row[-11] ),
    .C(net946),
    .A(\i_coord.y_inc_row[-10] ),
    .Y(_3162_),
    .D(net947));
 sg13g2_inv_1 _3887_ (.Y(_3163_),
    .A(_3162_));
 sg13g2_nor2_1 _3888_ (.A(_3155_),
    .B(_3162_),
    .Y(_3164_));
 sg13g2_nand2_1 _3889_ (.Y(_3165_),
    .A(\i_coord.y_inc_row[-7] ),
    .B(_3164_));
 sg13g2_xor2_1 _3890_ (.B(_3165_),
    .A(net945),
    .X(_3166_));
 sg13g2_and2_1 _3891_ (.A(_3160_),
    .B(_3166_),
    .X(_3167_));
 sg13g2_nand2_2 _3892_ (.Y(_3168_),
    .A(_3160_),
    .B(_3166_));
 sg13g2_nand3b_1 _3893_ (.B(net947),
    .C(_3160_),
    .Y(_3169_),
    .A_N(_3166_));
 sg13g2_o21ai_1 _3894_ (.B1(_3169_),
    .Y(_3170_),
    .A1(net947),
    .A2(_3168_));
 sg13g2_inv_1 _3895_ (.Y(_3171_),
    .A(_3170_));
 sg13g2_a21oi_1 _3896_ (.A1(net939),
    .A2(_3171_),
    .Y(\i_coord.l_xip.genblk2[2].state.D ),
    .B1(_3154_));
 sg13g2_xor2_1 _3897_ (.B(net947),
    .A(net946),
    .X(_3172_));
 sg13g2_nand2_1 _3898_ (.Y(_3173_),
    .A(net938),
    .B(_3172_));
 sg13g2_nor2_2 _3899_ (.A(_3097_),
    .B(net959),
    .Y(\i_coord.l_xir.genblk2[3].state.D ));
 sg13g2_o21ai_1 _3900_ (.B1(net964),
    .Y(_3174_),
    .A1(net939),
    .A2(net7));
 sg13g2_nor2_1 _3901_ (.A(net880),
    .B(_3168_),
    .Y(_3175_));
 sg13g2_nand2_1 _3902_ (.Y(_3176_),
    .A(net938),
    .B(_3167_));
 sg13g2_nor2_1 _3903_ (.A(_3172_),
    .B(_3175_),
    .Y(_3177_));
 sg13g2_nand2_1 _3904_ (.Y(_3178_),
    .A(net938),
    .B(_3168_));
 sg13g2_a21oi_1 _3905_ (.A1(_3172_),
    .A2(_3178_),
    .Y(_3179_),
    .B1(_3177_));
 sg13g2_nor2_1 _3906_ (.A(_3174_),
    .B(_3179_),
    .Y(\i_coord.l_xip.genblk2[3].state.D ));
 sg13g2_xor2_1 _3907_ (.B(_3157_),
    .A(\i_coord.y_inc_row[-11] ),
    .X(_3180_));
 sg13g2_and2_1 _3908_ (.A(net938),
    .B(_3180_),
    .X(_3181_));
 sg13g2_a221oi_1 _3909_ (.B2(_3181_),
    .C1(net958),
    .B1(_3168_),
    .A1(net881),
    .Y(_3182_),
    .A2(net8));
 sg13g2_o21ai_1 _3910_ (.B1(_3182_),
    .Y(\i_coord.l_xip.genblk2[4].state.D ),
    .A1(_3176_),
    .A2(_3180_));
 sg13g2_xor2_1 _3911_ (.B(_3161_),
    .A(\i_coord.y_inc_row[-10] ),
    .X(_3183_));
 sg13g2_nand3_1 _3912_ (.B(_3160_),
    .C(_3183_),
    .A(net939),
    .Y(_3184_));
 sg13g2_a22oi_1 _3913_ (.Y(_3185_),
    .B1(_3184_),
    .B2(_3176_),
    .A2(_3183_),
    .A1(_3167_));
 sg13g2_nand2_2 _3914_ (.Y(_3186_),
    .A(net880),
    .B(net9));
 sg13g2_nand3b_1 _3915_ (.B(_3186_),
    .C(net964),
    .Y(\i_coord.l_xip.genblk2[5].state.D ),
    .A_N(_3185_));
 sg13g2_xor2_1 _3916_ (.B(_3162_),
    .A(\i_coord.y_inc_row[-9] ),
    .X(_3187_));
 sg13g2_nor2_1 _3917_ (.A(_3159_),
    .B(_3187_),
    .Y(_3188_));
 sg13g2_nand2_1 _3918_ (.Y(_3189_),
    .A(net938),
    .B(_3188_));
 sg13g2_nand2_1 _3919_ (.Y(_3190_),
    .A(net880),
    .B(net10));
 sg13g2_a221oi_1 _3920_ (.B2(_3188_),
    .C1(net958),
    .B1(_3175_),
    .A1(net880),
    .Y(_3191_),
    .A2(net10));
 sg13g2_o21ai_1 _3921_ (.B1(_3191_),
    .Y(\i_coord.l_xip.genblk2[6].state.D ),
    .A1(_3178_),
    .A2(_3188_));
 sg13g2_a21oi_1 _3922_ (.A1(\i_coord.y_inc_row[-9] ),
    .A2(_3163_),
    .Y(_3192_),
    .B1(net308));
 sg13g2_nor3_2 _3923_ (.A(_3159_),
    .B(_3164_),
    .C(_3192_),
    .Y(_3193_));
 sg13g2_nand2_1 _3924_ (.Y(_3194_),
    .A(net938),
    .B(_3193_));
 sg13g2_a221oi_1 _3925_ (.B2(_3193_),
    .C1(net958),
    .B1(_3175_),
    .A1(net880),
    .Y(_3195_),
    .A2(net11));
 sg13g2_o21ai_1 _3926_ (.B1(_3195_),
    .Y(\i_coord.l_xip.genblk2[7].state.D ),
    .A1(_3178_),
    .A2(_3193_));
 sg13g2_and2_1 _3927_ (.A(net967),
    .B(net12),
    .X(\i_coord.l_xl.genblk2[11].state.D ));
 sg13g2_o21ai_1 _3928_ (.B1(net964),
    .Y(_3196_),
    .A1(net939),
    .A2(net12));
 sg13g2_or2_1 _3929_ (.X(_3197_),
    .B(_3164_),
    .A(\i_coord.y_inc_row[-7] ));
 sg13g2_a21o_1 _3930_ (.A2(_3197_),
    .A1(_3165_),
    .B1(_3159_),
    .X(_3198_));
 sg13g2_o21ai_1 _3931_ (.B1(net938),
    .Y(_3199_),
    .A1(_3166_),
    .A2(_3198_));
 sg13g2_a21oi_1 _3932_ (.A1(_3167_),
    .A2(_3198_),
    .Y(_3200_),
    .B1(_3199_));
 sg13g2_nor2_1 _3933_ (.A(_3196_),
    .B(_3200_),
    .Y(\i_coord.l_xip.genblk2[8].state.D ));
 sg13g2_and2_1 _3934_ (.A(net967),
    .B(net13),
    .X(\i_coord.l_xl.genblk2[12].state.D ));
 sg13g2_and2_2 _3935_ (.A(net880),
    .B(\i_coord.l_xl.genblk2[12].state.D ),
    .X(\i_coord.l_xip.genblk2[9].state.D ));
 sg13g2_nand3b_1 _3936_ (.B(_3160_),
    .C(net965),
    .Y(_3201_),
    .A_N(_0027_));
 sg13g2_nor2_1 _3937_ (.A(net333),
    .B(_3201_),
    .Y(\i_coord.l_yt.genblk2[0].state.D ));
 sg13g2_nor2_1 _3938_ (.A(net335),
    .B(_3201_),
    .Y(\i_coord.l_yt.genblk2[1].state.D ));
 sg13g2_nor3_2 _3939_ (.A(net881),
    .B(net958),
    .C(_3159_),
    .Y(_3202_));
 sg13g2_a21oi_1 _3940_ (.A1(\i_coord.y0[-11] ),
    .A2(net802),
    .Y(_3203_),
    .B1(\i_coord.l_xip.genblk2[0].state.D ));
 sg13g2_inv_1 _3941_ (.Y(\i_coord.l_yt.genblk2[2].state.D ),
    .A(_3203_));
 sg13g2_a21oi_1 _3942_ (.A1(\i_coord.y0[-10] ),
    .A2(net802),
    .Y(_3204_),
    .B1(\i_coord.l_xip.genblk2[1].state.D ));
 sg13g2_inv_1 _3943_ (.Y(\i_coord.l_yt.genblk2[3].state.D ),
    .A(_3204_));
 sg13g2_a21oi_1 _3944_ (.A1(_3119_),
    .A2(_3160_),
    .Y(_3205_),
    .B1(net882));
 sg13g2_nor2_1 _3945_ (.A(_3154_),
    .B(_3205_),
    .Y(\i_coord.l_yt.genblk2[4].state.D ));
 sg13g2_nand2_2 _3946_ (.Y(_3206_),
    .A(\i_coord.y0[-9] ),
    .B(net937));
 sg13g2_nand2_1 _3947_ (.Y(_3207_),
    .A(_3119_),
    .B(_3120_));
 sg13g2_nand3_1 _3948_ (.B(_3206_),
    .C(_3207_),
    .A(_3160_),
    .Y(_3208_));
 sg13g2_a21oi_1 _3949_ (.A1(net940),
    .A2(_3208_),
    .Y(\i_coord.l_yt.genblk2[5].state.D ),
    .B1(_3174_));
 sg13g2_xor2_1 _3950_ (.B(_3206_),
    .A(_0024_),
    .X(_3209_));
 sg13g2_and2_1 _3951_ (.A(net802),
    .B(_3209_),
    .X(_3210_));
 sg13g2_and2_2 _3952_ (.A(net8),
    .B(net964),
    .X(\i_coord.l_xir.genblk2[4].state.D ));
 sg13g2_a21o_1 _3953_ (.A2(\i_coord.l_xir.genblk2[4].state.D ),
    .A1(net882),
    .B1(_3210_),
    .X(\i_coord.l_yt.genblk2[6].state.D ));
 sg13g2_and2_1 _3954_ (.A(net9),
    .B(net964),
    .X(\i_coord.l_xir.genblk2[5].state.D ));
 sg13g2_nand4_1 _3955_ (.B(net937),
    .C(\i_coord.y0[-7] ),
    .A(\i_coord.y0[-9] ),
    .Y(_3211_),
    .D(\i_coord.y0[-6] ));
 sg13g2_o21ai_1 _3956_ (.B1(_3122_),
    .Y(_3212_),
    .A1(_3121_),
    .A2(_3206_));
 sg13g2_nand3_1 _3957_ (.B(_3211_),
    .C(_3212_),
    .A(_3202_),
    .Y(_3213_));
 sg13g2_o21ai_1 _3958_ (.B1(_3213_),
    .Y(\i_coord.l_yt.genblk2[7].state.D ),
    .A1(net959),
    .A2(_3186_));
 sg13g2_and2_1 _3959_ (.A(_3123_),
    .B(_3211_),
    .X(_3214_));
 sg13g2_nor2_1 _3960_ (.A(_3123_),
    .B(_3211_),
    .Y(_3215_));
 sg13g2_o21ai_1 _3961_ (.B1(_3202_),
    .Y(_3216_),
    .A1(_3214_),
    .A2(_3215_));
 sg13g2_nand2_2 _3962_ (.Y(_3217_),
    .A(net10),
    .B(net964));
 sg13g2_inv_1 _3963_ (.Y(\i_coord.l_xir.genblk2[6].state.D ),
    .A(_3217_));
 sg13g2_o21ai_1 _3964_ (.B1(_3216_),
    .Y(\i_coord.l_yt.genblk2[8].state.D ),
    .A1(net940),
    .A2(_3217_));
 sg13g2_and2_1 _3965_ (.A(_3124_),
    .B(_3214_),
    .X(_3218_));
 sg13g2_nor2_1 _3966_ (.A(_3124_),
    .B(_3214_),
    .Y(_3219_));
 sg13g2_o21ai_1 _3967_ (.B1(net802),
    .Y(_3220_),
    .A1(_3218_),
    .A2(_3219_));
 sg13g2_nand2_2 _3968_ (.Y(_3221_),
    .A(net11),
    .B(net964));
 sg13g2_inv_1 _3969_ (.Y(\i_coord.l_xir.genblk2[7].state.D ),
    .A(_3221_));
 sg13g2_o21ai_1 _3970_ (.B1(_3220_),
    .Y(\i_coord.l_yt.genblk2[9].state.D ),
    .A1(net940),
    .A2(_3221_));
 sg13g2_xnor2_1 _3971_ (.Y(_3222_),
    .A(_0023_),
    .B(_3218_));
 sg13g2_a21oi_1 _3972_ (.A1(_3160_),
    .A2(_3222_),
    .Y(_3223_),
    .B1(net882));
 sg13g2_nor2_1 _3973_ (.A(_3196_),
    .B(_3223_),
    .Y(\i_coord.l_yt.genblk2[10].state.D ));
 sg13g2_nor2b_1 _3974_ (.A(\i_coord.y0[-3] ),
    .B_N(_3218_),
    .Y(_3224_));
 sg13g2_xnor2_1 _3975_ (.Y(_3225_),
    .A(_0022_),
    .B(_3224_));
 sg13g2_a21oi_1 _3976_ (.A1(net802),
    .A2(_3225_),
    .Y(_3226_),
    .B1(\i_coord.l_xip.genblk2[9].state.D ));
 sg13g2_inv_1 _3977_ (.Y(\i_coord.l_yt.genblk2[11].state.D ),
    .A(_3226_));
 sg13g2_nor2b_1 _3978_ (.A(\i_coord.y0[-2] ),
    .B_N(_3224_),
    .Y(_3227_));
 sg13g2_nand2_1 _3979_ (.Y(_3228_),
    .A(net363),
    .B(_3227_));
 sg13g2_o21ai_1 _3980_ (.B1(net802),
    .Y(_3229_),
    .A1(_0021_),
    .A2(_3227_));
 sg13g2_inv_1 _3981_ (.Y(_3230_),
    .A(_3229_));
 sg13g2_a22oi_1 _3982_ (.Y(\i_coord.l_yt.genblk2[12].state.D ),
    .B1(_3228_),
    .B2(_3230_),
    .A2(_3153_),
    .A1(_3126_));
 sg13g2_nand2_1 _3983_ (.Y(\i_coord.l_xl.genblk2[14].state.D ),
    .A(net963),
    .B(_3128_));
 sg13g2_xnor2_1 _3984_ (.Y(_3231_),
    .A(_3127_),
    .B(_3228_));
 sg13g2_a22oi_1 _3985_ (.Y(\i_coord.l_yt.genblk2[13].state.D ),
    .B1(_3202_),
    .B2(_3231_),
    .A2(_3153_),
    .A1(_3128_));
 sg13g2_nand2_1 _3986_ (.Y(_3232_),
    .A(net16),
    .B(_3153_));
 sg13g2_and3_1 _3987_ (.X(_3233_),
    .A(_3125_),
    .B(_3127_),
    .C(_3227_));
 sg13g2_and2_1 _3988_ (.A(_3130_),
    .B(_3233_),
    .X(_3234_));
 sg13g2_o21ai_1 _3989_ (.B1(net802),
    .Y(_3235_),
    .A1(_3130_),
    .A2(_3233_));
 sg13g2_o21ai_1 _3990_ (.B1(_3232_),
    .Y(\i_coord.l_yt.genblk2[14].state.D ),
    .A1(_3234_),
    .A2(_3235_));
 sg13g2_nor2_1 _3991_ (.A(net960),
    .B(_3126_),
    .Y(\i_coord.l_xl.genblk2[13].state.D ));
 sg13g2_nand2b_1 _3992_ (.Y(\i_coord.l_xl.genblk2[15].state.D ),
    .B(net963),
    .A_N(net16));
 sg13g2_nor2b_1 _3993_ (.A(\step[2] ),
    .B_N(\step[1] ),
    .Y(_3236_));
 sg13g2_and3_1 _3994_ (.X(_3237_),
    .A(\step[3] ),
    .B(\step[4] ),
    .C(_3236_));
 sg13g2_nand3_1 _3995_ (.B(\step[4] ),
    .C(_3236_),
    .A(\step[3] ),
    .Y(_3238_));
 sg13g2_and2_1 _3996_ (.A(net957),
    .B(\step[1] ),
    .X(_3239_));
 sg13g2_nand2_2 _3997_ (.Y(_3240_),
    .A(net949),
    .B(net214));
 sg13g2_and2_1 _3998_ (.A(net278),
    .B(net866),
    .X(_3241_));
 sg13g2_nand2_2 _3999_ (.Y(_3242_),
    .A(net278),
    .B(net866));
 sg13g2_nand3_1 _4000_ (.B(\i_vga.timing_hor.counter[1] ),
    .C(_3241_),
    .A(net196),
    .Y(_3243_));
 sg13g2_or2_1 _4001_ (.X(_3244_),
    .B(_3243_),
    .A(_3085_));
 sg13g2_or2_1 _4002_ (.X(_3245_),
    .B(_3244_),
    .A(net241));
 sg13g2_nand4_1 _4003_ (.B(\i_vga.timing_hor.counter[9] ),
    .C(\i_vga.timing_hor.counter[7] ),
    .A(_3084_),
    .Y(_3246_),
    .D(\i_vga.timing_hor.counter[6] ));
 sg13g2_nor4_2 _4004_ (.A(\i_vga.timing_hor.counter[8] ),
    .B(\i_vga.timing_hor.counter[5] ),
    .C(_3245_),
    .Y(_3247_),
    .D(_3246_));
 sg13g2_or4_1 _4005_ (.A(\i_vga.timing_hor.counter[8] ),
    .B(\i_vga.timing_hor.counter[5] ),
    .C(_3245_),
    .D(_3246_),
    .X(_3248_));
 sg13g2_nand3_1 _4006_ (.B(\i_vga.timing_ver.counter[2] ),
    .C(\i_vga.timing_ver.counter[1] ),
    .A(\i_vga.timing_ver.counter[3] ),
    .Y(_3249_));
 sg13g2_nor4_2 _4007_ (.A(\i_vga.timing_ver.counter[0] ),
    .B(_3148_),
    .C(_3248_),
    .Y(_3250_),
    .D(_3249_));
 sg13g2_or4_1 _4008_ (.A(\i_vga.timing_ver.counter[0] ),
    .B(_3148_),
    .C(_3248_),
    .D(_3249_),
    .X(_3251_));
 sg13g2_nor2_1 _4009_ (.A(net254),
    .B(net264),
    .Y(_3252_));
 sg13g2_nand2b_1 _4010_ (.Y(_3253_),
    .B(\i_vga.timing_hor.counter[5] ),
    .A_N(\i_vga.timing_hor.counter[4] ));
 sg13g2_and2_1 _4011_ (.A(\i_vga.timing_hor.counter[9] ),
    .B(\i_vga.timing_hor.counter[8] ),
    .X(_3254_));
 sg13g2_nor3_1 _4012_ (.A(\i_vga.timing_hor.counter[7] ),
    .B(_0032_),
    .C(_3253_),
    .Y(_3255_));
 sg13g2_nand3_1 _4013_ (.B(_3254_),
    .C(_3255_),
    .A(net941),
    .Y(_3256_));
 sg13g2_nand3b_1 _4014_ (.B(_3086_),
    .C(\i_vga.timing_hor.counter[3] ),
    .Y(_3257_),
    .A_N(\i_vga.timing_hor.counter[2] ));
 sg13g2_nor4_2 _4015_ (.A(\i_vga.vblank ),
    .B(_3242_),
    .C(_3256_),
    .Y(_3258_),
    .D(_3257_));
 sg13g2_or4_2 _4016_ (.A(\i_vga.vblank ),
    .B(_3242_),
    .C(_3256_),
    .D(_3257_),
    .X(_3259_));
 sg13g2_nor2_1 _4017_ (.A(net778),
    .B(net801),
    .Y(_3260_));
 sg13g2_nand2_2 _4018_ (.Y(_3261_),
    .A(net770),
    .B(net794));
 sg13g2_or4_2 _4019_ (.A(\i_vga.timing_ver.counter[0] ),
    .B(_3148_),
    .C(_3248_),
    .D(_3249_),
    .X(_3262_));
 sg13g2_nor4_2 _4020_ (.A(\i_vga.vblank ),
    .B(_3242_),
    .C(_3256_),
    .Y(_3263_),
    .D(_3257_));
 sg13g2_or4_1 _4021_ (.A(\i_vga.vblank ),
    .B(_3242_),
    .C(_3256_),
    .D(_3257_),
    .X(_3264_));
 sg13g2_and2_1 _4022_ (.A(_3262_),
    .B(net791),
    .X(_3265_));
 sg13g2_nand2_2 _4023_ (.Y(_3266_),
    .A(_3262_),
    .B(net791));
 sg13g2_nand2_2 _4024_ (.Y(_3267_),
    .A(net949),
    .B(net765));
 sg13g2_nand2_2 _4025_ (.Y(_3268_),
    .A(net949),
    .B(net838));
 sg13g2_nor2_2 _4026_ (.A(net763),
    .B(_3268_),
    .Y(_3269_));
 sg13g2_or2_1 _4027_ (.X(_3270_),
    .B(_3268_),
    .A(net763));
 sg13g2_nor2b_1 _4028_ (.A(net950),
    .B_N(_0014_),
    .Y(_3271_));
 sg13g2_a21oi_2 _4029_ (.B1(_3271_),
    .Y(_3272_),
    .A2(_0007_),
    .A1(net950));
 sg13g2_mux2_1 _4030_ (.A0(_0014_),
    .A1(_0007_),
    .S(net950),
    .X(_3273_));
 sg13g2_mux2_1 _4031_ (.A0(net929),
    .A1(net902),
    .S(net955),
    .X(_3274_));
 sg13g2_nor2b_2 _4032_ (.A(net865),
    .B_N(net858),
    .Y(_3275_));
 sg13g2_mux2_2 _4033_ (.A0(net934),
    .A1(net906),
    .S(net955),
    .X(_3276_));
 sg13g2_mux2_2 _4034_ (.A0(\i_mandel.i_xy.x[-7] ),
    .A1(net904),
    .S(net955),
    .X(_3277_));
 sg13g2_and2_1 _4035_ (.A(net855),
    .B(net854),
    .X(_3278_));
 sg13g2_nand2_2 _4036_ (.Y(_3279_),
    .A(_3276_),
    .B(net854));
 sg13g2_nand2_1 _4037_ (.Y(_3280_),
    .A(net830),
    .B(net828));
 sg13g2_nor2_1 _4038_ (.A(_0016_),
    .B(net954),
    .Y(_3281_));
 sg13g2_nand2b_1 _4039_ (.Y(_3282_),
    .B(net952),
    .A_N(_0009_));
 sg13g2_nor2b_2 _4040_ (.A(_3281_),
    .B_N(_3282_),
    .Y(_3283_));
 sg13g2_nand2b_1 _4041_ (.Y(_3284_),
    .B(_3282_),
    .A_N(_3281_));
 sg13g2_nor2b_1 _4042_ (.A(net951),
    .B_N(_0015_),
    .Y(_3285_));
 sg13g2_a21oi_2 _4043_ (.B1(_3285_),
    .Y(_3286_),
    .A2(_0008_),
    .A1(net951));
 sg13g2_mux2_1 _4044_ (.A0(_0015_),
    .A1(_0008_),
    .S(net951),
    .X(_3287_));
 sg13g2_mux2_2 _4045_ (.A0(net916),
    .A1(net889),
    .S(net956),
    .X(_3288_));
 sg13g2_nor2b_2 _4046_ (.A(net852),
    .B_N(net849),
    .Y(_3289_));
 sg13g2_nand2_2 _4047_ (.Y(_3290_),
    .A(net824),
    .B(net850));
 sg13g2_nand2b_1 _4048_ (.Y(_3291_),
    .B(net950),
    .A_N(\i_mandel.i_xy.y[-3] ));
 sg13g2_mux2_2 _4049_ (.A0(net922),
    .A1(\i_mandel.i_xy.y[-3] ),
    .S(net950),
    .X(_3292_));
 sg13g2_o21ai_1 _4050_ (.B1(_3291_),
    .Y(_3293_),
    .A1(net950),
    .A2(net922));
 sg13g2_nor2b_2 _4051_ (.A(net864),
    .B_N(_3292_),
    .Y(_3294_));
 sg13g2_nand2b_2 _4052_ (.Y(_3295_),
    .B(net848),
    .A_N(net864));
 sg13g2_nand2b_1 _4053_ (.Y(_3296_),
    .B(net955),
    .A_N(\i_mandel.i_xy.y[-4] ));
 sg13g2_mux2_2 _4054_ (.A0(net925),
    .A1(\i_mandel.i_xy.y[-4] ),
    .S(net950),
    .X(_3297_));
 sg13g2_o21ai_1 _4055_ (.B1(_3296_),
    .Y(_3298_),
    .A1(net956),
    .A2(net925));
 sg13g2_nand2_1 _4056_ (.Y(_3299_),
    .A(net860),
    .B(net846));
 sg13g2_mux2_2 _4057_ (.A0(\i_mandel.i_xy.x[-5] ),
    .A1(net899),
    .S(net955),
    .X(_3300_));
 sg13g2_and2_2 _4058_ (.A(net846),
    .B(net843),
    .X(_3301_));
 sg13g2_nand2_2 _4059_ (.Y(_3302_),
    .A(net846),
    .B(net843));
 sg13g2_and3_2 _4060_ (.X(_3303_),
    .A(net860),
    .B(_3297_),
    .C(net843));
 sg13g2_nand3_1 _4061_ (.B(_3297_),
    .C(net843),
    .A(net857),
    .Y(_3304_));
 sg13g2_nand2_2 _4062_ (.Y(_3305_),
    .A(_3294_),
    .B(_3303_));
 sg13g2_nand3_1 _4063_ (.B(_3294_),
    .C(_3303_),
    .A(_3289_),
    .Y(_3306_));
 sg13g2_nor3_1 _4064_ (.A(net852),
    .B(_3295_),
    .C(_3304_),
    .Y(_3307_));
 sg13g2_nand3_1 _4065_ (.B(_3294_),
    .C(_3303_),
    .A(net824),
    .Y(_3308_));
 sg13g2_xnor2_1 _4066_ (.Y(_3309_),
    .A(_3288_),
    .B(_3308_));
 sg13g2_xnor2_1 _4067_ (.Y(_3310_),
    .A(_3288_),
    .B(_3307_));
 sg13g2_nand2_1 _4068_ (.Y(_3311_),
    .A(net826),
    .B(_3309_));
 sg13g2_nor2_1 _4069_ (.A(net954),
    .B(_0017_),
    .Y(_3312_));
 sg13g2_nand2b_1 _4070_ (.Y(_3313_),
    .B(net954),
    .A_N(_0010_));
 sg13g2_nor2b_2 _4071_ (.A(_3312_),
    .B_N(_3313_),
    .Y(_3314_));
 sg13g2_nand2b_2 _4072_ (.Y(_3315_),
    .B(_3313_),
    .A_N(_3312_));
 sg13g2_o21ai_1 _4073_ (.B1(net852),
    .Y(_3316_),
    .A1(_3295_),
    .A2(_3304_));
 sg13g2_and2_1 _4074_ (.A(_3308_),
    .B(_3316_),
    .X(_3317_));
 sg13g2_nand2_2 _4075_ (.Y(_3318_),
    .A(_3308_),
    .B(_3316_));
 sg13g2_nand3_1 _4076_ (.B(_3315_),
    .C(_3316_),
    .A(_3308_),
    .Y(_3319_));
 sg13g2_nor3_2 _4077_ (.A(_3283_),
    .B(_3310_),
    .C(_3319_),
    .Y(_3320_));
 sg13g2_nor2_1 _4078_ (.A(net950),
    .B(\i_mandel.i_xy.x[0] ),
    .Y(_3321_));
 sg13g2_nand2b_1 _4079_ (.Y(_3322_),
    .B(net951),
    .A_N(\i_mandel.i_xy.y[0] ));
 sg13g2_nor2b_1 _4080_ (.A(_3321_),
    .B_N(_3322_),
    .Y(_3323_));
 sg13g2_nand2b_2 _4081_ (.Y(_3324_),
    .B(_3322_),
    .A_N(_3321_));
 sg13g2_nand2_2 _4082_ (.Y(_3325_),
    .A(net824),
    .B(net820));
 sg13g2_inv_1 _4083_ (.Y(_3326_),
    .A(_3325_));
 sg13g2_nand2_1 _4084_ (.Y(_3327_),
    .A(_3289_),
    .B(net820));
 sg13g2_and2_1 _4085_ (.A(net850),
    .B(net821),
    .X(_3328_));
 sg13g2_nand2_2 _4086_ (.Y(_3329_),
    .A(net850),
    .B(net821));
 sg13g2_nor2_1 _4087_ (.A(_3308_),
    .B(_3329_),
    .Y(_3330_));
 sg13g2_a22oi_1 _4088_ (.Y(_3331_),
    .B1(_3328_),
    .B2(_3307_),
    .A2(_3324_),
    .A1(_3306_));
 sg13g2_nand2_1 _4089_ (.Y(_3332_),
    .A(net826),
    .B(net790));
 sg13g2_and2_1 _4090_ (.A(_3315_),
    .B(net790),
    .X(_3333_));
 sg13g2_nand2b_1 _4091_ (.Y(_3334_),
    .B(_3333_),
    .A_N(_3311_));
 sg13g2_xor2_1 _4092_ (.B(_3333_),
    .A(_3311_),
    .X(_3335_));
 sg13g2_nor3_1 _4093_ (.A(_3311_),
    .B(_3319_),
    .C(_3333_),
    .Y(_3336_));
 sg13g2_nor2_1 _4094_ (.A(net954),
    .B(_0018_),
    .Y(_3337_));
 sg13g2_nand2b_1 _4095_ (.Y(_3338_),
    .B(net952),
    .A_N(_0011_));
 sg13g2_nor2b_2 _4096_ (.A(_3337_),
    .B_N(_3338_),
    .Y(_3339_));
 sg13g2_nand2b_2 _4097_ (.Y(_3340_),
    .B(_3338_),
    .A_N(_3337_));
 sg13g2_nor2_1 _4098_ (.A(net956),
    .B(net913),
    .Y(_3341_));
 sg13g2_a21oi_2 _4099_ (.B1(_3341_),
    .Y(_3342_),
    .A2(_3132_),
    .A1(net956));
 sg13g2_and2_1 _4100_ (.A(net821),
    .B(net817),
    .X(_3343_));
 sg13g2_nand2_2 _4101_ (.Y(_3344_),
    .A(net820),
    .B(net817));
 sg13g2_xnor2_1 _4102_ (.Y(_3345_),
    .A(_3330_),
    .B(net819));
 sg13g2_nor2_1 _4103_ (.A(_3339_),
    .B(net787),
    .Y(_3346_));
 sg13g2_xnor2_1 _4104_ (.Y(_3347_),
    .A(_3320_),
    .B(_3335_));
 sg13g2_a21oi_1 _4105_ (.A1(_3346_),
    .A2(_3347_),
    .Y(_3348_),
    .B1(_3336_));
 sg13g2_nand2_1 _4106_ (.Y(_3349_),
    .A(net824),
    .B(net819));
 sg13g2_nand2_2 _4107_ (.Y(_3350_),
    .A(net857),
    .B(net848));
 sg13g2_nand2_1 _4108_ (.Y(_3351_),
    .A(net847),
    .B(net844));
 sg13g2_nor4_2 _4109_ (.A(_3290_),
    .B(_3302_),
    .C(_3344_),
    .Y(_3352_),
    .D(_3350_));
 sg13g2_nor2_2 _4110_ (.A(net864),
    .B(_3352_),
    .Y(_3353_));
 sg13g2_nand2b_2 _4111_ (.Y(_3354_),
    .B(net830),
    .A_N(_3352_));
 sg13g2_nor2_2 _4112_ (.A(_3339_),
    .B(net786),
    .Y(_3355_));
 sg13g2_inv_1 _4113_ (.Y(_3356_),
    .A(_3355_));
 sg13g2_nor2_1 _4114_ (.A(_3314_),
    .B(net787),
    .Y(_3357_));
 sg13g2_a21oi_1 _4115_ (.A1(_3309_),
    .A2(_3315_),
    .Y(_3358_),
    .B1(_3332_));
 sg13g2_xor2_1 _4116_ (.B(_3358_),
    .A(_3357_),
    .X(_3359_));
 sg13g2_nand2_1 _4117_ (.Y(_3360_),
    .A(_3355_),
    .B(_3359_));
 sg13g2_xnor2_1 _4118_ (.Y(_3361_),
    .A(_3355_),
    .B(_3359_));
 sg13g2_nor2_1 _4119_ (.A(_3348_),
    .B(_3361_),
    .Y(_3362_));
 sg13g2_nor2_1 _4120_ (.A(net953),
    .B(_0019_),
    .Y(_3363_));
 sg13g2_nand2b_1 _4121_ (.Y(_3364_),
    .B(net953),
    .A_N(_0012_));
 sg13g2_nor2b_2 _4122_ (.A(_3363_),
    .B_N(_3364_),
    .Y(_3365_));
 sg13g2_nand2b_2 _4123_ (.Y(_3366_),
    .B(_3364_),
    .A_N(_3363_));
 sg13g2_nor2_2 _4124_ (.A(net786),
    .B(_3365_),
    .Y(_3367_));
 sg13g2_nand2_2 _4125_ (.Y(_3368_),
    .A(_3353_),
    .B(_3366_));
 sg13g2_xor2_1 _4126_ (.B(_3361_),
    .A(_3348_),
    .X(_3369_));
 sg13g2_a21oi_1 _4127_ (.A1(_3367_),
    .A2(_3369_),
    .Y(_3370_),
    .B1(_3362_));
 sg13g2_o21ai_1 _4128_ (.B1(_3360_),
    .Y(_3371_),
    .A1(_3334_),
    .A2(_3357_));
 sg13g2_nor2_1 _4129_ (.A(_3314_),
    .B(net786),
    .Y(_3372_));
 sg13g2_nor3_1 _4130_ (.A(_3283_),
    .B(_3333_),
    .C(net787),
    .Y(_3373_));
 sg13g2_xnor2_1 _4131_ (.Y(_3374_),
    .A(_3372_),
    .B(_3373_));
 sg13g2_xnor2_1 _4132_ (.Y(_3375_),
    .A(_3355_),
    .B(_3374_));
 sg13g2_and2_1 _4133_ (.A(_3371_),
    .B(_3375_),
    .X(_3376_));
 sg13g2_xor2_1 _4134_ (.B(_3375_),
    .A(_3371_),
    .X(_3377_));
 sg13g2_xnor2_1 _4135_ (.Y(_3378_),
    .A(_3367_),
    .B(_3377_));
 sg13g2_or2_1 _4136_ (.X(_3379_),
    .B(_3378_),
    .A(_3370_));
 sg13g2_xnor2_1 _4137_ (.Y(_3380_),
    .A(_3370_),
    .B(_3378_));
 sg13g2_a21o_2 _4138_ (.A2(net823),
    .A1(_3275_),
    .B1(net848),
    .X(_3381_));
 sg13g2_and2_2 _4139_ (.A(_3305_),
    .B(_3381_),
    .X(_3382_));
 sg13g2_nand2_1 _4140_ (.Y(_3383_),
    .A(_3305_),
    .B(_3381_));
 sg13g2_nand3_1 _4141_ (.B(_3315_),
    .C(_3381_),
    .A(_3305_),
    .Y(_3384_));
 sg13g2_and4_1 _4142_ (.A(net826),
    .B(_3308_),
    .C(_3315_),
    .D(_3316_),
    .X(_3385_));
 sg13g2_nand2_1 _4143_ (.Y(_3386_),
    .A(_3382_),
    .B(_3385_));
 sg13g2_a22oi_1 _4144_ (.Y(_3387_),
    .B1(_3317_),
    .B2(net826),
    .A2(_3315_),
    .A1(_3309_));
 sg13g2_or3_1 _4145_ (.A(_3320_),
    .B(_3386_),
    .C(_3387_),
    .X(_3388_));
 sg13g2_and2_1 _4146_ (.A(net790),
    .B(_3340_),
    .X(_3389_));
 sg13g2_o21ai_1 _4147_ (.B1(_3386_),
    .Y(_3390_),
    .A1(_3320_),
    .A2(_3387_));
 sg13g2_nand3_1 _4148_ (.B(_3389_),
    .C(_3390_),
    .A(_3388_),
    .Y(_3391_));
 sg13g2_nand2_1 _4149_ (.Y(_3392_),
    .A(_3388_),
    .B(_3391_));
 sg13g2_xnor2_1 _4150_ (.Y(_3393_),
    .A(_3346_),
    .B(_3347_));
 sg13g2_nor2b_1 _4151_ (.A(_3393_),
    .B_N(_3392_),
    .Y(_3394_));
 sg13g2_xor2_1 _4152_ (.B(_3393_),
    .A(_3392_),
    .X(_3395_));
 sg13g2_nor2_1 _4153_ (.A(_3368_),
    .B(_3395_),
    .Y(_3396_));
 sg13g2_xnor2_1 _4154_ (.Y(_3397_),
    .A(_3368_),
    .B(_3369_));
 sg13g2_o21ai_1 _4155_ (.B1(_3397_),
    .Y(_3398_),
    .A1(_3394_),
    .A2(_3396_));
 sg13g2_or3_1 _4156_ (.A(_3394_),
    .B(_3396_),
    .C(_3397_),
    .X(_3399_));
 sg13g2_xnor2_1 _4157_ (.Y(_3400_),
    .A(_3368_),
    .B(_3395_));
 sg13g2_nand3_1 _4158_ (.B(_3305_),
    .C(_3381_),
    .A(net826),
    .Y(_3401_));
 sg13g2_nand3b_1 _4159_ (.B(net859),
    .C(net844),
    .Y(_3402_),
    .A_N(net865));
 sg13g2_a22oi_1 _4160_ (.Y(_3403_),
    .B1(_3402_),
    .B2(_3298_),
    .A2(net823),
    .A1(_3275_));
 sg13g2_a221oi_1 _4161_ (.B2(_3298_),
    .C1(_3314_),
    .B1(_3402_),
    .A1(_3275_),
    .Y(_3404_),
    .A2(_3301_));
 sg13g2_and4_1 _4162_ (.A(net827),
    .B(_3305_),
    .C(_3381_),
    .D(_3404_),
    .X(_3405_));
 sg13g2_a22oi_1 _4163_ (.Y(_3406_),
    .B1(_3401_),
    .B2(_3319_),
    .A2(_3385_),
    .A1(_3382_));
 sg13g2_and2_1 _4164_ (.A(_3405_),
    .B(_3406_),
    .X(_3407_));
 sg13g2_nor2_1 _4165_ (.A(_3310_),
    .B(_3339_),
    .Y(_3408_));
 sg13g2_xor2_1 _4166_ (.B(_3406_),
    .A(_3405_),
    .X(_3409_));
 sg13g2_a21o_1 _4167_ (.A2(_3409_),
    .A1(_3408_),
    .B1(_3407_),
    .X(_3410_));
 sg13g2_a21o_1 _4168_ (.A2(_3390_),
    .A1(_3388_),
    .B1(_3389_),
    .X(_3411_));
 sg13g2_nand3_1 _4169_ (.B(_3410_),
    .C(_3411_),
    .A(_3391_),
    .Y(_3412_));
 sg13g2_nor2_1 _4170_ (.A(net787),
    .B(_3365_),
    .Y(_3413_));
 sg13g2_a21o_1 _4171_ (.A2(_3411_),
    .A1(_3391_),
    .B1(_3410_),
    .X(_3414_));
 sg13g2_nand3_1 _4172_ (.B(_3413_),
    .C(_3414_),
    .A(_3412_),
    .Y(_3415_));
 sg13g2_and2_1 _4173_ (.A(_3412_),
    .B(_3415_),
    .X(_3416_));
 sg13g2_nor2_1 _4174_ (.A(_3400_),
    .B(_3416_),
    .Y(_3417_));
 sg13g2_xnor2_1 _4175_ (.Y(_3418_),
    .A(_3400_),
    .B(_3416_));
 sg13g2_nand2_1 _4176_ (.Y(_3419_),
    .A(net827),
    .B(_3403_));
 sg13g2_xor2_1 _4177_ (.B(net844),
    .A(_3275_),
    .X(_3420_));
 sg13g2_xnor2_1 _4178_ (.Y(_3421_),
    .A(_3275_),
    .B(net844));
 sg13g2_nor2_1 _4179_ (.A(_3314_),
    .B(_3421_),
    .Y(_3422_));
 sg13g2_and3_1 _4180_ (.X(_3423_),
    .A(net827),
    .B(_3404_),
    .C(net809));
 sg13g2_a21oi_1 _4181_ (.A1(_3384_),
    .A2(_3419_),
    .Y(_3424_),
    .B1(_3405_));
 sg13g2_nand2_1 _4182_ (.Y(_3425_),
    .A(_3423_),
    .B(_3424_));
 sg13g2_nand2_1 _4183_ (.Y(_3426_),
    .A(_3317_),
    .B(_3340_));
 sg13g2_xnor2_1 _4184_ (.Y(_3427_),
    .A(_3423_),
    .B(_3424_));
 sg13g2_o21ai_1 _4185_ (.B1(_3425_),
    .Y(_3428_),
    .A1(_3426_),
    .A2(_3427_));
 sg13g2_xnor2_1 _4186_ (.Y(_3429_),
    .A(_3408_),
    .B(_3409_));
 sg13g2_nand2b_1 _4187_ (.Y(_3430_),
    .B(_3428_),
    .A_N(_3429_));
 sg13g2_nand2_1 _4188_ (.Y(_3431_),
    .A(net790),
    .B(_3366_));
 sg13g2_xor2_1 _4189_ (.B(_3429_),
    .A(_3428_),
    .X(_3432_));
 sg13g2_or2_1 _4190_ (.X(_3433_),
    .B(_3432_),
    .A(_3431_));
 sg13g2_and2_1 _4191_ (.A(_3430_),
    .B(_3433_),
    .X(_3434_));
 sg13g2_o21ai_1 _4192_ (.B1(_3430_),
    .Y(_3435_),
    .A1(_3431_),
    .A2(_3432_));
 sg13g2_a21o_1 _4193_ (.A2(_3414_),
    .A1(_3412_),
    .B1(_3413_),
    .X(_3436_));
 sg13g2_nand2_1 _4194_ (.Y(_3437_),
    .A(_3415_),
    .B(_3436_));
 sg13g2_nand2_1 _4195_ (.Y(_3438_),
    .A(_3340_),
    .B(_3403_));
 sg13g2_nor2_1 _4196_ (.A(net863),
    .B(net857),
    .Y(_3439_));
 sg13g2_xor2_1 _4197_ (.B(net859),
    .A(net865),
    .X(_3440_));
 sg13g2_xnor2_1 _4198_ (.Y(_3441_),
    .A(net865),
    .B(net859));
 sg13g2_nor2_1 _4199_ (.A(_3314_),
    .B(_3440_),
    .Y(_3442_));
 sg13g2_nand3_1 _4200_ (.B(net809),
    .C(_3442_),
    .A(net827),
    .Y(_3443_));
 sg13g2_nand2_1 _4201_ (.Y(_3444_),
    .A(net827),
    .B(_3441_));
 sg13g2_o21ai_1 _4202_ (.B1(_3444_),
    .Y(_3445_),
    .A1(_3314_),
    .A2(_3421_));
 sg13g2_and2_1 _4203_ (.A(_3443_),
    .B(_3445_),
    .X(_3446_));
 sg13g2_nand2b_1 _4204_ (.Y(_3447_),
    .B(_3446_),
    .A_N(_3438_));
 sg13g2_nor2_1 _4205_ (.A(_3339_),
    .B(_3383_),
    .Y(_3448_));
 sg13g2_a21oi_1 _4206_ (.A1(net826),
    .A2(net809),
    .Y(_3449_),
    .B1(_3404_));
 sg13g2_or3_1 _4207_ (.A(_3423_),
    .B(_3443_),
    .C(_3449_),
    .X(_3450_));
 sg13g2_inv_1 _4208_ (.Y(_3451_),
    .A(_3450_));
 sg13g2_o21ai_1 _4209_ (.B1(_3443_),
    .Y(_3452_),
    .A1(_3423_),
    .A2(_3449_));
 sg13g2_and3_1 _4210_ (.X(_3453_),
    .A(_3448_),
    .B(_3450_),
    .C(_3452_));
 sg13g2_a21oi_1 _4211_ (.A1(_3450_),
    .A2(_3452_),
    .Y(_3454_),
    .B1(_3448_));
 sg13g2_or3_1 _4212_ (.A(_3447_),
    .B(_3453_),
    .C(_3454_),
    .X(_3455_));
 sg13g2_nor2_1 _4213_ (.A(_3318_),
    .B(_3365_),
    .Y(_3456_));
 sg13g2_o21ai_1 _4214_ (.B1(_3447_),
    .Y(_3457_),
    .A1(_3453_),
    .A2(_3454_));
 sg13g2_nand3_1 _4215_ (.B(_3456_),
    .C(_3457_),
    .A(_3455_),
    .Y(_3458_));
 sg13g2_nand2_1 _4216_ (.Y(_3459_),
    .A(_3455_),
    .B(_3458_));
 sg13g2_nor2_1 _4217_ (.A(_3310_),
    .B(_3365_),
    .Y(_3460_));
 sg13g2_nor2_1 _4218_ (.A(_3451_),
    .B(_3453_),
    .Y(_3461_));
 sg13g2_xnor2_1 _4219_ (.Y(_3462_),
    .A(_3426_),
    .B(_3427_));
 sg13g2_nor2_1 _4220_ (.A(_3461_),
    .B(_3462_),
    .Y(_3463_));
 sg13g2_xor2_1 _4221_ (.B(_3462_),
    .A(_3461_),
    .X(_3464_));
 sg13g2_xor2_1 _4222_ (.B(_3464_),
    .A(_3460_),
    .X(_3465_));
 sg13g2_nor2_1 _4223_ (.A(_3459_),
    .B(_3465_),
    .Y(_3466_));
 sg13g2_a21o_1 _4224_ (.A2(_3457_),
    .A1(_3455_),
    .B1(_3456_),
    .X(_3467_));
 sg13g2_xnor2_1 _4225_ (.Y(_3468_),
    .A(_3438_),
    .B(_3446_));
 sg13g2_nor2_1 _4226_ (.A(_3339_),
    .B(_3440_),
    .Y(_3469_));
 sg13g2_nand2_1 _4227_ (.Y(_3470_),
    .A(_3422_),
    .B(_3469_));
 sg13g2_nand3_1 _4228_ (.B(_3468_),
    .C(_3469_),
    .A(_3422_),
    .Y(_3471_));
 sg13g2_nand2_1 _4229_ (.Y(_3472_),
    .A(_3366_),
    .B(_3382_));
 sg13g2_xor2_1 _4230_ (.B(_3470_),
    .A(_3468_),
    .X(_3473_));
 sg13g2_o21ai_1 _4231_ (.B1(_3471_),
    .Y(_3474_),
    .A1(_3472_),
    .A2(_3473_));
 sg13g2_and3_1 _4232_ (.X(_3475_),
    .A(_3458_),
    .B(_3467_),
    .C(_3474_));
 sg13g2_nand3_1 _4233_ (.B(_3467_),
    .C(_3474_),
    .A(_3458_),
    .Y(_3476_));
 sg13g2_a21oi_1 _4234_ (.A1(_3458_),
    .A2(_3467_),
    .Y(_3477_),
    .B1(_3474_));
 sg13g2_a21o_1 _4235_ (.A2(_3467_),
    .A1(_3458_),
    .B1(_3474_),
    .X(_3478_));
 sg13g2_xnor2_1 _4236_ (.Y(_3479_),
    .A(_3472_),
    .B(_3473_));
 sg13g2_nand2_1 _4237_ (.Y(_3480_),
    .A(_3366_),
    .B(_3403_));
 sg13g2_nor2_1 _4238_ (.A(_3339_),
    .B(_3421_),
    .Y(_3481_));
 sg13g2_o21ai_1 _4239_ (.B1(_3470_),
    .Y(_3482_),
    .A1(_3442_),
    .A2(_3481_));
 sg13g2_nor2_1 _4240_ (.A(_3480_),
    .B(_3482_),
    .Y(_3483_));
 sg13g2_nand3_1 _4241_ (.B(net809),
    .C(_3469_),
    .A(_3366_),
    .Y(_3484_));
 sg13g2_inv_1 _4242_ (.Y(_3485_),
    .A(_3484_));
 sg13g2_xor2_1 _4243_ (.B(_3482_),
    .A(_3480_),
    .X(_3486_));
 sg13g2_a21oi_2 _4244_ (.B1(_3483_),
    .Y(_3487_),
    .A2(_3486_),
    .A1(_3485_));
 sg13g2_nor2_2 _4245_ (.A(_3479_),
    .B(_3487_),
    .Y(_3488_));
 sg13g2_or2_1 _4246_ (.X(_3489_),
    .B(_3487_),
    .A(_3479_));
 sg13g2_nor3_1 _4247_ (.A(_3475_),
    .B(_3477_),
    .C(_3489_),
    .Y(_3490_));
 sg13g2_nand3_1 _4248_ (.B(_3478_),
    .C(_3488_),
    .A(_3476_),
    .Y(_3491_));
 sg13g2_a21oi_1 _4249_ (.A1(_3478_),
    .A2(_3488_),
    .Y(_3492_),
    .B1(_3475_));
 sg13g2_a221oi_1 _4250_ (.B2(_3488_),
    .C1(_3475_),
    .B1(_3478_),
    .A1(_3459_),
    .Y(_3493_),
    .A2(_3465_));
 sg13g2_xor2_1 _4251_ (.B(_3432_),
    .A(_3431_),
    .X(_3494_));
 sg13g2_a21oi_1 _4252_ (.A1(_3460_),
    .A2(_3464_),
    .Y(_3495_),
    .B1(_3463_));
 sg13g2_nand2b_1 _4253_ (.Y(_3496_),
    .B(_3494_),
    .A_N(_3495_));
 sg13g2_xor2_1 _4254_ (.B(_3495_),
    .A(_3494_),
    .X(_3497_));
 sg13g2_or3_2 _4255_ (.A(_3466_),
    .B(_3493_),
    .C(_3497_),
    .X(_3498_));
 sg13g2_nand3_1 _4256_ (.B(_3435_),
    .C(_3436_),
    .A(_3415_),
    .Y(_3499_));
 sg13g2_and2_1 _4257_ (.A(_3496_),
    .B(_3499_),
    .X(_3500_));
 sg13g2_xnor2_1 _4258_ (.Y(_3501_),
    .A(_3434_),
    .B(_3437_));
 sg13g2_a22oi_1 _4259_ (.Y(_3502_),
    .B1(_3498_),
    .B2(_3500_),
    .A2(_3437_),
    .A1(_3434_));
 sg13g2_a221oi_1 _4260_ (.B2(_3500_),
    .C1(_3418_),
    .B1(_3498_),
    .A1(_3434_),
    .Y(_3503_),
    .A2(_3437_));
 sg13g2_nor2_1 _4261_ (.A(_3417_),
    .B(_3503_),
    .Y(_3504_));
 sg13g2_o21ai_1 _4262_ (.B1(_3398_),
    .Y(_3505_),
    .A1(_3400_),
    .A2(_3416_));
 sg13g2_o21ai_1 _4263_ (.B1(_3399_),
    .Y(_3506_),
    .A1(_3503_),
    .A2(_3505_));
 sg13g2_o21ai_1 _4264_ (.B1(_3379_),
    .Y(_3507_),
    .A1(_3380_),
    .A2(_3506_));
 sg13g2_a21o_1 _4265_ (.A2(_3377_),
    .A1(_3367_),
    .B1(_3376_),
    .X(_3508_));
 sg13g2_nand4_1 _4266_ (.B(net790),
    .C(net786),
    .A(net826),
    .Y(_3509_),
    .D(_3357_));
 sg13g2_o21ai_1 _4267_ (.B1(_3509_),
    .Y(_3510_),
    .A1(_3356_),
    .A2(_3374_));
 sg13g2_a21oi_1 _4268_ (.A1(_3283_),
    .A2(_3314_),
    .Y(_3511_),
    .B1(net786));
 sg13g2_nand4_1 _4269_ (.B(_3315_),
    .C(net787),
    .A(net826),
    .Y(_3512_),
    .D(_3353_));
 sg13g2_nand2_1 _4270_ (.Y(_3513_),
    .A(_3511_),
    .B(_3512_));
 sg13g2_nand2_1 _4271_ (.Y(_3514_),
    .A(_3355_),
    .B(_3513_));
 sg13g2_o21ai_1 _4272_ (.B1(_3514_),
    .Y(_3515_),
    .A1(_3340_),
    .A2(_3513_));
 sg13g2_xnor2_1 _4273_ (.Y(_3516_),
    .A(_3510_),
    .B(_3515_));
 sg13g2_nand2_1 _4274_ (.Y(_3517_),
    .A(_3367_),
    .B(_3516_));
 sg13g2_xnor2_1 _4275_ (.Y(_3518_),
    .A(_3367_),
    .B(_3516_));
 sg13g2_xor2_1 _4276_ (.B(_3518_),
    .A(_3508_),
    .X(_3519_));
 sg13g2_nor2_1 _4277_ (.A(_3355_),
    .B(_3511_),
    .Y(_3520_));
 sg13g2_xor2_1 _4278_ (.B(_3520_),
    .A(_3517_),
    .X(_3521_));
 sg13g2_a21o_1 _4279_ (.A2(_3518_),
    .A1(_3508_),
    .B1(_3521_),
    .X(_3522_));
 sg13g2_a21oi_2 _4280_ (.B1(_3522_),
    .Y(_3523_),
    .A2(_3519_),
    .A1(_3507_));
 sg13g2_nand2_2 _4281_ (.Y(_3524_),
    .A(net856),
    .B(net818));
 sg13g2_nand2_1 _4282_ (.Y(_3525_),
    .A(net853),
    .B(net818));
 sg13g2_nor2b_1 _4283_ (.A(_3280_),
    .B_N(net819),
    .Y(_3526_));
 sg13g2_a22oi_1 _4284_ (.Y(_3527_),
    .B1(net853),
    .B2(net818),
    .A2(net856),
    .A1(net830));
 sg13g2_nor2_1 _4285_ (.A(_3526_),
    .B(_3527_),
    .Y(_3528_));
 sg13g2_nor2_1 _4286_ (.A(net856),
    .B(net853),
    .Y(_3529_));
 sg13g2_nor2_1 _4287_ (.A(net863),
    .B(_3529_),
    .Y(_3530_));
 sg13g2_nor3_1 _4288_ (.A(net863),
    .B(net828),
    .C(_3529_),
    .Y(_0173_));
 sg13g2_nor2_1 _4289_ (.A(_3280_),
    .B(_3523_),
    .Y(_0174_));
 sg13g2_inv_1 _4290_ (.Y(_0175_),
    .A(_0174_));
 sg13g2_mux2_1 _4291_ (.A0(_3280_),
    .A1(_3530_),
    .S(_3523_),
    .X(_0176_));
 sg13g2_xnor2_1 _4292_ (.Y(_0177_),
    .A(_3275_),
    .B(_0176_));
 sg13g2_nand2_2 _4293_ (.Y(_0178_),
    .A(net847),
    .B(net816));
 sg13g2_xor2_1 _4294_ (.B(_3325_),
    .A(net850),
    .X(_0179_));
 sg13g2_o21ai_1 _4295_ (.B1(_3327_),
    .Y(_0180_),
    .A1(_0178_),
    .A2(_0179_));
 sg13g2_xnor2_1 _4296_ (.Y(_0181_),
    .A(net845),
    .B(net842));
 sg13g2_nor2_1 _4297_ (.A(net936),
    .B(net955),
    .Y(_0182_));
 sg13g2_nand2b_1 _4298_ (.Y(_0183_),
    .B(net955),
    .A_N(net907));
 sg13g2_nor2b_2 _4299_ (.A(_0182_),
    .B_N(_0183_),
    .Y(_0184_));
 sg13g2_nand2b_2 _4300_ (.Y(_0185_),
    .B(_0183_),
    .A_N(_0182_));
 sg13g2_nor2_2 _4301_ (.A(net862),
    .B(net815),
    .Y(_0186_));
 sg13g2_nor2_1 _4302_ (.A(net862),
    .B(_0185_),
    .Y(_0187_));
 sg13g2_mux2_2 _4303_ (.A0(_0186_),
    .A1(net807),
    .S(_0181_),
    .X(_0188_));
 sg13g2_inv_2 _4304_ (.Y(_0189_),
    .A(_0188_));
 sg13g2_and2_1 _4305_ (.A(_0180_),
    .B(_0188_),
    .X(_0190_));
 sg13g2_xnor2_1 _4306_ (.Y(_0191_),
    .A(_0180_),
    .B(_0189_));
 sg13g2_nor2_1 _4307_ (.A(net861),
    .B(_3302_),
    .Y(_0192_));
 sg13g2_o21ai_1 _4308_ (.B1(net807),
    .Y(_0193_),
    .A1(net845),
    .A2(net842));
 sg13g2_nand2b_2 _4309_ (.Y(_0194_),
    .B(_0193_),
    .A_N(_0192_));
 sg13g2_a21oi_1 _4310_ (.A1(_0191_),
    .A2(_0194_),
    .Y(_0195_),
    .B1(_0190_));
 sg13g2_nor2_1 _4311_ (.A(net739),
    .B(_0195_),
    .Y(_0196_));
 sg13g2_a21oi_2 _4312_ (.B1(_0174_),
    .Y(_0197_),
    .A2(_0176_),
    .A1(_3275_));
 sg13g2_inv_2 _4313_ (.Y(_0198_),
    .A(_0197_));
 sg13g2_xor2_1 _4314_ (.B(_0195_),
    .A(net739),
    .X(_0199_));
 sg13g2_a21oi_1 _4315_ (.A1(_0198_),
    .A2(_0199_),
    .Y(_0200_),
    .B1(_0196_));
 sg13g2_inv_1 _4316_ (.Y(_0201_),
    .A(_0200_));
 sg13g2_nor2_1 _4317_ (.A(net861),
    .B(net845),
    .Y(_0202_));
 sg13g2_nor2b_1 _4318_ (.A(_0178_),
    .B_N(_0202_),
    .Y(_0203_));
 sg13g2_xnor2_1 _4319_ (.Y(_0204_),
    .A(_0178_),
    .B(_0202_));
 sg13g2_xnor2_1 _4320_ (.Y(_0205_),
    .A(_3325_),
    .B(_0204_));
 sg13g2_nand2_1 _4321_ (.Y(_0206_),
    .A(net845),
    .B(net816));
 sg13g2_o21ai_1 _4322_ (.B1(_0206_),
    .Y(_0207_),
    .A1(net861),
    .A2(net842));
 sg13g2_or3_1 _4323_ (.A(net861),
    .B(net842),
    .C(_0206_),
    .X(_0208_));
 sg13g2_nor2_2 _4324_ (.A(_3293_),
    .B(_3324_),
    .Y(_0209_));
 sg13g2_nand2_1 _4325_ (.Y(_0210_),
    .A(_0207_),
    .B(_0209_));
 sg13g2_nand2_1 _4326_ (.Y(_0211_),
    .A(_0208_),
    .B(_0210_));
 sg13g2_nand2_1 _4327_ (.Y(_0212_),
    .A(_0205_),
    .B(_0211_));
 sg13g2_xor2_1 _4328_ (.B(_0179_),
    .A(_0178_),
    .X(_0213_));
 sg13g2_xor2_1 _4329_ (.B(_0211_),
    .A(_0205_),
    .X(_0214_));
 sg13g2_nand2_1 _4330_ (.Y(_0215_),
    .A(_0213_),
    .B(_0214_));
 sg13g2_nand2_1 _4331_ (.Y(_0216_),
    .A(_0212_),
    .B(_0215_));
 sg13g2_xnor2_1 _4332_ (.Y(_0217_),
    .A(_3328_),
    .B(_3349_));
 sg13g2_xnor2_1 _4333_ (.Y(_0218_),
    .A(_3294_),
    .B(_0217_));
 sg13g2_a21oi_1 _4334_ (.A1(_3326_),
    .A2(_0204_),
    .Y(_0219_),
    .B1(_0203_));
 sg13g2_nor3_1 _4335_ (.A(net864),
    .B(net847),
    .C(_3349_),
    .Y(_0220_));
 sg13g2_o21ai_1 _4336_ (.B1(_3349_),
    .Y(_0221_),
    .A1(net864),
    .A2(net847));
 sg13g2_nor2b_1 _4337_ (.A(_0220_),
    .B_N(_0221_),
    .Y(_0222_));
 sg13g2_xnor2_1 _4338_ (.Y(_0223_),
    .A(_3329_),
    .B(_0222_));
 sg13g2_nand2b_1 _4339_ (.Y(_0224_),
    .B(_0223_),
    .A_N(_0219_));
 sg13g2_nor2b_1 _4340_ (.A(_0223_),
    .B_N(_0219_),
    .Y(_0225_));
 sg13g2_xnor2_1 _4341_ (.Y(_0226_),
    .A(net861),
    .B(_0219_));
 sg13g2_a21oi_1 _4342_ (.A1(_0212_),
    .A2(_0215_),
    .Y(_0227_),
    .B1(_0226_));
 sg13g2_xor2_1 _4343_ (.B(_0194_),
    .A(_0191_),
    .X(_0228_));
 sg13g2_xor2_1 _4344_ (.B(_0226_),
    .A(_0216_),
    .X(_0229_));
 sg13g2_inv_1 _4345_ (.Y(_0230_),
    .A(_0229_));
 sg13g2_a21oi_1 _4346_ (.A1(_0228_),
    .A2(_0230_),
    .Y(_0231_),
    .B1(_0227_));
 sg13g2_a22oi_1 _4347_ (.Y(_0232_),
    .B1(_0217_),
    .B2(_3294_),
    .A2(_3343_),
    .A1(_3289_));
 sg13g2_nor2_1 _4348_ (.A(_0189_),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_xnor2_1 _4349_ (.Y(_0234_),
    .A(_0188_),
    .B(_0232_));
 sg13g2_xnor2_1 _4350_ (.Y(_0235_),
    .A(_0194_),
    .B(_0234_));
 sg13g2_o21ai_1 _4351_ (.B1(_0224_),
    .Y(_0236_),
    .A1(_0218_),
    .A2(_0225_));
 sg13g2_nor2_2 _4352_ (.A(net864),
    .B(net852),
    .Y(_0237_));
 sg13g2_nand2_1 _4353_ (.Y(_0238_),
    .A(net849),
    .B(net819));
 sg13g2_nand3_1 _4354_ (.B(net819),
    .C(_0237_),
    .A(net849),
    .Y(_0239_));
 sg13g2_xor2_1 _4355_ (.B(_0238_),
    .A(_0237_),
    .X(_0240_));
 sg13g2_xnor2_1 _4356_ (.Y(_0241_),
    .A(_3295_),
    .B(_0240_));
 sg13g2_a21o_1 _4357_ (.A2(_0222_),
    .A1(_3328_),
    .B1(_0220_),
    .X(_0242_));
 sg13g2_nor3_1 _4358_ (.A(net865),
    .B(net824),
    .C(_0238_),
    .Y(_0243_));
 sg13g2_a22oi_1 _4359_ (.Y(_0244_),
    .B1(net849),
    .B2(net819),
    .A2(net852),
    .A1(_3272_));
 sg13g2_nor2_1 _4360_ (.A(_0243_),
    .B(_0244_),
    .Y(_0245_));
 sg13g2_xnor2_1 _4361_ (.Y(_0246_),
    .A(net820),
    .B(_0245_));
 sg13g2_nand2b_1 _4362_ (.Y(_0247_),
    .B(_0242_),
    .A_N(_0246_));
 sg13g2_xor2_1 _4363_ (.B(_0246_),
    .A(_0242_),
    .X(_0248_));
 sg13g2_xor2_1 _4364_ (.B(_0248_),
    .A(_0241_),
    .X(_0249_));
 sg13g2_nand2_1 _4365_ (.Y(_0250_),
    .A(_0236_),
    .B(_0249_));
 sg13g2_xnor2_1 _4366_ (.Y(_0251_),
    .A(_0236_),
    .B(_0249_));
 sg13g2_xor2_1 _4367_ (.B(_0251_),
    .A(_0235_),
    .X(_0252_));
 sg13g2_nor2b_1 _4368_ (.A(_0231_),
    .B_N(_0252_),
    .Y(_0253_));
 sg13g2_xnor2_1 _4369_ (.Y(_0254_),
    .A(_0197_),
    .B(_0199_));
 sg13g2_xnor2_1 _4370_ (.Y(_0255_),
    .A(_0231_),
    .B(_0252_));
 sg13g2_a21oi_1 _4371_ (.A1(_0254_),
    .A2(_0255_),
    .Y(_0256_),
    .B1(_0253_));
 sg13g2_a21oi_1 _4372_ (.A1(_0194_),
    .A2(_0234_),
    .Y(_0257_),
    .B1(_0233_));
 sg13g2_nor2_1 _4373_ (.A(net739),
    .B(_0257_),
    .Y(_0258_));
 sg13g2_xor2_1 _4374_ (.B(_0257_),
    .A(net739),
    .X(_0259_));
 sg13g2_xnor2_1 _4375_ (.Y(_0260_),
    .A(_0197_),
    .B(_0259_));
 sg13g2_inv_1 _4376_ (.Y(_0261_),
    .A(_0260_));
 sg13g2_o21ai_1 _4377_ (.B1(_0250_),
    .Y(_0262_),
    .A1(_0235_),
    .A2(_0251_));
 sg13g2_o21ai_1 _4378_ (.B1(_0239_),
    .Y(_0263_),
    .A1(_3295_),
    .A2(_0240_));
 sg13g2_and2_1 _4379_ (.A(_0188_),
    .B(_0263_),
    .X(_0264_));
 sg13g2_xnor2_1 _4380_ (.Y(_0265_),
    .A(_0189_),
    .B(_0263_));
 sg13g2_xnor2_1 _4381_ (.Y(_0266_),
    .A(_0194_),
    .B(_0265_));
 sg13g2_o21ai_1 _4382_ (.B1(_0247_),
    .Y(_0267_),
    .A1(_0241_),
    .A2(_0248_));
 sg13g2_o21ai_1 _4383_ (.B1(net830),
    .Y(_0268_),
    .A1(net824),
    .A2(net849));
 sg13g2_a21oi_1 _4384_ (.A1(net849),
    .A2(_0237_),
    .Y(_0269_),
    .B1(_0268_));
 sg13g2_xnor2_1 _4385_ (.Y(_0270_),
    .A(_3294_),
    .B(_0269_));
 sg13g2_inv_1 _4386_ (.Y(_0271_),
    .A(_0270_));
 sg13g2_nor2_1 _4387_ (.A(net862),
    .B(net849),
    .Y(_0272_));
 sg13g2_a21oi_1 _4388_ (.A1(net820),
    .A2(_0245_),
    .Y(_0273_),
    .B1(_0243_));
 sg13g2_nor2b_1 _4389_ (.A(_0273_),
    .B_N(_0272_),
    .Y(_0274_));
 sg13g2_xnor2_1 _4390_ (.Y(_0275_),
    .A(_0272_),
    .B(_0273_));
 sg13g2_xnor2_1 _4391_ (.Y(_0276_),
    .A(_0270_),
    .B(_0275_));
 sg13g2_nand2_1 _4392_ (.Y(_0277_),
    .A(_0267_),
    .B(_0276_));
 sg13g2_xnor2_1 _4393_ (.Y(_0278_),
    .A(_0267_),
    .B(_0276_));
 sg13g2_xor2_1 _4394_ (.B(_0278_),
    .A(_0266_),
    .X(_0279_));
 sg13g2_nand2_1 _4395_ (.Y(_0280_),
    .A(_0262_),
    .B(_0279_));
 sg13g2_xnor2_1 _4396_ (.Y(_0281_),
    .A(_0262_),
    .B(_0279_));
 sg13g2_xor2_1 _4397_ (.B(_0281_),
    .A(_0260_),
    .X(_0282_));
 sg13g2_nor2_1 _4398_ (.A(_0256_),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_xor2_1 _4399_ (.B(_0282_),
    .A(_0256_),
    .X(_0284_));
 sg13g2_xnor2_1 _4400_ (.Y(_0285_),
    .A(_0200_),
    .B(_0284_));
 sg13g2_nand2_1 _4401_ (.Y(_0286_),
    .A(_0207_),
    .B(_0208_));
 sg13g2_nand2_1 _4402_ (.Y(_0287_),
    .A(net842),
    .B(net816));
 sg13g2_nand3_1 _4403_ (.B(net816),
    .C(_3439_),
    .A(net842),
    .Y(_0288_));
 sg13g2_nand2_1 _4404_ (.Y(_0289_),
    .A(net845),
    .B(net820));
 sg13g2_xor2_1 _4405_ (.B(_0287_),
    .A(_3439_),
    .X(_0290_));
 sg13g2_o21ai_1 _4406_ (.B1(_0288_),
    .Y(_0291_),
    .A1(_0289_),
    .A2(_0290_));
 sg13g2_mux2_1 _4407_ (.A0(_0291_),
    .A1(_0209_),
    .S(_0286_),
    .X(_0292_));
 sg13g2_xnor2_1 _4408_ (.Y(_0293_),
    .A(_0213_),
    .B(_0214_));
 sg13g2_nor2b_1 _4409_ (.A(_0293_),
    .B_N(_0292_),
    .Y(_0294_));
 sg13g2_a22oi_1 _4410_ (.Y(_0295_),
    .B1(net816),
    .B2(net845),
    .A2(net842),
    .A1(net830));
 sg13g2_a21oi_1 _4411_ (.A1(net816),
    .A2(_0192_),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_a22oi_1 _4412_ (.Y(_0297_),
    .B1(_0296_),
    .B2(net807),
    .A2(_0192_),
    .A1(net816));
 sg13g2_xnor2_1 _4413_ (.Y(_0298_),
    .A(_3290_),
    .B(_0188_));
 sg13g2_nand2b_1 _4414_ (.Y(_0299_),
    .B(_0298_),
    .A_N(_0297_));
 sg13g2_xnor2_1 _4415_ (.Y(_0300_),
    .A(_0297_),
    .B(_0298_));
 sg13g2_xnor2_1 _4416_ (.Y(_0301_),
    .A(_0292_),
    .B(_0293_));
 sg13g2_a21oi_1 _4417_ (.A1(_0300_),
    .A2(_0301_),
    .Y(_0302_),
    .B1(_0294_));
 sg13g2_xor2_1 _4418_ (.B(_0229_),
    .A(_0228_),
    .X(_0303_));
 sg13g2_nor2_1 _4419_ (.A(_0302_),
    .B(_0303_),
    .Y(_0304_));
 sg13g2_o21ai_1 _4420_ (.B1(_0299_),
    .Y(_0305_),
    .A1(_3290_),
    .A2(_0189_));
 sg13g2_nand2b_1 _4421_ (.Y(_0306_),
    .B(_0305_),
    .A_N(net739));
 sg13g2_xnor2_1 _4422_ (.Y(_0307_),
    .A(net739),
    .B(_0305_));
 sg13g2_nand2_1 _4423_ (.Y(_0308_),
    .A(_0198_),
    .B(_0307_));
 sg13g2_xnor2_1 _4424_ (.Y(_0309_),
    .A(_0197_),
    .B(_0307_));
 sg13g2_xor2_1 _4425_ (.B(_0303_),
    .A(_0302_),
    .X(_0310_));
 sg13g2_a21oi_1 _4426_ (.A1(_0309_),
    .A2(_0310_),
    .Y(_0311_),
    .B1(_0304_));
 sg13g2_xnor2_1 _4427_ (.Y(_0312_),
    .A(_0254_),
    .B(_0255_));
 sg13g2_nor2_1 _4428_ (.A(_0311_),
    .B(_0312_),
    .Y(_0313_));
 sg13g2_nand2_1 _4429_ (.Y(_0314_),
    .A(_0306_),
    .B(_0308_));
 sg13g2_xor2_1 _4430_ (.B(_0312_),
    .A(_0311_),
    .X(_0315_));
 sg13g2_and2_1 _4431_ (.A(_0314_),
    .B(_0315_),
    .X(_0316_));
 sg13g2_o21ai_1 _4432_ (.B1(_0285_),
    .Y(_0317_),
    .A1(_0313_),
    .A2(_0316_));
 sg13g2_a21oi_1 _4433_ (.A1(_0198_),
    .A2(_0259_),
    .Y(_0318_),
    .B1(_0258_));
 sg13g2_o21ai_1 _4434_ (.B1(_0280_),
    .Y(_0319_),
    .A1(_0261_),
    .A2(_0281_));
 sg13g2_a21oi_1 _4435_ (.A1(_0194_),
    .A2(_0265_),
    .Y(_0320_),
    .B1(_0264_));
 sg13g2_nor2_1 _4436_ (.A(net740),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_xor2_1 _4437_ (.B(_0320_),
    .A(net740),
    .X(_0322_));
 sg13g2_xnor2_1 _4438_ (.Y(_0323_),
    .A(_0197_),
    .B(_0322_));
 sg13g2_inv_1 _4439_ (.Y(_0324_),
    .A(_0323_));
 sg13g2_o21ai_1 _4440_ (.B1(_0277_),
    .Y(_0325_),
    .A1(_0266_),
    .A2(_0278_));
 sg13g2_a22oi_1 _4441_ (.Y(_0326_),
    .B1(_0269_),
    .B2(_3294_),
    .A2(_0237_),
    .A1(net849));
 sg13g2_nor2_1 _4442_ (.A(_0189_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_xnor2_1 _4443_ (.Y(_0328_),
    .A(_0188_),
    .B(_0326_));
 sg13g2_xor2_1 _4444_ (.B(_0328_),
    .A(_0194_),
    .X(_0329_));
 sg13g2_a21oi_1 _4445_ (.A1(_0271_),
    .A2(_0275_),
    .Y(_0330_),
    .B1(_0274_));
 sg13g2_o21ai_1 _4446_ (.B1(net817),
    .Y(_0331_),
    .A1(net862),
    .A2(net821));
 sg13g2_o21ai_1 _4447_ (.B1(_0331_),
    .Y(_0332_),
    .A1(net862),
    .A2(net817));
 sg13g2_o21ai_1 _4448_ (.B1(_0332_),
    .Y(_0333_),
    .A1(net830),
    .A2(_3344_));
 sg13g2_nor2_1 _4449_ (.A(_0270_),
    .B(_0333_),
    .Y(_0334_));
 sg13g2_xor2_1 _4450_ (.B(_0333_),
    .A(_0270_),
    .X(_0335_));
 sg13g2_nor2b_1 _4451_ (.A(_0330_),
    .B_N(_0335_),
    .Y(_0336_));
 sg13g2_xnor2_1 _4452_ (.Y(_0337_),
    .A(_0330_),
    .B(_0335_));
 sg13g2_xor2_1 _4453_ (.B(_0337_),
    .A(_0329_),
    .X(_0338_));
 sg13g2_nand2_1 _4454_ (.Y(_0339_),
    .A(_0325_),
    .B(_0338_));
 sg13g2_xnor2_1 _4455_ (.Y(_0340_),
    .A(_0325_),
    .B(_0338_));
 sg13g2_xor2_1 _4456_ (.B(_0340_),
    .A(_0323_),
    .X(_0341_));
 sg13g2_nand2b_1 _4457_ (.Y(_0342_),
    .B(_0319_),
    .A_N(_0341_));
 sg13g2_xor2_1 _4458_ (.B(_0341_),
    .A(_0319_),
    .X(_0343_));
 sg13g2_xor2_1 _4459_ (.B(_0343_),
    .A(_0318_),
    .X(_0344_));
 sg13g2_a21oi_2 _4460_ (.B1(_0283_),
    .Y(_0345_),
    .A2(_0284_),
    .A1(_0201_));
 sg13g2_nor2b_1 _4461_ (.A(_0345_),
    .B_N(_0344_),
    .Y(_0346_));
 sg13g2_xor2_1 _4462_ (.B(_0345_),
    .A(_0344_),
    .X(_0347_));
 sg13g2_nor2_1 _4463_ (.A(_0317_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_or3_1 _4464_ (.A(_0285_),
    .B(_0313_),
    .C(_0316_),
    .X(_0349_));
 sg13g2_and2_1 _4465_ (.A(_0317_),
    .B(_0349_),
    .X(_0350_));
 sg13g2_xnor2_1 _4466_ (.Y(_0351_),
    .A(_0314_),
    .B(_0315_));
 sg13g2_nor2_1 _4467_ (.A(net863),
    .B(net853),
    .Y(_0352_));
 sg13g2_nand2_1 _4468_ (.Y(_0353_),
    .A(net857),
    .B(net818));
 sg13g2_nand3_1 _4469_ (.B(net819),
    .C(_0352_),
    .A(net857),
    .Y(_0354_));
 sg13g2_nand2_2 _4470_ (.Y(_0355_),
    .A(net842),
    .B(net820));
 sg13g2_xor2_1 _4471_ (.B(_0353_),
    .A(_0352_),
    .X(_0356_));
 sg13g2_o21ai_1 _4472_ (.B1(_0354_),
    .Y(_0357_),
    .A1(_0355_),
    .A2(_0356_));
 sg13g2_xor2_1 _4473_ (.B(_0290_),
    .A(_0289_),
    .X(_0358_));
 sg13g2_nand2_1 _4474_ (.Y(_0359_),
    .A(_0357_),
    .B(_0358_));
 sg13g2_xnor2_1 _4475_ (.Y(_0360_),
    .A(_0357_),
    .B(_0358_));
 sg13g2_o21ai_1 _4476_ (.B1(_0359_),
    .Y(_0361_),
    .A1(net852),
    .A2(_0360_));
 sg13g2_xor2_1 _4477_ (.B(_0291_),
    .A(_0286_),
    .X(_0362_));
 sg13g2_inv_1 _4478_ (.Y(_0363_),
    .A(_0362_));
 sg13g2_a22oi_1 _4479_ (.Y(_0364_),
    .B1(_0287_),
    .B2(_0289_),
    .A2(_3343_),
    .A1(net823));
 sg13g2_nand2_1 _4480_ (.Y(_0365_),
    .A(net807),
    .B(_0364_));
 sg13g2_o21ai_1 _4481_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_3302_),
    .A2(_3344_));
 sg13g2_and2_1 _4482_ (.A(net850),
    .B(net847),
    .X(_0367_));
 sg13g2_xor2_1 _4483_ (.B(_0296_),
    .A(net807),
    .X(_0368_));
 sg13g2_xor2_1 _4484_ (.B(_0368_),
    .A(_0367_),
    .X(_0369_));
 sg13g2_and2_1 _4485_ (.A(_0366_),
    .B(_0369_),
    .X(_0370_));
 sg13g2_xnor2_1 _4486_ (.Y(_0371_),
    .A(_0366_),
    .B(_0369_));
 sg13g2_xnor2_1 _4487_ (.Y(_0372_),
    .A(_0361_),
    .B(_0362_));
 sg13g2_nor2b_1 _4488_ (.A(_0371_),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_a21oi_1 _4489_ (.A1(_0361_),
    .A2(_0363_),
    .Y(_0374_),
    .B1(_0373_));
 sg13g2_xnor2_1 _4490_ (.Y(_0375_),
    .A(_0300_),
    .B(_0301_));
 sg13g2_nor2_1 _4491_ (.A(_0374_),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_a21oi_1 _4492_ (.A1(_0367_),
    .A2(_0368_),
    .Y(_0377_),
    .B1(_0370_));
 sg13g2_nor2_1 _4493_ (.A(_0177_),
    .B(_0377_),
    .Y(_0378_));
 sg13g2_xor2_1 _4494_ (.B(_0377_),
    .A(net740),
    .X(_0379_));
 sg13g2_xnor2_1 _4495_ (.Y(_0380_),
    .A(_0197_),
    .B(_0379_));
 sg13g2_xor2_1 _4496_ (.B(_0375_),
    .A(_0374_),
    .X(_0381_));
 sg13g2_a21oi_1 _4497_ (.A1(_0380_),
    .A2(_0381_),
    .Y(_0382_),
    .B1(_0376_));
 sg13g2_xnor2_1 _4498_ (.Y(_0383_),
    .A(_0309_),
    .B(_0310_));
 sg13g2_nor2_1 _4499_ (.A(_0382_),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_a21oi_1 _4500_ (.A1(_0198_),
    .A2(_0379_),
    .Y(_0385_),
    .B1(_0378_));
 sg13g2_inv_1 _4501_ (.Y(_0386_),
    .A(_0385_));
 sg13g2_xor2_1 _4502_ (.B(_0383_),
    .A(_0382_),
    .X(_0387_));
 sg13g2_a21oi_1 _4503_ (.A1(_0386_),
    .A2(_0387_),
    .Y(_0388_),
    .B1(_0384_));
 sg13g2_nor2_1 _4504_ (.A(_0351_),
    .B(_0388_),
    .Y(_0389_));
 sg13g2_nand2_1 _4505_ (.Y(_0390_),
    .A(_0350_),
    .B(_0389_));
 sg13g2_xnor2_1 _4506_ (.Y(_0391_),
    .A(_0351_),
    .B(_0388_));
 sg13g2_xnor2_1 _4507_ (.Y(_0392_),
    .A(_0385_),
    .B(_0387_));
 sg13g2_nor2_1 _4508_ (.A(net862),
    .B(net856),
    .Y(_0393_));
 sg13g2_nand3_1 _4509_ (.B(net818),
    .C(_0393_),
    .A(net853),
    .Y(_0394_));
 sg13g2_nand2_2 _4510_ (.Y(_0395_),
    .A(net857),
    .B(net822));
 sg13g2_xnor2_1 _4511_ (.Y(_0396_),
    .A(_3525_),
    .B(_0393_));
 sg13g2_nand2b_1 _4512_ (.Y(_0397_),
    .B(_0396_),
    .A_N(_0395_));
 sg13g2_nand2_1 _4513_ (.Y(_0398_),
    .A(_0394_),
    .B(_0397_));
 sg13g2_xor2_1 _4514_ (.B(_0356_),
    .A(_0355_),
    .X(_0399_));
 sg13g2_nand2_1 _4515_ (.Y(_0400_),
    .A(_0398_),
    .B(_0399_));
 sg13g2_nand2_1 _4516_ (.Y(_0401_),
    .A(net850),
    .B(net845));
 sg13g2_xnor2_1 _4517_ (.Y(_0402_),
    .A(_0398_),
    .B(_0399_));
 sg13g2_o21ai_1 _4518_ (.B1(_0400_),
    .Y(_0403_),
    .A1(_0401_),
    .A2(_0402_));
 sg13g2_xnor2_1 _4519_ (.Y(_0404_),
    .A(net824),
    .B(_0360_));
 sg13g2_nand2_1 _4520_ (.Y(_0405_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_xor2_1 _4521_ (.B(_0401_),
    .A(_0355_),
    .X(_0406_));
 sg13g2_nand2_1 _4522_ (.Y(_0407_),
    .A(net807),
    .B(_0406_));
 sg13g2_o21ai_1 _4523_ (.B1(_0407_),
    .Y(_0408_),
    .A1(_3302_),
    .A2(_3329_));
 sg13g2_nor2_2 _4524_ (.A(net852),
    .B(_3293_),
    .Y(_0409_));
 sg13g2_xor2_1 _4525_ (.B(_0364_),
    .A(net807),
    .X(_0410_));
 sg13g2_xnor2_1 _4526_ (.Y(_0411_),
    .A(_0409_),
    .B(_0410_));
 sg13g2_nor2b_1 _4527_ (.A(_0411_),
    .B_N(_0408_),
    .Y(_0412_));
 sg13g2_xor2_1 _4528_ (.B(_0411_),
    .A(_0408_),
    .X(_0413_));
 sg13g2_xnor2_1 _4529_ (.Y(_0414_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_o21ai_1 _4530_ (.B1(_0405_),
    .Y(_0415_),
    .A1(_0413_),
    .A2(_0414_));
 sg13g2_xnor2_1 _4531_ (.Y(_0416_),
    .A(_0371_),
    .B(_0372_));
 sg13g2_nand2_1 _4532_ (.Y(_0417_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_a21o_1 _4533_ (.A2(_0410_),
    .A1(_0409_),
    .B1(_0412_),
    .X(_0418_));
 sg13g2_nor2b_1 _4534_ (.A(net740),
    .B_N(_0418_),
    .Y(_0419_));
 sg13g2_xnor2_1 _4535_ (.Y(_0420_),
    .A(net740),
    .B(_0418_));
 sg13g2_xnor2_1 _4536_ (.Y(_0421_),
    .A(_0197_),
    .B(_0420_));
 sg13g2_inv_1 _4537_ (.Y(_0422_),
    .A(_0421_));
 sg13g2_xnor2_1 _4538_ (.Y(_0423_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_o21ai_1 _4539_ (.B1(_0417_),
    .Y(_0424_),
    .A1(_0422_),
    .A2(_0423_));
 sg13g2_xnor2_1 _4540_ (.Y(_0425_),
    .A(_0380_),
    .B(_0381_));
 sg13g2_nor2b_1 _4541_ (.A(_0425_),
    .B_N(_0424_),
    .Y(_0426_));
 sg13g2_a21o_1 _4542_ (.A2(_0420_),
    .A1(_0198_),
    .B1(_0419_),
    .X(_0427_));
 sg13g2_xor2_1 _4543_ (.B(_0425_),
    .A(_0424_),
    .X(_0428_));
 sg13g2_nor2b_1 _4544_ (.A(_0428_),
    .B_N(_0427_),
    .Y(_0429_));
 sg13g2_nor2_1 _4545_ (.A(_0426_),
    .B(_0429_),
    .Y(_0430_));
 sg13g2_nor2b_1 _4546_ (.A(_0430_),
    .B_N(_0392_),
    .Y(_0431_));
 sg13g2_nor2b_1 _4547_ (.A(_0391_),
    .B_N(_0431_),
    .Y(_0432_));
 sg13g2_nand2_2 _4548_ (.Y(_0433_),
    .A(net822),
    .B(net815));
 sg13g2_and2_2 _4549_ (.A(net855),
    .B(_0184_),
    .X(_0434_));
 sg13g2_nand2_1 _4550_ (.Y(_0435_),
    .A(_3276_),
    .B(_0184_));
 sg13g2_nor2_2 _4551_ (.A(_3287_),
    .B(_0185_),
    .Y(_0436_));
 sg13g2_nand2_1 _4552_ (.Y(_0437_),
    .A(net854),
    .B(net848));
 sg13g2_inv_1 _4553_ (.Y(_0438_),
    .A(_0437_));
 sg13g2_nand2_1 _4554_ (.Y(_0439_),
    .A(net856),
    .B(net825));
 sg13g2_nand2_2 _4555_ (.Y(_0440_),
    .A(net851),
    .B(net815));
 sg13g2_a22oi_1 _4556_ (.Y(_0441_),
    .B1(_0439_),
    .B2(_0440_),
    .A2(_0434_),
    .A1(_3289_));
 sg13g2_a22oi_1 _4557_ (.Y(_0442_),
    .B1(_0438_),
    .B2(_0441_),
    .A2(_0434_),
    .A1(_3289_));
 sg13g2_nor2_1 _4558_ (.A(_0433_),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_xnor2_1 _4559_ (.Y(_0444_),
    .A(_0433_),
    .B(_0442_));
 sg13g2_inv_1 _4560_ (.Y(_0445_),
    .A(_0444_));
 sg13g2_a21oi_1 _4561_ (.A1(net860),
    .A2(net846),
    .Y(_0446_),
    .B1(net843));
 sg13g2_nor3_1 _4562_ (.A(_3303_),
    .B(_0440_),
    .C(_0446_),
    .Y(_0447_));
 sg13g2_o21ai_1 _4563_ (.B1(_3304_),
    .Y(_0448_),
    .A1(_0440_),
    .A2(_0446_));
 sg13g2_xor2_1 _4564_ (.B(_0448_),
    .A(_0444_),
    .X(_0449_));
 sg13g2_nand2_1 _4565_ (.Y(_0450_),
    .A(net828),
    .B(_3289_));
 sg13g2_a22oi_1 _4566_ (.Y(_0451_),
    .B1(net851),
    .B2(net856),
    .A2(net824),
    .A1(net853));
 sg13g2_a21oi_2 _4567_ (.B1(_0451_),
    .Y(_0452_),
    .A2(_3289_),
    .A1(net828));
 sg13g2_xnor2_1 _4568_ (.Y(_0453_),
    .A(_3350_),
    .B(_0452_));
 sg13g2_nand2b_1 _4569_ (.Y(_0454_),
    .B(_0453_),
    .A_N(_0433_));
 sg13g2_xnor2_1 _4570_ (.Y(_0455_),
    .A(_0433_),
    .B(_0453_));
 sg13g2_nor2b_1 _4571_ (.A(_0449_),
    .B_N(_0455_),
    .Y(_0456_));
 sg13g2_nand2_2 _4572_ (.Y(_0457_),
    .A(net858),
    .B(net854));
 sg13g2_nand2_2 _4573_ (.Y(_0458_),
    .A(net857),
    .B(net851));
 sg13g2_nor2_1 _4574_ (.A(_3290_),
    .B(_0457_),
    .Y(_0459_));
 sg13g2_nand2_1 _4575_ (.Y(_0460_),
    .A(net857),
    .B(net825));
 sg13g2_nand2_1 _4576_ (.Y(_0461_),
    .A(net853),
    .B(net851));
 sg13g2_a21oi_1 _4577_ (.A1(_0460_),
    .A2(_0461_),
    .Y(_0462_),
    .B1(_0459_));
 sg13g2_nor2b_1 _4578_ (.A(_3351_),
    .B_N(_0462_),
    .Y(_0463_));
 sg13g2_xnor2_1 _4579_ (.Y(_0464_),
    .A(_3351_),
    .B(_0462_));
 sg13g2_nand2_2 _4580_ (.Y(_0465_),
    .A(net818),
    .B(net815));
 sg13g2_nand2_1 _4581_ (.Y(_0466_),
    .A(net856),
    .B(net822));
 sg13g2_nor2_1 _4582_ (.A(_3524_),
    .B(_0433_),
    .Y(_0467_));
 sg13g2_xor2_1 _4583_ (.B(_0466_),
    .A(_0465_),
    .X(_0468_));
 sg13g2_nand2_1 _4584_ (.Y(_0469_),
    .A(_0464_),
    .B(_0468_));
 sg13g2_xnor2_1 _4585_ (.Y(_0470_),
    .A(_0464_),
    .B(_0468_));
 sg13g2_xnor2_1 _4586_ (.Y(_0471_),
    .A(_0454_),
    .B(_0470_));
 sg13g2_o21ai_1 _4587_ (.B1(_0450_),
    .Y(_0472_),
    .A1(_3350_),
    .A2(_0451_));
 sg13g2_nor2_2 _4588_ (.A(_3293_),
    .B(_3298_),
    .Y(_0473_));
 sg13g2_nand2_1 _4589_ (.Y(_0474_),
    .A(net847),
    .B(net846));
 sg13g2_a22oi_1 _4590_ (.Y(_0475_),
    .B1(_3351_),
    .B2(_3298_),
    .A2(net823),
    .A1(net847));
 sg13g2_nand2b_1 _4591_ (.Y(_0476_),
    .B(_0475_),
    .A_N(_0465_));
 sg13g2_xnor2_1 _4592_ (.Y(_0477_),
    .A(_0465_),
    .B(_0475_));
 sg13g2_nand2_1 _4593_ (.Y(_0478_),
    .A(_0472_),
    .B(_0477_));
 sg13g2_xnor2_1 _4594_ (.Y(_0479_),
    .A(_0472_),
    .B(_0477_));
 sg13g2_xnor2_1 _4595_ (.Y(_0480_),
    .A(net823),
    .B(_0479_));
 sg13g2_nand2b_1 _4596_ (.Y(_0481_),
    .B(_0480_),
    .A_N(_0471_));
 sg13g2_xnor2_1 _4597_ (.Y(_0482_),
    .A(_0471_),
    .B(_0480_));
 sg13g2_nand2_1 _4598_ (.Y(_0483_),
    .A(_0456_),
    .B(_0482_));
 sg13g2_xnor2_1 _4599_ (.Y(_0484_),
    .A(_0456_),
    .B(_0482_));
 sg13g2_nand2_2 _4600_ (.Y(_0485_),
    .A(net856),
    .B(net848));
 sg13g2_xnor2_1 _4601_ (.Y(_0486_),
    .A(_3418_),
    .B(_3502_));
 sg13g2_xnor2_1 _4602_ (.Y(_0487_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_a22oi_1 _4603_ (.Y(_0488_),
    .B1(_0486_),
    .B2(_0487_),
    .A2(_0409_),
    .A1(net828));
 sg13g2_and2_1 _4604_ (.A(_3398_),
    .B(_3399_),
    .X(_0489_));
 sg13g2_xnor2_1 _4605_ (.Y(_0490_),
    .A(_3504_),
    .B(_0489_));
 sg13g2_xnor2_1 _4606_ (.Y(_0491_),
    .A(_0452_),
    .B(_0490_));
 sg13g2_xor2_1 _4607_ (.B(_0491_),
    .A(_0488_),
    .X(_0492_));
 sg13g2_nand2b_1 _4608_ (.Y(_0493_),
    .B(_0492_),
    .A_N(_3350_));
 sg13g2_o21ai_1 _4609_ (.B1(_0493_),
    .Y(_0494_),
    .A1(_0488_),
    .A2(_0491_));
 sg13g2_a21oi_1 _4610_ (.A1(_0445_),
    .A2(_0448_),
    .Y(_0495_),
    .B1(_0443_));
 sg13g2_a22oi_1 _4611_ (.Y(_0496_),
    .B1(_0452_),
    .B2(_0490_),
    .A2(_3289_),
    .A1(net828));
 sg13g2_nand2_1 _4612_ (.Y(_0497_),
    .A(net853),
    .B(net822));
 sg13g2_nor2_1 _4613_ (.A(_3279_),
    .B(_3329_),
    .Y(_0498_));
 sg13g2_a21oi_1 _4614_ (.A1(_0461_),
    .A2(_0466_),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_xor2_1 _4615_ (.B(_3506_),
    .A(_3380_),
    .X(_0500_));
 sg13g2_xnor2_1 _4616_ (.Y(_0501_),
    .A(_0499_),
    .B(_0500_));
 sg13g2_nor2_1 _4617_ (.A(_0496_),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_xor2_1 _4618_ (.B(_0501_),
    .A(_0496_),
    .X(_0503_));
 sg13g2_nor2b_1 _4619_ (.A(_0460_),
    .B_N(_0503_),
    .Y(_0504_));
 sg13g2_xor2_1 _4620_ (.B(_0503_),
    .A(_0460_),
    .X(_0505_));
 sg13g2_nor2_1 _4621_ (.A(_0495_),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_xor2_1 _4622_ (.B(_0505_),
    .A(_0495_),
    .X(_0507_));
 sg13g2_xnor2_1 _4623_ (.Y(_0508_),
    .A(_0494_),
    .B(_0507_));
 sg13g2_o21ai_1 _4624_ (.B1(_0483_),
    .Y(_0509_),
    .A1(_0484_),
    .A2(_0508_));
 sg13g2_o21ai_1 _4625_ (.B1(_0481_),
    .Y(_0510_),
    .A1(_0454_),
    .A2(_0470_));
 sg13g2_o21ai_1 _4626_ (.B1(_0476_),
    .Y(_0511_),
    .A1(_3293_),
    .A2(_3302_));
 sg13g2_nor2_1 _4627_ (.A(_0459_),
    .B(_0463_),
    .Y(_0512_));
 sg13g2_nand2_1 _4628_ (.Y(_0513_),
    .A(net825),
    .B(net844));
 sg13g2_xnor2_1 _4629_ (.Y(_0514_),
    .A(_0473_),
    .B(_0513_));
 sg13g2_xor2_1 _4630_ (.B(_0514_),
    .A(net808),
    .X(_0515_));
 sg13g2_o21ai_1 _4631_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_0459_),
    .A2(_0463_));
 sg13g2_xnor2_1 _4632_ (.Y(_0517_),
    .A(_0512_),
    .B(_0515_));
 sg13g2_nand2_1 _4633_ (.Y(_0518_),
    .A(_0511_),
    .B(_0517_));
 sg13g2_xnor2_1 _4634_ (.Y(_0519_),
    .A(_0511_),
    .B(_0517_));
 sg13g2_nand2b_1 _4635_ (.Y(_0520_),
    .B(_0186_),
    .A_N(_3524_));
 sg13g2_xnor2_1 _4636_ (.Y(_0521_),
    .A(_3524_),
    .B(_0186_));
 sg13g2_nand2b_1 _4637_ (.Y(_0522_),
    .B(_0521_),
    .A_N(_0497_));
 sg13g2_xnor2_1 _4638_ (.Y(_0523_),
    .A(_0497_),
    .B(_0521_));
 sg13g2_xor2_1 _4639_ (.B(_0523_),
    .A(_0467_),
    .X(_0524_));
 sg13g2_nor2_1 _4640_ (.A(_0458_),
    .B(_0513_),
    .Y(_0525_));
 sg13g2_xor2_1 _4641_ (.B(_0513_),
    .A(_0458_),
    .X(_0526_));
 sg13g2_xnor2_1 _4642_ (.Y(_0527_),
    .A(_0474_),
    .B(_0526_));
 sg13g2_and2_1 _4643_ (.A(_0524_),
    .B(_0527_),
    .X(_0528_));
 sg13g2_xnor2_1 _4644_ (.Y(_0529_),
    .A(_0524_),
    .B(_0527_));
 sg13g2_xor2_1 _4645_ (.B(_0529_),
    .A(_0469_),
    .X(_0530_));
 sg13g2_nand2b_1 _4646_ (.Y(_0531_),
    .B(_0530_),
    .A_N(_0519_));
 sg13g2_xnor2_1 _4647_ (.Y(_0532_),
    .A(_0519_),
    .B(_0530_));
 sg13g2_and2_1 _4648_ (.A(_0510_),
    .B(_0532_),
    .X(_0533_));
 sg13g2_xor2_1 _4649_ (.B(_0532_),
    .A(_0510_),
    .X(_0534_));
 sg13g2_nor2_1 _4650_ (.A(_0502_),
    .B(_0504_),
    .Y(_0535_));
 sg13g2_o21ai_1 _4651_ (.B1(_0478_),
    .Y(_0536_),
    .A1(_3302_),
    .A2(_0479_));
 sg13g2_a21o_1 _4652_ (.A2(_0500_),
    .A1(_0499_),
    .B1(_0498_),
    .X(_0537_));
 sg13g2_xor2_1 _4653_ (.B(_0497_),
    .A(_3524_),
    .X(_0538_));
 sg13g2_nand2_1 _4654_ (.Y(_0539_),
    .A(net830),
    .B(_0538_));
 sg13g2_xnor2_1 _4655_ (.Y(_0540_),
    .A(net862),
    .B(_0538_));
 sg13g2_nand2_1 _4656_ (.Y(_0541_),
    .A(_0537_),
    .B(_0540_));
 sg13g2_xnor2_1 _4657_ (.Y(_0542_),
    .A(_0537_),
    .B(_0540_));
 sg13g2_xnor2_1 _4658_ (.Y(_0543_),
    .A(_3507_),
    .B(_3519_));
 sg13g2_xor2_1 _4659_ (.B(_0543_),
    .A(_0542_),
    .X(_0544_));
 sg13g2_nand2_1 _4660_ (.Y(_0545_),
    .A(_0536_),
    .B(_0544_));
 sg13g2_xnor2_1 _4661_ (.Y(_0546_),
    .A(_0536_),
    .B(_0544_));
 sg13g2_xor2_1 _4662_ (.B(_0546_),
    .A(_0535_),
    .X(_0547_));
 sg13g2_xnor2_1 _4663_ (.Y(_0548_),
    .A(_0534_),
    .B(_0547_));
 sg13g2_nor2b_1 _4664_ (.A(_0548_),
    .B_N(_0509_),
    .Y(_0549_));
 sg13g2_a21oi_2 _4665_ (.B1(_0506_),
    .Y(_0550_),
    .A2(_0507_),
    .A1(_0494_));
 sg13g2_xor2_1 _4666_ (.B(_0548_),
    .A(_0509_),
    .X(_0551_));
 sg13g2_nor2_1 _4667_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_nor2_1 _4668_ (.A(_0549_),
    .B(_0552_),
    .Y(_0553_));
 sg13g2_o21ai_1 _4669_ (.B1(_0545_),
    .Y(_0554_),
    .A1(_0535_),
    .A2(_0546_));
 sg13g2_a21o_1 _4670_ (.A2(_0547_),
    .A1(_0534_),
    .B1(_0533_),
    .X(_0555_));
 sg13g2_o21ai_1 _4671_ (.B1(_0531_),
    .Y(_0556_),
    .A1(_0469_),
    .A2(_0529_));
 sg13g2_a22oi_1 _4672_ (.Y(_0557_),
    .B1(_0514_),
    .B2(net808),
    .A2(_0409_),
    .A1(net823));
 sg13g2_inv_1 _4673_ (.Y(_0558_),
    .A(_0557_));
 sg13g2_a21oi_2 _4674_ (.B1(_0525_),
    .Y(_0559_),
    .A2(_0526_),
    .A1(_0473_));
 sg13g2_nor2_1 _4675_ (.A(_3290_),
    .B(_3302_),
    .Y(_0560_));
 sg13g2_a22oi_1 _4676_ (.Y(_0561_),
    .B1(net843),
    .B2(net850),
    .A2(net845),
    .A1(net825));
 sg13g2_nor2_2 _4677_ (.A(_0560_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_xnor2_1 _4678_ (.Y(_0563_),
    .A(net808),
    .B(_0562_));
 sg13g2_nor2_1 _4679_ (.A(_0559_),
    .B(_0563_),
    .Y(_0564_));
 sg13g2_xor2_1 _4680_ (.B(_0563_),
    .A(_0559_),
    .X(_0565_));
 sg13g2_xnor2_1 _4681_ (.Y(_0566_),
    .A(_0557_),
    .B(_0565_));
 sg13g2_a21oi_1 _4682_ (.A1(_0467_),
    .A2(_0523_),
    .Y(_0567_),
    .B1(_0528_));
 sg13g2_xnor2_1 _4683_ (.Y(_0568_),
    .A(net848),
    .B(_0562_));
 sg13g2_nand2_1 _4684_ (.Y(_0569_),
    .A(_0520_),
    .B(_0522_));
 sg13g2_xnor2_1 _4685_ (.Y(_0570_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_nand2_1 _4686_ (.Y(_0571_),
    .A(_0569_),
    .B(_0570_));
 sg13g2_xnor2_1 _4687_ (.Y(_0572_),
    .A(_0569_),
    .B(_0570_));
 sg13g2_xor2_1 _4688_ (.B(_0572_),
    .A(_0568_),
    .X(_0573_));
 sg13g2_nor2b_1 _4689_ (.A(_0567_),
    .B_N(_0573_),
    .Y(_0574_));
 sg13g2_xnor2_1 _4690_ (.Y(_0575_),
    .A(_0567_),
    .B(_0573_));
 sg13g2_xnor2_1 _4691_ (.Y(_0576_),
    .A(_0566_),
    .B(_0575_));
 sg13g2_nand2b_1 _4692_ (.Y(_0577_),
    .B(_0556_),
    .A_N(_0576_));
 sg13g2_xor2_1 _4693_ (.B(_0576_),
    .A(_0556_),
    .X(_0578_));
 sg13g2_o21ai_1 _4694_ (.B1(_0541_),
    .Y(_0579_),
    .A1(_0542_),
    .A2(_0543_));
 sg13g2_and2_1 _4695_ (.A(_0516_),
    .B(_0518_),
    .X(_0580_));
 sg13g2_o21ai_1 _4696_ (.B1(_0539_),
    .Y(_0581_),
    .A1(_3279_),
    .A2(_3344_));
 sg13g2_xnor2_1 _4697_ (.Y(_0582_),
    .A(_3523_),
    .B(_3528_));
 sg13g2_xor2_1 _4698_ (.B(_0582_),
    .A(_0581_),
    .X(_0583_));
 sg13g2_nor2b_1 _4699_ (.A(_0395_),
    .B_N(_0583_),
    .Y(_0584_));
 sg13g2_xnor2_1 _4700_ (.Y(_0585_),
    .A(_0395_),
    .B(_0583_));
 sg13g2_nor2b_1 _4701_ (.A(_0580_),
    .B_N(_0585_),
    .Y(_0586_));
 sg13g2_xnor2_1 _4702_ (.Y(_0587_),
    .A(_0580_),
    .B(_0585_));
 sg13g2_xnor2_1 _4703_ (.Y(_0588_),
    .A(_0579_),
    .B(_0587_));
 sg13g2_xor2_1 _4704_ (.B(_0588_),
    .A(_0578_),
    .X(_0589_));
 sg13g2_xnor2_1 _4705_ (.Y(_0590_),
    .A(_0555_),
    .B(_0589_));
 sg13g2_nor2b_1 _4706_ (.A(_0590_),
    .B_N(_0554_),
    .Y(_0591_));
 sg13g2_xnor2_1 _4707_ (.Y(_0592_),
    .A(_0554_),
    .B(_0590_));
 sg13g2_nand2b_1 _4708_ (.Y(_0593_),
    .B(_0592_),
    .A_N(_0553_));
 sg13g2_a21o_1 _4709_ (.A2(_0589_),
    .A1(_0555_),
    .B1(_0591_),
    .X(_0594_));
 sg13g2_a21oi_1 _4710_ (.A1(_0579_),
    .A2(_0587_),
    .Y(_0595_),
    .B1(_0586_));
 sg13g2_o21ai_1 _4711_ (.B1(_0577_),
    .Y(_0596_),
    .A1(_0578_),
    .A2(_0588_));
 sg13g2_a21oi_1 _4712_ (.A1(_0566_),
    .A2(_0575_),
    .Y(_0597_),
    .B1(_0574_));
 sg13g2_a21oi_1 _4713_ (.A1(net808),
    .A2(_0562_),
    .Y(_0598_),
    .B1(_0560_));
 sg13g2_inv_1 _4714_ (.Y(_0599_),
    .A(_0598_));
 sg13g2_a21oi_1 _4715_ (.A1(net847),
    .A2(_0562_),
    .Y(_0600_),
    .B1(_0560_));
 sg13g2_xnor2_1 _4716_ (.Y(_0601_),
    .A(net807),
    .B(_0406_));
 sg13g2_nor2_1 _4717_ (.A(_0600_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_xor2_1 _4718_ (.B(_0601_),
    .A(_0600_),
    .X(_0603_));
 sg13g2_xnor2_1 _4719_ (.Y(_0604_),
    .A(_0598_),
    .B(_0603_));
 sg13g2_inv_1 _4720_ (.Y(_0605_),
    .A(_0604_));
 sg13g2_o21ai_1 _4721_ (.B1(_0571_),
    .Y(_0606_),
    .A1(_0568_),
    .A2(_0572_));
 sg13g2_xor2_1 _4722_ (.B(_0402_),
    .A(_0401_),
    .X(_0607_));
 sg13g2_xnor2_1 _4723_ (.Y(_0608_),
    .A(_0606_),
    .B(_0607_));
 sg13g2_nor2_1 _4724_ (.A(_0605_),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_xnor2_1 _4725_ (.Y(_0610_),
    .A(_0605_),
    .B(_0608_));
 sg13g2_nor2_1 _4726_ (.A(_0597_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_xor2_1 _4727_ (.B(_0610_),
    .A(_0597_),
    .X(_0612_));
 sg13g2_a21o_1 _4728_ (.A2(_0582_),
    .A1(_0581_),
    .B1(_0584_),
    .X(_0613_));
 sg13g2_a21oi_1 _4729_ (.A1(_0558_),
    .A2(_0565_),
    .Y(_0614_),
    .B1(_0564_));
 sg13g2_mux2_1 _4730_ (.A0(_3527_),
    .A1(_3526_),
    .S(_3523_),
    .X(_0615_));
 sg13g2_xnor2_1 _4731_ (.Y(_0616_),
    .A(_0173_),
    .B(_0615_));
 sg13g2_xnor2_1 _4732_ (.Y(_0617_),
    .A(_0353_),
    .B(_0616_));
 sg13g2_nor2_1 _4733_ (.A(_0614_),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_xor2_1 _4734_ (.B(_0617_),
    .A(_0614_),
    .X(_0619_));
 sg13g2_xor2_1 _4735_ (.B(_0619_),
    .A(_0613_),
    .X(_0620_));
 sg13g2_xnor2_1 _4736_ (.Y(_0621_),
    .A(_0612_),
    .B(_0620_));
 sg13g2_nand2b_1 _4737_ (.Y(_0622_),
    .B(_0596_),
    .A_N(_0621_));
 sg13g2_xor2_1 _4738_ (.B(_0621_),
    .A(_0596_),
    .X(_0623_));
 sg13g2_xor2_1 _4739_ (.B(_0623_),
    .A(_0595_),
    .X(_0624_));
 sg13g2_nand2_1 _4740_ (.Y(_0625_),
    .A(_0594_),
    .B(_0624_));
 sg13g2_xnor2_1 _4741_ (.Y(_0626_),
    .A(_0594_),
    .B(_0624_));
 sg13g2_nor2_1 _4742_ (.A(_0593_),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_nand2_1 _4743_ (.Y(_0628_),
    .A(_0593_),
    .B(_0626_));
 sg13g2_xor2_1 _4744_ (.B(_0592_),
    .A(_0553_),
    .X(_0629_));
 sg13g2_xor2_1 _4745_ (.B(_0455_),
    .A(_0449_),
    .X(_0630_));
 sg13g2_and2_1 _4746_ (.A(net858),
    .B(_3300_),
    .X(_0631_));
 sg13g2_nand2_1 _4747_ (.Y(_0632_),
    .A(net854),
    .B(_3297_));
 sg13g2_xnor2_1 _4748_ (.Y(_0633_),
    .A(_0631_),
    .B(_0632_));
 sg13g2_nand2_1 _4749_ (.Y(_0634_),
    .A(_0436_),
    .B(_0633_));
 sg13g2_o21ai_1 _4750_ (.B1(_0634_),
    .Y(_0635_),
    .A1(_3302_),
    .A2(_0457_));
 sg13g2_nor3_1 _4751_ (.A(net852),
    .B(_0185_),
    .C(_0485_),
    .Y(_0636_));
 sg13g2_o21ai_1 _4752_ (.B1(_0440_),
    .Y(_0637_),
    .A1(_3303_),
    .A2(_0446_));
 sg13g2_nor2b_1 _4753_ (.A(_0447_),
    .B_N(_0637_),
    .Y(_0638_));
 sg13g2_xnor2_1 _4754_ (.Y(_0639_),
    .A(_0636_),
    .B(_0638_));
 sg13g2_nor2b_1 _4755_ (.A(_0639_),
    .B_N(_0635_),
    .Y(_0640_));
 sg13g2_xor2_1 _4756_ (.B(_0639_),
    .A(_0635_),
    .X(_0641_));
 sg13g2_xnor2_1 _4757_ (.Y(_0642_),
    .A(_0437_),
    .B(_0441_));
 sg13g2_nand2b_1 _4758_ (.Y(_0643_),
    .B(_0642_),
    .A_N(_0641_));
 sg13g2_nor2_1 _4759_ (.A(_0630_),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_a22oi_1 _4760_ (.Y(_0645_),
    .B1(_0485_),
    .B2(_0632_),
    .A2(_0473_),
    .A1(net829));
 sg13g2_nand3_1 _4761_ (.B(_3498_),
    .C(_3501_),
    .A(_3496_),
    .Y(_0646_));
 sg13g2_a21o_1 _4762_ (.A2(_3498_),
    .A1(_3496_),
    .B1(_3501_),
    .X(_0647_));
 sg13g2_nand3_1 _4763_ (.B(_0646_),
    .C(_0647_),
    .A(_0645_),
    .Y(_0648_));
 sg13g2_o21ai_1 _4764_ (.B1(_0648_),
    .Y(_0649_),
    .A1(_3279_),
    .A2(_0474_));
 sg13g2_xnor2_1 _4765_ (.Y(_0650_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_nor2b_1 _4766_ (.A(_0650_),
    .B_N(_0649_),
    .Y(_0651_));
 sg13g2_xnor2_1 _4767_ (.Y(_0652_),
    .A(_0649_),
    .B(_0650_));
 sg13g2_nor2b_1 _4768_ (.A(_3299_),
    .B_N(_0652_),
    .Y(_0653_));
 sg13g2_nor2_1 _4769_ (.A(_0651_),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_a21oi_1 _4770_ (.A1(_0636_),
    .A2(_0638_),
    .Y(_0655_),
    .B1(_0640_));
 sg13g2_xor2_1 _4771_ (.B(_0492_),
    .A(_3350_),
    .X(_0656_));
 sg13g2_or2_1 _4772_ (.X(_0657_),
    .B(_0656_),
    .A(_0655_));
 sg13g2_xnor2_1 _4773_ (.Y(_0658_),
    .A(_0655_),
    .B(_0656_));
 sg13g2_xor2_1 _4774_ (.B(_0658_),
    .A(_0654_),
    .X(_0659_));
 sg13g2_xor2_1 _4775_ (.B(_0643_),
    .A(_0630_),
    .X(_0660_));
 sg13g2_a21oi_1 _4776_ (.A1(_0659_),
    .A2(_0660_),
    .Y(_0661_),
    .B1(_0644_));
 sg13g2_xor2_1 _4777_ (.B(_0508_),
    .A(_0484_),
    .X(_0662_));
 sg13g2_nor2b_1 _4778_ (.A(_0661_),
    .B_N(_0662_),
    .Y(_0663_));
 sg13g2_o21ai_1 _4779_ (.B1(_0657_),
    .Y(_0664_),
    .A1(_0654_),
    .A2(_0658_));
 sg13g2_xnor2_1 _4780_ (.Y(_0665_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_a21oi_1 _4781_ (.A1(_0664_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(_0663_));
 sg13g2_xor2_1 _4782_ (.B(_0551_),
    .A(_0550_),
    .X(_0667_));
 sg13g2_nand2b_1 _4783_ (.Y(_0668_),
    .B(_0667_),
    .A_N(_0666_));
 sg13g2_xnor2_1 _4784_ (.Y(_0669_),
    .A(_0666_),
    .B(_0667_));
 sg13g2_nand2b_1 _4785_ (.Y(_0670_),
    .B(_0669_),
    .A_N(_0458_));
 sg13g2_nand2_1 _4786_ (.Y(_0671_),
    .A(_0668_),
    .B(_0670_));
 sg13g2_a21oi_2 _4787_ (.B1(_0629_),
    .Y(_0672_),
    .A2(_0670_),
    .A1(_0668_));
 sg13g2_inv_1 _4788_ (.Y(_0673_),
    .A(_0672_));
 sg13g2_xor2_1 _4789_ (.B(_0671_),
    .A(_0629_),
    .X(_0674_));
 sg13g2_xor2_1 _4790_ (.B(_0633_),
    .A(_0436_),
    .X(_0675_));
 sg13g2_nand2_1 _4791_ (.Y(_0676_),
    .A(net829),
    .B(net823));
 sg13g2_a22oi_1 _4792_ (.Y(_0677_),
    .B1(_3300_),
    .B2(net854),
    .A2(net846),
    .A1(net855));
 sg13g2_a21oi_2 _4793_ (.B1(_0677_),
    .Y(_0678_),
    .A2(_3301_),
    .A1(net829));
 sg13g2_inv_1 _4794_ (.Y(_0679_),
    .A(_0678_));
 sg13g2_nand2_1 _4795_ (.Y(_0680_),
    .A(net848),
    .B(_0184_));
 sg13g2_inv_1 _4796_ (.Y(_0681_),
    .A(_0680_));
 sg13g2_a22oi_1 _4797_ (.Y(_0682_),
    .B1(_0678_),
    .B2(_0681_),
    .A2(_3301_),
    .A1(net829));
 sg13g2_nand2b_1 _4798_ (.Y(_0683_),
    .B(_0675_),
    .A_N(_0682_));
 sg13g2_xor2_1 _4799_ (.B(_0682_),
    .A(_0675_),
    .X(_0684_));
 sg13g2_xnor2_1 _4800_ (.Y(_0685_),
    .A(_0436_),
    .B(_0485_));
 sg13g2_nor2b_1 _4801_ (.A(_0684_),
    .B_N(_0685_),
    .Y(_0686_));
 sg13g2_xnor2_1 _4802_ (.Y(_0687_),
    .A(_0641_),
    .B(_0642_));
 sg13g2_nand2_1 _4803_ (.Y(_0688_),
    .A(_0686_),
    .B(_0687_));
 sg13g2_xnor2_1 _4804_ (.Y(_0689_),
    .A(_0686_),
    .B(_0687_));
 sg13g2_o21ai_1 _4805_ (.B1(_3497_),
    .Y(_0690_),
    .A1(_3466_),
    .A2(_3493_));
 sg13g2_nand2_1 _4806_ (.Y(_0691_),
    .A(_3498_),
    .B(_0690_));
 sg13g2_o21ai_1 _4807_ (.B1(_0676_),
    .Y(_0692_),
    .A1(_0679_),
    .A2(_0691_));
 sg13g2_a21o_1 _4808_ (.A2(_0647_),
    .A1(_0646_),
    .B1(_0645_),
    .X(_0693_));
 sg13g2_nand3_1 _4809_ (.B(_0692_),
    .C(_0693_),
    .A(_0648_),
    .Y(_0694_));
 sg13g2_a21o_1 _4810_ (.A2(_0693_),
    .A1(_0648_),
    .B1(_0692_),
    .X(_0695_));
 sg13g2_nand3_1 _4811_ (.B(_0694_),
    .C(_0695_),
    .A(_0631_),
    .Y(_0696_));
 sg13g2_nand2_1 _4812_ (.Y(_0697_),
    .A(_0694_),
    .B(_0696_));
 sg13g2_xnor2_1 _4813_ (.Y(_0698_),
    .A(_3299_),
    .B(_0652_));
 sg13g2_nor2b_1 _4814_ (.A(_0683_),
    .B_N(_0698_),
    .Y(_0699_));
 sg13g2_xnor2_1 _4815_ (.Y(_0700_),
    .A(_0683_),
    .B(_0698_));
 sg13g2_xnor2_1 _4816_ (.Y(_0701_),
    .A(_0697_),
    .B(_0700_));
 sg13g2_o21ai_1 _4817_ (.B1(_0688_),
    .Y(_0702_),
    .A1(_0689_),
    .A2(_0701_));
 sg13g2_xnor2_1 _4818_ (.Y(_0703_),
    .A(_0659_),
    .B(_0660_));
 sg13g2_nor2b_1 _4819_ (.A(_0703_),
    .B_N(_0702_),
    .Y(_0704_));
 sg13g2_a21o_1 _4820_ (.A2(_0700_),
    .A1(_0697_),
    .B1(_0699_),
    .X(_0705_));
 sg13g2_xnor2_1 _4821_ (.Y(_0706_),
    .A(_0702_),
    .B(_0703_));
 sg13g2_a21oi_2 _4822_ (.B1(_0704_),
    .Y(_0707_),
    .A2(_0706_),
    .A1(_0705_));
 sg13g2_xnor2_1 _4823_ (.Y(_0708_),
    .A(_0664_),
    .B(_0665_));
 sg13g2_nor2_1 _4824_ (.A(_0707_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_xnor2_1 _4825_ (.Y(_0710_),
    .A(_0458_),
    .B(_0669_));
 sg13g2_xor2_1 _4826_ (.B(_0710_),
    .A(_0709_),
    .X(_0711_));
 sg13g2_nand2_2 _4827_ (.Y(_0712_),
    .A(net858),
    .B(net855));
 sg13g2_and3_1 _4828_ (.X(_0713_),
    .A(net858),
    .B(net855),
    .C(_3277_));
 sg13g2_xnor2_1 _4829_ (.Y(_0714_),
    .A(_3277_),
    .B(_0712_));
 sg13g2_xor2_1 _4830_ (.B(_0712_),
    .A(_3277_),
    .X(_0715_));
 sg13g2_a21oi_1 _4831_ (.A1(_3476_),
    .A2(_3478_),
    .Y(_0716_),
    .B1(_3488_));
 sg13g2_o21ai_1 _4832_ (.B1(_3489_),
    .Y(_0717_),
    .A1(_3475_),
    .A2(_3477_));
 sg13g2_nor3_1 _4833_ (.A(_3490_),
    .B(_0715_),
    .C(_0716_),
    .Y(_0718_));
 sg13g2_or2_1 _4834_ (.X(_0719_),
    .B(_0718_),
    .A(_0713_));
 sg13g2_nand2_1 _4835_ (.Y(_0720_),
    .A(net828),
    .B(_0631_));
 sg13g2_nand2_1 _4836_ (.Y(_0721_),
    .A(net855),
    .B(_3300_));
 sg13g2_nand2_1 _4837_ (.Y(_0722_),
    .A(_0457_),
    .B(_0721_));
 sg13g2_nand2_1 _4838_ (.Y(_0723_),
    .A(_0720_),
    .B(_0722_));
 sg13g2_xnor2_1 _4839_ (.Y(_0724_),
    .A(_3459_),
    .B(_3465_));
 sg13g2_xnor2_1 _4840_ (.Y(_0725_),
    .A(_3492_),
    .B(_0724_));
 sg13g2_xnor2_1 _4841_ (.Y(_0726_),
    .A(_0723_),
    .B(_0725_));
 sg13g2_nand2b_1 _4842_ (.Y(_0727_),
    .B(_0719_),
    .A_N(_0726_));
 sg13g2_xor2_1 _4843_ (.B(_0726_),
    .A(_0719_),
    .X(_0728_));
 sg13g2_o21ai_1 _4844_ (.B1(_0727_),
    .Y(_0729_),
    .A1(_0457_),
    .A2(_0728_));
 sg13g2_nand2_1 _4845_ (.Y(_0730_),
    .A(net844),
    .B(_0434_));
 sg13g2_o21ai_1 _4846_ (.B1(_0720_),
    .Y(_0731_),
    .A1(_0723_),
    .A2(_0725_));
 sg13g2_xnor2_1 _4847_ (.Y(_0732_),
    .A(_0679_),
    .B(_0691_));
 sg13g2_nor2b_1 _4848_ (.A(_0732_),
    .B_N(_0731_),
    .Y(_0733_));
 sg13g2_xnor2_1 _4849_ (.Y(_0734_),
    .A(_0731_),
    .B(_0732_));
 sg13g2_xnor2_1 _4850_ (.Y(_0735_),
    .A(net858),
    .B(_0734_));
 sg13g2_nor2_1 _4851_ (.A(_0730_),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_xor2_1 _4852_ (.B(_0735_),
    .A(_0730_),
    .X(_0737_));
 sg13g2_xnor2_1 _4853_ (.Y(_0738_),
    .A(_0729_),
    .B(_0737_));
 sg13g2_nand2_1 _4854_ (.Y(_0739_),
    .A(net846),
    .B(net815));
 sg13g2_xor2_1 _4855_ (.B(_0680_),
    .A(_0678_),
    .X(_0740_));
 sg13g2_nor2_1 _4856_ (.A(_0739_),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_and2_1 _4857_ (.A(_0739_),
    .B(_0740_),
    .X(_0742_));
 sg13g2_nor3_1 _4858_ (.A(_0680_),
    .B(_0741_),
    .C(_0742_),
    .Y(_0743_));
 sg13g2_inv_1 _4859_ (.Y(_0744_),
    .A(_0743_));
 sg13g2_xor2_1 _4860_ (.B(_0739_),
    .A(_0678_),
    .X(_0745_));
 sg13g2_nor2_1 _4861_ (.A(_0738_),
    .B(_0745_),
    .Y(_0746_));
 sg13g2_xor2_1 _4862_ (.B(_0685_),
    .A(_0684_),
    .X(_0747_));
 sg13g2_xnor2_1 _4863_ (.Y(_0748_),
    .A(_0743_),
    .B(_0747_));
 sg13g2_a21oi_1 _4864_ (.A1(net858),
    .A2(_0734_),
    .Y(_0749_),
    .B1(_0733_));
 sg13g2_a21o_1 _4865_ (.A2(_0695_),
    .A1(_0694_),
    .B1(_0631_),
    .X(_0750_));
 sg13g2_and3_1 _4866_ (.X(_0751_),
    .A(_0696_),
    .B(_0741_),
    .C(_0750_));
 sg13g2_a21oi_1 _4867_ (.A1(_0696_),
    .A2(_0750_),
    .Y(_0752_),
    .B1(_0741_));
 sg13g2_or3_1 _4868_ (.A(_0749_),
    .B(_0751_),
    .C(_0752_),
    .X(_0753_));
 sg13g2_o21ai_1 _4869_ (.B1(_0749_),
    .Y(_0754_),
    .A1(_0751_),
    .A2(_0752_));
 sg13g2_nand3_1 _4870_ (.B(_0753_),
    .C(_0754_),
    .A(_0748_),
    .Y(_0755_));
 sg13g2_a21o_1 _4871_ (.A2(_0754_),
    .A1(_0753_),
    .B1(_0748_),
    .X(_0756_));
 sg13g2_nand3_1 _4872_ (.B(_0755_),
    .C(_0756_),
    .A(_0746_),
    .Y(_0757_));
 sg13g2_a21oi_1 _4873_ (.A1(_0729_),
    .A2(_0737_),
    .Y(_0758_),
    .B1(_0736_));
 sg13g2_inv_1 _4874_ (.Y(_0759_),
    .A(_0758_));
 sg13g2_a21o_1 _4875_ (.A2(_0756_),
    .A1(_0755_),
    .B1(_0746_),
    .X(_0760_));
 sg13g2_nand3_1 _4876_ (.B(_0759_),
    .C(_0760_),
    .A(_0757_),
    .Y(_0761_));
 sg13g2_nand2_1 _4877_ (.Y(_0762_),
    .A(_0757_),
    .B(_0761_));
 sg13g2_nand2b_1 _4878_ (.Y(_0763_),
    .B(_0753_),
    .A_N(_0751_));
 sg13g2_o21ai_1 _4879_ (.B1(_0755_),
    .Y(_0764_),
    .A1(_0744_),
    .A2(_0747_));
 sg13g2_xor2_1 _4880_ (.B(_0701_),
    .A(_0689_),
    .X(_0765_));
 sg13g2_xnor2_1 _4881_ (.Y(_0766_),
    .A(_0764_),
    .B(_0765_));
 sg13g2_nor2b_1 _4882_ (.A(_0766_),
    .B_N(_0763_),
    .Y(_0767_));
 sg13g2_xor2_1 _4883_ (.B(_0766_),
    .A(_0763_),
    .X(_0768_));
 sg13g2_nand2b_1 _4884_ (.Y(_0769_),
    .B(_0762_),
    .A_N(_0768_));
 sg13g2_a21oi_1 _4885_ (.A1(_0764_),
    .A2(_0765_),
    .Y(_0770_),
    .B1(_0767_));
 sg13g2_xnor2_1 _4886_ (.Y(_0771_),
    .A(_0705_),
    .B(_0706_));
 sg13g2_nor2_1 _4887_ (.A(_0770_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_xor2_1 _4888_ (.B(_0771_),
    .A(_0770_),
    .X(_0773_));
 sg13g2_nor2b_1 _4889_ (.A(_0769_),
    .B_N(_0773_),
    .Y(_0774_));
 sg13g2_xnor2_1 _4890_ (.Y(_0775_),
    .A(_0762_),
    .B(_0768_));
 sg13g2_a21o_1 _4891_ (.A2(_0760_),
    .A1(_0757_),
    .B1(_0759_),
    .X(_0776_));
 sg13g2_xnor2_1 _4892_ (.Y(_0777_),
    .A(_0738_),
    .B(_0745_));
 sg13g2_xor2_1 _4893_ (.B(_0728_),
    .A(_0457_),
    .X(_0778_));
 sg13g2_a21oi_1 _4894_ (.A1(_3491_),
    .A2(_0717_),
    .Y(_0779_),
    .B1(_0714_));
 sg13g2_nor3_1 _4895_ (.A(_3490_),
    .B(_0714_),
    .C(_0716_),
    .Y(_0780_));
 sg13g2_a21oi_1 _4896_ (.A1(_3491_),
    .A2(_0717_),
    .Y(_0781_),
    .B1(_0715_));
 sg13g2_nor3_1 _4897_ (.A(_3279_),
    .B(_0718_),
    .C(_0779_),
    .Y(_0782_));
 sg13g2_a21oi_1 _4898_ (.A1(_3491_),
    .A2(_0717_),
    .Y(_0783_),
    .B1(_0712_));
 sg13g2_inv_1 _4899_ (.Y(_0784_),
    .A(_0783_));
 sg13g2_nor2_1 _4900_ (.A(_0782_),
    .B(_0783_),
    .Y(_0785_));
 sg13g2_nor2b_1 _4901_ (.A(_0785_),
    .B_N(_0778_),
    .Y(_0786_));
 sg13g2_xnor2_1 _4902_ (.Y(_0787_),
    .A(_0778_),
    .B(_0785_));
 sg13g2_nand2b_1 _4903_ (.Y(_0788_),
    .B(_0185_),
    .A_N(net855));
 sg13g2_nand3_1 _4904_ (.B(_0435_),
    .C(_0788_),
    .A(net844),
    .Y(_0789_));
 sg13g2_inv_1 _4905_ (.Y(_0790_),
    .A(_0789_));
 sg13g2_a21oi_1 _4906_ (.A1(_0787_),
    .A2(_0790_),
    .Y(_0791_),
    .B1(_0786_));
 sg13g2_nor2_1 _4907_ (.A(_0777_),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_nand3_1 _4908_ (.B(_0776_),
    .C(_0792_),
    .A(_0761_),
    .Y(_0793_));
 sg13g2_nand4_1 _4909_ (.B(_0775_),
    .C(_0776_),
    .A(_0761_),
    .Y(_0794_),
    .D(_0792_));
 sg13g2_xnor2_1 _4910_ (.Y(_0795_),
    .A(_0777_),
    .B(_0791_));
 sg13g2_nand2_1 _4911_ (.Y(_0796_),
    .A(net854),
    .B(net815));
 sg13g2_xor2_1 _4912_ (.B(_0796_),
    .A(net855),
    .X(_0797_));
 sg13g2_xnor2_1 _4913_ (.Y(_0798_),
    .A(_3484_),
    .B(_3486_));
 sg13g2_nand2b_1 _4914_ (.Y(_0799_),
    .B(_0798_),
    .A_N(_0797_));
 sg13g2_o21ai_1 _4915_ (.B1(_0799_),
    .Y(_0800_),
    .A1(_3279_),
    .A2(_0185_));
 sg13g2_xnor2_1 _4916_ (.Y(_0801_),
    .A(_3479_),
    .B(_3487_));
 sg13g2_nand2b_1 _4917_ (.Y(_0802_),
    .B(_0800_),
    .A_N(_0801_));
 sg13g2_nand2_2 _4918_ (.Y(_0803_),
    .A(net859),
    .B(net815));
 sg13g2_xor2_1 _4919_ (.B(_0801_),
    .A(_0800_),
    .X(_0804_));
 sg13g2_o21ai_1 _4920_ (.B1(_0802_),
    .Y(_0805_),
    .A1(_0803_),
    .A2(_0804_));
 sg13g2_nor3_1 _4921_ (.A(net828),
    .B(_0780_),
    .C(_0781_),
    .Y(_0806_));
 sg13g2_o21ai_1 _4922_ (.B1(_0712_),
    .Y(_0807_),
    .A1(_0782_),
    .A2(_0806_));
 sg13g2_and3_1 _4923_ (.X(_0808_),
    .A(_0784_),
    .B(_0805_),
    .C(_0807_));
 sg13g2_nand3_1 _4924_ (.B(_0805_),
    .C(_0807_),
    .A(_0784_),
    .Y(_0809_));
 sg13g2_xnor2_1 _4925_ (.Y(_0810_),
    .A(_0787_),
    .B(_0789_));
 sg13g2_and2_1 _4926_ (.A(_0808_),
    .B(_0810_),
    .X(_0811_));
 sg13g2_nor2b_1 _4927_ (.A(_0795_),
    .B_N(_0811_),
    .Y(_0812_));
 sg13g2_a21o_1 _4928_ (.A2(_0776_),
    .A1(_0761_),
    .B1(_0792_),
    .X(_0813_));
 sg13g2_and3_1 _4929_ (.X(_0814_),
    .A(_0793_),
    .B(_0812_),
    .C(_0813_));
 sg13g2_nand3_1 _4930_ (.B(_0812_),
    .C(_0813_),
    .A(_0793_),
    .Y(_0815_));
 sg13g2_xnor2_1 _4931_ (.Y(_0816_),
    .A(_0808_),
    .B(_0810_));
 sg13g2_xor2_1 _4932_ (.B(_0804_),
    .A(_0803_),
    .X(_0817_));
 sg13g2_a21oi_1 _4933_ (.A1(_3366_),
    .A2(net809),
    .Y(_0818_),
    .B1(_3469_));
 sg13g2_nor2_1 _4934_ (.A(_3485_),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_xnor2_1 _4935_ (.Y(_0820_),
    .A(_0797_),
    .B(_0798_));
 sg13g2_and3_1 _4936_ (.X(_0821_),
    .A(_0434_),
    .B(_0819_),
    .C(_0820_));
 sg13g2_nand2_1 _4937_ (.Y(_0822_),
    .A(_0817_),
    .B(_0821_));
 sg13g2_xor2_1 _4938_ (.B(_0821_),
    .A(_0817_),
    .X(_0823_));
 sg13g2_nor2b_1 _4939_ (.A(_0803_),
    .B_N(_0823_),
    .Y(_0824_));
 sg13g2_a21o_1 _4940_ (.A2(_0807_),
    .A1(_0784_),
    .B1(_0805_),
    .X(_0825_));
 sg13g2_and3_1 _4941_ (.X(_0826_),
    .A(_0809_),
    .B(_0824_),
    .C(_0825_));
 sg13g2_a21oi_1 _4942_ (.A1(_0809_),
    .A2(_0825_),
    .Y(_0827_),
    .B1(_0824_));
 sg13g2_or3_1 _4943_ (.A(_0822_),
    .B(_0826_),
    .C(_0827_),
    .X(_0828_));
 sg13g2_nand2b_1 _4944_ (.Y(_0829_),
    .B(_0828_),
    .A_N(_0826_));
 sg13g2_nand2b_1 _4945_ (.Y(_0830_),
    .B(_0829_),
    .A_N(_0816_));
 sg13g2_xnor2_1 _4946_ (.Y(_0831_),
    .A(_0795_),
    .B(_0811_));
 sg13g2_nor2_1 _4947_ (.A(_0795_),
    .B(_0830_),
    .Y(_0832_));
 sg13g2_xor2_1 _4948_ (.B(_0829_),
    .A(_0816_),
    .X(_0833_));
 sg13g2_o21ai_1 _4949_ (.B1(_0822_),
    .Y(_0834_),
    .A1(_0826_),
    .A2(_0827_));
 sg13g2_a21oi_1 _4950_ (.A1(_0434_),
    .A2(_0819_),
    .Y(_0835_),
    .B1(_0820_));
 sg13g2_nor4_2 _4951_ (.A(_0796_),
    .B(_0804_),
    .C(_0821_),
    .Y(_0836_),
    .D(_0835_));
 sg13g2_and3_1 _4952_ (.X(_0837_),
    .A(_0828_),
    .B(_0834_),
    .C(_0836_));
 sg13g2_nand3_1 _4953_ (.B(_0834_),
    .C(_0836_),
    .A(_0828_),
    .Y(_0838_));
 sg13g2_a21oi_1 _4954_ (.A1(_0828_),
    .A2(_0834_),
    .Y(_0839_),
    .B1(_0836_));
 sg13g2_or4_1 _4955_ (.A(_0435_),
    .B(_0798_),
    .C(_0804_),
    .D(_0819_),
    .X(_0840_));
 sg13g2_nor3_1 _4956_ (.A(_0837_),
    .B(_0839_),
    .C(_0840_),
    .Y(_0841_));
 sg13g2_a21oi_1 _4957_ (.A1(net858),
    .A2(net815),
    .Y(_0842_),
    .B1(_0823_));
 sg13g2_nor3_1 _4958_ (.A(_3365_),
    .B(_3440_),
    .C(_0185_),
    .Y(_0843_));
 sg13g2_nand3_1 _4959_ (.B(_0819_),
    .C(_0843_),
    .A(_3486_),
    .Y(_0844_));
 sg13g2_nor3_1 _4960_ (.A(_0824_),
    .B(_0842_),
    .C(_0844_),
    .Y(_0845_));
 sg13g2_o21ai_1 _4961_ (.B1(_0840_),
    .Y(_0846_),
    .A1(_0837_),
    .A2(_0839_));
 sg13g2_nand2b_1 _4962_ (.Y(_0847_),
    .B(_0846_),
    .A_N(_0841_));
 sg13g2_a21o_1 _4963_ (.A2(_0846_),
    .A1(_0845_),
    .B1(_0841_),
    .X(_0848_));
 sg13g2_xnor2_1 _4964_ (.Y(_0849_),
    .A(_0833_),
    .B(_0837_));
 sg13g2_nand2_1 _4965_ (.Y(_0850_),
    .A(_0848_),
    .B(_0849_));
 sg13g2_o21ai_1 _4966_ (.B1(_0850_),
    .Y(_0851_),
    .A1(_0833_),
    .A2(_0838_));
 sg13g2_xnor2_1 _4967_ (.Y(_0852_),
    .A(_0830_),
    .B(_0831_));
 sg13g2_a21o_1 _4968_ (.A2(_0852_),
    .A1(_0851_),
    .B1(_0832_),
    .X(_0853_));
 sg13g2_a21o_1 _4969_ (.A2(_0813_),
    .A1(_0793_),
    .B1(_0812_),
    .X(_0854_));
 sg13g2_and3_1 _4970_ (.X(_0855_),
    .A(_0815_),
    .B(_0853_),
    .C(_0854_));
 sg13g2_a21oi_1 _4971_ (.A1(_0853_),
    .A2(_0854_),
    .Y(_0856_),
    .B1(_0814_));
 sg13g2_xor2_1 _4972_ (.B(_0793_),
    .A(_0775_),
    .X(_0857_));
 sg13g2_o21ai_1 _4973_ (.B1(_0794_),
    .Y(_0858_),
    .A1(_0856_),
    .A2(_0857_));
 sg13g2_xnor2_1 _4974_ (.Y(_0859_),
    .A(_0769_),
    .B(_0773_));
 sg13g2_a21o_1 _4975_ (.A2(_0859_),
    .A1(_0858_),
    .B1(_0774_),
    .X(_0860_));
 sg13g2_xor2_1 _4976_ (.B(_0708_),
    .A(_0707_),
    .X(_0861_));
 sg13g2_and2_1 _4977_ (.A(_0772_),
    .B(_0861_),
    .X(_0862_));
 sg13g2_xnor2_1 _4978_ (.Y(_0863_),
    .A(_0772_),
    .B(_0861_));
 sg13g2_inv_1 _4979_ (.Y(_0864_),
    .A(_0863_));
 sg13g2_nand3_1 _4980_ (.B(_0860_),
    .C(_0864_),
    .A(_0711_),
    .Y(_0865_));
 sg13g2_o21ai_1 _4981_ (.B1(_0710_),
    .Y(_0866_),
    .A1(_0709_),
    .A2(_0862_));
 sg13g2_a21oi_1 _4982_ (.A1(_0865_),
    .A2(_0866_),
    .Y(_0867_),
    .B1(_0674_));
 sg13g2_a21o_2 _4983_ (.A2(_0866_),
    .A1(_0865_),
    .B1(_0674_),
    .X(_0868_));
 sg13g2_nor2b_1 _4984_ (.A(_0627_),
    .B_N(_0628_),
    .Y(_0869_));
 sg13g2_nand2b_1 _4985_ (.Y(_0870_),
    .B(_0628_),
    .A_N(_0627_));
 sg13g2_a21oi_1 _4986_ (.A1(_0673_),
    .A2(_0868_),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_nor2_1 _4987_ (.A(_0627_),
    .B(_0672_),
    .Y(_0872_));
 sg13g2_a22oi_1 _4988_ (.Y(_0873_),
    .B1(_0868_),
    .B2(_0872_),
    .A2(_0626_),
    .A1(_0593_));
 sg13g2_o21ai_1 _4989_ (.B1(_0622_),
    .Y(_0874_),
    .A1(_0595_),
    .A2(_0623_));
 sg13g2_a21oi_1 _4990_ (.A1(_0613_),
    .A2(_0619_),
    .Y(_0875_),
    .B1(_0618_));
 sg13g2_a21oi_1 _4991_ (.A1(_0612_),
    .A2(_0620_),
    .Y(_0876_),
    .B1(_0611_));
 sg13g2_a21oi_1 _4992_ (.A1(_0606_),
    .A2(_0607_),
    .Y(_0877_),
    .B1(_0609_));
 sg13g2_xor2_1 _4993_ (.B(_0414_),
    .A(_0413_),
    .X(_0878_));
 sg13g2_nor2b_1 _4994_ (.A(_0877_),
    .B_N(_0878_),
    .Y(_0879_));
 sg13g2_xnor2_1 _4995_ (.Y(_0880_),
    .A(_0877_),
    .B(_0878_));
 sg13g2_o21ai_1 _4996_ (.B1(_0175_),
    .Y(_0881_),
    .A1(_0353_),
    .A2(_0616_));
 sg13g2_a21oi_1 _4997_ (.A1(_0599_),
    .A2(_0603_),
    .Y(_0882_),
    .B1(_0602_));
 sg13g2_nor2_1 _4998_ (.A(net740),
    .B(_0882_),
    .Y(_0883_));
 sg13g2_nand2_1 _4999_ (.Y(_0884_),
    .A(net740),
    .B(_0882_));
 sg13g2_nand2b_1 _5000_ (.Y(_0885_),
    .B(_0884_),
    .A_N(_0883_));
 sg13g2_xnor2_1 _5001_ (.Y(_0886_),
    .A(_0881_),
    .B(_0885_));
 sg13g2_xnor2_1 _5002_ (.Y(_0887_),
    .A(_0880_),
    .B(_0886_));
 sg13g2_nor2_1 _5003_ (.A(_0876_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_xor2_1 _5004_ (.B(_0887_),
    .A(_0876_),
    .X(_0889_));
 sg13g2_nor2b_1 _5005_ (.A(_0875_),
    .B_N(_0889_),
    .Y(_0890_));
 sg13g2_xnor2_1 _5006_ (.Y(_0891_),
    .A(_0875_),
    .B(_0889_));
 sg13g2_and2_1 _5007_ (.A(_0874_),
    .B(_0891_),
    .X(_0892_));
 sg13g2_xnor2_1 _5008_ (.Y(_0893_),
    .A(_0874_),
    .B(_0891_));
 sg13g2_nor2_1 _5009_ (.A(_0625_),
    .B(_0893_),
    .Y(_0894_));
 sg13g2_xor2_1 _5010_ (.B(_0893_),
    .A(_0625_),
    .X(_0895_));
 sg13g2_a21o_1 _5011_ (.A2(_0884_),
    .A1(_0881_),
    .B1(_0883_),
    .X(_0896_));
 sg13g2_a21oi_1 _5012_ (.A1(_0880_),
    .A2(_0886_),
    .Y(_0897_),
    .B1(_0879_));
 sg13g2_xor2_1 _5013_ (.B(_0423_),
    .A(_0421_),
    .X(_0898_));
 sg13g2_nor2_1 _5014_ (.A(_0897_),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_xor2_1 _5015_ (.B(_0898_),
    .A(_0897_),
    .X(_0900_));
 sg13g2_xnor2_1 _5016_ (.Y(_0901_),
    .A(_0896_),
    .B(_0900_));
 sg13g2_nor2_1 _5017_ (.A(_0888_),
    .B(_0890_),
    .Y(_0902_));
 sg13g2_nor2_1 _5018_ (.A(_0901_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_xor2_1 _5019_ (.B(_0902_),
    .A(_0901_),
    .X(_0904_));
 sg13g2_nand2_1 _5020_ (.Y(_0905_),
    .A(_0892_),
    .B(_0904_));
 sg13g2_xor2_1 _5021_ (.B(_0904_),
    .A(_0892_),
    .X(_0906_));
 sg13g2_nand2_1 _5022_ (.Y(_0907_),
    .A(_0895_),
    .B(_0906_));
 sg13g2_a221oi_1 _5023_ (.B2(_0872_),
    .C1(_0907_),
    .B1(_0868_),
    .A1(_0593_),
    .Y(_0908_),
    .A2(_0626_));
 sg13g2_o21ai_1 _5024_ (.B1(_0894_),
    .Y(_0909_),
    .A1(_0892_),
    .A2(_0904_));
 sg13g2_nand2_1 _5025_ (.Y(_0910_),
    .A(_0905_),
    .B(_0909_));
 sg13g2_nor2_1 _5026_ (.A(_0908_),
    .B(_0910_),
    .Y(_0911_));
 sg13g2_xor2_1 _5027_ (.B(_0428_),
    .A(_0427_),
    .X(_0912_));
 sg13g2_a21oi_1 _5028_ (.A1(_0896_),
    .A2(_0900_),
    .Y(_0913_),
    .B1(_0899_));
 sg13g2_nor2_1 _5029_ (.A(_0912_),
    .B(_0913_),
    .Y(_0914_));
 sg13g2_xor2_1 _5030_ (.B(_0913_),
    .A(_0912_),
    .X(_0915_));
 sg13g2_nand2_1 _5031_ (.Y(_0916_),
    .A(_0903_),
    .B(_0915_));
 sg13g2_xnor2_1 _5032_ (.Y(_0917_),
    .A(_0903_),
    .B(_0915_));
 sg13g2_inv_1 _5033_ (.Y(_0918_),
    .A(_0917_));
 sg13g2_xnor2_1 _5034_ (.Y(_0919_),
    .A(_0392_),
    .B(_0430_));
 sg13g2_nor2_1 _5035_ (.A(_0914_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_xor2_1 _5036_ (.B(_0919_),
    .A(_0914_),
    .X(_0921_));
 sg13g2_nor2b_1 _5037_ (.A(_0917_),
    .B_N(_0921_),
    .Y(_0922_));
 sg13g2_o21ai_1 _5038_ (.B1(_0922_),
    .Y(_0923_),
    .A1(_0908_),
    .A2(_0910_));
 sg13g2_nor2_1 _5039_ (.A(_0916_),
    .B(_0920_),
    .Y(_0924_));
 sg13g2_a21oi_1 _5040_ (.A1(_0914_),
    .A2(_0919_),
    .Y(_0925_),
    .B1(_0924_));
 sg13g2_xor2_1 _5041_ (.B(_0431_),
    .A(_0391_),
    .X(_0926_));
 sg13g2_a21oi_1 _5042_ (.A1(_0923_),
    .A2(_0925_),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_xor2_1 _5043_ (.B(_0389_),
    .A(_0350_),
    .X(_0928_));
 sg13g2_o21ai_1 _5044_ (.B1(_0928_),
    .Y(_0929_),
    .A1(_0432_),
    .A2(_0927_));
 sg13g2_xnor2_1 _5045_ (.Y(_0930_),
    .A(_0317_),
    .B(_0347_));
 sg13g2_a21oi_1 _5046_ (.A1(_0390_),
    .A2(_0929_),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_a21oi_1 _5047_ (.A1(_0198_),
    .A2(_0322_),
    .Y(_0932_),
    .B1(_0321_));
 sg13g2_o21ai_1 _5048_ (.B1(_0339_),
    .Y(_0933_),
    .A1(_0324_),
    .A2(_0340_));
 sg13g2_a21oi_1 _5049_ (.A1(_0194_),
    .A2(_0328_),
    .Y(_0934_),
    .B1(_0327_));
 sg13g2_nor2_1 _5050_ (.A(net739),
    .B(_0934_),
    .Y(_0935_));
 sg13g2_xor2_1 _5051_ (.B(_0934_),
    .A(net739),
    .X(_0936_));
 sg13g2_nor2_1 _5052_ (.A(_0198_),
    .B(_0936_),
    .Y(_0937_));
 sg13g2_xnor2_1 _5053_ (.Y(_0938_),
    .A(_0197_),
    .B(_0936_));
 sg13g2_inv_1 _5054_ (.Y(_0939_),
    .A(_0938_));
 sg13g2_a21o_1 _5055_ (.A2(_0337_),
    .A1(_0329_),
    .B1(_0336_),
    .X(_0940_));
 sg13g2_a21oi_2 _5056_ (.B1(_0334_),
    .Y(_0941_),
    .A2(_3343_),
    .A1(net861));
 sg13g2_or2_1 _5057_ (.X(_0942_),
    .B(net816),
    .A(net820));
 sg13g2_a21oi_1 _5058_ (.A1(_3344_),
    .A2(_0942_),
    .Y(_0943_),
    .B1(net861));
 sg13g2_xor2_1 _5059_ (.B(_0943_),
    .A(_0270_),
    .X(_0944_));
 sg13g2_xnor2_1 _5060_ (.Y(_0945_),
    .A(_0941_),
    .B(_0944_));
 sg13g2_xnor2_1 _5061_ (.Y(_0946_),
    .A(_0329_),
    .B(_0945_));
 sg13g2_nand2_1 _5062_ (.Y(_0947_),
    .A(_0940_),
    .B(_0946_));
 sg13g2_xnor2_1 _5063_ (.Y(_0948_),
    .A(_0940_),
    .B(_0946_));
 sg13g2_xor2_1 _5064_ (.B(_0948_),
    .A(_0938_),
    .X(_0949_));
 sg13g2_inv_1 _5065_ (.Y(_0950_),
    .A(_0949_));
 sg13g2_xnor2_1 _5066_ (.Y(_0951_),
    .A(_0933_),
    .B(_0950_));
 sg13g2_nor2_1 _5067_ (.A(_0932_),
    .B(_0951_),
    .Y(_0952_));
 sg13g2_xor2_1 _5068_ (.B(_0951_),
    .A(_0932_),
    .X(_0953_));
 sg13g2_o21ai_1 _5069_ (.B1(_0342_),
    .Y(_0954_),
    .A1(_0318_),
    .A2(_0343_));
 sg13g2_xor2_1 _5070_ (.B(_0954_),
    .A(_0953_),
    .X(_0955_));
 sg13g2_nand2_1 _5071_ (.Y(_0956_),
    .A(_0346_),
    .B(_0955_));
 sg13g2_xor2_1 _5072_ (.B(_0955_),
    .A(_0346_),
    .X(_0957_));
 sg13g2_o21ai_1 _5073_ (.B1(_0957_),
    .Y(_0958_),
    .A1(_0348_),
    .A2(_0931_));
 sg13g2_or3_1 _5074_ (.A(_0348_),
    .B(_0931_),
    .C(_0957_),
    .X(_0959_));
 sg13g2_and2_1 _5075_ (.A(_0958_),
    .B(_0959_),
    .X(\i_mandel.l_sq.genblk2[17].state.D ));
 sg13g2_and2_1 _5076_ (.A(\i_mandel.l_sq.genblk2[17].state.Q ),
    .B(\i_mandel.l_sq.genblk2[17].state.D ),
    .X(_0960_));
 sg13g2_xor2_1 _5077_ (.B(\i_mandel.l_sq.genblk2[17].state.D ),
    .A(\i_mandel.l_sq.genblk2[17].state.Q ),
    .X(_0961_));
 sg13g2_nand3_1 _5078_ (.B(_0929_),
    .C(_0930_),
    .A(_0390_),
    .Y(_0962_));
 sg13g2_nor2b_1 _5079_ (.A(_0931_),
    .B_N(_0962_),
    .Y(\i_mandel.l_sq.genblk2[16].state.D ));
 sg13g2_nand2_1 _5080_ (.Y(_0963_),
    .A(\i_mandel.l_sq.genblk2[16].state.Q ),
    .B(\i_mandel.l_sq.genblk2[16].state.D ));
 sg13g2_a21oi_1 _5081_ (.A1(_0873_),
    .A2(_0895_),
    .Y(_0964_),
    .B1(_0894_));
 sg13g2_xor2_1 _5082_ (.B(_0964_),
    .A(_0906_),
    .X(_0965_));
 sg13g2_inv_1 _5083_ (.Y(\i_mandel.l_sq.genblk2[11].state.D ),
    .A(_0965_));
 sg13g2_nor2_1 _5084_ (.A(\i_mandel.l_sq.genblk2[11].state.Q ),
    .B(\i_mandel.l_sq.genblk2[11].state.D ),
    .Y(_0966_));
 sg13g2_xor2_1 _5085_ (.B(_0895_),
    .A(_0873_),
    .X(\i_mandel.l_sq.genblk2[10].state.D ));
 sg13g2_xnor2_1 _5086_ (.Y(_0967_),
    .A(\i_mandel.l_sq.genblk2[10].state.Q ),
    .B(\i_mandel.l_sq.genblk2[10].state.D ));
 sg13g2_nor3_1 _5087_ (.A(_0672_),
    .B(_0867_),
    .C(_0869_),
    .Y(_0968_));
 sg13g2_a21oi_1 _5088_ (.A1(_0673_),
    .A2(_0868_),
    .Y(_0969_),
    .B1(_0869_));
 sg13g2_nor3_2 _5089_ (.A(_0672_),
    .B(_0867_),
    .C(_0870_),
    .Y(_0970_));
 sg13g2_nor2_1 _5090_ (.A(_0969_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_inv_1 _5091_ (.Y(\i_mandel.l_sq.genblk2[9].state.D ),
    .A(_0971_));
 sg13g2_nor3_2 _5092_ (.A(_3091_),
    .B(_0871_),
    .C(_0968_),
    .Y(_0972_));
 sg13g2_o21ai_1 _5093_ (.B1(\i_mandel.l_sq.genblk2[9].state.Q ),
    .Y(_0973_),
    .A1(_0969_),
    .A2(_0970_));
 sg13g2_a21oi_1 _5094_ (.A1(_0860_),
    .A2(_0864_),
    .Y(_0974_),
    .B1(_0862_));
 sg13g2_xor2_1 _5095_ (.B(_0974_),
    .A(_0711_),
    .X(_0975_));
 sg13g2_inv_1 _5096_ (.Y(\i_mandel.l_sq.genblk2[7].state.D ),
    .A(_0975_));
 sg13g2_nor2_1 _5097_ (.A(_3092_),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_xnor2_1 _5098_ (.Y(\i_mandel.l_sq.genblk2[6].state.D ),
    .A(_0860_),
    .B(_0863_));
 sg13g2_and2_1 _5099_ (.A(\i_mandel.l_sq.genblk2[6].state.Q ),
    .B(\i_mandel.l_sq.genblk2[6].state.D ),
    .X(_0977_));
 sg13g2_xor2_1 _5100_ (.B(_0859_),
    .A(_0858_),
    .X(\i_mandel.l_sq.genblk2[5].state.D ));
 sg13g2_nand2_1 _5101_ (.Y(_0978_),
    .A(\i_mandel.l_sq.genblk2[5].state.Q ),
    .B(\i_mandel.l_sq.genblk2[5].state.D ));
 sg13g2_xnor2_1 _5102_ (.Y(_0979_),
    .A(\i_mandel.l_sq.genblk2[5].state.Q ),
    .B(\i_mandel.l_sq.genblk2[5].state.D ));
 sg13g2_xor2_1 _5103_ (.B(_0857_),
    .A(_0856_),
    .X(\i_mandel.l_sq.genblk2[4].state.D ));
 sg13g2_and2_1 _5104_ (.A(\i_mandel.l_sq.genblk2[4].state.Q ),
    .B(\i_mandel.l_sq.genblk2[4].state.D ),
    .X(_0980_));
 sg13g2_inv_1 _5105_ (.Y(_0981_),
    .A(_0980_));
 sg13g2_o21ai_1 _5106_ (.B1(_0978_),
    .Y(_0982_),
    .A1(_0979_),
    .A2(_0981_));
 sg13g2_xor2_1 _5107_ (.B(\i_mandel.l_sq.genblk2[6].state.D ),
    .A(\i_mandel.l_sq.genblk2[6].state.Q ),
    .X(_0983_));
 sg13g2_a21o_1 _5108_ (.A2(_0983_),
    .A1(_0982_),
    .B1(_0977_),
    .X(_0984_));
 sg13g2_xnor2_1 _5109_ (.Y(_0985_),
    .A(\i_mandel.l_sq.genblk2[7].state.Q ),
    .B(_0975_));
 sg13g2_a21oi_1 _5110_ (.A1(_0984_),
    .A2(_0985_),
    .Y(_0986_),
    .B1(_0976_));
 sg13g2_nand3_1 _5111_ (.B(_0865_),
    .C(_0866_),
    .A(_0674_),
    .Y(_0987_));
 sg13g2_and2_2 _5112_ (.A(_0868_),
    .B(_0987_),
    .X(\i_mandel.l_sq.genblk2[8].state.D ));
 sg13g2_and2_1 _5113_ (.A(\i_mandel.l_sq.genblk2[8].state.Q ),
    .B(\i_mandel.l_sq.genblk2[8].state.D ),
    .X(_0988_));
 sg13g2_a221oi_1 _5114_ (.B2(\i_mandel.l_sq.genblk2[8].state.Q ),
    .C1(_0976_),
    .B1(\i_mandel.l_sq.genblk2[8].state.D ),
    .A1(_0984_),
    .Y(_0989_),
    .A2(_0985_));
 sg13g2_nor3_1 _5115_ (.A(\i_mandel.l_sq.genblk2[9].state.Q ),
    .B(_0969_),
    .C(_0970_),
    .Y(_0990_));
 sg13g2_nor2_1 _5116_ (.A(\i_mandel.l_sq.genblk2[8].state.Q ),
    .B(\i_mandel.l_sq.genblk2[8].state.D ),
    .Y(_0991_));
 sg13g2_nor4_1 _5117_ (.A(_0972_),
    .B(_0988_),
    .C(_0990_),
    .D(_0991_),
    .Y(_0992_));
 sg13g2_or4_2 _5118_ (.A(_0972_),
    .B(_0989_),
    .C(_0990_),
    .D(_0991_),
    .X(_0993_));
 sg13g2_a21oi_1 _5119_ (.A1(_0973_),
    .A2(_0993_),
    .Y(_0994_),
    .B1(_0967_));
 sg13g2_a21o_1 _5120_ (.A2(_0993_),
    .A1(_0973_),
    .B1(_0967_),
    .X(_0995_));
 sg13g2_a21o_1 _5121_ (.A2(\i_mandel.l_sq.genblk2[10].state.D ),
    .A1(\i_mandel.l_sq.genblk2[10].state.Q ),
    .B1(_0994_),
    .X(_0996_));
 sg13g2_a22oi_1 _5122_ (.Y(_0997_),
    .B1(\i_mandel.l_sq.genblk2[10].state.D ),
    .B2(\i_mandel.l_sq.genblk2[10].state.Q ),
    .A2(\i_mandel.l_sq.genblk2[11].state.D ),
    .A1(\i_mandel.l_sq.genblk2[11].state.Q ));
 sg13g2_a21o_1 _5123_ (.A2(_0997_),
    .A1(_0995_),
    .B1(_0966_),
    .X(_0998_));
 sg13g2_o21ai_1 _5124_ (.B1(_0918_),
    .Y(_0999_),
    .A1(_0908_),
    .A2(_0910_));
 sg13g2_a21o_1 _5125_ (.A2(_0999_),
    .A1(_0916_),
    .B1(_0921_),
    .X(_1000_));
 sg13g2_nand3_1 _5126_ (.B(_0921_),
    .C(_0999_),
    .A(_0916_),
    .Y(_1001_));
 sg13g2_and2_1 _5127_ (.A(_1000_),
    .B(_1001_),
    .X(_1002_));
 sg13g2_inv_1 _5128_ (.Y(\i_mandel.l_sq.genblk2[13].state.D ),
    .A(_1002_));
 sg13g2_a21oi_1 _5129_ (.A1(_1000_),
    .A2(_1001_),
    .Y(_1003_),
    .B1(_3090_));
 sg13g2_nand3_1 _5130_ (.B(_1000_),
    .C(_1001_),
    .A(_3090_),
    .Y(_1004_));
 sg13g2_nand2b_1 _5131_ (.Y(_1005_),
    .B(_1004_),
    .A_N(_1003_));
 sg13g2_xnor2_1 _5132_ (.Y(\i_mandel.l_sq.genblk2[12].state.D ),
    .A(_0911_),
    .B(_0918_));
 sg13g2_and2_1 _5133_ (.A(\i_mandel.l_sq.genblk2[12].state.Q ),
    .B(\i_mandel.l_sq.genblk2[12].state.D ),
    .X(_1006_));
 sg13g2_nor2_1 _5134_ (.A(\i_mandel.l_sq.genblk2[12].state.Q ),
    .B(\i_mandel.l_sq.genblk2[12].state.D ),
    .Y(_1007_));
 sg13g2_xor2_1 _5135_ (.B(\i_mandel.l_sq.genblk2[12].state.D ),
    .A(\i_mandel.l_sq.genblk2[12].state.Q ),
    .X(_1008_));
 sg13g2_nand3b_1 _5136_ (.B(_1004_),
    .C(_1008_),
    .Y(_1009_),
    .A_N(_1003_));
 sg13g2_nor2_1 _5137_ (.A(_0998_),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_a21oi_1 _5138_ (.A1(_1004_),
    .A2(_1006_),
    .Y(_1011_),
    .B1(_1003_));
 sg13g2_o21ai_1 _5139_ (.B1(_1011_),
    .Y(_1012_),
    .A1(_0998_),
    .A2(_1009_));
 sg13g2_or3_1 _5140_ (.A(_0432_),
    .B(_0927_),
    .C(_0928_),
    .X(_1013_));
 sg13g2_and2_2 _5141_ (.A(_0929_),
    .B(_1013_),
    .X(\i_mandel.l_sq.genblk2[15].state.D ));
 sg13g2_a21oi_1 _5142_ (.A1(_0929_),
    .A2(_1013_),
    .Y(_1014_),
    .B1(\i_mandel.l_sq.genblk2[15].state.Q ));
 sg13g2_and3_1 _5143_ (.X(_1015_),
    .A(\i_mandel.l_sq.genblk2[15].state.Q ),
    .B(_0929_),
    .C(_1013_));
 sg13g2_or2_1 _5144_ (.X(_1016_),
    .B(_1015_),
    .A(_1014_));
 sg13g2_nand3_1 _5145_ (.B(_0925_),
    .C(_0926_),
    .A(_0923_),
    .Y(_1017_));
 sg13g2_nand2b_2 _5146_ (.Y(_1018_),
    .B(_1017_),
    .A_N(_0927_));
 sg13g2_inv_1 _5147_ (.Y(\i_mandel.l_sq.genblk2[14].state.D ),
    .A(_1018_));
 sg13g2_nor2_1 _5148_ (.A(_3089_),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_and2_1 _5149_ (.A(_3089_),
    .B(_1018_),
    .X(_1020_));
 sg13g2_nor2_1 _5150_ (.A(_1019_),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_nor4_1 _5151_ (.A(_1014_),
    .B(_1015_),
    .C(_1019_),
    .D(_1020_),
    .Y(_1022_));
 sg13g2_nor2b_1 _5152_ (.A(_1014_),
    .B_N(_1019_),
    .Y(_1023_));
 sg13g2_a221oi_1 _5153_ (.B2(_1012_),
    .C1(_1023_),
    .B1(_1022_),
    .A1(\i_mandel.l_sq.genblk2[15].state.Q ),
    .Y(_1024_),
    .A2(\i_mandel.l_sq.genblk2[15].state.D ));
 sg13g2_xnor2_1 _5154_ (.Y(_1025_),
    .A(\i_mandel.l_sq.genblk2[16].state.Q ),
    .B(\i_mandel.l_sq.genblk2[16].state.D ));
 sg13g2_o21ai_1 _5155_ (.B1(_0963_),
    .Y(_1026_),
    .A1(_1024_),
    .A2(_1025_));
 sg13g2_a21oi_1 _5156_ (.A1(_0961_),
    .A2(_1026_),
    .Y(_1027_),
    .B1(_0960_));
 sg13g2_nand2_1 _5157_ (.Y(_1028_),
    .A(_0956_),
    .B(_0958_));
 sg13g2_a21oi_1 _5158_ (.A1(_0933_),
    .A2(_0950_),
    .Y(_1029_),
    .B1(_0952_));
 sg13g2_o21ai_1 _5159_ (.B1(_0947_),
    .Y(_1030_),
    .A1(_0939_),
    .A2(_0948_));
 sg13g2_nor2_1 _5160_ (.A(net861),
    .B(_0942_),
    .Y(_1031_));
 sg13g2_nand2_1 _5161_ (.Y(_1032_),
    .A(net830),
    .B(_3343_));
 sg13g2_a21oi_1 _5162_ (.A1(_0270_),
    .A2(_1032_),
    .Y(_1033_),
    .B1(_1031_));
 sg13g2_a21oi_1 _5163_ (.A1(_0941_),
    .A2(_0944_),
    .Y(_1034_),
    .B1(_1033_));
 sg13g2_o21ai_1 _5164_ (.B1(_1033_),
    .Y(_1035_),
    .A1(_0941_),
    .A2(_0944_));
 sg13g2_nand2b_1 _5165_ (.Y(_1036_),
    .B(_1035_),
    .A_N(_0329_));
 sg13g2_nand2b_1 _5166_ (.Y(_1037_),
    .B(_1036_),
    .A_N(_1034_));
 sg13g2_xor2_1 _5167_ (.B(_1037_),
    .A(_0935_),
    .X(_1038_));
 sg13g2_xnor2_1 _5168_ (.Y(_1039_),
    .A(_0937_),
    .B(_1038_));
 sg13g2_xor2_1 _5169_ (.B(_1039_),
    .A(_1030_),
    .X(_1040_));
 sg13g2_a22oi_1 _5170_ (.Y(_1041_),
    .B1(_1029_),
    .B2(_1040_),
    .A2(_0954_),
    .A1(_0953_));
 sg13g2_o21ai_1 _5171_ (.B1(_1041_),
    .Y(_1042_),
    .A1(_1029_),
    .A2(_1040_));
 sg13g2_xnor2_1 _5172_ (.Y(\i_mandel.l_sq.genblk2[18].state.D ),
    .A(_1028_),
    .B(_1042_));
 sg13g2_xor2_1 _5173_ (.B(\i_mandel.l_sq.genblk2[18].state.D ),
    .A(\i_mandel.l_sq.genblk2[18].state.Q ),
    .X(_1043_));
 sg13g2_xnor2_1 _5174_ (.Y(_1044_),
    .A(_1027_),
    .B(_1043_));
 sg13g2_xnor2_1 _5175_ (.Y(_1045_),
    .A(_0961_),
    .B(_1026_));
 sg13g2_xnor2_1 _5176_ (.Y(_1046_),
    .A(_1024_),
    .B(_1025_));
 sg13g2_a21oi_1 _5177_ (.A1(_1012_),
    .A2(_1021_),
    .Y(_1047_),
    .B1(_1019_));
 sg13g2_xnor2_1 _5178_ (.Y(_1048_),
    .A(_1012_),
    .B(_1021_));
 sg13g2_mux2_1 _5179_ (.A0(_1006_),
    .A1(_1007_),
    .S(_1005_),
    .X(_1049_));
 sg13g2_a21o_1 _5180_ (.A2(_1049_),
    .A1(_0998_),
    .B1(_1010_),
    .X(_1050_));
 sg13g2_xnor2_1 _5181_ (.Y(_1051_),
    .A(\i_mandel.l_sq.genblk2[11].state.Q ),
    .B(\i_mandel.l_sq.genblk2[11].state.D ));
 sg13g2_nand2_1 _5182_ (.Y(_1052_),
    .A(_0996_),
    .B(_1051_));
 sg13g2_nor2_1 _5183_ (.A(_0996_),
    .B(_1051_),
    .Y(_1053_));
 sg13g2_and3_1 _5184_ (.X(_1054_),
    .A(_0967_),
    .B(_0973_),
    .C(_0993_));
 sg13g2_nor2_1 _5185_ (.A(_0986_),
    .B(_0992_),
    .Y(_1055_));
 sg13g2_xnor2_1 _5186_ (.Y(_1056_),
    .A(_0984_),
    .B(_0985_));
 sg13g2_xnor2_1 _5187_ (.Y(_1057_),
    .A(_0982_),
    .B(_0983_));
 sg13g2_nor2_1 _5188_ (.A(\i_mandel.l_sq.genblk2[4].state.Q ),
    .B(\i_mandel.l_sq.genblk2[4].state.D ),
    .Y(_1058_));
 sg13g2_nand2_1 _5189_ (.Y(_1059_),
    .A(_0979_),
    .B(_1058_));
 sg13g2_o21ai_1 _5190_ (.B1(_1059_),
    .Y(_1060_),
    .A1(_0979_),
    .A2(_0981_));
 sg13g2_nand3_1 _5191_ (.B(_1057_),
    .C(_1060_),
    .A(_1056_),
    .Y(_1061_));
 sg13g2_nor2_1 _5192_ (.A(_1055_),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_o21ai_1 _5193_ (.B1(_0991_),
    .Y(_1063_),
    .A1(_0972_),
    .A2(_0990_));
 sg13g2_and2_1 _5194_ (.A(_0993_),
    .B(_1063_),
    .X(_1064_));
 sg13g2_o21ai_1 _5195_ (.B1(_1062_),
    .Y(_1065_),
    .A1(_0994_),
    .A2(_1054_));
 sg13g2_nor3_1 _5196_ (.A(_1053_),
    .B(_1064_),
    .C(_1065_),
    .Y(_1066_));
 sg13g2_nand4_1 _5197_ (.B(_1050_),
    .C(_1052_),
    .A(_1048_),
    .Y(_1067_),
    .D(_1066_));
 sg13g2_xnor2_1 _5198_ (.Y(_1068_),
    .A(_1016_),
    .B(_1047_));
 sg13g2_nor2b_1 _5199_ (.A(_1067_),
    .B_N(_1068_),
    .Y(_1069_));
 sg13g2_o21ai_1 _5200_ (.B1(_1045_),
    .Y(_1070_),
    .A1(_1046_),
    .A2(_1069_));
 sg13g2_nor2_1 _5201_ (.A(_1044_),
    .B(_1070_),
    .Y(_1071_));
 sg13g2_nor3_2 _5202_ (.A(_3094_),
    .B(_1044_),
    .C(_1070_),
    .Y(_1072_));
 sg13g2_nor4_2 _5203_ (.A(_3094_),
    .B(_0013_),
    .C(_1044_),
    .Y(_1073_),
    .D(_1070_));
 sg13g2_xnor2_1 _5204_ (.Y(_1074_),
    .A(net212),
    .B(_1073_));
 sg13g2_nand2_1 _5205_ (.Y(_1075_),
    .A(net754),
    .B(_1074_));
 sg13g2_nor2_1 _5206_ (.A(net353),
    .B(net754),
    .Y(_1076_));
 sg13g2_nand2b_1 _5207_ (.Y(_1077_),
    .B(_3270_),
    .A_N(\last_iter[2] ));
 sg13g2_a21o_2 _5208_ (.A2(_1074_),
    .A1(net754),
    .B1(_1076_),
    .X(_1078_));
 sg13g2_inv_1 _5209_ (.Y(_0168_),
    .A(_1078_));
 sg13g2_xnor2_1 _5210_ (.Y(_1079_),
    .A(net205),
    .B(_1071_));
 sg13g2_nor2_1 _5211_ (.A(net357),
    .B(_3269_),
    .Y(_1080_));
 sg13g2_a21o_1 _5212_ (.A2(_1079_),
    .A1(_3269_),
    .B1(_1080_),
    .X(_1081_));
 sg13g2_inv_2 _5213_ (.Y(_0166_),
    .A(_1081_));
 sg13g2_a21o_1 _5214_ (.A2(_1073_),
    .A1(\iter[2] ),
    .B1(_3137_),
    .X(_1082_));
 sg13g2_nand3_1 _5215_ (.B(_3137_),
    .C(_1073_),
    .A(\iter[2] ),
    .Y(_1083_));
 sg13g2_and2_1 _5216_ (.A(_1082_),
    .B(_1083_),
    .X(_1084_));
 sg13g2_and3_1 _5217_ (.X(_1085_),
    .A(net754),
    .B(_1082_),
    .C(_1083_));
 sg13g2_nand3_1 _5218_ (.B(_1082_),
    .C(_1083_),
    .A(_3269_),
    .Y(_1086_));
 sg13g2_nand2_1 _5219_ (.Y(_1087_),
    .A(_3138_),
    .B(_3270_));
 sg13g2_and2_2 _5220_ (.A(_1086_),
    .B(_1087_),
    .X(_0169_));
 sg13g2_a221oi_1 _5221_ (.B2(_1087_),
    .C1(_0166_),
    .B1(_1086_),
    .A1(_1075_),
    .Y(_1088_),
    .A2(_1077_));
 sg13g2_xnor2_1 _5222_ (.Y(_1089_),
    .A(_0013_),
    .B(_1072_));
 sg13g2_mux2_1 _5223_ (.A0(_3146_),
    .A1(_1089_),
    .S(net754),
    .X(_1090_));
 sg13g2_nand2_1 _5224_ (.Y(_1091_),
    .A(_0168_),
    .B(_1090_));
 sg13g2_a221oi_1 _5225_ (.B2(_1081_),
    .C1(_1085_),
    .B1(_1078_),
    .A1(_3138_),
    .Y(_1092_),
    .A2(_3270_));
 sg13g2_a21o_1 _5226_ (.A2(_1092_),
    .A1(_1091_),
    .B1(_1088_),
    .X(_0000_));
 sg13g2_nor2_1 _5227_ (.A(_0168_),
    .B(_1090_),
    .Y(_1093_));
 sg13g2_mux2_1 _5228_ (.A0(net299),
    .A1(_1074_),
    .S(net754),
    .X(_1094_));
 sg13g2_xnor2_1 _5229_ (.Y(_1095_),
    .A(_1090_),
    .B(_1094_));
 sg13g2_mux2_1 _5230_ (.A0(_1093_),
    .A1(_1095_),
    .S(_0169_),
    .X(_0001_));
 sg13g2_nor2_1 _5231_ (.A(net342),
    .B(net754),
    .Y(_1096_));
 sg13g2_xnor2_1 _5232_ (.Y(_1097_),
    .A(net192),
    .B(_1072_));
 sg13g2_a21o_2 _5233_ (.A2(_1097_),
    .A1(net754),
    .B1(_1096_),
    .X(_1098_));
 sg13g2_inv_1 _5234_ (.Y(_0167_),
    .A(_1098_));
 sg13g2_a221oi_1 _5235_ (.B2(_0166_),
    .C1(_1078_),
    .B1(_1098_),
    .A1(_1086_),
    .Y(_1099_),
    .A2(_1087_));
 sg13g2_a21oi_1 _5236_ (.A1(_1081_),
    .A2(_1098_),
    .Y(_1100_),
    .B1(_1078_));
 sg13g2_o21ai_1 _5237_ (.B1(_0168_),
    .Y(_1101_),
    .A1(_0166_),
    .A2(_0167_));
 sg13g2_a221oi_1 _5238_ (.B2(_0167_),
    .C1(_1085_),
    .B1(_0166_),
    .A1(_3138_),
    .Y(_1102_),
    .A2(_3270_));
 sg13g2_a21o_1 _5239_ (.A2(_1102_),
    .A1(_1101_),
    .B1(_1099_),
    .X(_0002_));
 sg13g2_mux2_1 _5240_ (.A0(_1100_),
    .A1(_1094_),
    .S(_0169_),
    .X(_0003_));
 sg13g2_or2_1 _5241_ (.X(_1103_),
    .B(_3257_),
    .A(net366));
 sg13g2_nor2_1 _5242_ (.A(_3253_),
    .B(_1103_),
    .Y(_1104_));
 sg13g2_nor2_1 _5243_ (.A(\i_vga.timing_hor.counter[3] ),
    .B(_3253_),
    .Y(_1105_));
 sg13g2_nor2_1 _5244_ (.A(net229),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_nand2_1 _5245_ (.Y(_1107_),
    .A(net941),
    .B(_1106_));
 sg13g2_nor2_1 _5246_ (.A(_1104_),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_o21ai_1 _5247_ (.B1(_3254_),
    .Y(_1109_),
    .A1(net254),
    .A2(_1108_));
 sg13g2_o21ai_1 _5248_ (.B1(_1109_),
    .Y(_1110_),
    .A1(_3256_),
    .A2(_1103_));
 sg13g2_nor4_1 _5249_ (.A(net941),
    .B(net264),
    .C(_1104_),
    .D(_1106_),
    .Y(_1111_));
 sg13g2_o21ai_1 _5250_ (.B1(_1110_),
    .Y(_0004_),
    .A1(_3252_),
    .A2(_1111_));
 sg13g2_xnor2_1 _5251_ (.Y(\i_mandel.l_sq.genblk2[0].state.D ),
    .A(_0845_),
    .B(_0847_));
 sg13g2_xor2_1 _5252_ (.B(_0849_),
    .A(_0848_),
    .X(\i_mandel.l_sq.genblk2[1].state.D ));
 sg13g2_xor2_1 _5253_ (.B(_0852_),
    .A(_0851_),
    .X(\i_mandel.l_sq.genblk2[2].state.D ));
 sg13g2_a21oi_2 _5254_ (.B1(_0853_),
    .Y(_1112_),
    .A2(_0854_),
    .A1(_0815_));
 sg13g2_nor2_1 _5255_ (.A(_0855_),
    .B(_1112_),
    .Y(\i_mandel.l_sq.genblk2[3].state.D ));
 sg13g2_nor2b_1 _5256_ (.A(net1),
    .B_N(net2),
    .Y(_1113_));
 sg13g2_nand2_1 _5257_ (.Y(_1114_),
    .A(net3),
    .B(_1113_));
 sg13g2_a21oi_1 _5258_ (.A1(net965),
    .A2(_1114_),
    .Y(\i_coord.l_xir.gated_clk ),
    .B1(clknet_1_1__leaf_clk));
 sg13g2_nand2b_1 _5259_ (.Y(_1115_),
    .B(net1),
    .A_N(net2));
 sg13g2_or2_1 _5260_ (.X(_1116_),
    .B(_1115_),
    .A(_3093_));
 sg13g2_a21oi_1 _5261_ (.A1(net965),
    .A2(_1116_),
    .Y(\i_coord.l_yip.gated_clk ),
    .B1(clknet_1_1__leaf_clk));
 sg13g2_nor2_1 _5262_ (.A(net1),
    .B(net2),
    .Y(_1117_));
 sg13g2_nand2_1 _5263_ (.Y(_1118_),
    .A(net965),
    .B(_0027_));
 sg13g2_a21oi_1 _5264_ (.A1(net3),
    .A2(_1117_),
    .Y(_1119_),
    .B1(_1118_));
 sg13g2_nor2_1 _5265_ (.A(clknet_1_0__leaf_clk),
    .B(_1119_),
    .Y(\i_coord.l_xip.gated_clk ));
 sg13g2_a21oi_1 _5266_ (.A1(_3093_),
    .A2(_1113_),
    .Y(_1120_),
    .B1(_1118_));
 sg13g2_nor2_1 _5267_ (.A(clknet_1_1__leaf_clk),
    .B(_1120_),
    .Y(\i_coord.l_yt.gated_clk ));
 sg13g2_o21ai_1 _5268_ (.B1(net965),
    .Y(_1121_),
    .A1(net3),
    .A2(_1115_));
 sg13g2_nor2b_1 _5269_ (.A(clknet_1_0__leaf_clk),
    .B_N(_1121_),
    .Y(\i_coord.l_xl.gated_clk ));
 sg13g2_nor2_1 _5270_ (.A(net949),
    .B(clknet_1_0__leaf_clk),
    .Y(\i_mandel.i_xy.hc.gated_clk ));
 sg13g2_nor2_1 _5271_ (.A(net953),
    .B(_0012_),
    .Y(_1122_));
 sg13g2_nand2b_1 _5272_ (.Y(_1123_),
    .B(net953),
    .A_N(_0019_));
 sg13g2_nor2b_2 _5273_ (.A(_1122_),
    .B_N(_1123_),
    .Y(_1124_));
 sg13g2_nand2b_2 _5274_ (.Y(_1125_),
    .B(_1123_),
    .A_N(_1122_));
 sg13g2_nor2_1 _5275_ (.A(_3421_),
    .B(_1124_),
    .Y(_1126_));
 sg13g2_nor2_1 _5276_ (.A(net952),
    .B(_0011_),
    .Y(_1127_));
 sg13g2_nand2b_1 _5277_ (.Y(_1128_),
    .B(net952),
    .A_N(_0018_));
 sg13g2_nor2b_2 _5278_ (.A(_1127_),
    .B_N(_1128_),
    .Y(_1129_));
 sg13g2_nand2b_2 _5279_ (.Y(_1130_),
    .B(_1128_),
    .A_N(_1127_));
 sg13g2_nor2_1 _5280_ (.A(_3440_),
    .B(_1129_),
    .Y(_1131_));
 sg13g2_and2_1 _5281_ (.A(_1126_),
    .B(_1131_),
    .X(_1132_));
 sg13g2_xor2_1 _5282_ (.B(_1131_),
    .A(_1126_),
    .X(\i_mandel.i_xy.hc.genblk2[0].state.D ));
 sg13g2_nand2_1 _5283_ (.Y(_1133_),
    .A(_3403_),
    .B(_1125_));
 sg13g2_nor2_1 _5284_ (.A(net952),
    .B(_0010_),
    .Y(_1134_));
 sg13g2_nand2b_1 _5285_ (.Y(_1135_),
    .B(net952),
    .A_N(_0017_));
 sg13g2_nor2b_1 _5286_ (.A(_1134_),
    .B_N(_1135_),
    .Y(_1136_));
 sg13g2_nand2b_1 _5287_ (.Y(_1137_),
    .B(_1135_),
    .A_N(_1134_));
 sg13g2_nor2_1 _5288_ (.A(_3421_),
    .B(_1129_),
    .Y(_1138_));
 sg13g2_nand3_1 _5289_ (.B(_1131_),
    .C(net812),
    .A(_3420_),
    .Y(_1139_));
 sg13g2_nor2_1 _5290_ (.A(_3440_),
    .B(net813),
    .Y(_1140_));
 sg13g2_o21ai_1 _5291_ (.B1(_1139_),
    .Y(_1141_),
    .A1(_1138_),
    .A2(_1140_));
 sg13g2_or2_1 _5292_ (.X(_1142_),
    .B(_1141_),
    .A(_1133_));
 sg13g2_xor2_1 _5293_ (.B(_1141_),
    .A(_1133_),
    .X(_1143_));
 sg13g2_and2_1 _5294_ (.A(_1132_),
    .B(_1143_),
    .X(_1144_));
 sg13g2_xor2_1 _5295_ (.B(_1143_),
    .A(_1132_),
    .X(\i_mandel.i_xy.hc.genblk2[1].state.D ));
 sg13g2_nor2_1 _5296_ (.A(_0009_),
    .B(net952),
    .Y(_1145_));
 sg13g2_nand2b_1 _5297_ (.Y(_1146_),
    .B(net952),
    .A_N(_0016_));
 sg13g2_nor2b_1 _5298_ (.A(_1145_),
    .B_N(_1146_),
    .Y(_1147_));
 sg13g2_nand2b_1 _5299_ (.Y(_1148_),
    .B(_1146_),
    .A_N(_1145_));
 sg13g2_nor4_1 _5300_ (.A(_3421_),
    .B(_3440_),
    .C(net813),
    .D(_1147_),
    .Y(_1149_));
 sg13g2_nand3_1 _5301_ (.B(_1140_),
    .C(net810),
    .A(net809),
    .Y(_1150_));
 sg13g2_nand2_1 _5302_ (.Y(_1151_),
    .A(_3441_),
    .B(net810));
 sg13g2_o21ai_1 _5303_ (.B1(_1151_),
    .Y(_1152_),
    .A1(_3421_),
    .A2(net814));
 sg13g2_and4_2 _5304_ (.A(_3403_),
    .B(_1130_),
    .C(_1150_),
    .D(_1152_),
    .X(_1153_));
 sg13g2_a22oi_1 _5305_ (.Y(_1154_),
    .B1(_1150_),
    .B2(_1152_),
    .A2(_1130_),
    .A1(_3403_));
 sg13g2_nor3_1 _5306_ (.A(_1139_),
    .B(_1153_),
    .C(_1154_),
    .Y(_1155_));
 sg13g2_or3_1 _5307_ (.A(_1139_),
    .B(_1153_),
    .C(_1154_),
    .X(_1156_));
 sg13g2_o21ai_1 _5308_ (.B1(_1139_),
    .Y(_1157_),
    .A1(_1153_),
    .A2(_1154_));
 sg13g2_and4_1 _5309_ (.A(_3382_),
    .B(_1125_),
    .C(_1156_),
    .D(_1157_),
    .X(_1158_));
 sg13g2_a22oi_1 _5310_ (.Y(_1159_),
    .B1(_1156_),
    .B2(_1157_),
    .A2(_1125_),
    .A1(_3382_));
 sg13g2_nor3_1 _5311_ (.A(_1142_),
    .B(_1158_),
    .C(_1159_),
    .Y(_1160_));
 sg13g2_o21ai_1 _5312_ (.B1(_1142_),
    .Y(_1161_),
    .A1(_1158_),
    .A2(_1159_));
 sg13g2_nand2b_1 _5313_ (.Y(_1162_),
    .B(_1161_),
    .A_N(_1160_));
 sg13g2_xnor2_1 _5314_ (.Y(\i_mandel.i_xy.hc.genblk2[2].state.D ),
    .A(_1144_),
    .B(_1162_));
 sg13g2_a21oi_1 _5315_ (.A1(_1144_),
    .A2(_1161_),
    .Y(_1163_),
    .B1(_1160_));
 sg13g2_or2_1 _5316_ (.X(_1164_),
    .B(_1158_),
    .A(_1155_));
 sg13g2_nor2_1 _5317_ (.A(_3318_),
    .B(_1124_),
    .Y(_1165_));
 sg13g2_nand2_1 _5318_ (.Y(_1166_),
    .A(_3382_),
    .B(_1130_));
 sg13g2_nand2_1 _5319_ (.Y(_1167_),
    .A(_3403_),
    .B(net810));
 sg13g2_nor3_1 _5320_ (.A(_3421_),
    .B(net813),
    .C(_1167_),
    .Y(_1168_));
 sg13g2_nand4_1 _5321_ (.B(net809),
    .C(net812),
    .A(_3403_),
    .Y(_1169_),
    .D(net810));
 sg13g2_a221oi_1 _5322_ (.B2(_3298_),
    .C1(net814),
    .B1(_3402_),
    .A1(_3275_),
    .Y(_1170_),
    .A2(net823));
 sg13g2_a21o_1 _5323_ (.A2(net810),
    .A1(net809),
    .B1(_1170_),
    .X(_1171_));
 sg13g2_and3_1 _5324_ (.X(_1172_),
    .A(_1149_),
    .B(_1169_),
    .C(_1171_));
 sg13g2_a21oi_1 _5325_ (.A1(_1169_),
    .A2(_1171_),
    .Y(_1173_),
    .B1(_1149_));
 sg13g2_or3_1 _5326_ (.A(_1166_),
    .B(_1172_),
    .C(_1173_),
    .X(_1174_));
 sg13g2_o21ai_1 _5327_ (.B1(_1166_),
    .Y(_1175_),
    .A1(_1172_),
    .A2(_1173_));
 sg13g2_nand3_1 _5328_ (.B(_1174_),
    .C(_1175_),
    .A(_1153_),
    .Y(_1176_));
 sg13g2_a21o_1 _5329_ (.A2(_1175_),
    .A1(_1174_),
    .B1(_1153_),
    .X(_1177_));
 sg13g2_nand3_1 _5330_ (.B(_1176_),
    .C(_1177_),
    .A(_1165_),
    .Y(_1178_));
 sg13g2_a21o_1 _5331_ (.A2(_1177_),
    .A1(_1176_),
    .B1(_1165_),
    .X(_1179_));
 sg13g2_and3_1 _5332_ (.X(_1180_),
    .A(_1164_),
    .B(_1178_),
    .C(_1179_));
 sg13g2_nand3_1 _5333_ (.B(_1178_),
    .C(_1179_),
    .A(_1164_),
    .Y(_1181_));
 sg13g2_a21oi_1 _5334_ (.A1(_1178_),
    .A2(_1179_),
    .Y(_1182_),
    .B1(_1164_));
 sg13g2_nor3_1 _5335_ (.A(_1163_),
    .B(_1180_),
    .C(_1182_),
    .Y(_1183_));
 sg13g2_o21ai_1 _5336_ (.B1(_1163_),
    .Y(_1184_),
    .A1(_1180_),
    .A2(_1182_));
 sg13g2_nor2b_2 _5337_ (.A(_1183_),
    .B_N(_1184_),
    .Y(\i_mandel.i_xy.hc.genblk2[3].state.D ));
 sg13g2_o21ai_1 _5338_ (.B1(_1181_),
    .Y(_1185_),
    .A1(_1163_),
    .A2(_1182_));
 sg13g2_nand2_1 _5339_ (.Y(_1186_),
    .A(_1176_),
    .B(_1178_));
 sg13g2_nor2_1 _5340_ (.A(_3310_),
    .B(_1124_),
    .Y(_1187_));
 sg13g2_nor2b_1 _5341_ (.A(_1172_),
    .B_N(_1174_),
    .Y(_1188_));
 sg13g2_nor2_1 _5342_ (.A(_3318_),
    .B(_1129_),
    .Y(_1189_));
 sg13g2_nor2_1 _5343_ (.A(_3383_),
    .B(_1147_),
    .Y(_1190_));
 sg13g2_and4_1 _5344_ (.A(_3305_),
    .B(_3381_),
    .C(net810),
    .D(_1170_),
    .X(_1191_));
 sg13g2_nand3_1 _5345_ (.B(_3381_),
    .C(net812),
    .A(_3305_),
    .Y(_1192_));
 sg13g2_a21oi_1 _5346_ (.A1(_1167_),
    .A2(_1192_),
    .Y(_1193_),
    .B1(_1191_));
 sg13g2_xnor2_1 _5347_ (.Y(_1194_),
    .A(_1168_),
    .B(_1193_));
 sg13g2_nor3_1 _5348_ (.A(_3318_),
    .B(_1129_),
    .C(_1194_),
    .Y(_1195_));
 sg13g2_xnor2_1 _5349_ (.Y(_1196_),
    .A(_1189_),
    .B(_1194_));
 sg13g2_nor2b_1 _5350_ (.A(_1188_),
    .B_N(_1196_),
    .Y(_1197_));
 sg13g2_xnor2_1 _5351_ (.Y(_1198_),
    .A(_1188_),
    .B(_1196_));
 sg13g2_xnor2_1 _5352_ (.Y(_1199_),
    .A(_1187_),
    .B(_1198_));
 sg13g2_nor2b_1 _5353_ (.A(_1199_),
    .B_N(_1186_),
    .Y(_1200_));
 sg13g2_nand2b_1 _5354_ (.Y(_1201_),
    .B(_1199_),
    .A_N(_1186_));
 sg13g2_nand2b_1 _5355_ (.Y(_1202_),
    .B(_1201_),
    .A_N(_1200_));
 sg13g2_xnor2_1 _5356_ (.Y(\i_mandel.i_xy.hc.genblk2[4].state.D ),
    .A(_1185_),
    .B(_1202_));
 sg13g2_a21oi_1 _5357_ (.A1(_1185_),
    .A2(_1201_),
    .Y(_1203_),
    .B1(_1200_));
 sg13g2_a21o_1 _5358_ (.A2(_1198_),
    .A1(_1187_),
    .B1(_1197_),
    .X(_1204_));
 sg13g2_and2_1 _5359_ (.A(net790),
    .B(_1125_),
    .X(_1205_));
 sg13g2_a21o_1 _5360_ (.A2(_1193_),
    .A1(_1168_),
    .B1(_1195_),
    .X(_1206_));
 sg13g2_nor2_1 _5361_ (.A(_3310_),
    .B(_1129_),
    .Y(_1207_));
 sg13g2_nor2_1 _5362_ (.A(_3318_),
    .B(_1147_),
    .Y(_1208_));
 sg13g2_nand4_1 _5363_ (.B(_3382_),
    .C(net812),
    .A(_3317_),
    .Y(_1209_),
    .D(net810));
 sg13g2_nor2_1 _5364_ (.A(_3318_),
    .B(net813),
    .Y(_1210_));
 sg13g2_o21ai_1 _5365_ (.B1(_1209_),
    .Y(_1211_),
    .A1(_1190_),
    .A2(_1210_));
 sg13g2_nor4_1 _5366_ (.A(_3383_),
    .B(net813),
    .C(_1167_),
    .D(_1211_),
    .Y(_1212_));
 sg13g2_xnor2_1 _5367_ (.Y(_1213_),
    .A(_1191_),
    .B(_1211_));
 sg13g2_xnor2_1 _5368_ (.Y(_1214_),
    .A(_1207_),
    .B(_1213_));
 sg13g2_nor2b_1 _5369_ (.A(_1214_),
    .B_N(_1206_),
    .Y(_1215_));
 sg13g2_xnor2_1 _5370_ (.Y(_1216_),
    .A(_1206_),
    .B(_1214_));
 sg13g2_xor2_1 _5371_ (.B(_1216_),
    .A(_1205_),
    .X(_1217_));
 sg13g2_nand2_1 _5372_ (.Y(_1218_),
    .A(_1204_),
    .B(_1217_));
 sg13g2_xnor2_1 _5373_ (.Y(_1219_),
    .A(_1204_),
    .B(_1217_));
 sg13g2_xor2_1 _5374_ (.B(_1219_),
    .A(_1203_),
    .X(\i_mandel.i_xy.hc.genblk2[5].state.D ));
 sg13g2_o21ai_1 _5375_ (.B1(_1218_),
    .Y(_1220_),
    .A1(_1203_),
    .A2(_1219_));
 sg13g2_a21oi_1 _5376_ (.A1(_1205_),
    .A2(_1216_),
    .Y(_1221_),
    .B1(_1215_));
 sg13g2_nand2b_1 _5377_ (.Y(_1222_),
    .B(_1125_),
    .A_N(_3345_));
 sg13g2_a21oi_1 _5378_ (.A1(_1207_),
    .A2(_1213_),
    .Y(_1223_),
    .B1(_1212_));
 sg13g2_nand2_1 _5379_ (.Y(_1224_),
    .A(net790),
    .B(_1130_));
 sg13g2_nand2_1 _5380_ (.Y(_1225_),
    .A(_3309_),
    .B(net811));
 sg13g2_nand3_1 _5381_ (.B(_1137_),
    .C(_1208_),
    .A(_3309_),
    .Y(_1226_));
 sg13g2_nor2_1 _5382_ (.A(_3310_),
    .B(net814),
    .Y(_1227_));
 sg13g2_o21ai_1 _5383_ (.B1(_1226_),
    .Y(_1228_),
    .A1(_1208_),
    .A2(_1227_));
 sg13g2_xor2_1 _5384_ (.B(_1228_),
    .A(_1209_),
    .X(_1229_));
 sg13g2_nand2b_1 _5385_ (.Y(_1230_),
    .B(_1229_),
    .A_N(_1224_));
 sg13g2_xnor2_1 _5386_ (.Y(_1231_),
    .A(_1224_),
    .B(_1229_));
 sg13g2_nand2b_1 _5387_ (.Y(_1232_),
    .B(_1231_),
    .A_N(_1223_));
 sg13g2_xor2_1 _5388_ (.B(_1231_),
    .A(_1223_),
    .X(_1233_));
 sg13g2_xnor2_1 _5389_ (.Y(_1234_),
    .A(_1222_),
    .B(_1233_));
 sg13g2_nor2_1 _5390_ (.A(_1221_),
    .B(_1234_),
    .Y(_1235_));
 sg13g2_xor2_1 _5391_ (.B(_1234_),
    .A(_1221_),
    .X(_1236_));
 sg13g2_xor2_1 _5392_ (.B(_1236_),
    .A(_1220_),
    .X(\i_mandel.i_xy.hc.genblk2[6].state.D ));
 sg13g2_a21oi_1 _5393_ (.A1(_1220_),
    .A2(_1236_),
    .Y(_1237_),
    .B1(_1235_));
 sg13g2_o21ai_1 _5394_ (.B1(_1232_),
    .Y(_1238_),
    .A1(_1222_),
    .A2(_1233_));
 sg13g2_nor2_2 _5395_ (.A(_3354_),
    .B(_1124_),
    .Y(_1239_));
 sg13g2_nand2_2 _5396_ (.Y(_1240_),
    .A(_3353_),
    .B(_1125_));
 sg13g2_o21ai_1 _5397_ (.B1(_1230_),
    .Y(_1241_),
    .A1(_1209_),
    .A2(_1228_));
 sg13g2_nor2_1 _5398_ (.A(_3345_),
    .B(_1129_),
    .Y(_1242_));
 sg13g2_and2_1 _5399_ (.A(_3331_),
    .B(net811),
    .X(_1243_));
 sg13g2_nand2_1 _5400_ (.Y(_1244_),
    .A(net790),
    .B(net812));
 sg13g2_xnor2_1 _5401_ (.Y(_1245_),
    .A(_1225_),
    .B(_1244_));
 sg13g2_nor2_1 _5402_ (.A(_1226_),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_nand2_1 _5403_ (.Y(_1247_),
    .A(_1226_),
    .B(_1245_));
 sg13g2_nand2b_1 _5404_ (.Y(_1248_),
    .B(_1247_),
    .A_N(_1246_));
 sg13g2_xnor2_1 _5405_ (.Y(_1249_),
    .A(_1242_),
    .B(_1248_));
 sg13g2_nand2_1 _5406_ (.Y(_1250_),
    .A(_1241_),
    .B(_1249_));
 sg13g2_xnor2_1 _5407_ (.Y(_1251_),
    .A(_1241_),
    .B(_1249_));
 sg13g2_xnor2_1 _5408_ (.Y(_1252_),
    .A(_1239_),
    .B(_1251_));
 sg13g2_nand2_1 _5409_ (.Y(_1253_),
    .A(_1238_),
    .B(_1252_));
 sg13g2_xnor2_1 _5410_ (.Y(_1254_),
    .A(_1238_),
    .B(_1252_));
 sg13g2_xor2_1 _5411_ (.B(_1254_),
    .A(_1237_),
    .X(\i_mandel.i_xy.hc.genblk2[7].state.D ));
 sg13g2_o21ai_1 _5412_ (.B1(_1253_),
    .Y(_1255_),
    .A1(_1237_),
    .A2(_1254_));
 sg13g2_o21ai_1 _5413_ (.B1(_1250_),
    .Y(_1256_),
    .A1(_1240_),
    .A2(_1251_));
 sg13g2_a21oi_1 _5414_ (.A1(_1242_),
    .A2(_1247_),
    .Y(_1257_),
    .B1(_1246_));
 sg13g2_nor2_1 _5415_ (.A(_3354_),
    .B(_1129_),
    .Y(_1258_));
 sg13g2_nand2_2 _5416_ (.Y(_1259_),
    .A(_3353_),
    .B(_1130_));
 sg13g2_nor2_1 _5417_ (.A(_3345_),
    .B(net813),
    .Y(_1260_));
 sg13g2_nand2b_1 _5418_ (.Y(_1261_),
    .B(_1243_),
    .A_N(_1227_));
 sg13g2_nand4_1 _5419_ (.B(net787),
    .C(net812),
    .A(_3309_),
    .Y(_1262_),
    .D(_1243_));
 sg13g2_xor2_1 _5420_ (.B(_1261_),
    .A(_1260_),
    .X(_1263_));
 sg13g2_xnor2_1 _5421_ (.Y(_1264_),
    .A(_1259_),
    .B(_1263_));
 sg13g2_nor2_1 _5422_ (.A(_1257_),
    .B(_1264_),
    .Y(_1265_));
 sg13g2_xnor2_1 _5423_ (.Y(_1266_),
    .A(_1257_),
    .B(_1264_));
 sg13g2_nor2_1 _5424_ (.A(_1240_),
    .B(_1266_),
    .Y(_1267_));
 sg13g2_xnor2_1 _5425_ (.Y(_1268_),
    .A(_1240_),
    .B(_1266_));
 sg13g2_nor2b_1 _5426_ (.A(_1268_),
    .B_N(_1256_),
    .Y(_1269_));
 sg13g2_xor2_1 _5427_ (.B(_1268_),
    .A(_1256_),
    .X(_1270_));
 sg13g2_inv_1 _5428_ (.Y(_1271_),
    .A(_1270_));
 sg13g2_xnor2_1 _5429_ (.Y(\i_mandel.i_xy.hc.genblk2[8].state.D ),
    .A(_1255_),
    .B(_1270_));
 sg13g2_o21ai_1 _5430_ (.B1(_1262_),
    .Y(_1272_),
    .A1(_1259_),
    .A2(_1263_));
 sg13g2_nor2_1 _5431_ (.A(net786),
    .B(net813),
    .Y(_1273_));
 sg13g2_nand3b_1 _5432_ (.B(net811),
    .C(_1244_),
    .Y(_1274_),
    .A_N(net787));
 sg13g2_xor2_1 _5433_ (.B(_1274_),
    .A(_1273_),
    .X(_1275_));
 sg13g2_xnor2_1 _5434_ (.Y(_1276_),
    .A(_1259_),
    .B(_1275_));
 sg13g2_nand2b_1 _5435_ (.Y(_1277_),
    .B(_1272_),
    .A_N(_1276_));
 sg13g2_xor2_1 _5436_ (.B(_1276_),
    .A(_1272_),
    .X(_1278_));
 sg13g2_or2_1 _5437_ (.X(_1279_),
    .B(_1278_),
    .A(_1240_));
 sg13g2_xnor2_1 _5438_ (.Y(_1280_),
    .A(_1239_),
    .B(_1278_));
 sg13g2_o21ai_1 _5439_ (.B1(_1280_),
    .Y(_1281_),
    .A1(_1265_),
    .A2(_1267_));
 sg13g2_or3_1 _5440_ (.A(_1265_),
    .B(_1267_),
    .C(_1280_),
    .X(_1282_));
 sg13g2_nand2_1 _5441_ (.Y(_1283_),
    .A(_1281_),
    .B(_1282_));
 sg13g2_a21oi_1 _5442_ (.A1(_1255_),
    .A2(_1271_),
    .Y(_1284_),
    .B1(_1269_));
 sg13g2_xor2_1 _5443_ (.B(_1284_),
    .A(_1283_),
    .X(\i_mandel.i_xy.hc.genblk2[9].state.D ));
 sg13g2_nand3_1 _5444_ (.B(_1243_),
    .C(_1260_),
    .A(net786),
    .Y(_1285_));
 sg13g2_o21ai_1 _5445_ (.B1(_1285_),
    .Y(_1286_),
    .A1(_1259_),
    .A2(_1275_));
 sg13g2_nand3_1 _5446_ (.B(net812),
    .C(net811),
    .A(net787),
    .Y(_1287_));
 sg13g2_o21ai_1 _5447_ (.B1(_1287_),
    .Y(_1288_),
    .A1(net812),
    .A2(net810));
 sg13g2_nor2_1 _5448_ (.A(net786),
    .B(_1288_),
    .Y(_1289_));
 sg13g2_xnor2_1 _5449_ (.Y(_1290_),
    .A(_1258_),
    .B(_1289_));
 sg13g2_inv_1 _5450_ (.Y(_1291_),
    .A(_1290_));
 sg13g2_xnor2_1 _5451_ (.Y(_1292_),
    .A(_1286_),
    .B(_1290_));
 sg13g2_xnor2_1 _5452_ (.Y(_1293_),
    .A(_1239_),
    .B(_1292_));
 sg13g2_nand3_1 _5453_ (.B(_1279_),
    .C(_1293_),
    .A(_1277_),
    .Y(_1294_));
 sg13g2_a21o_1 _5454_ (.A2(_1279_),
    .A1(_1277_),
    .B1(_1293_),
    .X(_1295_));
 sg13g2_nand2_1 _5455_ (.Y(_1296_),
    .A(_1294_),
    .B(_1295_));
 sg13g2_o21ai_1 _5456_ (.B1(_1281_),
    .Y(_1297_),
    .A1(_1283_),
    .A2(_1284_));
 sg13g2_xnor2_1 _5457_ (.Y(\i_mandel.i_xy.hc.genblk2[10].state.D ),
    .A(_1296_),
    .B(_1297_));
 sg13g2_a221oi_1 _5458_ (.B2(_1129_),
    .C1(_1289_),
    .B1(_1273_),
    .A1(net813),
    .Y(_1298_),
    .A2(_1258_));
 sg13g2_nor3_1 _5459_ (.A(_1240_),
    .B(_1286_),
    .C(_1291_),
    .Y(_1299_));
 sg13g2_nand3_1 _5460_ (.B(_1286_),
    .C(_1291_),
    .A(_1240_),
    .Y(_1300_));
 sg13g2_nand2b_1 _5461_ (.Y(_1301_),
    .B(_1300_),
    .A_N(_1299_));
 sg13g2_xnor2_1 _5462_ (.Y(_1302_),
    .A(_1298_),
    .B(_1301_));
 sg13g2_nand2_1 _5463_ (.Y(_1303_),
    .A(_1281_),
    .B(_1295_));
 sg13g2_a21oi_2 _5464_ (.B1(_1302_),
    .Y(_1304_),
    .A2(_1303_),
    .A1(_1294_));
 sg13g2_inv_1 _5465_ (.Y(\i_mandel.i_xy.hc.genblk2[11].state.D ),
    .A(_1304_));
 sg13g2_nand2_2 _5466_ (.Y(_1305_),
    .A(net963),
    .B(_3268_));
 sg13g2_and3_1 _5467_ (.X(_0033_),
    .A(net184),
    .B(net963),
    .C(_3268_));
 sg13g2_nor2_1 _5468_ (.A(net949),
    .B(net214),
    .Y(_1306_));
 sg13g2_nor3_1 _5469_ (.A(net867),
    .B(_1305_),
    .C(_1306_),
    .Y(_0034_));
 sg13g2_xnor2_1 _5470_ (.Y(_1307_),
    .A(net227),
    .B(net867));
 sg13g2_nor2_1 _5471_ (.A(_1305_),
    .B(_1307_),
    .Y(_0035_));
 sg13g2_and3_1 _5472_ (.X(_1308_),
    .A(\step[2] ),
    .B(net193),
    .C(net867));
 sg13g2_a21oi_1 _5473_ (.A1(\step[2] ),
    .A2(net867),
    .Y(_1309_),
    .B1(net193));
 sg13g2_nor3_1 _5474_ (.A(_1305_),
    .B(_1308_),
    .C(net194),
    .Y(_0036_));
 sg13g2_xnor2_1 _5475_ (.Y(_1310_),
    .A(net219),
    .B(_1308_));
 sg13g2_nor2_1 _5476_ (.A(_1305_),
    .B(net220),
    .Y(_0037_));
 sg13g2_and2_1 _5477_ (.A(\i_coord.l_xir.genblk2[2].state.Q ),
    .B(\i_coord.x_row_start[-11] ),
    .X(_1311_));
 sg13g2_or2_1 _5478_ (.X(_1312_),
    .B(\i_coord.x_row_start[-11] ),
    .A(\i_coord.l_xir.genblk2[2].state.Q ));
 sg13g2_nand2b_1 _5479_ (.Y(_1313_),
    .B(_1312_),
    .A_N(_1311_));
 sg13g2_nand2_1 _5480_ (.Y(_1314_),
    .A(\i_coord.l_xir.genblk2[0].state.Q ),
    .B(net206));
 sg13g2_xor2_1 _5481_ (.B(net271),
    .A(\i_coord.l_xir.genblk2[1].state.Q ),
    .X(_1315_));
 sg13g2_nor2b_1 _5482_ (.A(_1314_),
    .B_N(_1315_),
    .Y(_1316_));
 sg13g2_a21o_1 _5483_ (.A2(\i_coord.x_row_start[-12] ),
    .A1(\i_coord.l_xir.genblk2[1].state.Q ),
    .B1(_1316_),
    .X(_1317_));
 sg13g2_a21oi_1 _5484_ (.A1(_1312_),
    .A2(_1317_),
    .Y(_1318_),
    .B1(_1311_));
 sg13g2_nand2_1 _5485_ (.Y(_1319_),
    .A(\i_coord.l_xir.genblk2[3].state.Q ),
    .B(\i_coord.x_row_start[-10] ));
 sg13g2_xnor2_1 _5486_ (.Y(_1320_),
    .A(\i_coord.l_xir.genblk2[3].state.Q ),
    .B(\i_coord.x_row_start[-10] ));
 sg13g2_or2_1 _5487_ (.X(_1321_),
    .B(_1320_),
    .A(_1318_));
 sg13g2_xor2_1 _5488_ (.B(_1320_),
    .A(_1318_),
    .X(_1322_));
 sg13g2_nand2_1 _5489_ (.Y(_1323_),
    .A(\i_coord.l_xl.genblk2[3].state.Q ),
    .B(net780));
 sg13g2_o21ai_1 _5490_ (.B1(net770),
    .Y(_1324_),
    .A1(net794),
    .A2(_1322_));
 sg13g2_a22oi_1 _5491_ (.Y(_0038_),
    .B1(_1323_),
    .B2(_1324_),
    .A2(net761),
    .A1(_3098_));
 sg13g2_xnor2_1 _5492_ (.Y(_1325_),
    .A(\i_coord.l_xir.genblk2[4].state.Q ),
    .B(\i_coord.x_row_start[-9] ));
 sg13g2_a21oi_1 _5493_ (.A1(_1319_),
    .A2(_1321_),
    .Y(_1326_),
    .B1(_1325_));
 sg13g2_and3_1 _5494_ (.X(_1327_),
    .A(_1319_),
    .B(_1321_),
    .C(_1325_));
 sg13g2_or3_1 _5495_ (.A(net779),
    .B(_1326_),
    .C(_1327_),
    .X(_1328_));
 sg13g2_a21oi_1 _5496_ (.A1(\i_coord.l_xl.genblk2[4].state.Q ),
    .A2(net780),
    .Y(_1329_),
    .B1(net765));
 sg13g2_a22oi_1 _5497_ (.Y(_0039_),
    .B1(_1328_),
    .B2(_1329_),
    .A2(net761),
    .A1(_3099_));
 sg13g2_a21o_1 _5498_ (.A2(\i_coord.x_row_start[-9] ),
    .A1(\i_coord.l_xir.genblk2[4].state.Q ),
    .B1(_1326_),
    .X(_1330_));
 sg13g2_nand2_1 _5499_ (.Y(_1331_),
    .A(\i_coord.l_xir.genblk2[5].state.Q ),
    .B(\i_coord.x_row_start[-8] ));
 sg13g2_xor2_1 _5500_ (.B(\i_coord.x_row_start[-8] ),
    .A(\i_coord.l_xir.genblk2[5].state.Q ),
    .X(_1332_));
 sg13g2_o21ai_1 _5501_ (.B1(net770),
    .Y(_1333_),
    .A1(_1330_),
    .A2(_1332_));
 sg13g2_a21o_1 _5502_ (.A2(_1332_),
    .A1(_1330_),
    .B1(_1333_),
    .X(_1334_));
 sg13g2_a21oi_1 _5503_ (.A1(\i_coord.l_xl.genblk2[5].state.Q ),
    .A2(net780),
    .Y(_1335_),
    .B1(net765));
 sg13g2_a22oi_1 _5504_ (.Y(_0040_),
    .B1(_1334_),
    .B2(_1335_),
    .A2(net761),
    .A1(_3100_));
 sg13g2_nand2_1 _5505_ (.Y(_1336_),
    .A(\i_coord.l_xir.genblk2[6].state.Q ),
    .B(\i_coord.x_row_start[-7] ));
 sg13g2_xnor2_1 _5506_ (.Y(_1337_),
    .A(\i_coord.l_xir.genblk2[6].state.Q ),
    .B(\i_coord.x_row_start[-7] ));
 sg13g2_o21ai_1 _5507_ (.B1(_1330_),
    .Y(_1338_),
    .A1(\i_coord.l_xir.genblk2[5].state.Q ),
    .A2(\i_coord.x_row_start[-8] ));
 sg13g2_nand3_1 _5508_ (.B(_1337_),
    .C(_1338_),
    .A(_1331_),
    .Y(_1339_));
 sg13g2_a21o_1 _5509_ (.A2(_1338_),
    .A1(_1331_),
    .B1(_1337_),
    .X(_1340_));
 sg13g2_nand3_1 _5510_ (.B(_1339_),
    .C(_1340_),
    .A(net770),
    .Y(_1341_));
 sg13g2_a21oi_1 _5511_ (.A1(\i_coord.l_xl.genblk2[6].state.Q ),
    .A2(net779),
    .Y(_1342_),
    .B1(net765));
 sg13g2_a22oi_1 _5512_ (.Y(_0041_),
    .B1(_1341_),
    .B2(_1342_),
    .A2(net759),
    .A1(_3101_));
 sg13g2_nand2_1 _5513_ (.Y(_1343_),
    .A(net805),
    .B(net218));
 sg13g2_xnor2_1 _5514_ (.Y(_1344_),
    .A(net805),
    .B(\i_coord.x_row_start[-6] ));
 sg13g2_a21o_1 _5515_ (.A2(_1340_),
    .A1(_1336_),
    .B1(_1344_),
    .X(_1345_));
 sg13g2_nand3_1 _5516_ (.B(_1340_),
    .C(_1344_),
    .A(_1336_),
    .Y(_1346_));
 sg13g2_and2_1 _5517_ (.A(_1345_),
    .B(_1346_),
    .X(_1347_));
 sg13g2_a221oi_1 _5518_ (.B2(_1347_),
    .C1(net764),
    .B1(_3262_),
    .A1(\i_coord.l_xl.genblk2[7].state.Q ),
    .Y(_1348_),
    .A2(net779));
 sg13g2_a21oi_1 _5519_ (.A1(_3103_),
    .A2(net759),
    .Y(_0042_),
    .B1(_1348_));
 sg13g2_xnor2_1 _5520_ (.Y(_1349_),
    .A(net805),
    .B(\i_coord.x_row_start[-5] ));
 sg13g2_nand3_1 _5521_ (.B(_1345_),
    .C(_1349_),
    .A(_1343_),
    .Y(_1350_));
 sg13g2_a21oi_1 _5522_ (.A1(_1343_),
    .A2(_1345_),
    .Y(_1351_),
    .B1(_1349_));
 sg13g2_nor2_1 _5523_ (.A(net777),
    .B(_1351_),
    .Y(_1352_));
 sg13g2_nand2_1 _5524_ (.Y(_1353_),
    .A(_1350_),
    .B(_1352_));
 sg13g2_a21oi_1 _5525_ (.A1(\i_coord.l_xl.genblk2[8].state.Q ),
    .A2(net779),
    .Y(_1354_),
    .B1(net765));
 sg13g2_a22oi_1 _5526_ (.Y(_0043_),
    .B1(_1353_),
    .B2(_1354_),
    .A2(net759),
    .A1(_3104_));
 sg13g2_xor2_1 _5527_ (.B(\i_coord.x_row_start[-4] ),
    .A(net805),
    .X(_1355_));
 sg13g2_a21o_1 _5528_ (.A2(\i_coord.x_row_start[-5] ),
    .A1(\i_coord.l_xir.genblk2[7].state.Q ),
    .B1(_1351_),
    .X(_1356_));
 sg13g2_a21oi_1 _5529_ (.A1(_1355_),
    .A2(_1356_),
    .Y(_1357_),
    .B1(net777));
 sg13g2_o21ai_1 _5530_ (.B1(_1357_),
    .Y(_1358_),
    .A1(_1355_),
    .A2(_1356_));
 sg13g2_a21oi_1 _5531_ (.A1(\i_coord.l_xl.genblk2[9].state.Q ),
    .A2(net777),
    .Y(_1359_),
    .B1(net764));
 sg13g2_a22oi_1 _5532_ (.Y(_0044_),
    .B1(_1358_),
    .B2(_1359_),
    .A2(net759),
    .A1(_3105_));
 sg13g2_xnor2_1 _5533_ (.Y(_1360_),
    .A(net805),
    .B(\i_coord.x_row_start[-3] ));
 sg13g2_nand2_1 _5534_ (.Y(_1361_),
    .A(_1351_),
    .B(_1355_));
 sg13g2_o21ai_1 _5535_ (.B1(net805),
    .Y(_1362_),
    .A1(\i_coord.x_row_start[-5] ),
    .A2(\i_coord.x_row_start[-4] ));
 sg13g2_a21oi_1 _5536_ (.A1(_1361_),
    .A2(_1362_),
    .Y(_1363_),
    .B1(_1360_));
 sg13g2_nand3_1 _5537_ (.B(_1361_),
    .C(_1362_),
    .A(_1360_),
    .Y(_1364_));
 sg13g2_nor2b_1 _5538_ (.A(_1363_),
    .B_N(_1364_),
    .Y(_1365_));
 sg13g2_a221oi_1 _5539_ (.B2(_1365_),
    .C1(net764),
    .B1(_3262_),
    .A1(\i_coord.l_xl.genblk2[10].state.Q ),
    .Y(_1366_),
    .A2(net777));
 sg13g2_a21oi_1 _5540_ (.A1(_3106_),
    .A2(net758),
    .Y(_0045_),
    .B1(_1366_));
 sg13g2_xnor2_1 _5541_ (.Y(_1367_),
    .A(net806),
    .B(\i_coord.x_row_start[-2] ));
 sg13g2_a21oi_1 _5542_ (.A1(net805),
    .A2(\i_coord.x_row_start[-3] ),
    .Y(_1368_),
    .B1(_1363_));
 sg13g2_o21ai_1 _5543_ (.B1(net769),
    .Y(_1369_),
    .A1(_1367_),
    .A2(_1368_));
 sg13g2_a21o_1 _5544_ (.A2(_1368_),
    .A1(_1367_),
    .B1(_1369_),
    .X(_1370_));
 sg13g2_a21oi_1 _5545_ (.A1(\i_coord.l_xl.genblk2[11].state.Q ),
    .A2(net778),
    .Y(_1371_),
    .B1(net764));
 sg13g2_a22oi_1 _5546_ (.Y(_0046_),
    .B1(_1370_),
    .B2(_1371_),
    .A2(net758),
    .A1(_3107_));
 sg13g2_xnor2_1 _5547_ (.Y(_1372_),
    .A(net806),
    .B(\i_coord.x_row_start[-1] ));
 sg13g2_nor3_1 _5548_ (.A(_1360_),
    .B(_1361_),
    .C(_1367_),
    .Y(_1373_));
 sg13g2_o21ai_1 _5549_ (.B1(net805),
    .Y(_1374_),
    .A1(\i_coord.x_row_start[-3] ),
    .A2(\i_coord.x_row_start[-2] ));
 sg13g2_nand3b_1 _5550_ (.B(_1374_),
    .C(_1362_),
    .Y(_1375_),
    .A_N(_1373_));
 sg13g2_nand2b_1 _5551_ (.Y(_1376_),
    .B(_1375_),
    .A_N(_1372_));
 sg13g2_xnor2_1 _5552_ (.Y(_1377_),
    .A(_1372_),
    .B(_1375_));
 sg13g2_a221oi_1 _5553_ (.B2(_1377_),
    .C1(net764),
    .B1(_3262_),
    .A1(\i_coord.l_xl.genblk2[12].state.Q ),
    .Y(_1378_),
    .A2(net776));
 sg13g2_a21oi_1 _5554_ (.A1(_3108_),
    .A2(net758),
    .Y(_0047_),
    .B1(_1378_));
 sg13g2_xnor2_1 _5555_ (.Y(_1379_),
    .A(net806),
    .B(\i_coord.x_row_start[0] ));
 sg13g2_o21ai_1 _5556_ (.B1(_1376_),
    .Y(_1380_),
    .A1(_3102_),
    .A2(_3108_));
 sg13g2_xnor2_1 _5557_ (.Y(_1381_),
    .A(_1379_),
    .B(_1380_));
 sg13g2_nand2_1 _5558_ (.Y(_1382_),
    .A(_3262_),
    .B(_1381_));
 sg13g2_a21oi_1 _5559_ (.A1(\i_coord.l_xl.genblk2[13].state.Q ),
    .A2(net775),
    .Y(_1383_),
    .B1(net764));
 sg13g2_a22oi_1 _5560_ (.Y(_0048_),
    .B1(_1382_),
    .B2(_1383_),
    .A2(net758),
    .A1(_3109_));
 sg13g2_xnor2_1 _5561_ (.Y(_1384_),
    .A(net806),
    .B(\i_coord.x_row_start[1] ));
 sg13g2_or2_1 _5562_ (.X(_1385_),
    .B(_1379_),
    .A(_1376_));
 sg13g2_o21ai_1 _5563_ (.B1(net806),
    .Y(_1386_),
    .A1(\i_coord.x_row_start[-1] ),
    .A2(\i_coord.x_row_start[0] ));
 sg13g2_a21oi_1 _5564_ (.A1(_1385_),
    .A2(_1386_),
    .Y(_1387_),
    .B1(_1384_));
 sg13g2_and3_1 _5565_ (.X(_1388_),
    .A(_1384_),
    .B(_1385_),
    .C(_1386_));
 sg13g2_or3_1 _5566_ (.A(net775),
    .B(_1387_),
    .C(_1388_),
    .X(_1389_));
 sg13g2_a21oi_1 _5567_ (.A1(\i_coord.l_xl.genblk2[14].state.Q ),
    .A2(net775),
    .Y(_1390_),
    .B1(net764));
 sg13g2_a22oi_1 _5568_ (.Y(_0049_),
    .B1(_1389_),
    .B2(_1390_),
    .A2(net757),
    .A1(_3110_));
 sg13g2_a21oi_1 _5569_ (.A1(net806),
    .A2(\i_coord.x_row_start[1] ),
    .Y(_1391_),
    .B1(_1387_));
 sg13g2_xnor2_1 _5570_ (.Y(_1392_),
    .A(net806),
    .B(net225));
 sg13g2_a21oi_1 _5571_ (.A1(_1391_),
    .A2(_1392_),
    .Y(_1393_),
    .B1(net775));
 sg13g2_o21ai_1 _5572_ (.B1(_1393_),
    .Y(_1394_),
    .A1(_1391_),
    .A2(_1392_));
 sg13g2_a21oi_2 _5573_ (.B1(net764),
    .Y(_1395_),
    .A2(net775),
    .A1(\i_coord.l_xl.genblk2[15].state.Q ));
 sg13g2_a22oi_1 _5574_ (.Y(_0050_),
    .B1(_1394_),
    .B2(_1395_),
    .A2(net757),
    .A1(_3111_));
 sg13g2_nand3_1 _5575_ (.B(net2),
    .C(net3),
    .A(net1),
    .Y(_1396_));
 sg13g2_and2_2 _5576_ (.A(net880),
    .B(_1396_),
    .X(_1397_));
 sg13g2_nand2_1 _5577_ (.Y(_1398_),
    .A(net881),
    .B(_1396_));
 sg13g2_nor2_2 _5578_ (.A(net939),
    .B(_1396_),
    .Y(_1399_));
 sg13g2_nand2b_1 _5579_ (.Y(_1400_),
    .B(_1399_),
    .A_N(net4));
 sg13g2_o21ai_1 _5580_ (.B1(_1400_),
    .Y(_1401_),
    .A1(net948),
    .A2(_1398_));
 sg13g2_a22oi_1 _5581_ (.Y(_0051_),
    .B1(_1401_),
    .B2(net966),
    .A2(net802),
    .A1(net948));
 sg13g2_a22oi_1 _5582_ (.Y(_1402_),
    .B1(_1399_),
    .B2(net5),
    .A2(_1397_),
    .A1(net946));
 sg13g2_a21oi_1 _5583_ (.A1(_3173_),
    .A2(_1402_),
    .Y(_0052_),
    .B1(net958));
 sg13g2_a21oi_1 _5584_ (.A1(_3096_),
    .A2(_1399_),
    .Y(_1403_),
    .B1(_3181_));
 sg13g2_o21ai_1 _5585_ (.B1(_1403_),
    .Y(_1404_),
    .A1(net345),
    .A2(_1398_));
 sg13g2_nand2_1 _5586_ (.Y(_0053_),
    .A(net966),
    .B(_1404_));
 sg13g2_o21ai_1 _5587_ (.B1(net880),
    .Y(_1405_),
    .A1(_3097_),
    .A2(_1396_));
 sg13g2_a22oi_1 _5588_ (.Y(_1406_),
    .B1(_1405_),
    .B2(_3184_),
    .A2(_1397_),
    .A1(net326));
 sg13g2_nand2_1 _5589_ (.Y(_0054_),
    .A(net966),
    .B(_1406_));
 sg13g2_a22oi_1 _5590_ (.Y(_1407_),
    .B1(_1399_),
    .B2(net8),
    .A2(_1397_),
    .A1(net339));
 sg13g2_a21oi_1 _5591_ (.A1(_3189_),
    .A2(_1407_),
    .Y(_0055_),
    .B1(net958));
 sg13g2_a22oi_1 _5592_ (.Y(_1408_),
    .B1(_1399_),
    .B2(net9),
    .A2(_1397_),
    .A1(net308));
 sg13g2_a21oi_1 _5593_ (.A1(_3194_),
    .A2(_1408_),
    .Y(_0056_),
    .B1(net958));
 sg13g2_o21ai_1 _5594_ (.B1(net966),
    .Y(_1409_),
    .A1(_3190_),
    .A2(_1396_));
 sg13g2_a221oi_1 _5595_ (.B2(net343),
    .C1(_1409_),
    .B1(_1397_),
    .A1(net939),
    .Y(_1410_),
    .A2(_3198_));
 sg13g2_inv_1 _5596_ (.Y(_0057_),
    .A(_1410_));
 sg13g2_a22oi_1 _5597_ (.Y(_1411_),
    .B1(_1399_),
    .B2(net11),
    .A2(_1397_),
    .A1(net945));
 sg13g2_nand3_1 _5598_ (.B(_3178_),
    .C(_1411_),
    .A(net967),
    .Y(_0058_));
 sg13g2_nor2_2 _5599_ (.A(net940),
    .B(net783),
    .Y(_1412_));
 sg13g2_nand2_1 _5600_ (.Y(_1413_),
    .A(net882),
    .B(net771));
 sg13g2_nand2_1 _5601_ (.Y(_1414_),
    .A(\i_coord.l_yt.genblk2[0].state.Q ),
    .B(net755));
 sg13g2_nand2_1 _5602_ (.Y(_1415_),
    .A(net948),
    .B(net799));
 sg13g2_xor2_1 _5603_ (.B(_1415_),
    .A(net276),
    .X(_1416_));
 sg13g2_o21ai_1 _5604_ (.B1(_1414_),
    .Y(_0059_),
    .A1(net755),
    .A2(_1416_));
 sg13g2_nor2_2 _5605_ (.A(net797),
    .B(net756),
    .Y(_1417_));
 sg13g2_nand2_2 _5606_ (.Y(_1418_),
    .A(_3258_),
    .B(_1412_));
 sg13g2_nand2_1 _5607_ (.Y(_1419_),
    .A(net948),
    .B(\i_coord.y_row_start[-13] ));
 sg13g2_nand2_1 _5608_ (.Y(_1420_),
    .A(\i_coord.y_inc_row[-12] ),
    .B(net233));
 sg13g2_xor2_1 _5609_ (.B(\i_coord.y_row_start[-12] ),
    .A(net946),
    .X(_1421_));
 sg13g2_nand2b_1 _5610_ (.Y(_1422_),
    .B(_1421_),
    .A_N(_1419_));
 sg13g2_xor2_1 _5611_ (.B(_1421_),
    .A(_1419_),
    .X(_1423_));
 sg13g2_nor2_2 _5612_ (.A(net940),
    .B(net762),
    .Y(_1424_));
 sg13g2_nand2_2 _5613_ (.Y(_1425_),
    .A(net882),
    .B(net766));
 sg13g2_a22oi_1 _5614_ (.Y(_1426_),
    .B1(_1424_),
    .B2(net233),
    .A2(net755),
    .A1(\i_coord.l_yt.genblk2[1].state.Q ));
 sg13g2_nor2_2 _5615_ (.A(net792),
    .B(net755),
    .Y(_1427_));
 sg13g2_o21ai_1 _5616_ (.B1(_1426_),
    .Y(_0060_),
    .A1(_1418_),
    .A2(_1423_));
 sg13g2_nand2_1 _5617_ (.Y(_1428_),
    .A(\i_coord.y_inc_row[-11] ),
    .B(net292));
 sg13g2_xnor2_1 _5618_ (.Y(_1429_),
    .A(\i_coord.y_inc_row[-11] ),
    .B(\i_coord.y_row_start[-11] ));
 sg13g2_nand3_1 _5619_ (.B(_1422_),
    .C(_1429_),
    .A(_1420_),
    .Y(_1430_));
 sg13g2_a21o_1 _5620_ (.A2(_1422_),
    .A1(_1420_),
    .B1(_1429_),
    .X(_1431_));
 sg13g2_nand2_1 _5621_ (.Y(_1432_),
    .A(_1430_),
    .B(_1431_));
 sg13g2_nand2b_1 _5622_ (.Y(_1433_),
    .B(net755),
    .A_N(\i_coord.l_yt.genblk2[2].state.Q ));
 sg13g2_o21ai_1 _5623_ (.B1(_1433_),
    .Y(_1434_),
    .A1(net292),
    .A2(_1425_));
 sg13g2_a21oi_1 _5624_ (.A1(_1417_),
    .A2(_1432_),
    .Y(_0061_),
    .B1(_1434_));
 sg13g2_nand2_1 _5625_ (.Y(_1435_),
    .A(\i_coord.y_inc_row[-10] ),
    .B(\i_coord.y_row_start[-10] ));
 sg13g2_xnor2_1 _5626_ (.Y(_1436_),
    .A(\i_coord.y_inc_row[-10] ),
    .B(\i_coord.y_row_start[-10] ));
 sg13g2_nand3_1 _5627_ (.B(_1431_),
    .C(_1436_),
    .A(_1428_),
    .Y(_1437_));
 sg13g2_a21o_1 _5628_ (.A2(_1431_),
    .A1(_1428_),
    .B1(_1436_),
    .X(_1438_));
 sg13g2_nand2_1 _5629_ (.Y(_1439_),
    .A(_1437_),
    .B(_1438_));
 sg13g2_nand2b_1 _5630_ (.Y(_1440_),
    .B(net755),
    .A_N(\i_coord.l_yt.genblk2[3].state.Q ));
 sg13g2_o21ai_1 _5631_ (.B1(_1440_),
    .Y(_1441_),
    .A1(net298),
    .A2(_1425_));
 sg13g2_a21oi_1 _5632_ (.A1(_1417_),
    .A2(_1439_),
    .Y(_0062_),
    .B1(_1441_));
 sg13g2_a22oi_1 _5633_ (.Y(_1442_),
    .B1(_1424_),
    .B2(net282),
    .A2(net755),
    .A1(\i_coord.l_yt.genblk2[4].state.Q ));
 sg13g2_xnor2_1 _5634_ (.Y(_1443_),
    .A(\i_coord.y_inc_row[-9] ),
    .B(\i_coord.y_row_start[-9] ));
 sg13g2_a21oi_1 _5635_ (.A1(_1435_),
    .A2(_1438_),
    .Y(_1444_),
    .B1(_1443_));
 sg13g2_nand3_1 _5636_ (.B(_1438_),
    .C(_1443_),
    .A(_1435_),
    .Y(_1445_));
 sg13g2_nand2_1 _5637_ (.Y(_1446_),
    .A(_1417_),
    .B(_1445_));
 sg13g2_o21ai_1 _5638_ (.B1(_1442_),
    .Y(_0063_),
    .A1(_1444_),
    .A2(_1446_));
 sg13g2_a22oi_1 _5639_ (.Y(_1447_),
    .B1(_1424_),
    .B2(net244),
    .A2(net755),
    .A1(\i_coord.l_yt.genblk2[5].state.Q ));
 sg13g2_a21o_1 _5640_ (.A2(\i_coord.y_row_start[-9] ),
    .A1(\i_coord.y_inc_row[-9] ),
    .B1(_1444_),
    .X(_1448_));
 sg13g2_or2_1 _5641_ (.X(_1449_),
    .B(\i_coord.y_row_start[-8] ),
    .A(\i_coord.y_inc_row[-8] ));
 sg13g2_nand2_1 _5642_ (.Y(_1450_),
    .A(\i_coord.y_inc_row[-8] ),
    .B(\i_coord.y_row_start[-8] ));
 sg13g2_nand2_1 _5643_ (.Y(_1451_),
    .A(_1449_),
    .B(_1450_));
 sg13g2_xnor2_1 _5644_ (.Y(_1452_),
    .A(_1448_),
    .B(_1451_));
 sg13g2_nand2_1 _5645_ (.Y(_1453_),
    .A(_1427_),
    .B(_1452_));
 sg13g2_nand2_1 _5646_ (.Y(_0064_),
    .A(_1447_),
    .B(_1453_));
 sg13g2_nand2_1 _5647_ (.Y(_1454_),
    .A(\i_coord.y_inc_row[-7] ),
    .B(\i_coord.y_row_start[-7] ));
 sg13g2_xnor2_1 _5648_ (.Y(_1455_),
    .A(\i_coord.y_inc_row[-7] ),
    .B(\i_coord.y_row_start[-7] ));
 sg13g2_nand2b_1 _5649_ (.Y(_1456_),
    .B(_1450_),
    .A_N(_1448_));
 sg13g2_nand2_1 _5650_ (.Y(_1457_),
    .A(_1449_),
    .B(_1456_));
 sg13g2_nand2_1 _5651_ (.Y(_1458_),
    .A(_1455_),
    .B(_1457_));
 sg13g2_or2_1 _5652_ (.X(_1459_),
    .B(_1457_),
    .A(_1455_));
 sg13g2_a21oi_1 _5653_ (.A1(_1458_),
    .A2(_1459_),
    .Y(_1460_),
    .B1(_1418_));
 sg13g2_nor2_1 _5654_ (.A(\i_coord.l_yt.genblk2[6].state.Q ),
    .B(_1412_),
    .Y(_1461_));
 sg13g2_nor2_1 _5655_ (.A(net249),
    .B(_1425_),
    .Y(_1462_));
 sg13g2_nor3_1 _5656_ (.A(_1460_),
    .B(_1461_),
    .C(_1462_),
    .Y(_0065_));
 sg13g2_nand2_1 _5657_ (.Y(_1463_),
    .A(net944),
    .B(net252));
 sg13g2_xnor2_1 _5658_ (.Y(_1464_),
    .A(net944),
    .B(\i_coord.y_row_start[-6] ));
 sg13g2_nand3_1 _5659_ (.B(_1459_),
    .C(_1464_),
    .A(_1454_),
    .Y(_1465_));
 sg13g2_a21o_1 _5660_ (.A2(_1459_),
    .A1(_1454_),
    .B1(_1464_),
    .X(_1466_));
 sg13g2_a21oi_1 _5661_ (.A1(_1465_),
    .A2(_1466_),
    .Y(_1467_),
    .B1(_1418_));
 sg13g2_nor2_1 _5662_ (.A(net252),
    .B(_1425_),
    .Y(_1468_));
 sg13g2_nor2_1 _5663_ (.A(\i_coord.l_yt.genblk2[7].state.Q ),
    .B(_1412_),
    .Y(_1469_));
 sg13g2_nor3_1 _5664_ (.A(_1467_),
    .B(_1468_),
    .C(_1469_),
    .Y(_0066_));
 sg13g2_a22oi_1 _5665_ (.Y(_1470_),
    .B1(_1424_),
    .B2(net279),
    .A2(net756),
    .A1(\i_coord.l_yt.genblk2[8].state.Q ));
 sg13g2_nand2_1 _5666_ (.Y(_1471_),
    .A(net943),
    .B(\i_coord.y_row_start[-5] ));
 sg13g2_xnor2_1 _5667_ (.Y(_1472_),
    .A(net944),
    .B(\i_coord.y_row_start[-5] ));
 sg13g2_a21o_1 _5668_ (.A2(_1466_),
    .A1(_1463_),
    .B1(_1472_),
    .X(_1473_));
 sg13g2_nand3_1 _5669_ (.B(_1466_),
    .C(_1472_),
    .A(_1463_),
    .Y(_1474_));
 sg13g2_nand3_1 _5670_ (.B(_1473_),
    .C(_1474_),
    .A(_1427_),
    .Y(_1475_));
 sg13g2_nand2_1 _5671_ (.Y(_0067_),
    .A(_1470_),
    .B(_1475_));
 sg13g2_xor2_1 _5672_ (.B(net270),
    .A(net943),
    .X(_1476_));
 sg13g2_nand2_1 _5673_ (.Y(_1477_),
    .A(_1471_),
    .B(_1473_));
 sg13g2_nor2_1 _5674_ (.A(\i_coord.l_yt.genblk2[9].state.Q ),
    .B(_1412_),
    .Y(_1478_));
 sg13g2_xnor2_1 _5675_ (.Y(_1479_),
    .A(_1476_),
    .B(_1477_));
 sg13g2_a221oi_1 _5676_ (.B2(_1417_),
    .C1(_1478_),
    .B1(_1479_),
    .A1(_3112_),
    .Y(_0068_),
    .A2(_1424_));
 sg13g2_and2_1 _5677_ (.A(net942),
    .B(\i_coord.y_row_start[-3] ),
    .X(_1480_));
 sg13g2_xor2_1 _5678_ (.B(\i_coord.y_row_start[-3] ),
    .A(net942),
    .X(_1481_));
 sg13g2_nor2b_1 _5679_ (.A(_1473_),
    .B_N(_1476_),
    .Y(_1482_));
 sg13g2_o21ai_1 _5680_ (.B1(net943),
    .Y(_1483_),
    .A1(\i_coord.y_row_start[-5] ),
    .A2(\i_coord.y_row_start[-4] ));
 sg13g2_nand2b_1 _5681_ (.Y(_1484_),
    .B(_1483_),
    .A_N(_1482_));
 sg13g2_xor2_1 _5682_ (.B(_1484_),
    .A(_1481_),
    .X(_1485_));
 sg13g2_a22oi_1 _5683_ (.Y(_1486_),
    .B1(_1427_),
    .B2(_1485_),
    .A2(net756),
    .A1(\i_coord.l_yt.genblk2[10].state.Q ));
 sg13g2_o21ai_1 _5684_ (.B1(_1486_),
    .Y(_0069_),
    .A1(_3113_),
    .A2(_1425_));
 sg13g2_a21oi_1 _5685_ (.A1(_1481_),
    .A2(_1484_),
    .Y(_1487_),
    .B1(_1480_));
 sg13g2_xor2_1 _5686_ (.B(\i_coord.y_row_start[-2] ),
    .A(net943),
    .X(_1488_));
 sg13g2_nand2_1 _5687_ (.Y(_1489_),
    .A(\i_coord.l_yt.genblk2[11].state.Q ),
    .B(net756));
 sg13g2_xor2_1 _5688_ (.B(_1488_),
    .A(_1487_),
    .X(_1490_));
 sg13g2_a22oi_1 _5689_ (.Y(_1491_),
    .B1(_1490_),
    .B2(_1412_),
    .A2(_1489_),
    .A1(_1418_));
 sg13g2_a21o_1 _5690_ (.A2(_1424_),
    .A1(net245),
    .B1(_1491_),
    .X(_0070_));
 sg13g2_a22oi_1 _5691_ (.Y(_1492_),
    .B1(_1424_),
    .B2(net275),
    .A2(net756),
    .A1(\i_coord.l_yt.genblk2[12].state.Q ));
 sg13g2_xnor2_1 _5692_ (.Y(_1493_),
    .A(net942),
    .B(\i_coord.y_row_start[-1] ));
 sg13g2_and2_1 _5693_ (.A(_1481_),
    .B(_1488_),
    .X(_1494_));
 sg13g2_a221oi_1 _5694_ (.B2(_1494_),
    .C1(_1480_),
    .B1(_1482_),
    .A1(net942),
    .Y(_1495_),
    .A2(\i_coord.y_row_start[-2] ));
 sg13g2_nand3_1 _5695_ (.B(_1493_),
    .C(_1495_),
    .A(_1483_),
    .Y(_1496_));
 sg13g2_a21oi_1 _5696_ (.A1(_1483_),
    .A2(_1495_),
    .Y(_1497_),
    .B1(_1493_));
 sg13g2_nand2_1 _5697_ (.Y(_1498_),
    .A(_1417_),
    .B(_1496_));
 sg13g2_o21ai_1 _5698_ (.B1(_1492_),
    .Y(_0071_),
    .A1(_1497_),
    .A2(_1498_));
 sg13g2_and2_1 _5699_ (.A(net942),
    .B(\i_coord.y_row_start[0] ),
    .X(_1499_));
 sg13g2_xor2_1 _5700_ (.B(\i_coord.y_row_start[0] ),
    .A(net943),
    .X(_1500_));
 sg13g2_a21o_1 _5701_ (.A2(\i_coord.y_row_start[-1] ),
    .A1(net942),
    .B1(_1497_),
    .X(_1501_));
 sg13g2_and2_1 _5702_ (.A(_1500_),
    .B(_1501_),
    .X(_1502_));
 sg13g2_o21ai_1 _5703_ (.B1(_1417_),
    .Y(_1503_),
    .A1(_1500_),
    .A2(_1501_));
 sg13g2_a22oi_1 _5704_ (.Y(_1504_),
    .B1(_1424_),
    .B2(net263),
    .A2(net756),
    .A1(\i_coord.l_yt.genblk2[13].state.Q ));
 sg13g2_o21ai_1 _5705_ (.B1(_1504_),
    .Y(_0072_),
    .A1(_1502_),
    .A2(_1503_));
 sg13g2_a221oi_1 _5706_ (.B2(_1500_),
    .C1(_1499_),
    .B1(_1497_),
    .A1(net942),
    .Y(_1505_),
    .A2(\i_coord.y_row_start[-1] ));
 sg13g2_xnor2_1 _5707_ (.Y(_1506_),
    .A(net942),
    .B(net210));
 sg13g2_nor2_1 _5708_ (.A(net210),
    .B(_1425_),
    .Y(_1507_));
 sg13g2_xnor2_1 _5709_ (.Y(_1508_),
    .A(_1505_),
    .B(_1506_));
 sg13g2_a221oi_1 _5710_ (.B2(_1508_),
    .C1(_1507_),
    .B1(_1427_),
    .A1(_3114_),
    .Y(_0073_),
    .A2(net756));
 sg13g2_o21ai_1 _5711_ (.B1(net967),
    .Y(_1509_),
    .A1(\i_coord.demo_update_delay ),
    .A2(net781));
 sg13g2_a21oi_1 _5712_ (.A1(_3088_),
    .A2(net781),
    .Y(_0074_),
    .B1(_1509_));
 sg13g2_nor3_1 _5713_ (.A(_0168_),
    .B(_0166_),
    .C(_0167_),
    .Y(_1510_));
 sg13g2_nor3_1 _5714_ (.A(_1078_),
    .B(_0166_),
    .C(_1098_),
    .Y(_1511_));
 sg13g2_nor3_1 _5715_ (.A(_0169_),
    .B(_1510_),
    .C(_1511_),
    .Y(_0075_));
 sg13g2_nor3_1 _5716_ (.A(_1078_),
    .B(_1081_),
    .C(_1098_),
    .Y(_1512_));
 sg13g2_nor2_1 _5717_ (.A(_0169_),
    .B(_1512_),
    .Y(_0076_));
 sg13g2_nor2_1 _5718_ (.A(\i_vga.timing_ver.counter[9] ),
    .B(net242),
    .Y(_1513_));
 sg13g2_nand3_1 _5719_ (.B(_3147_),
    .C(_1513_),
    .A(net284),
    .Y(_1514_));
 sg13g2_nand3_1 _5720_ (.B(net315),
    .C(_3247_),
    .A(net208),
    .Y(_1515_));
 sg13g2_nor2_1 _5721_ (.A(_3087_),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_nand2_1 _5722_ (.Y(_1517_),
    .A(net365),
    .B(_1516_));
 sg13g2_inv_1 _5723_ (.Y(_1518_),
    .A(_1517_));
 sg13g2_o21ai_1 _5724_ (.B1(net962),
    .Y(_1519_),
    .A1(_1514_),
    .A2(_1517_));
 sg13g2_xnor2_1 _5725_ (.Y(_1520_),
    .A(net315),
    .B(_3247_));
 sg13g2_nand2b_1 _5726_ (.Y(_0077_),
    .B(net316),
    .A_N(_1519_));
 sg13g2_a21oi_1 _5727_ (.A1(\i_vga.timing_ver.counter[0] ),
    .A2(_3247_),
    .Y(_1521_),
    .B1(net208));
 sg13g2_nand2_1 _5728_ (.Y(_1522_),
    .A(net961),
    .B(_1515_));
 sg13g2_nor2_1 _5729_ (.A(net209),
    .B(_1522_),
    .Y(_0078_));
 sg13g2_xnor2_1 _5730_ (.Y(_1523_),
    .A(_3087_),
    .B(_1515_));
 sg13g2_nand2b_1 _5731_ (.Y(_0079_),
    .B(_1523_),
    .A_N(_1519_));
 sg13g2_nor2_1 _5732_ (.A(net331),
    .B(_1516_),
    .Y(_1524_));
 sg13g2_a21o_1 _5733_ (.A2(_1518_),
    .A1(_1514_),
    .B1(_1524_),
    .X(_1525_));
 sg13g2_nand2_1 _5734_ (.Y(_0080_),
    .A(net962),
    .B(net332));
 sg13g2_xor2_1 _5735_ (.B(_1517_),
    .A(net284),
    .X(_1526_));
 sg13g2_nor2_1 _5736_ (.A(net960),
    .B(net285),
    .Y(_0081_));
 sg13g2_a21oi_1 _5737_ (.A1(\i_vga.timing_ver.counter[4] ),
    .A2(_1518_),
    .Y(_1527_),
    .B1(net242));
 sg13g2_and3_1 _5738_ (.X(_1528_),
    .A(net242),
    .B(net364),
    .C(_1518_));
 sg13g2_o21ai_1 _5739_ (.B1(net962),
    .Y(_0082_),
    .A1(net243),
    .A2(_1528_));
 sg13g2_xnor2_1 _5740_ (.Y(_1529_),
    .A(net266),
    .B(_1528_));
 sg13g2_nand2_1 _5741_ (.Y(_0083_),
    .A(net962),
    .B(_1529_));
 sg13g2_a21oi_1 _5742_ (.A1(\i_vga.timing_ver.counter[6] ),
    .A2(_1528_),
    .Y(_1530_),
    .B1(net221));
 sg13g2_nand3_1 _5743_ (.B(\i_vga.timing_ver.counter[6] ),
    .C(_1528_),
    .A(net221),
    .Y(_1531_));
 sg13g2_inv_1 _5744_ (.Y(_1532_),
    .A(_1531_));
 sg13g2_o21ai_1 _5745_ (.B1(net962),
    .Y(_0084_),
    .A1(net222),
    .A2(_1532_));
 sg13g2_xor2_1 _5746_ (.B(_1531_),
    .A(net261),
    .X(_1533_));
 sg13g2_nand2_1 _5747_ (.Y(_0085_),
    .A(net961),
    .B(net262));
 sg13g2_nor2_1 _5748_ (.A(net216),
    .B(_1531_),
    .Y(_1534_));
 sg13g2_xnor2_1 _5749_ (.Y(_1535_),
    .A(net204),
    .B(net217));
 sg13g2_nand2b_1 _5750_ (.Y(_0086_),
    .B(_1535_),
    .A_N(_1519_));
 sg13g2_o21ai_1 _5751_ (.B1(net961),
    .Y(_1536_),
    .A1(net278),
    .A2(net866));
 sg13g2_nor2_1 _5752_ (.A(_3241_),
    .B(_1536_),
    .Y(_0087_));
 sg13g2_o21ai_1 _5753_ (.B1(net961),
    .Y(_1537_),
    .A1(_3086_),
    .A2(_3242_));
 sg13g2_a21oi_1 _5754_ (.A1(_3086_),
    .A2(_3242_),
    .Y(_0088_),
    .B1(_1537_));
 sg13g2_a21oi_1 _5755_ (.A1(\i_vga.timing_hor.counter[1] ),
    .A2(_3241_),
    .Y(_1538_),
    .B1(net196));
 sg13g2_nand2_1 _5756_ (.Y(_1539_),
    .A(net961),
    .B(_3243_));
 sg13g2_nor2_1 _5757_ (.A(net197),
    .B(_1539_),
    .Y(_0089_));
 sg13g2_nand2_1 _5758_ (.Y(_1540_),
    .A(net961),
    .B(_3244_));
 sg13g2_a21oi_1 _5759_ (.A1(_3085_),
    .A2(_3243_),
    .Y(_0090_),
    .B1(_1540_));
 sg13g2_a21oi_1 _5760_ (.A1(net241),
    .A2(_3244_),
    .Y(_1541_),
    .B1(net960));
 sg13g2_nand2_1 _5761_ (.Y(_0091_),
    .A(_3245_),
    .B(_1541_));
 sg13g2_nor2_1 _5762_ (.A(_3240_),
    .B(_3247_),
    .Y(_1542_));
 sg13g2_nand3_1 _5763_ (.B(\i_vga.timing_hor.counter[2] ),
    .C(\i_vga.timing_hor.counter[0] ),
    .A(\i_vga.timing_hor.counter[4] ),
    .Y(_1543_));
 sg13g2_nor3_1 _5764_ (.A(_3085_),
    .B(_3086_),
    .C(_1543_),
    .Y(_1544_));
 sg13g2_xnor2_1 _5765_ (.Y(_1545_),
    .A(net229),
    .B(_1544_));
 sg13g2_a22oi_1 _5766_ (.Y(_1546_),
    .B1(_1542_),
    .B2(net230),
    .A2(_3240_),
    .A1(\i_vga.timing_hor.counter[5] ));
 sg13g2_nor2_1 _5767_ (.A(net960),
    .B(net231),
    .Y(_0092_));
 sg13g2_and2_1 _5768_ (.A(\i_vga.timing_hor.counter[5] ),
    .B(_1544_),
    .X(_1547_));
 sg13g2_nand2_1 _5769_ (.Y(_1548_),
    .A(net866),
    .B(_1547_));
 sg13g2_a21oi_1 _5770_ (.A1(net941),
    .A2(_1548_),
    .Y(_1549_),
    .B1(net960));
 sg13g2_o21ai_1 _5771_ (.B1(_1549_),
    .Y(_0093_),
    .A1(net941),
    .A2(_1548_));
 sg13g2_and3_1 _5772_ (.X(_1550_),
    .A(\i_vga.timing_hor.counter[7] ),
    .B(net941),
    .C(_1547_));
 sg13g2_nand3_1 _5773_ (.B(net941),
    .C(_1547_),
    .A(\i_vga.timing_hor.counter[7] ),
    .Y(_1551_));
 sg13g2_a22oi_1 _5774_ (.Y(_1552_),
    .B1(_1542_),
    .B2(_1551_),
    .A2(_3240_),
    .A1(net254));
 sg13g2_a21oi_1 _5775_ (.A1(net941),
    .A2(_1547_),
    .Y(_1553_),
    .B1(net254));
 sg13g2_nor3_1 _5776_ (.A(net960),
    .B(_1552_),
    .C(net255),
    .Y(_0094_));
 sg13g2_nor2_1 _5777_ (.A(net305),
    .B(_1551_),
    .Y(_1554_));
 sg13g2_o21ai_1 _5778_ (.B1(net866),
    .Y(_1555_),
    .A1(_3247_),
    .A2(_1554_));
 sg13g2_nand3_1 _5779_ (.B(net866),
    .C(_1550_),
    .A(net305),
    .Y(_1556_));
 sg13g2_nand2_1 _5780_ (.Y(_1557_),
    .A(net305),
    .B(_1556_));
 sg13g2_nand3_1 _5781_ (.B(_1555_),
    .C(_1557_),
    .A(net961),
    .Y(_0095_));
 sg13g2_nand4_1 _5782_ (.B(\i_vga.timing_hor.counter[8] ),
    .C(net866),
    .A(\i_vga.timing_hor.counter[9] ),
    .Y(_1558_),
    .D(_1550_));
 sg13g2_xor2_1 _5783_ (.B(_1556_),
    .A(net295),
    .X(_1559_));
 sg13g2_nand2_1 _5784_ (.Y(_0096_),
    .A(net962),
    .B(net296));
 sg13g2_and3_1 _5785_ (.X(_1560_),
    .A(_3084_),
    .B(_3254_),
    .C(_1550_));
 sg13g2_o21ai_1 _5786_ (.B1(net866),
    .Y(_1561_),
    .A1(_3247_),
    .A2(_1560_));
 sg13g2_a21oi_1 _5787_ (.A1(net290),
    .A2(_1558_),
    .Y(_1562_),
    .B1(net960));
 sg13g2_nand2_1 _5788_ (.Y(_0097_),
    .A(_1561_),
    .B(net291));
 sg13g2_nor3_1 _5789_ (.A(net224),
    .B(net3),
    .C(net958),
    .Y(_1563_));
 sg13g2_and3_1 _5790_ (.X(_0098_),
    .A(net785),
    .B(_1117_),
    .C(_1563_));
 sg13g2_nand3_1 _5791_ (.B(net833),
    .C(net760),
    .A(net949),
    .Y(_1564_));
 sg13g2_and2_1 _5792_ (.A(net949),
    .B(_1564_),
    .X(_1565_));
 sg13g2_nand2_1 _5793_ (.Y(_1566_),
    .A(net949),
    .B(_1564_));
 sg13g2_nor2_1 _5794_ (.A(net206),
    .B(net795),
    .Y(_1567_));
 sg13g2_nor2_2 _5795_ (.A(net869),
    .B(net782),
    .Y(_1568_));
 sg13g2_nand2_1 _5796_ (.Y(_1569_),
    .A(\i_coord.l_xip.genblk2[0].state.Q ),
    .B(\i_coord.x0[-13] ));
 sg13g2_xnor2_1 _5797_ (.Y(_1570_),
    .A(\i_coord.l_xip.genblk2[0].state.Q ),
    .B(\i_coord.x0[-13] ));
 sg13g2_a21oi_1 _5798_ (.A1(net795),
    .A2(_1570_),
    .Y(_1571_),
    .B1(_1567_));
 sg13g2_a22oi_1 _5799_ (.Y(_1572_),
    .B1(_1568_),
    .B2(_1571_),
    .A2(net869),
    .A1(\i_coord.x0[-13] ));
 sg13g2_a21oi_1 _5800_ (.A1(net795),
    .A2(_1572_),
    .Y(_1573_),
    .B1(_1567_));
 sg13g2_nand3_1 _5801_ (.B(net751),
    .C(_1573_),
    .A(net771),
    .Y(_1574_));
 sg13g2_o21ai_1 _5802_ (.B1(_1574_),
    .Y(_0099_),
    .A1(_3139_),
    .A2(net751));
 sg13g2_nand2_1 _5803_ (.Y(_1575_),
    .A(net271),
    .B(net799));
 sg13g2_xor2_1 _5804_ (.B(\i_coord.x0[-12] ),
    .A(\i_coord.l_xip.genblk2[1].state.Q ),
    .X(_1576_));
 sg13g2_nor2b_1 _5805_ (.A(_1569_),
    .B_N(_1576_),
    .Y(_1577_));
 sg13g2_xor2_1 _5806_ (.B(_1576_),
    .A(_1569_),
    .X(_1578_));
 sg13g2_o21ai_1 _5807_ (.B1(_1575_),
    .Y(_1579_),
    .A1(net799),
    .A2(_1578_));
 sg13g2_a22oi_1 _5808_ (.Y(_1580_),
    .B1(_1568_),
    .B2(_1579_),
    .A2(net869),
    .A1(\i_coord.x0[-12] ));
 sg13g2_o21ai_1 _5809_ (.B1(_1575_),
    .Y(_1581_),
    .A1(net799),
    .A2(_1580_));
 sg13g2_nand3_1 _5810_ (.B(net750),
    .C(_1581_),
    .A(net771),
    .Y(_1582_));
 sg13g2_o21ai_1 _5811_ (.B1(_1582_),
    .Y(_0100_),
    .A1(_3141_),
    .A2(net750));
 sg13g2_nand2_1 _5812_ (.Y(_1583_),
    .A(\i_coord.x_row_start[-11] ),
    .B(net798));
 sg13g2_xnor2_1 _5813_ (.Y(_1584_),
    .A(\i_coord.l_xip.genblk2[2].state.Q ),
    .B(\i_coord.x0[-11] ));
 sg13g2_a21oi_1 _5814_ (.A1(\i_coord.l_xip.genblk2[1].state.Q ),
    .A2(\i_coord.x0[-12] ),
    .Y(_1585_),
    .B1(_1577_));
 sg13g2_nor2_1 _5815_ (.A(_1584_),
    .B(_1585_),
    .Y(_1586_));
 sg13g2_a21o_1 _5816_ (.A2(_1585_),
    .A1(_1584_),
    .B1(net798),
    .X(_1587_));
 sg13g2_o21ai_1 _5817_ (.B1(_1583_),
    .Y(_1588_),
    .A1(_1586_),
    .A2(_1587_));
 sg13g2_nand2_1 _5818_ (.Y(_1589_),
    .A(_1568_),
    .B(_1588_));
 sg13g2_o21ai_1 _5819_ (.B1(_1589_),
    .Y(_1590_),
    .A1(_3142_),
    .A2(net875));
 sg13g2_mux2_1 _5820_ (.A0(net247),
    .A1(_1590_),
    .S(net795),
    .X(_1591_));
 sg13g2_nand3_1 _5821_ (.B(net750),
    .C(_1591_),
    .A(net771),
    .Y(_1592_));
 sg13g2_o21ai_1 _5822_ (.B1(_1592_),
    .Y(_0101_),
    .A1(_3142_),
    .A2(net750));
 sg13g2_a21oi_1 _5823_ (.A1(\i_coord.l_xip.genblk2[2].state.Q ),
    .A2(\i_coord.x0[-11] ),
    .Y(_1593_),
    .B1(_1586_));
 sg13g2_nand2_1 _5824_ (.Y(_1594_),
    .A(\i_coord.l_xip.genblk2[3].state.Q ),
    .B(\i_coord.x0[-10] ));
 sg13g2_xnor2_1 _5825_ (.Y(_1595_),
    .A(\i_coord.l_xip.genblk2[3].state.Q ),
    .B(\i_coord.x0[-10] ));
 sg13g2_xnor2_1 _5826_ (.Y(_1596_),
    .A(_1593_),
    .B(_1595_));
 sg13g2_a221oi_1 _5827_ (.B2(_1596_),
    .C1(net780),
    .B1(net792),
    .A1(_3098_),
    .Y(_1597_),
    .A2(net798));
 sg13g2_a21oi_1 _5828_ (.A1(\i_coord.l_xl.genblk2[3].state.Q ),
    .A2(net782),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_nor2_1 _5829_ (.A(\i_coord.x0[-10] ),
    .B(net878),
    .Y(_1599_));
 sg13g2_a21oi_1 _5830_ (.A1(net873),
    .A2(_1598_),
    .Y(_1600_),
    .B1(_1599_));
 sg13g2_a21oi_1 _5831_ (.A1(net763),
    .A2(_1598_),
    .Y(_1601_),
    .B1(net748));
 sg13g2_o21ai_1 _5832_ (.B1(_1601_),
    .Y(_1602_),
    .A1(net763),
    .A2(_1600_));
 sg13g2_o21ai_1 _5833_ (.B1(_1602_),
    .Y(_0102_),
    .A1(_3143_),
    .A2(net753));
 sg13g2_o21ai_1 _5834_ (.B1(_1594_),
    .Y(_1603_),
    .A1(_1593_),
    .A2(_1595_));
 sg13g2_and2_1 _5835_ (.A(\i_coord.l_xip.genblk2[4].state.Q ),
    .B(\i_coord.x0[-9] ),
    .X(_1604_));
 sg13g2_xor2_1 _5836_ (.B(\i_coord.x0[-9] ),
    .A(\i_coord.l_xip.genblk2[4].state.Q ),
    .X(_1605_));
 sg13g2_xnor2_1 _5837_ (.Y(_1606_),
    .A(_1603_),
    .B(_1605_));
 sg13g2_o21ai_1 _5838_ (.B1(net769),
    .Y(_1607_),
    .A1(\i_coord.x_row_start[-9] ),
    .A2(net794));
 sg13g2_a21o_1 _5839_ (.A2(_1606_),
    .A1(net791),
    .B1(_1607_),
    .X(_1608_));
 sg13g2_a21oi_1 _5840_ (.A1(\i_coord.l_xl.genblk2[4].state.Q ),
    .A2(net780),
    .Y(_1609_),
    .B1(net869));
 sg13g2_nand2_1 _5841_ (.Y(_1610_),
    .A(_1608_),
    .B(_1609_));
 sg13g2_o21ai_1 _5842_ (.B1(_1610_),
    .Y(_1611_),
    .A1(\i_coord.x0[-9] ),
    .A2(net873));
 sg13g2_a221oi_1 _5843_ (.B2(net761),
    .C1(net746),
    .B1(_1611_),
    .A1(_1329_),
    .Y(_1612_),
    .A2(_1608_));
 sg13g2_a21o_1 _5844_ (.A2(net746),
    .A1(net287),
    .B1(_1612_),
    .X(_0103_));
 sg13g2_a21o_1 _5845_ (.A2(_1605_),
    .A1(_1603_),
    .B1(_1604_),
    .X(_1613_));
 sg13g2_nand2_1 _5846_ (.Y(_1614_),
    .A(\i_coord.l_xip.genblk2[5].state.Q ),
    .B(\i_coord.x0[-8] ));
 sg13g2_xor2_1 _5847_ (.B(\i_coord.x0[-8] ),
    .A(\i_coord.l_xip.genblk2[5].state.Q ),
    .X(_1615_));
 sg13g2_xnor2_1 _5848_ (.Y(_1616_),
    .A(_1613_),
    .B(_1615_));
 sg13g2_o21ai_1 _5849_ (.B1(net769),
    .Y(_1617_),
    .A1(\i_coord.x_row_start[-8] ),
    .A2(net793));
 sg13g2_a21o_1 _5850_ (.A2(_1616_),
    .A1(net794),
    .B1(_1617_),
    .X(_1618_));
 sg13g2_a21oi_1 _5851_ (.A1(\i_coord.l_xl.genblk2[5].state.Q ),
    .A2(net780),
    .Y(_1619_),
    .B1(net868));
 sg13g2_nand2_1 _5852_ (.Y(_1620_),
    .A(_1618_),
    .B(_1619_));
 sg13g2_o21ai_1 _5853_ (.B1(_1620_),
    .Y(_1621_),
    .A1(\i_coord.x0[-8] ),
    .A2(net873));
 sg13g2_a221oi_1 _5854_ (.B2(net761),
    .C1(net746),
    .B1(_1621_),
    .A1(_1335_),
    .Y(_1622_),
    .A2(_1618_));
 sg13g2_a21o_1 _5855_ (.A2(net746),
    .A1(net306),
    .B1(_1622_),
    .X(_0104_));
 sg13g2_xnor2_1 _5856_ (.Y(_1623_),
    .A(\i_coord.l_xip.genblk2[6].state.Q ),
    .B(\i_coord.x0[-7] ));
 sg13g2_o21ai_1 _5857_ (.B1(_1613_),
    .Y(_1624_),
    .A1(\i_coord.l_xip.genblk2[5].state.Q ),
    .A2(\i_coord.x0[-8] ));
 sg13g2_and3_1 _5858_ (.X(_1625_),
    .A(_1614_),
    .B(_1623_),
    .C(_1624_));
 sg13g2_a21oi_1 _5859_ (.A1(_1614_),
    .A2(_1624_),
    .Y(_1626_),
    .B1(_1623_));
 sg13g2_or2_1 _5860_ (.X(_1627_),
    .B(_1626_),
    .A(_1625_));
 sg13g2_o21ai_1 _5861_ (.B1(net769),
    .Y(_1628_),
    .A1(\i_coord.x_row_start[-7] ),
    .A2(net793));
 sg13g2_a21o_1 _5862_ (.A2(_1627_),
    .A1(net791),
    .B1(_1628_),
    .X(_1629_));
 sg13g2_a21oi_1 _5863_ (.A1(\i_coord.l_xl.genblk2[6].state.Q ),
    .A2(net779),
    .Y(_1630_),
    .B1(net868));
 sg13g2_nand2_1 _5864_ (.Y(_1631_),
    .A(_1629_),
    .B(_1630_));
 sg13g2_o21ai_1 _5865_ (.B1(_1631_),
    .Y(_1632_),
    .A1(\i_coord.x0[-7] ),
    .A2(net873));
 sg13g2_a221oi_1 _5866_ (.B2(net759),
    .C1(net746),
    .B1(_1632_),
    .A1(_1342_),
    .Y(_1633_),
    .A2(_1629_));
 sg13g2_a21o_1 _5867_ (.A2(net746),
    .A1(net303),
    .B1(_1633_),
    .X(_0105_));
 sg13g2_nand2_1 _5868_ (.Y(_1634_),
    .A(net240),
    .B(net749));
 sg13g2_a21oi_1 _5869_ (.A1(\i_coord.l_xip.genblk2[6].state.Q ),
    .A2(\i_coord.x0[-7] ),
    .Y(_1635_),
    .B1(_1626_));
 sg13g2_nand2_1 _5870_ (.Y(_1636_),
    .A(\i_coord.l_xip.genblk2[7].state.Q ),
    .B(\i_coord.x0[-6] ));
 sg13g2_xnor2_1 _5871_ (.Y(_1637_),
    .A(\i_coord.l_xip.genblk2[7].state.Q ),
    .B(\i_coord.x0[-6] ));
 sg13g2_xnor2_1 _5872_ (.Y(_1638_),
    .A(_1635_),
    .B(_1637_));
 sg13g2_a221oi_1 _5873_ (.B2(_1638_),
    .C1(net779),
    .B1(net792),
    .A1(_3103_),
    .Y(_1639_),
    .A2(net801));
 sg13g2_a21o_1 _5874_ (.A2(net779),
    .A1(\i_coord.l_xl.genblk2[7].state.Q ),
    .B1(_1639_),
    .X(_1640_));
 sg13g2_nor2_1 _5875_ (.A(net868),
    .B(_1640_),
    .Y(_1641_));
 sg13g2_a21oi_1 _5876_ (.A1(_3144_),
    .A2(net868),
    .Y(_1642_),
    .B1(_1641_));
 sg13g2_nand2_1 _5877_ (.Y(_1643_),
    .A(net841),
    .B(_1642_));
 sg13g2_nor2_1 _5878_ (.A(net759),
    .B(_1640_),
    .Y(_1644_));
 sg13g2_o21ai_1 _5879_ (.B1(net753),
    .Y(_1645_),
    .A1(net763),
    .A2(_1642_));
 sg13g2_o21ai_1 _5880_ (.B1(_1634_),
    .Y(_0106_),
    .A1(_1644_),
    .A2(_1645_));
 sg13g2_and2_1 _5881_ (.A(\i_coord.l_xip.genblk2[8].state.Q ),
    .B(\i_coord.x0[-5] ),
    .X(_1646_));
 sg13g2_xor2_1 _5882_ (.B(\i_coord.x0[-5] ),
    .A(\i_coord.l_xip.genblk2[8].state.Q ),
    .X(_1647_));
 sg13g2_o21ai_1 _5883_ (.B1(_1636_),
    .Y(_1648_),
    .A1(_1635_),
    .A2(_1637_));
 sg13g2_xnor2_1 _5884_ (.Y(_1649_),
    .A(_1647_),
    .B(_1648_));
 sg13g2_o21ai_1 _5885_ (.B1(net769),
    .Y(_1650_),
    .A1(\i_coord.x_row_start[-5] ),
    .A2(net793));
 sg13g2_a21o_1 _5886_ (.A2(_1649_),
    .A1(net791),
    .B1(_1650_),
    .X(_1651_));
 sg13g2_a21oi_1 _5887_ (.A1(\i_coord.l_xl.genblk2[8].state.Q ),
    .A2(net779),
    .Y(_1652_),
    .B1(net868));
 sg13g2_nand2_1 _5888_ (.Y(_1653_),
    .A(_1651_),
    .B(_1652_));
 sg13g2_o21ai_1 _5889_ (.B1(_1653_),
    .Y(_1654_),
    .A1(\i_coord.x0[-5] ),
    .A2(net871));
 sg13g2_a221oi_1 _5890_ (.B2(net759),
    .C1(net744),
    .B1(_1654_),
    .A1(_1354_),
    .Y(_1655_),
    .A2(_1651_));
 sg13g2_a21o_1 _5891_ (.A2(net745),
    .A1(net301),
    .B1(_1655_),
    .X(_0107_));
 sg13g2_xnor2_1 _5892_ (.Y(_1656_),
    .A(net789),
    .B(\i_coord.x0[-4] ));
 sg13g2_a21o_1 _5893_ (.A2(_1648_),
    .A1(_1647_),
    .B1(_1646_),
    .X(_1657_));
 sg13g2_o21ai_1 _5894_ (.B1(net793),
    .Y(_1658_),
    .A1(_1656_),
    .A2(_1657_));
 sg13g2_a21oi_1 _5895_ (.A1(_1656_),
    .A2(_1657_),
    .Y(_1659_),
    .B1(_1658_));
 sg13g2_o21ai_1 _5896_ (.B1(net769),
    .Y(_1660_),
    .A1(\i_coord.x_row_start[-4] ),
    .A2(net793));
 sg13g2_nor2_1 _5897_ (.A(_1659_),
    .B(_1660_),
    .Y(_1661_));
 sg13g2_inv_1 _5898_ (.Y(_1662_),
    .A(_1661_));
 sg13g2_a21oi_1 _5899_ (.A1(\i_coord.l_xl.genblk2[9].state.Q ),
    .A2(net777),
    .Y(_1663_),
    .B1(_1661_));
 sg13g2_nand2_1 _5900_ (.Y(_1664_),
    .A(net871),
    .B(_1663_));
 sg13g2_o21ai_1 _5901_ (.B1(_1664_),
    .Y(_1665_),
    .A1(\i_coord.x0[-4] ),
    .A2(net871));
 sg13g2_a221oi_1 _5902_ (.B2(net759),
    .C1(net745),
    .B1(_1665_),
    .A1(_1359_),
    .Y(_1666_),
    .A2(_1662_));
 sg13g2_a21o_1 _5903_ (.A2(net745),
    .A1(net312),
    .B1(_1666_),
    .X(_0108_));
 sg13g2_nand2_1 _5904_ (.Y(_1667_),
    .A(net789),
    .B(\i_coord.x0[-3] ));
 sg13g2_xor2_1 _5905_ (.B(\i_coord.x0[-3] ),
    .A(net789),
    .X(_1668_));
 sg13g2_o21ai_1 _5906_ (.B1(_1657_),
    .Y(_1669_),
    .A1(net789),
    .A2(\i_coord.x0[-4] ));
 sg13g2_inv_1 _5907_ (.Y(_1670_),
    .A(_1669_));
 sg13g2_a21oi_1 _5908_ (.A1(net789),
    .A2(\i_coord.x0[-4] ),
    .Y(_1671_),
    .B1(_1670_));
 sg13g2_nand2b_1 _5909_ (.Y(_1672_),
    .B(_1668_),
    .A_N(_1671_));
 sg13g2_xor2_1 _5910_ (.B(_1671_),
    .A(_1668_),
    .X(_1673_));
 sg13g2_a221oi_1 _5911_ (.B2(_1673_),
    .C1(net778),
    .B1(net791),
    .A1(_3106_),
    .Y(_1674_),
    .A2(net801));
 sg13g2_a21oi_1 _5912_ (.A1(\i_coord.l_xl.genblk2[10].state.Q ),
    .A2(net777),
    .Y(_1675_),
    .B1(_1674_));
 sg13g2_nand2_1 _5913_ (.Y(_1676_),
    .A(net871),
    .B(_1675_));
 sg13g2_o21ai_1 _5914_ (.B1(_1676_),
    .Y(_1677_),
    .A1(\i_coord.x0[-3] ),
    .A2(net870));
 sg13g2_nand2_1 _5915_ (.Y(_1678_),
    .A(net757),
    .B(_1677_));
 sg13g2_a21oi_1 _5916_ (.A1(_3266_),
    .A2(_1675_),
    .Y(_1679_),
    .B1(net745));
 sg13g2_a22oi_1 _5917_ (.Y(_1680_),
    .B1(_1678_),
    .B2(_1679_),
    .A2(net745),
    .A1(net310));
 sg13g2_inv_1 _5918_ (.Y(_0109_),
    .A(_1680_));
 sg13g2_nor2_1 _5919_ (.A(net789),
    .B(\i_coord.x0[-2] ),
    .Y(_1681_));
 sg13g2_xor2_1 _5920_ (.B(\i_coord.x0[-2] ),
    .A(net788),
    .X(_1682_));
 sg13g2_nand3_1 _5921_ (.B(_1672_),
    .C(_1682_),
    .A(_1667_),
    .Y(_1683_));
 sg13g2_a21oi_1 _5922_ (.A1(_1667_),
    .A2(_1672_),
    .Y(_1684_),
    .B1(_1682_));
 sg13g2_nor2_1 _5923_ (.A(net801),
    .B(_1684_),
    .Y(_1685_));
 sg13g2_a221oi_1 _5924_ (.B2(_1685_),
    .C1(net776),
    .B1(_1683_),
    .A1(_3107_),
    .Y(_1686_),
    .A2(_3263_));
 sg13g2_inv_1 _5925_ (.Y(_1687_),
    .A(_1686_));
 sg13g2_a21oi_1 _5926_ (.A1(\i_coord.l_xl.genblk2[11].state.Q ),
    .A2(net777),
    .Y(_1688_),
    .B1(_1686_));
 sg13g2_nand2_1 _5927_ (.Y(_1689_),
    .A(net870),
    .B(_1688_));
 sg13g2_o21ai_1 _5928_ (.B1(_1689_),
    .Y(_1690_),
    .A1(\i_coord.x0[-2] ),
    .A2(net870));
 sg13g2_a221oi_1 _5929_ (.B2(net758),
    .C1(net744),
    .B1(_1690_),
    .A1(_1371_),
    .Y(_1691_),
    .A2(_1687_));
 sg13g2_a21o_1 _5930_ (.A2(net744),
    .A1(net311),
    .B1(_1691_),
    .X(_0110_));
 sg13g2_xor2_1 _5931_ (.B(\i_coord.x0[-1] ),
    .A(net788),
    .X(_1692_));
 sg13g2_o21ai_1 _5932_ (.B1(net789),
    .Y(_1693_),
    .A1(\i_coord.x0[-3] ),
    .A2(\i_coord.x0[-2] ));
 sg13g2_o21ai_1 _5933_ (.B1(_1693_),
    .Y(_1694_),
    .A1(_1672_),
    .A2(_1681_));
 sg13g2_and2_1 _5934_ (.A(_1692_),
    .B(_1694_),
    .X(_1695_));
 sg13g2_xnor2_1 _5935_ (.Y(_1696_),
    .A(_1692_),
    .B(_1694_));
 sg13g2_a221oi_1 _5936_ (.B2(_1696_),
    .C1(net776),
    .B1(net791),
    .A1(_3108_),
    .Y(_1697_),
    .A2(net801));
 sg13g2_a21o_1 _5937_ (.A2(net776),
    .A1(\i_coord.l_xl.genblk2[12].state.Q ),
    .B1(_1697_),
    .X(_1698_));
 sg13g2_nand2b_1 _5938_ (.Y(_1699_),
    .B(net868),
    .A_N(\i_coord.x0[-1] ));
 sg13g2_o21ai_1 _5939_ (.B1(_1699_),
    .Y(_1700_),
    .A1(net868),
    .A2(_1698_));
 sg13g2_o21ai_1 _5940_ (.B1(net753),
    .Y(_1701_),
    .A1(net757),
    .A2(_1698_));
 sg13g2_a21oi_1 _5941_ (.A1(net757),
    .A2(_1700_),
    .Y(_1702_),
    .B1(_1701_));
 sg13g2_a21o_1 _5942_ (.A2(net744),
    .A1(net313),
    .B1(_1702_),
    .X(_0111_));
 sg13g2_xor2_1 _5943_ (.B(\i_coord.x0[0] ),
    .A(net788),
    .X(_1703_));
 sg13g2_a21oi_1 _5944_ (.A1(net788),
    .A2(\i_coord.x0[-1] ),
    .Y(_1704_),
    .B1(_1695_));
 sg13g2_o21ai_1 _5945_ (.B1(net793),
    .Y(_1705_),
    .A1(_1703_),
    .A2(_1704_));
 sg13g2_a21oi_1 _5946_ (.A1(_1703_),
    .A2(_1704_),
    .Y(_1706_),
    .B1(_1705_));
 sg13g2_o21ai_1 _5947_ (.B1(net769),
    .Y(_1707_),
    .A1(\i_coord.x_row_start[0] ),
    .A2(net793));
 sg13g2_nor2_1 _5948_ (.A(_1706_),
    .B(_1707_),
    .Y(_1708_));
 sg13g2_inv_1 _5949_ (.Y(_1709_),
    .A(_1708_));
 sg13g2_a21oi_1 _5950_ (.A1(\i_coord.l_xl.genblk2[13].state.Q ),
    .A2(net776),
    .Y(_1710_),
    .B1(_1708_));
 sg13g2_nand2_1 _5951_ (.Y(_1711_),
    .A(net870),
    .B(_1710_));
 sg13g2_o21ai_1 _5952_ (.B1(_1711_),
    .Y(_1712_),
    .A1(\i_coord.x0[0] ),
    .A2(net870));
 sg13g2_a221oi_1 _5953_ (.B2(net757),
    .C1(net744),
    .B1(_1712_),
    .A1(_1383_),
    .Y(_1713_),
    .A2(_1709_));
 sg13g2_a21o_1 _5954_ (.A2(net744),
    .A1(net302),
    .B1(_1713_),
    .X(_0112_));
 sg13g2_xnor2_1 _5955_ (.Y(_1714_),
    .A(net788),
    .B(\i_coord.x0[1] ));
 sg13g2_nand2_1 _5956_ (.Y(_1715_),
    .A(_1695_),
    .B(_1703_));
 sg13g2_o21ai_1 _5957_ (.B1(net788),
    .Y(_1716_),
    .A1(\i_coord.x0[-1] ),
    .A2(\i_coord.x0[0] ));
 sg13g2_and3_1 _5958_ (.X(_1717_),
    .A(_1714_),
    .B(_1715_),
    .C(_1716_));
 sg13g2_a21oi_1 _5959_ (.A1(_1715_),
    .A2(_1716_),
    .Y(_1718_),
    .B1(_1714_));
 sg13g2_or2_1 _5960_ (.X(_1719_),
    .B(_1718_),
    .A(_1717_));
 sg13g2_a221oi_1 _5961_ (.B2(_1719_),
    .C1(net775),
    .B1(net791),
    .A1(_3110_),
    .Y(_1720_),
    .A2(net801));
 sg13g2_inv_1 _5962_ (.Y(_1721_),
    .A(_1720_));
 sg13g2_a21oi_1 _5963_ (.A1(\i_coord.l_xl.genblk2[14].state.Q ),
    .A2(net775),
    .Y(_1722_),
    .B1(_1720_));
 sg13g2_nand2_1 _5964_ (.Y(_1723_),
    .A(net870),
    .B(_1722_));
 sg13g2_o21ai_1 _5965_ (.B1(_1723_),
    .Y(_1724_),
    .A1(\i_coord.x0[1] ),
    .A2(net870));
 sg13g2_nor2_1 _5966_ (.A(net831),
    .B(_1724_),
    .Y(_1725_));
 sg13g2_a221oi_1 _5967_ (.B2(net757),
    .C1(net744),
    .B1(_1724_),
    .A1(_1390_),
    .Y(_1726_),
    .A2(_1721_));
 sg13g2_a21o_1 _5968_ (.A2(net744),
    .A1(net297),
    .B1(_1726_),
    .X(_0113_));
 sg13g2_a21oi_1 _5969_ (.A1(net788),
    .A2(\i_coord.x0[1] ),
    .Y(_1727_),
    .B1(_1718_));
 sg13g2_xor2_1 _5970_ (.B(\i_coord.x0[2] ),
    .A(net788),
    .X(_1728_));
 sg13g2_a21oi_1 _5971_ (.A1(_1727_),
    .A2(_1728_),
    .Y(_1729_),
    .B1(net801));
 sg13g2_o21ai_1 _5972_ (.B1(_1729_),
    .Y(_1730_),
    .A1(_1727_),
    .A2(_1728_));
 sg13g2_o21ai_1 _5973_ (.B1(net769),
    .Y(_1731_),
    .A1(\i_coord.x_row_start[2] ),
    .A2(net793));
 sg13g2_nand2b_1 _5974_ (.Y(_1732_),
    .B(_1730_),
    .A_N(_1731_));
 sg13g2_a21oi_1 _5975_ (.A1(\i_coord.l_xl.genblk2[15].state.Q ),
    .A2(net775),
    .Y(_1733_),
    .B1(net868));
 sg13g2_nand2_1 _5976_ (.Y(_1734_),
    .A(_1732_),
    .B(_1733_));
 sg13g2_o21ai_1 _5977_ (.B1(_1734_),
    .Y(_1735_),
    .A1(\i_coord.x0[2] ),
    .A2(net870));
 sg13g2_a22oi_1 _5978_ (.Y(_1736_),
    .B1(_1735_),
    .B2(net757),
    .A2(_1732_),
    .A1(_1395_));
 sg13g2_mux2_1 _5979_ (.A0(net260),
    .A1(_1736_),
    .S(net753),
    .X(_0114_));
 sg13g2_nand2b_1 _5980_ (.Y(_1737_),
    .B(net799),
    .A_N(\i_coord.y_row_start[-13] ));
 sg13g2_nand2_1 _5981_ (.Y(_1738_),
    .A(\i_coord.y0[-13] ),
    .B(\i_coord.l_yip.genblk2[0].state.Q ));
 sg13g2_xnor2_1 _5982_ (.Y(_1739_),
    .A(\i_coord.y0[-13] ),
    .B(\i_coord.l_yip.genblk2[0].state.Q ));
 sg13g2_a21oi_1 _5983_ (.A1(net795),
    .A2(_1739_),
    .Y(_1740_),
    .B1(net782));
 sg13g2_a22oi_1 _5984_ (.Y(_1741_),
    .B1(_1737_),
    .B2(_1740_),
    .A2(net782),
    .A1(\i_coord.l_yt.genblk2[0].state.Q ));
 sg13g2_nor2_1 _5985_ (.A(net246),
    .B(net875),
    .Y(_1742_));
 sg13g2_a21oi_1 _5986_ (.A1(net874),
    .A2(_1741_),
    .Y(_1743_),
    .B1(_1742_));
 sg13g2_o21ai_1 _5987_ (.B1(net750),
    .Y(_1744_),
    .A1(net761),
    .A2(_1741_));
 sg13g2_a21oi_1 _5988_ (.A1(net766),
    .A2(_1743_),
    .Y(_1745_),
    .B1(_1744_));
 sg13g2_a21oi_1 _5989_ (.A1(_3116_),
    .A2(net748),
    .Y(_0115_),
    .B1(_1745_));
 sg13g2_nor2_1 _5990_ (.A(net250),
    .B(net874),
    .Y(_1746_));
 sg13g2_nand2_1 _5991_ (.Y(_1747_),
    .A(\i_coord.y0[-12] ),
    .B(\i_coord.l_yip.genblk2[1].state.Q ));
 sg13g2_xnor2_1 _5992_ (.Y(_1748_),
    .A(\i_coord.y0[-12] ),
    .B(\i_coord.l_yip.genblk2[1].state.Q ));
 sg13g2_or2_1 _5993_ (.X(_1749_),
    .B(_1748_),
    .A(_1738_));
 sg13g2_xnor2_1 _5994_ (.Y(_1750_),
    .A(_1738_),
    .B(_1748_));
 sg13g2_a21oi_1 _5995_ (.A1(\i_coord.y_row_start[-12] ),
    .A2(net800),
    .Y(_1751_),
    .B1(net785));
 sg13g2_o21ai_1 _5996_ (.B1(_1751_),
    .Y(_1752_),
    .A1(net800),
    .A2(_1750_));
 sg13g2_o21ai_1 _5997_ (.B1(_1752_),
    .Y(_1753_),
    .A1(\i_coord.l_yt.genblk2[1].state.Q ),
    .A2(net772));
 sg13g2_a21oi_1 _5998_ (.A1(net874),
    .A2(_1753_),
    .Y(_1754_),
    .B1(_1746_));
 sg13g2_o21ai_1 _5999_ (.B1(net750),
    .Y(_1755_),
    .A1(net766),
    .A2(_1753_));
 sg13g2_a21oi_1 _6000_ (.A1(net766),
    .A2(_1754_),
    .Y(_1756_),
    .B1(_1755_));
 sg13g2_a21oi_1 _6001_ (.A1(_3117_),
    .A2(net748),
    .Y(_0116_),
    .B1(_1756_));
 sg13g2_and2_1 _6002_ (.A(\i_coord.y0[-11] ),
    .B(\i_coord.l_yip.genblk2[2].state.Q ),
    .X(_1757_));
 sg13g2_xnor2_1 _6003_ (.Y(_1758_),
    .A(\i_coord.y0[-11] ),
    .B(\i_coord.l_yip.genblk2[2].state.Q ));
 sg13g2_and3_1 _6004_ (.X(_1759_),
    .A(_1747_),
    .B(_1749_),
    .C(_1758_));
 sg13g2_a21oi_1 _6005_ (.A1(_1747_),
    .A2(_1749_),
    .Y(_1760_),
    .B1(_1758_));
 sg13g2_or2_1 _6006_ (.X(_1761_),
    .B(_1760_),
    .A(_1759_));
 sg13g2_a21oi_1 _6007_ (.A1(\i_coord.y_row_start[-11] ),
    .A2(net799),
    .Y(_1762_),
    .B1(net785));
 sg13g2_o21ai_1 _6008_ (.B1(_1762_),
    .Y(_1763_),
    .A1(_3263_),
    .A2(_1761_));
 sg13g2_o21ai_1 _6009_ (.B1(_1763_),
    .Y(_1764_),
    .A1(\i_coord.l_yt.genblk2[2].state.Q ),
    .A2(net772));
 sg13g2_nand2_1 _6010_ (.Y(_1765_),
    .A(net874),
    .B(_1764_));
 sg13g2_o21ai_1 _6011_ (.B1(_1765_),
    .Y(_1766_),
    .A1(\i_coord.y0[-11] ),
    .A2(net874));
 sg13g2_nand2_1 _6012_ (.Y(_1767_),
    .A(net766),
    .B(_1766_));
 sg13g2_a21oi_1 _6013_ (.A1(net762),
    .A2(_1764_),
    .Y(_1768_),
    .B1(net748));
 sg13g2_a22oi_1 _6014_ (.Y(_1769_),
    .B1(_1767_),
    .B2(_1768_),
    .A2(net748),
    .A1(net325));
 sg13g2_inv_1 _6015_ (.Y(_0117_),
    .A(_1769_));
 sg13g2_nand2_1 _6016_ (.Y(_1770_),
    .A(\i_coord.y0[-10] ),
    .B(\i_coord.l_yip.genblk2[3].state.Q ));
 sg13g2_xor2_1 _6017_ (.B(\i_coord.l_yip.genblk2[3].state.Q ),
    .A(\i_coord.y0[-10] ),
    .X(_1771_));
 sg13g2_o21ai_1 _6018_ (.B1(_1771_),
    .Y(_1772_),
    .A1(_1757_),
    .A2(_1760_));
 sg13g2_or3_1 _6019_ (.A(_1757_),
    .B(_1760_),
    .C(_1771_),
    .X(_1773_));
 sg13g2_nand3_1 _6020_ (.B(_1772_),
    .C(_1773_),
    .A(net795),
    .Y(_1774_));
 sg13g2_nand2_1 _6021_ (.Y(_1775_),
    .A(\i_coord.y_row_start[-10] ),
    .B(net799));
 sg13g2_nand3_1 _6022_ (.B(_1774_),
    .C(_1775_),
    .A(net772),
    .Y(_1776_));
 sg13g2_o21ai_1 _6023_ (.B1(_1776_),
    .Y(_1777_),
    .A1(\i_coord.l_yt.genblk2[3].state.Q ),
    .A2(net771));
 sg13g2_nor2_1 _6024_ (.A(\i_coord.y0[-10] ),
    .B(net874),
    .Y(_1778_));
 sg13g2_a21oi_1 _6025_ (.A1(net874),
    .A2(_1777_),
    .Y(_1779_),
    .B1(_1778_));
 sg13g2_o21ai_1 _6026_ (.B1(net750),
    .Y(_1780_),
    .A1(net761),
    .A2(_1777_));
 sg13g2_a21oi_1 _6027_ (.A1(net766),
    .A2(_1779_),
    .Y(_1781_),
    .B1(_1780_));
 sg13g2_a21oi_1 _6028_ (.A1(_3118_),
    .A2(net748),
    .Y(_0118_),
    .B1(_1781_));
 sg13g2_nor2_1 _6029_ (.A(\i_coord.y0[-9] ),
    .B(net875),
    .Y(_1782_));
 sg13g2_xnor2_1 _6030_ (.Y(_1783_),
    .A(\i_coord.y0[-9] ),
    .B(\i_coord.l_yip.genblk2[4].state.Q ));
 sg13g2_a21oi_1 _6031_ (.A1(_1770_),
    .A2(_1772_),
    .Y(_1784_),
    .B1(_1783_));
 sg13g2_and3_1 _6032_ (.X(_1785_),
    .A(_1770_),
    .B(_1772_),
    .C(_1783_));
 sg13g2_o21ai_1 _6033_ (.B1(net797),
    .Y(_1786_),
    .A1(_1784_),
    .A2(_1785_));
 sg13g2_o21ai_1 _6034_ (.B1(_1786_),
    .Y(_1787_),
    .A1(\i_coord.y_row_start[-9] ),
    .A2(net795));
 sg13g2_nor2_1 _6035_ (.A(net782),
    .B(_1787_),
    .Y(_1788_));
 sg13g2_a21oi_2 _6036_ (.B1(_1788_),
    .Y(_1789_),
    .A2(net782),
    .A1(\i_coord.l_yt.genblk2[4].state.Q ));
 sg13g2_a21oi_1 _6037_ (.A1(net874),
    .A2(_1789_),
    .Y(_1790_),
    .B1(_1782_));
 sg13g2_o21ai_1 _6038_ (.B1(net750),
    .Y(_1791_),
    .A1(net767),
    .A2(_1789_));
 sg13g2_a21oi_1 _6039_ (.A1(net767),
    .A2(_1790_),
    .Y(_1792_),
    .B1(_1791_));
 sg13g2_a21oi_1 _6040_ (.A1(_3119_),
    .A2(net748),
    .Y(_0119_),
    .B1(_1792_));
 sg13g2_nor2_1 _6041_ (.A(net937),
    .B(net875),
    .Y(_1793_));
 sg13g2_a21o_1 _6042_ (.A2(\i_coord.l_yip.genblk2[4].state.Q ),
    .A1(\i_coord.y0[-9] ),
    .B1(_1784_),
    .X(_1794_));
 sg13g2_nand2_1 _6043_ (.Y(_1795_),
    .A(net937),
    .B(\i_coord.l_yip.genblk2[5].state.Q ));
 sg13g2_xor2_1 _6044_ (.B(\i_coord.l_yip.genblk2[5].state.Q ),
    .A(net937),
    .X(_1796_));
 sg13g2_o21ai_1 _6045_ (.B1(net797),
    .Y(_1797_),
    .A1(_1794_),
    .A2(_1796_));
 sg13g2_a21oi_1 _6046_ (.A1(_1794_),
    .A2(_1796_),
    .Y(_1798_),
    .B1(_1797_));
 sg13g2_a21oi_1 _6047_ (.A1(\i_coord.y_row_start[-8] ),
    .A2(net800),
    .Y(_1799_),
    .B1(net782));
 sg13g2_nand2b_1 _6048_ (.Y(_1800_),
    .B(_1799_),
    .A_N(_1798_));
 sg13g2_o21ai_1 _6049_ (.B1(_1800_),
    .Y(_1801_),
    .A1(\i_coord.l_yt.genblk2[5].state.Q ),
    .A2(net771));
 sg13g2_a21oi_1 _6050_ (.A1(net875),
    .A2(_1801_),
    .Y(_1802_),
    .B1(_1793_));
 sg13g2_o21ai_1 _6051_ (.B1(net751),
    .Y(_1803_),
    .A1(net767),
    .A2(_1801_));
 sg13g2_a21oi_1 _6052_ (.A1(net767),
    .A2(_1802_),
    .Y(_1804_),
    .B1(_1803_));
 sg13g2_a21oi_1 _6053_ (.A1(_3120_),
    .A2(net748),
    .Y(_0120_),
    .B1(_1804_));
 sg13g2_nor2_1 _6054_ (.A(\i_coord.l_yt.genblk2[6].state.Q ),
    .B(net773),
    .Y(_1805_));
 sg13g2_nand2_1 _6055_ (.Y(_1806_),
    .A(\i_coord.y0[-7] ),
    .B(\i_coord.l_yip.genblk2[6].state.Q ));
 sg13g2_xnor2_1 _6056_ (.Y(_1807_),
    .A(\i_coord.y0[-7] ),
    .B(\i_coord.l_yip.genblk2[6].state.Q ));
 sg13g2_o21ai_1 _6057_ (.B1(_1794_),
    .Y(_1808_),
    .A1(net937),
    .A2(\i_coord.l_yip.genblk2[5].state.Q ));
 sg13g2_a21o_1 _6058_ (.A2(_1808_),
    .A1(_1795_),
    .B1(_1807_),
    .X(_1809_));
 sg13g2_nand3_1 _6059_ (.B(_1807_),
    .C(_1808_),
    .A(_1795_),
    .Y(_1810_));
 sg13g2_nand3_1 _6060_ (.B(_1809_),
    .C(_1810_),
    .A(net796),
    .Y(_1811_));
 sg13g2_a21oi_1 _6061_ (.A1(\i_coord.y_row_start[-7] ),
    .A2(net800),
    .Y(_1812_),
    .B1(net783));
 sg13g2_a21o_1 _6062_ (.A2(_1812_),
    .A1(_1811_),
    .B1(_1805_),
    .X(_1813_));
 sg13g2_nand2_1 _6063_ (.Y(_1814_),
    .A(net876),
    .B(_1813_));
 sg13g2_o21ai_1 _6064_ (.B1(_1814_),
    .Y(_1815_),
    .A1(\i_coord.y0[-7] ),
    .A2(net876));
 sg13g2_nand2_1 _6065_ (.Y(_1816_),
    .A(net767),
    .B(_1815_));
 sg13g2_a21oi_1 _6066_ (.A1(net762),
    .A2(_1813_),
    .Y(_1817_),
    .B1(net747));
 sg13g2_a22oi_1 _6067_ (.Y(_1818_),
    .B1(_1816_),
    .B2(_1817_),
    .A2(net747),
    .A1(net272));
 sg13g2_inv_1 _6068_ (.Y(_0121_),
    .A(_1818_));
 sg13g2_and2_1 _6069_ (.A(_1806_),
    .B(_1809_),
    .X(_1819_));
 sg13g2_xnor2_1 _6070_ (.Y(_1820_),
    .A(\i_coord.y0[-6] ),
    .B(\i_coord.l_yip.genblk2[7].state.Q ));
 sg13g2_or2_1 _6071_ (.X(_1821_),
    .B(_1820_),
    .A(_1819_));
 sg13g2_a21oi_1 _6072_ (.A1(_1819_),
    .A2(_1820_),
    .Y(_1822_),
    .B1(_3258_));
 sg13g2_a22oi_1 _6073_ (.Y(_1823_),
    .B1(_1821_),
    .B2(_1822_),
    .A2(net800),
    .A1(\i_coord.y_row_start[-6] ));
 sg13g2_nand2_1 _6074_ (.Y(_1824_),
    .A(net773),
    .B(_1823_));
 sg13g2_o21ai_1 _6075_ (.B1(_1824_),
    .Y(_1825_),
    .A1(\i_coord.l_yt.genblk2[7].state.Q ),
    .A2(net772));
 sg13g2_nor2_1 _6076_ (.A(\i_coord.y0[-6] ),
    .B(net876),
    .Y(_1826_));
 sg13g2_a21oi_1 _6077_ (.A1(net876),
    .A2(_1825_),
    .Y(_1827_),
    .B1(_1826_));
 sg13g2_a21oi_1 _6078_ (.A1(net763),
    .A2(_1825_),
    .Y(_1828_),
    .B1(net747));
 sg13g2_o21ai_1 _6079_ (.B1(_1828_),
    .Y(_1829_),
    .A1(_3266_),
    .A2(_1827_));
 sg13g2_o21ai_1 _6080_ (.B1(_1829_),
    .Y(_0122_),
    .A1(_3122_),
    .A2(net752));
 sg13g2_and2_1 _6081_ (.A(\i_coord.y0[-5] ),
    .B(\i_coord.l_yip.genblk2[8].state.Q ),
    .X(_1830_));
 sg13g2_xor2_1 _6082_ (.B(\i_coord.l_yip.genblk2[8].state.Q ),
    .A(\i_coord.y0[-5] ),
    .X(_1831_));
 sg13g2_o21ai_1 _6083_ (.B1(_1821_),
    .Y(_1832_),
    .A1(_3122_),
    .A2(_3134_));
 sg13g2_xnor2_1 _6084_ (.Y(_1833_),
    .A(_1831_),
    .B(_1832_));
 sg13g2_o21ai_1 _6085_ (.B1(net773),
    .Y(_1834_),
    .A1(\i_coord.y_row_start[-5] ),
    .A2(net796));
 sg13g2_a21oi_1 _6086_ (.A1(net796),
    .A2(_1833_),
    .Y(_1835_),
    .B1(_1834_));
 sg13g2_a21oi_1 _6087_ (.A1(\i_coord.l_yt.genblk2[8].state.Q ),
    .A2(net783),
    .Y(_1836_),
    .B1(_1835_));
 sg13g2_nor2_1 _6088_ (.A(\i_coord.y0[-5] ),
    .B(net876),
    .Y(_1837_));
 sg13g2_a21oi_1 _6089_ (.A1(net876),
    .A2(_1836_),
    .Y(_1838_),
    .B1(_1837_));
 sg13g2_a21oi_1 _6090_ (.A1(_3261_),
    .A2(_1836_),
    .Y(_1839_),
    .B1(net747));
 sg13g2_o21ai_1 _6091_ (.B1(_1839_),
    .Y(_1840_),
    .A1(_3266_),
    .A2(_1838_));
 sg13g2_o21ai_1 _6092_ (.B1(_1840_),
    .Y(_0123_),
    .A1(_3123_),
    .A2(net752));
 sg13g2_xnor2_1 _6093_ (.Y(_1841_),
    .A(\i_coord.y0[-4] ),
    .B(net803));
 sg13g2_a21o_1 _6094_ (.A2(_1832_),
    .A1(_1831_),
    .B1(_1830_),
    .X(_1842_));
 sg13g2_a21oi_1 _6095_ (.A1(_1841_),
    .A2(_1842_),
    .Y(_1843_),
    .B1(_3258_));
 sg13g2_o21ai_1 _6096_ (.B1(_1843_),
    .Y(_1844_),
    .A1(_1841_),
    .A2(_1842_));
 sg13g2_a21oi_1 _6097_ (.A1(_3112_),
    .A2(net800),
    .Y(_1845_),
    .B1(net783));
 sg13g2_a22oi_1 _6098_ (.Y(_1846_),
    .B1(_1844_),
    .B2(_1845_),
    .A2(net783),
    .A1(\i_coord.l_yt.genblk2[9].state.Q ));
 sg13g2_nor2_1 _6099_ (.A(\i_coord.y0[-4] ),
    .B(net876),
    .Y(_1847_));
 sg13g2_a21oi_1 _6100_ (.A1(net876),
    .A2(_1846_),
    .Y(_1848_),
    .B1(_1847_));
 sg13g2_a21oi_1 _6101_ (.A1(net762),
    .A2(_1846_),
    .Y(_1849_),
    .B1(net749));
 sg13g2_o21ai_1 _6102_ (.B1(_1849_),
    .Y(_1850_),
    .A1(_3266_),
    .A2(_1848_));
 sg13g2_o21ai_1 _6103_ (.B1(_1850_),
    .Y(_0124_),
    .A1(_3124_),
    .A2(net752));
 sg13g2_nand2_1 _6104_ (.Y(_1851_),
    .A(net248),
    .B(net749));
 sg13g2_and2_1 _6105_ (.A(\i_coord.y0[-3] ),
    .B(net803),
    .X(_1852_));
 sg13g2_xor2_1 _6106_ (.B(net803),
    .A(\i_coord.y0[-3] ),
    .X(_1853_));
 sg13g2_o21ai_1 _6107_ (.B1(_1842_),
    .Y(_1854_),
    .A1(\i_coord.y0[-4] ),
    .A2(net803));
 sg13g2_o21ai_1 _6108_ (.B1(_1854_),
    .Y(_1855_),
    .A1(_3124_),
    .A2(_3136_));
 sg13g2_xnor2_1 _6109_ (.Y(_1856_),
    .A(_1853_),
    .B(_1855_));
 sg13g2_a221oi_1 _6110_ (.B2(_1856_),
    .C1(net784),
    .B1(net792),
    .A1(_3113_),
    .Y(_1857_),
    .A2(net800));
 sg13g2_a21o_1 _6111_ (.A2(net783),
    .A1(\i_coord.l_yt.genblk2[10].state.Q ),
    .B1(_1857_),
    .X(_1858_));
 sg13g2_mux2_1 _6112_ (.A0(\i_coord.y0[-3] ),
    .A1(_1858_),
    .S(net877),
    .X(_1859_));
 sg13g2_nor2_1 _6113_ (.A(net762),
    .B(_1859_),
    .Y(_1860_));
 sg13g2_o21ai_1 _6114_ (.B1(net752),
    .Y(_1861_),
    .A1(net766),
    .A2(_1858_));
 sg13g2_o21ai_1 _6115_ (.B1(_1851_),
    .Y(_0125_),
    .A1(_1860_),
    .A2(_1861_));
 sg13g2_nand2_1 _6116_ (.Y(_1862_),
    .A(net228),
    .B(net747));
 sg13g2_nor2_1 _6117_ (.A(\i_coord.y0[-2] ),
    .B(net804),
    .Y(_1863_));
 sg13g2_nand2_1 _6118_ (.Y(_1864_),
    .A(\i_coord.y0[-2] ),
    .B(net803));
 sg13g2_nor2b_1 _6119_ (.A(_1863_),
    .B_N(_1864_),
    .Y(_1865_));
 sg13g2_a21oi_1 _6120_ (.A1(_1853_),
    .A2(_1855_),
    .Y(_1866_),
    .B1(_1852_));
 sg13g2_o21ai_1 _6121_ (.B1(net792),
    .Y(_1867_),
    .A1(_1865_),
    .A2(_1866_));
 sg13g2_a21oi_1 _6122_ (.A1(_1865_),
    .A2(_1866_),
    .Y(_1868_),
    .B1(_1867_));
 sg13g2_o21ai_1 _6123_ (.B1(net773),
    .Y(_1869_),
    .A1(\i_coord.y_row_start[-2] ),
    .A2(net796));
 sg13g2_nand2_1 _6124_ (.Y(_1870_),
    .A(\i_coord.l_yt.genblk2[11].state.Q ),
    .B(net784));
 sg13g2_o21ai_1 _6125_ (.B1(_1870_),
    .Y(_1871_),
    .A1(_1868_),
    .A2(_1869_));
 sg13g2_mux2_1 _6126_ (.A0(\i_coord.y0[-2] ),
    .A1(_1871_),
    .S(net877),
    .X(_1872_));
 sg13g2_nor2_1 _6127_ (.A(net762),
    .B(_1872_),
    .Y(_1873_));
 sg13g2_o21ai_1 _6128_ (.B1(net751),
    .Y(_1874_),
    .A1(net766),
    .A2(_1871_));
 sg13g2_o21ai_1 _6129_ (.B1(_1862_),
    .Y(_0126_),
    .A1(_1873_),
    .A2(_1874_));
 sg13g2_and2_1 _6130_ (.A(\i_coord.y0[-1] ),
    .B(net804),
    .X(_1875_));
 sg13g2_xor2_1 _6131_ (.B(net804),
    .A(\i_coord.y0[-1] ),
    .X(_1876_));
 sg13g2_o21ai_1 _6132_ (.B1(_1864_),
    .Y(_1877_),
    .A1(_1863_),
    .A2(_1866_));
 sg13g2_xnor2_1 _6133_ (.Y(_1878_),
    .A(_1876_),
    .B(_1877_));
 sg13g2_o21ai_1 _6134_ (.B1(net772),
    .Y(_1879_),
    .A1(\i_coord.y_row_start[-1] ),
    .A2(net796));
 sg13g2_a21oi_1 _6135_ (.A1(net796),
    .A2(_1878_),
    .Y(_1880_),
    .B1(_1879_));
 sg13g2_a21oi_1 _6136_ (.A1(\i_coord.l_yt.genblk2[12].state.Q ),
    .A2(net783),
    .Y(_1881_),
    .B1(_1880_));
 sg13g2_nor2_1 _6137_ (.A(net307),
    .B(net877),
    .Y(_1882_));
 sg13g2_a21oi_1 _6138_ (.A1(net877),
    .A2(_1881_),
    .Y(_1883_),
    .B1(_1882_));
 sg13g2_a21oi_1 _6139_ (.A1(net762),
    .A2(_1881_),
    .Y(_1884_),
    .B1(net747));
 sg13g2_o21ai_1 _6140_ (.B1(_1884_),
    .Y(_1885_),
    .A1(_3266_),
    .A2(_1883_));
 sg13g2_o21ai_1 _6141_ (.B1(_1885_),
    .Y(_0127_),
    .A1(_3125_),
    .A2(net751));
 sg13g2_a21o_1 _6142_ (.A2(_1877_),
    .A1(_1876_),
    .B1(_1875_),
    .X(_1886_));
 sg13g2_xor2_1 _6143_ (.B(net804),
    .A(\i_coord.y0[0] ),
    .X(_1887_));
 sg13g2_xnor2_1 _6144_ (.Y(_1888_),
    .A(_1886_),
    .B(_1887_));
 sg13g2_o21ai_1 _6145_ (.B1(net772),
    .Y(_1889_),
    .A1(\i_coord.y_row_start[0] ),
    .A2(net796));
 sg13g2_a21oi_1 _6146_ (.A1(net792),
    .A2(_1888_),
    .Y(_1890_),
    .B1(_1889_));
 sg13g2_a21oi_1 _6147_ (.A1(\i_coord.l_yt.genblk2[13].state.Q ),
    .A2(net783),
    .Y(_1891_),
    .B1(_1890_));
 sg13g2_nor2_1 _6148_ (.A(\i_coord.y0[0] ),
    .B(net877),
    .Y(_1892_));
 sg13g2_a21oi_1 _6149_ (.A1(net877),
    .A2(_1891_),
    .Y(_1893_),
    .B1(_1892_));
 sg13g2_a21oi_1 _6150_ (.A1(net762),
    .A2(_1891_),
    .Y(_1894_),
    .B1(net747));
 sg13g2_o21ai_1 _6151_ (.B1(_1894_),
    .Y(_1895_),
    .A1(_3266_),
    .A2(_1893_));
 sg13g2_o21ai_1 _6152_ (.B1(_1895_),
    .Y(_0128_),
    .A1(_3127_),
    .A2(net751));
 sg13g2_nor2_1 _6153_ (.A(net803),
    .B(_1886_),
    .Y(_1896_));
 sg13g2_mux2_1 _6154_ (.A0(net803),
    .A1(_1886_),
    .S(_3127_),
    .X(_1897_));
 sg13g2_nor3_1 _6155_ (.A(\i_coord.y0[1] ),
    .B(_1896_),
    .C(_1897_),
    .Y(_1898_));
 sg13g2_o21ai_1 _6156_ (.B1(\i_coord.y0[1] ),
    .Y(_1899_),
    .A1(_1896_),
    .A2(_1897_));
 sg13g2_nor2_1 _6157_ (.A(_3263_),
    .B(_1898_),
    .Y(_1900_));
 sg13g2_o21ai_1 _6158_ (.B1(net772),
    .Y(_1901_),
    .A1(\i_coord.y_row_start[1] ),
    .A2(net796));
 sg13g2_a21oi_1 _6159_ (.A1(_1899_),
    .A2(_1900_),
    .Y(_1902_),
    .B1(_1901_));
 sg13g2_a21oi_2 _6160_ (.B1(_1902_),
    .Y(_1903_),
    .A2(net784),
    .A1(\i_coord.l_yt.genblk2[14].state.Q ));
 sg13g2_nor2_1 _6161_ (.A(\i_coord.y0[1] ),
    .B(net877),
    .Y(_1904_));
 sg13g2_a21oi_2 _6162_ (.B1(_1904_),
    .Y(_1905_),
    .A2(_1903_),
    .A1(net877));
 sg13g2_a21oi_1 _6163_ (.A1(_3261_),
    .A2(_1903_),
    .Y(_1906_),
    .B1(net747));
 sg13g2_o21ai_1 _6164_ (.B1(_1906_),
    .Y(_1907_),
    .A1(_3266_),
    .A2(_1905_));
 sg13g2_o21ai_1 _6165_ (.B1(_1907_),
    .Y(_0129_),
    .A1(_3129_),
    .A2(net751));
 sg13g2_nor2_1 _6166_ (.A(\i_mandel.i_xy.hc.genblk1.genblk1.CG.GATE ),
    .B(net763),
    .Y(_1908_));
 sg13g2_o21ai_1 _6167_ (.B1(_1908_),
    .Y(_1909_),
    .A1(net838),
    .A2(_1071_));
 sg13g2_xnor2_1 _6168_ (.Y(_1910_),
    .A(\i_coord.x0[-13] ),
    .B(\i_mandel.l_sq.genblk2[1].state.D ));
 sg13g2_nand2_1 _6169_ (.Y(_1911_),
    .A(\i_mandel.l_sq.genblk2[1].state.Q ),
    .B(_1910_));
 sg13g2_xnor2_1 _6170_ (.Y(_1912_),
    .A(\i_mandel.l_sq.genblk2[1].state.Q ),
    .B(_1910_));
 sg13g2_a21oi_2 _6171_ (.B1(_1912_),
    .Y(_1913_),
    .A2(\i_mandel.l_sq.genblk2[0].state.D ),
    .A1(_3140_));
 sg13g2_inv_1 _6172_ (.Y(_1914_),
    .A(_1913_));
 sg13g2_nand3_1 _6173_ (.B(\i_mandel.l_sq.genblk2[0].state.D ),
    .C(_1912_),
    .A(_3140_),
    .Y(_1915_));
 sg13g2_a21oi_1 _6174_ (.A1(_1914_),
    .A2(_1915_),
    .Y(_1916_),
    .B1(net839));
 sg13g2_a21oi_1 _6175_ (.A1(net839),
    .A2(_1572_),
    .Y(_1917_),
    .B1(_1916_));
 sg13g2_mux2_1 _6176_ (.A0(_1917_),
    .A1(net203),
    .S(net733),
    .X(_0130_));
 sg13g2_nor2_1 _6177_ (.A(_3141_),
    .B(\i_mandel.l_sq.genblk2[2].state.D ),
    .Y(_1918_));
 sg13g2_xnor2_1 _6178_ (.Y(_1919_),
    .A(\i_coord.x0[-12] ),
    .B(\i_mandel.l_sq.genblk2[2].state.D ));
 sg13g2_xnor2_1 _6179_ (.Y(_1920_),
    .A(\i_mandel.l_sq.genblk2[2].state.Q ),
    .B(_1919_));
 sg13g2_o21ai_1 _6180_ (.B1(_1911_),
    .Y(_1921_),
    .A1(_3139_),
    .A2(\i_mandel.l_sq.genblk2[1].state.D ));
 sg13g2_nor2b_1 _6181_ (.A(_1920_),
    .B_N(_1921_),
    .Y(_1922_));
 sg13g2_xnor2_1 _6182_ (.Y(_1923_),
    .A(_1920_),
    .B(_1921_));
 sg13g2_a21oi_1 _6183_ (.A1(_1913_),
    .A2(_1923_),
    .Y(_1924_),
    .B1(net839));
 sg13g2_o21ai_1 _6184_ (.B1(_1924_),
    .Y(_1925_),
    .A1(_1913_),
    .A2(_1923_));
 sg13g2_o21ai_1 _6185_ (.B1(_1925_),
    .Y(_1926_),
    .A1(net836),
    .A2(_1580_));
 sg13g2_mux2_1 _6186_ (.A0(_1926_),
    .A1(net199),
    .S(net733),
    .X(_0131_));
 sg13g2_a21o_1 _6187_ (.A2(_1923_),
    .A1(_1913_),
    .B1(_1922_),
    .X(_1927_));
 sg13g2_a21oi_1 _6188_ (.A1(\i_mandel.l_sq.genblk2[2].state.Q ),
    .A2(_1919_),
    .Y(_1928_),
    .B1(_1918_));
 sg13g2_nor2b_1 _6189_ (.A(\i_mandel.l_sq.genblk2[3].state.D ),
    .B_N(\i_coord.x0[-11] ),
    .Y(_1929_));
 sg13g2_o21ai_1 _6190_ (.B1(\i_coord.x0[-11] ),
    .Y(_1930_),
    .A1(_0855_),
    .A2(_1112_));
 sg13g2_or3_1 _6191_ (.A(\i_coord.x0[-11] ),
    .B(_0855_),
    .C(_1112_),
    .X(_1931_));
 sg13g2_and3_1 _6192_ (.X(_1932_),
    .A(\i_mandel.l_sq.genblk2[3].state.Q ),
    .B(_1930_),
    .C(_1931_));
 sg13g2_a21oi_1 _6193_ (.A1(_1930_),
    .A2(_1931_),
    .Y(_1933_),
    .B1(\i_mandel.l_sq.genblk2[3].state.Q ));
 sg13g2_nor3_1 _6194_ (.A(_1928_),
    .B(_1932_),
    .C(_1933_),
    .Y(_1934_));
 sg13g2_o21ai_1 _6195_ (.B1(_1928_),
    .Y(_1935_),
    .A1(_1932_),
    .A2(_1933_));
 sg13g2_nor2b_1 _6196_ (.A(_1934_),
    .B_N(_1935_),
    .Y(_1936_));
 sg13g2_xnor2_1 _6197_ (.Y(_1937_),
    .A(_1927_),
    .B(_1936_));
 sg13g2_nand2_1 _6198_ (.Y(_1938_),
    .A(net836),
    .B(_1937_));
 sg13g2_o21ai_1 _6199_ (.B1(_1938_),
    .Y(_1939_),
    .A1(net836),
    .A2(_1590_));
 sg13g2_nand2_1 _6200_ (.Y(_1940_),
    .A(net186),
    .B(net733));
 sg13g2_o21ai_1 _6201_ (.B1(_1940_),
    .Y(_0132_),
    .A1(net733),
    .A2(_1939_));
 sg13g2_a21oi_1 _6202_ (.A1(_1927_),
    .A2(_1935_),
    .Y(_1941_),
    .B1(_1934_));
 sg13g2_or2_1 _6203_ (.X(_1942_),
    .B(_1932_),
    .A(_1929_));
 sg13g2_nor2_1 _6204_ (.A(_3143_),
    .B(\i_mandel.l_sq.genblk2[4].state.D ),
    .Y(_1943_));
 sg13g2_xnor2_1 _6205_ (.Y(_1944_),
    .A(\i_coord.x0[-10] ),
    .B(\i_mandel.l_sq.genblk2[4].state.D ));
 sg13g2_xnor2_1 _6206_ (.Y(_1945_),
    .A(\i_mandel.l_sq.genblk2[4].state.Q ),
    .B(_1944_));
 sg13g2_nand2b_1 _6207_ (.Y(_1946_),
    .B(_1942_),
    .A_N(_1945_));
 sg13g2_xor2_1 _6208_ (.B(_1945_),
    .A(_1942_),
    .X(_1947_));
 sg13g2_xnor2_1 _6209_ (.Y(_1948_),
    .A(_1941_),
    .B(_1947_));
 sg13g2_nand2_1 _6210_ (.Y(_1949_),
    .A(net833),
    .B(_1948_));
 sg13g2_o21ai_1 _6211_ (.B1(_1949_),
    .Y(_1950_),
    .A1(net833),
    .A2(_1600_));
 sg13g2_nand2_1 _6212_ (.Y(_1951_),
    .A(net185),
    .B(net733));
 sg13g2_o21ai_1 _6213_ (.B1(_1951_),
    .Y(_0133_),
    .A1(net734),
    .A2(_1950_));
 sg13g2_o21ai_1 _6214_ (.B1(_1946_),
    .Y(_1952_),
    .A1(_1941_),
    .A2(_1947_));
 sg13g2_a21oi_1 _6215_ (.A1(\i_mandel.l_sq.genblk2[4].state.Q ),
    .A2(_1944_),
    .Y(_1953_),
    .B1(_1943_));
 sg13g2_nor2b_1 _6216_ (.A(\i_mandel.l_sq.genblk2[5].state.D ),
    .B_N(\i_coord.x0[-9] ),
    .Y(_1954_));
 sg13g2_xnor2_1 _6217_ (.Y(_1955_),
    .A(\i_coord.x0[-9] ),
    .B(\i_mandel.l_sq.genblk2[5].state.D ));
 sg13g2_xnor2_1 _6218_ (.Y(_1956_),
    .A(\i_mandel.l_sq.genblk2[5].state.Q ),
    .B(_1955_));
 sg13g2_nor2_1 _6219_ (.A(_1953_),
    .B(_1956_),
    .Y(_1957_));
 sg13g2_nand2_1 _6220_ (.Y(_1958_),
    .A(_1953_),
    .B(_1956_));
 sg13g2_nand2b_1 _6221_ (.Y(_1959_),
    .B(_1958_),
    .A_N(_1957_));
 sg13g2_xor2_1 _6222_ (.B(_1959_),
    .A(_1952_),
    .X(_1960_));
 sg13g2_or2_1 _6223_ (.X(_1961_),
    .B(_1611_),
    .A(net833));
 sg13g2_o21ai_1 _6224_ (.B1(_1961_),
    .Y(_1962_),
    .A1(net841),
    .A2(_1960_));
 sg13g2_mux2_1 _6225_ (.A0(_1962_),
    .A1(net936),
    .S(net734),
    .X(_0134_));
 sg13g2_and2_1 _6226_ (.A(net841),
    .B(_1621_),
    .X(_1963_));
 sg13g2_a21oi_1 _6227_ (.A1(_1952_),
    .A2(_1958_),
    .Y(_1964_),
    .B1(_1957_));
 sg13g2_nor2b_1 _6228_ (.A(\i_mandel.l_sq.genblk2[6].state.D ),
    .B_N(\i_coord.x0[-8] ),
    .Y(_1965_));
 sg13g2_xnor2_1 _6229_ (.Y(_1966_),
    .A(\i_coord.x0[-8] ),
    .B(\i_mandel.l_sq.genblk2[6].state.D ));
 sg13g2_xnor2_1 _6230_ (.Y(_1967_),
    .A(\i_mandel.l_sq.genblk2[6].state.Q ),
    .B(_1966_));
 sg13g2_a21oi_1 _6231_ (.A1(\i_mandel.l_sq.genblk2[5].state.Q ),
    .A2(_1955_),
    .Y(_1968_),
    .B1(_1954_));
 sg13g2_or2_1 _6232_ (.X(_1969_),
    .B(_1968_),
    .A(_1967_));
 sg13g2_xnor2_1 _6233_ (.Y(_1970_),
    .A(_1967_),
    .B(_1968_));
 sg13g2_xnor2_1 _6234_ (.Y(_1971_),
    .A(_1964_),
    .B(_1970_));
 sg13g2_a21oi_1 _6235_ (.A1(net833),
    .A2(_1971_),
    .Y(_1972_),
    .B1(_1963_));
 sg13g2_mux2_1 _6236_ (.A0(_1972_),
    .A1(net934),
    .S(net738),
    .X(_0135_));
 sg13g2_o21ai_1 _6237_ (.B1(_1969_),
    .Y(_1973_),
    .A1(_1964_),
    .A2(_1970_));
 sg13g2_and2_1 _6238_ (.A(\i_coord.x0[-7] ),
    .B(_0975_),
    .X(_1974_));
 sg13g2_xor2_1 _6239_ (.B(_0975_),
    .A(\i_coord.x0[-7] ),
    .X(_1975_));
 sg13g2_xnor2_1 _6240_ (.Y(_1976_),
    .A(\i_mandel.l_sq.genblk2[7].state.Q ),
    .B(_1975_));
 sg13g2_a21oi_1 _6241_ (.A1(\i_mandel.l_sq.genblk2[6].state.Q ),
    .A2(_1966_),
    .Y(_1977_),
    .B1(_1965_));
 sg13g2_nor2_1 _6242_ (.A(_1976_),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_nand2_1 _6243_ (.Y(_1979_),
    .A(_1976_),
    .B(_1977_));
 sg13g2_nand2b_1 _6244_ (.Y(_1980_),
    .B(_1979_),
    .A_N(_1978_));
 sg13g2_xnor2_1 _6245_ (.Y(_1981_),
    .A(_1973_),
    .B(_1980_));
 sg13g2_nand2_1 _6246_ (.Y(_1982_),
    .A(net833),
    .B(_1981_));
 sg13g2_o21ai_1 _6247_ (.B1(_1982_),
    .Y(_1983_),
    .A1(net833),
    .A2(_1632_));
 sg13g2_mux2_1 _6248_ (.A0(_1983_),
    .A1(net274),
    .S(net732),
    .X(_0136_));
 sg13g2_a21oi_1 _6249_ (.A1(_1973_),
    .A2(_1979_),
    .Y(_1984_),
    .B1(_1978_));
 sg13g2_xnor2_1 _6250_ (.Y(_1985_),
    .A(\i_coord.x0[-6] ),
    .B(\i_mandel.l_sq.genblk2[8].state.D ));
 sg13g2_nand2_1 _6251_ (.Y(_1986_),
    .A(\i_mandel.l_sq.genblk2[8].state.Q ),
    .B(_1985_));
 sg13g2_xnor2_1 _6252_ (.Y(_1987_),
    .A(\i_mandel.l_sq.genblk2[8].state.Q ),
    .B(_1985_));
 sg13g2_a21o_1 _6253_ (.A2(_1975_),
    .A1(\i_mandel.l_sq.genblk2[7].state.Q ),
    .B1(_1974_),
    .X(_1988_));
 sg13g2_nand2b_1 _6254_ (.Y(_1989_),
    .B(_1988_),
    .A_N(_1987_));
 sg13g2_nor2b_1 _6255_ (.A(_1988_),
    .B_N(_1987_),
    .Y(_1990_));
 sg13g2_xnor2_1 _6256_ (.Y(_1991_),
    .A(_1987_),
    .B(_1988_));
 sg13g2_xor2_1 _6257_ (.B(_1991_),
    .A(_1984_),
    .X(_1992_));
 sg13g2_o21ai_1 _6258_ (.B1(_1643_),
    .Y(_1993_),
    .A1(net838),
    .A2(_1992_));
 sg13g2_mux2_1 _6259_ (.A0(_1993_),
    .A1(net321),
    .S(net736),
    .X(_0137_));
 sg13g2_o21ai_1 _6260_ (.B1(_1989_),
    .Y(_1994_),
    .A1(_1984_),
    .A2(_1990_));
 sg13g2_o21ai_1 _6261_ (.B1(_1986_),
    .Y(_1995_),
    .A1(_3144_),
    .A2(\i_mandel.l_sq.genblk2[8].state.D ));
 sg13g2_and2_1 _6262_ (.A(\i_coord.x0[-5] ),
    .B(_0971_),
    .X(_1996_));
 sg13g2_xor2_1 _6263_ (.B(_0971_),
    .A(\i_coord.x0[-5] ),
    .X(_1997_));
 sg13g2_xnor2_1 _6264_ (.Y(_1998_),
    .A(\i_mandel.l_sq.genblk2[9].state.Q ),
    .B(_1997_));
 sg13g2_nor2b_1 _6265_ (.A(_1998_),
    .B_N(_1995_),
    .Y(_1999_));
 sg13g2_nand2b_1 _6266_ (.Y(_2000_),
    .B(_1998_),
    .A_N(_1995_));
 sg13g2_nand2b_1 _6267_ (.Y(_2001_),
    .B(_2000_),
    .A_N(_1999_));
 sg13g2_xnor2_1 _6268_ (.Y(_2002_),
    .A(_1994_),
    .B(_2001_));
 sg13g2_nor2_1 _6269_ (.A(net838),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_a21oi_2 _6270_ (.B1(_2003_),
    .Y(_2004_),
    .A2(_1654_),
    .A1(net838));
 sg13g2_mux2_1 _6271_ (.A0(_2004_),
    .A1(net267),
    .S(net734),
    .X(_0138_));
 sg13g2_a21oi_1 _6272_ (.A1(_1994_),
    .A2(_2000_),
    .Y(_2005_),
    .B1(_1999_));
 sg13g2_nor2b_1 _6273_ (.A(\i_mandel.l_sq.genblk2[10].state.D ),
    .B_N(\i_coord.x0[-4] ),
    .Y(_2006_));
 sg13g2_xnor2_1 _6274_ (.Y(_2007_),
    .A(\i_coord.x0[-4] ),
    .B(\i_mandel.l_sq.genblk2[10].state.D ));
 sg13g2_xnor2_1 _6275_ (.Y(_2008_),
    .A(\i_mandel.l_sq.genblk2[10].state.Q ),
    .B(_2007_));
 sg13g2_a21oi_1 _6276_ (.A1(\i_mandel.l_sq.genblk2[9].state.Q ),
    .A2(_1997_),
    .Y(_2009_),
    .B1(_1996_));
 sg13g2_or2_1 _6277_ (.X(_2010_),
    .B(_2009_),
    .A(_2008_));
 sg13g2_xnor2_1 _6278_ (.Y(_2011_),
    .A(_2008_),
    .B(_2009_));
 sg13g2_o21ai_1 _6279_ (.B1(net832),
    .Y(_2012_),
    .A1(_2005_),
    .A2(_2011_));
 sg13g2_a21o_1 _6280_ (.A2(_2011_),
    .A1(_2005_),
    .B1(_2012_),
    .X(_2013_));
 sg13g2_o21ai_1 _6281_ (.B1(_2013_),
    .Y(_2014_),
    .A1(net832),
    .A2(_1665_));
 sg13g2_mux2_1 _6282_ (.A0(_2014_),
    .A1(net925),
    .S(net732),
    .X(_0139_));
 sg13g2_o21ai_1 _6283_ (.B1(_2010_),
    .Y(_2015_),
    .A1(_2005_),
    .A2(_2011_));
 sg13g2_and2_1 _6284_ (.A(\i_coord.x0[-3] ),
    .B(_0965_),
    .X(_2016_));
 sg13g2_xnor2_1 _6285_ (.Y(_2017_),
    .A(\i_coord.x0[-3] ),
    .B(\i_mandel.l_sq.genblk2[11].state.D ));
 sg13g2_xnor2_1 _6286_ (.Y(_2018_),
    .A(\i_mandel.l_sq.genblk2[11].state.Q ),
    .B(_2017_));
 sg13g2_a21oi_1 _6287_ (.A1(\i_mandel.l_sq.genblk2[10].state.Q ),
    .A2(_2007_),
    .Y(_2019_),
    .B1(_2006_));
 sg13g2_nor2_1 _6288_ (.A(_2018_),
    .B(_2019_),
    .Y(_2020_));
 sg13g2_nand2_1 _6289_ (.Y(_2021_),
    .A(_2018_),
    .B(_2019_));
 sg13g2_nand2b_1 _6290_ (.Y(_2022_),
    .B(_2021_),
    .A_N(_2020_));
 sg13g2_xnor2_1 _6291_ (.Y(_2023_),
    .A(_2015_),
    .B(_2022_));
 sg13g2_nand2_1 _6292_ (.Y(_2024_),
    .A(net832),
    .B(_2023_));
 sg13g2_o21ai_1 _6293_ (.B1(_2024_),
    .Y(_2025_),
    .A1(net831),
    .A2(_1677_));
 sg13g2_mux2_1 _6294_ (.A0(_2025_),
    .A1(net922),
    .S(net732),
    .X(_0140_));
 sg13g2_a21oi_1 _6295_ (.A1(_2015_),
    .A2(_2021_),
    .Y(_2026_),
    .B1(_2020_));
 sg13g2_nor2b_1 _6296_ (.A(\i_mandel.l_sq.genblk2[12].state.D ),
    .B_N(\i_coord.x0[-2] ),
    .Y(_2027_));
 sg13g2_xnor2_1 _6297_ (.Y(_2028_),
    .A(\i_coord.x0[-2] ),
    .B(\i_mandel.l_sq.genblk2[12].state.D ));
 sg13g2_xnor2_1 _6298_ (.Y(_2029_),
    .A(\i_mandel.l_sq.genblk2[12].state.Q ),
    .B(_2028_));
 sg13g2_a21oi_1 _6299_ (.A1(\i_mandel.l_sq.genblk2[11].state.Q ),
    .A2(_2017_),
    .Y(_2030_),
    .B1(_2016_));
 sg13g2_or2_1 _6300_ (.X(_2031_),
    .B(_2030_),
    .A(_2029_));
 sg13g2_xor2_1 _6301_ (.B(_2030_),
    .A(_2029_),
    .X(_2032_));
 sg13g2_nand2b_1 _6302_ (.Y(_2033_),
    .B(_2032_),
    .A_N(_2026_));
 sg13g2_xnor2_1 _6303_ (.Y(_2034_),
    .A(_2026_),
    .B(_2032_));
 sg13g2_nand2_1 _6304_ (.Y(_2035_),
    .A(net831),
    .B(_2034_));
 sg13g2_o21ai_1 _6305_ (.B1(_2035_),
    .Y(_2036_),
    .A1(net831),
    .A2(_1690_));
 sg13g2_mux2_1 _6306_ (.A0(_2036_),
    .A1(net211),
    .S(net738),
    .X(_0141_));
 sg13g2_and2_1 _6307_ (.A(\i_coord.x0[-1] ),
    .B(_1002_),
    .X(_2037_));
 sg13g2_xor2_1 _6308_ (.B(_1002_),
    .A(\i_coord.x0[-1] ),
    .X(_2038_));
 sg13g2_xnor2_1 _6309_ (.Y(_2039_),
    .A(\i_mandel.l_sq.genblk2[13].state.Q ),
    .B(_2038_));
 sg13g2_a21oi_1 _6310_ (.A1(\i_mandel.l_sq.genblk2[12].state.Q ),
    .A2(_2028_),
    .Y(_2040_),
    .B1(_2027_));
 sg13g2_nor2_1 _6311_ (.A(_2039_),
    .B(_2040_),
    .Y(_2041_));
 sg13g2_xnor2_1 _6312_ (.Y(_2042_),
    .A(_2039_),
    .B(_2040_));
 sg13g2_a21oi_1 _6313_ (.A1(_2031_),
    .A2(_2033_),
    .Y(_2043_),
    .B1(_2042_));
 sg13g2_and3_1 _6314_ (.X(_2044_),
    .A(_2031_),
    .B(_2033_),
    .C(_2042_));
 sg13g2_or3_1 _6315_ (.A(net838),
    .B(_2043_),
    .C(_2044_),
    .X(_2045_));
 sg13g2_o21ai_1 _6316_ (.B1(_2045_),
    .Y(_2046_),
    .A1(net831),
    .A2(_1700_));
 sg13g2_mux2_1 _6317_ (.A0(_2046_),
    .A1(net347),
    .S(net733),
    .X(_0142_));
 sg13g2_or2_1 _6318_ (.X(_2047_),
    .B(_2043_),
    .A(_2041_));
 sg13g2_and2_1 _6319_ (.A(\i_coord.x0[0] ),
    .B(_1018_),
    .X(_2048_));
 sg13g2_xor2_1 _6320_ (.B(_1018_),
    .A(\i_coord.x0[0] ),
    .X(_2049_));
 sg13g2_xnor2_1 _6321_ (.Y(_2050_),
    .A(\i_mandel.l_sq.genblk2[14].state.Q ),
    .B(_2049_));
 sg13g2_a21o_1 _6322_ (.A2(_2038_),
    .A1(\i_mandel.l_sq.genblk2[13].state.Q ),
    .B1(_2037_),
    .X(_2051_));
 sg13g2_nand2b_1 _6323_ (.Y(_2052_),
    .B(_2051_),
    .A_N(_2050_));
 sg13g2_xnor2_1 _6324_ (.Y(_2053_),
    .A(_2050_),
    .B(_2051_));
 sg13g2_o21ai_1 _6325_ (.B1(_2053_),
    .Y(_2054_),
    .A1(_2041_),
    .A2(_2043_));
 sg13g2_o21ai_1 _6326_ (.B1(net831),
    .Y(_2055_),
    .A1(_2047_),
    .A2(_2053_));
 sg13g2_nand2b_1 _6327_ (.Y(_2056_),
    .B(_2054_),
    .A_N(_2055_));
 sg13g2_o21ai_1 _6328_ (.B1(_2056_),
    .Y(_2057_),
    .A1(net831),
    .A2(_1712_));
 sg13g2_mux2_1 _6329_ (.A0(_2057_),
    .A1(net286),
    .S(net732),
    .X(_0143_));
 sg13g2_xnor2_1 _6330_ (.Y(_2058_),
    .A(\i_coord.x0[1] ),
    .B(\i_mandel.l_sq.genblk2[15].state.D ));
 sg13g2_nand2_1 _6331_ (.Y(_2059_),
    .A(\i_mandel.l_sq.genblk2[15].state.Q ),
    .B(_2058_));
 sg13g2_xnor2_1 _6332_ (.Y(_2060_),
    .A(\i_mandel.l_sq.genblk2[15].state.Q ),
    .B(_2058_));
 sg13g2_a21oi_1 _6333_ (.A1(\i_mandel.l_sq.genblk2[14].state.Q ),
    .A2(_2049_),
    .Y(_2061_),
    .B1(_2048_));
 sg13g2_or2_1 _6334_ (.X(_2062_),
    .B(_2061_),
    .A(_2060_));
 sg13g2_xnor2_1 _6335_ (.Y(_2063_),
    .A(_2060_),
    .B(_2061_));
 sg13g2_nand3_1 _6336_ (.B(_2054_),
    .C(_2063_),
    .A(_2052_),
    .Y(_2064_));
 sg13g2_a21o_1 _6337_ (.A2(_2054_),
    .A1(_2052_),
    .B1(_2063_),
    .X(_2065_));
 sg13g2_nand3_1 _6338_ (.B(_2064_),
    .C(_2065_),
    .A(net831),
    .Y(_2066_));
 sg13g2_nor2_1 _6339_ (.A(_1725_),
    .B(net732),
    .Y(_2067_));
 sg13g2_a22oi_1 _6340_ (.Y(_0144_),
    .B1(_2066_),
    .B2(_2067_),
    .A2(net732),
    .A1(_3133_));
 sg13g2_nand2_1 _6341_ (.Y(_2068_),
    .A(net191),
    .B(net732));
 sg13g2_o21ai_1 _6342_ (.B1(_2059_),
    .Y(_2069_),
    .A1(_3145_),
    .A2(\i_mandel.l_sq.genblk2[15].state.D ));
 sg13g2_xnor2_1 _6343_ (.Y(_2070_),
    .A(\i_coord.x0[2] ),
    .B(_1025_));
 sg13g2_xnor2_1 _6344_ (.Y(_2071_),
    .A(_2069_),
    .B(_2070_));
 sg13g2_and3_1 _6345_ (.X(_2072_),
    .A(_2062_),
    .B(_2065_),
    .C(_2071_));
 sg13g2_a21oi_1 _6346_ (.A1(_2062_),
    .A2(_2065_),
    .Y(_2073_),
    .B1(_2071_));
 sg13g2_nor3_1 _6347_ (.A(net838),
    .B(_2072_),
    .C(_2073_),
    .Y(_2074_));
 sg13g2_a21o_1 _6348_ (.A2(_1735_),
    .A1(net838),
    .B1(net732),
    .X(_2075_));
 sg13g2_o21ai_1 _6349_ (.B1(_2068_),
    .Y(_0145_),
    .A1(_2074_),
    .A2(_2075_));
 sg13g2_nand2_1 _6350_ (.Y(_2076_),
    .A(net205),
    .B(_3267_));
 sg13g2_o21ai_1 _6351_ (.B1(_2076_),
    .Y(_0146_),
    .A1(_1079_),
    .A2(_1564_));
 sg13g2_nand2_1 _6352_ (.Y(_2077_),
    .A(net192),
    .B(_3267_));
 sg13g2_o21ai_1 _6353_ (.B1(_2077_),
    .Y(_0147_),
    .A1(_1097_),
    .A2(_1564_));
 sg13g2_nand2_1 _6354_ (.Y(_2078_),
    .A(net212),
    .B(_3267_));
 sg13g2_o21ai_1 _6355_ (.B1(_2078_),
    .Y(_0148_),
    .A1(_1074_),
    .A2(_1564_));
 sg13g2_nand2_1 _6356_ (.Y(_2079_),
    .A(net189),
    .B(_3267_));
 sg13g2_o21ai_1 _6357_ (.B1(_2079_),
    .Y(_0149_),
    .A1(_1084_),
    .A2(_1564_));
 sg13g2_and2_1 _6358_ (.A(\i_mandel.i_xy.hc.genblk2[2].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[2].state.D ),
    .X(_2080_));
 sg13g2_nand2_2 _6359_ (.Y(_2081_),
    .A(net935),
    .B(net902));
 sg13g2_nand2_1 _6360_ (.Y(_2082_),
    .A(\i_mandel.i_xy.hc.genblk2[3].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[3].state.D ));
 sg13g2_xnor2_1 _6361_ (.Y(_2083_),
    .A(\i_mandel.i_xy.hc.genblk2[3].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[3].state.D ));
 sg13g2_nand2_2 _6362_ (.Y(_2084_),
    .A(net932),
    .B(net906));
 sg13g2_nand2_1 _6363_ (.Y(_2085_),
    .A(net936),
    .B(net904));
 sg13g2_nand2_1 _6364_ (.Y(_2086_),
    .A(net931),
    .B(net907));
 sg13g2_xor2_1 _6365_ (.B(_2085_),
    .A(_2084_),
    .X(_2087_));
 sg13g2_nand2b_1 _6366_ (.Y(_2088_),
    .B(_2087_),
    .A_N(_2086_));
 sg13g2_o21ai_1 _6367_ (.B1(_2088_),
    .Y(_2089_),
    .A1(_2084_),
    .A2(_2085_));
 sg13g2_nand2_1 _6368_ (.Y(_2090_),
    .A(net929),
    .B(net907));
 sg13g2_nand2_2 _6369_ (.Y(_2091_),
    .A(net904),
    .B(net931));
 sg13g2_nor2_1 _6370_ (.A(_2084_),
    .B(_2091_),
    .Y(_2092_));
 sg13g2_a22oi_1 _6371_ (.Y(_2093_),
    .B1(net931),
    .B2(net906),
    .A2(net904),
    .A1(net932));
 sg13g2_nor2_1 _6372_ (.A(_2092_),
    .B(_2093_),
    .Y(_2094_));
 sg13g2_nand2b_1 _6373_ (.Y(_2095_),
    .B(_2094_),
    .A_N(_2090_));
 sg13g2_xnor2_1 _6374_ (.Y(_2096_),
    .A(_2090_),
    .B(_2094_));
 sg13g2_nand2_1 _6375_ (.Y(_2097_),
    .A(_2089_),
    .B(_2096_));
 sg13g2_xnor2_1 _6376_ (.Y(_2098_),
    .A(_2089_),
    .B(_2096_));
 sg13g2_xor2_1 _6377_ (.B(_2098_),
    .A(_2083_),
    .X(_2099_));
 sg13g2_nand2_1 _6378_ (.Y(_2100_),
    .A(net936),
    .B(net907));
 sg13g2_nor2_1 _6379_ (.A(_2084_),
    .B(_2100_),
    .Y(_2101_));
 sg13g2_xnor2_1 _6380_ (.Y(_2102_),
    .A(_2086_),
    .B(_2087_));
 sg13g2_xnor2_1 _6381_ (.Y(_2103_),
    .A(_2101_),
    .B(_2102_));
 sg13g2_xnor2_1 _6382_ (.Y(_2104_),
    .A(\i_mandel.i_xy.hc.genblk2[2].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[2].state.D ));
 sg13g2_nor2_1 _6383_ (.A(_2103_),
    .B(_2104_),
    .Y(_2105_));
 sg13g2_a21oi_1 _6384_ (.A1(_2101_),
    .A2(_2102_),
    .Y(_2106_),
    .B1(_2105_));
 sg13g2_nand2b_1 _6385_ (.Y(_2107_),
    .B(_2099_),
    .A_N(_2106_));
 sg13g2_xnor2_1 _6386_ (.Y(_2108_),
    .A(_2099_),
    .B(_2106_));
 sg13g2_nand2b_1 _6387_ (.Y(_2109_),
    .B(_2108_),
    .A_N(_2081_));
 sg13g2_xnor2_1 _6388_ (.Y(_2110_),
    .A(_2081_),
    .B(_2108_));
 sg13g2_nand2_1 _6389_ (.Y(_2111_),
    .A(\i_mandel.i_xy.hc.genblk2[1].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[1].state.D ));
 sg13g2_xnor2_1 _6390_ (.Y(_2112_),
    .A(\i_mandel.i_xy.hc.genblk2[1].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[1].state.D ));
 sg13g2_a22oi_1 _6391_ (.Y(_2113_),
    .B1(net907),
    .B2(net932),
    .A2(net906),
    .A1(net936));
 sg13g2_nor2_1 _6392_ (.A(_2101_),
    .B(_2113_),
    .Y(_2114_));
 sg13g2_nand2b_1 _6393_ (.Y(_2115_),
    .B(_2114_),
    .A_N(_2112_));
 sg13g2_xnor2_1 _6394_ (.Y(_2116_),
    .A(_2103_),
    .B(_2104_));
 sg13g2_nor2_1 _6395_ (.A(_2115_),
    .B(_2116_),
    .Y(_2117_));
 sg13g2_nand2_1 _6396_ (.Y(_2118_),
    .A(_2110_),
    .B(_2117_));
 sg13g2_xnor2_1 _6397_ (.Y(_2119_),
    .A(_2112_),
    .B(_2114_));
 sg13g2_nor2_1 _6398_ (.A(\i_mandel.i_xy.hc.genblk2[0].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[0].state.D ),
    .Y(_2120_));
 sg13g2_and2_1 _6399_ (.A(\i_mandel.i_xy.hc.genblk2[0].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[0].state.D ),
    .X(_2121_));
 sg13g2_nor3_1 _6400_ (.A(_2100_),
    .B(_2120_),
    .C(_2121_),
    .Y(_2122_));
 sg13g2_xor2_1 _6401_ (.B(_2116_),
    .A(_2115_),
    .X(_2123_));
 sg13g2_and3_1 _6402_ (.X(_2124_),
    .A(_2119_),
    .B(_2122_),
    .C(_2123_));
 sg13g2_nor2_1 _6403_ (.A(_2117_),
    .B(_2124_),
    .Y(_2125_));
 sg13g2_xnor2_1 _6404_ (.Y(_2126_),
    .A(_2110_),
    .B(_2125_));
 sg13g2_nand2_1 _6405_ (.Y(_2127_),
    .A(_2119_),
    .B(_2121_));
 sg13g2_a21oi_1 _6406_ (.A1(_2119_),
    .A2(_2122_),
    .Y(_2128_),
    .B1(_2123_));
 sg13g2_a21oi_1 _6407_ (.A1(_2111_),
    .A2(_2127_),
    .Y(_2129_),
    .B1(_2128_));
 sg13g2_nand2b_1 _6408_ (.Y(_2130_),
    .B(_2129_),
    .A_N(_2124_));
 sg13g2_o21ai_1 _6409_ (.B1(_2130_),
    .Y(_2131_),
    .A1(_2111_),
    .A2(_2127_));
 sg13g2_o21ai_1 _6410_ (.B1(_2131_),
    .Y(_2132_),
    .A1(_2080_),
    .A2(_2126_));
 sg13g2_a21o_1 _6411_ (.A2(_2126_),
    .A1(_2080_),
    .B1(_2132_),
    .X(_2133_));
 sg13g2_a22oi_1 _6412_ (.Y(_2134_),
    .B1(_2126_),
    .B2(_2080_),
    .A2(_2124_),
    .A1(_2110_));
 sg13g2_nand2_1 _6413_ (.Y(_2135_),
    .A(net898),
    .B(net933));
 sg13g2_nor2_1 _6414_ (.A(_2081_),
    .B(_2135_),
    .Y(_2136_));
 sg13g2_a22oi_1 _6415_ (.Y(_2137_),
    .B1(net902),
    .B2(net932),
    .A2(net935),
    .A1(net899));
 sg13g2_nor2_1 _6416_ (.A(_2136_),
    .B(_2137_),
    .Y(_2138_));
 sg13g2_o21ai_1 _6417_ (.B1(_2095_),
    .Y(_2139_),
    .A1(_2084_),
    .A2(_2091_));
 sg13g2_nand2_1 _6418_ (.Y(_2140_),
    .A(net927),
    .B(net907));
 sg13g2_nand2_1 _6419_ (.Y(_2141_),
    .A(net904),
    .B(net929));
 sg13g2_nand2_1 _6420_ (.Y(_2142_),
    .A(net929),
    .B(net906));
 sg13g2_xor2_1 _6421_ (.B(_2142_),
    .A(_2091_),
    .X(_2143_));
 sg13g2_nand2b_1 _6422_ (.Y(_2144_),
    .B(_2143_),
    .A_N(_2140_));
 sg13g2_xnor2_1 _6423_ (.Y(_2145_),
    .A(_2140_),
    .B(_2143_));
 sg13g2_xnor2_1 _6424_ (.Y(_2146_),
    .A(_2139_),
    .B(_2145_));
 sg13g2_nand2_1 _6425_ (.Y(_2147_),
    .A(\i_mandel.i_xy.hc.genblk2[4].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[4].state.D ));
 sg13g2_xnor2_1 _6426_ (.Y(_2148_),
    .A(\i_mandel.i_xy.hc.genblk2[4].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[4].state.D ));
 sg13g2_nor2_1 _6427_ (.A(_2146_),
    .B(_2148_),
    .Y(_2149_));
 sg13g2_xor2_1 _6428_ (.B(_2148_),
    .A(_2146_),
    .X(_2150_));
 sg13g2_o21ai_1 _6429_ (.B1(_2097_),
    .Y(_2151_),
    .A1(_2083_),
    .A2(_2098_));
 sg13g2_and2_1 _6430_ (.A(_2150_),
    .B(_2151_),
    .X(_2152_));
 sg13g2_xor2_1 _6431_ (.B(_2151_),
    .A(_2150_),
    .X(_2153_));
 sg13g2_xnor2_1 _6432_ (.Y(_2154_),
    .A(_2138_),
    .B(_2153_));
 sg13g2_nand2_1 _6433_ (.Y(_2155_),
    .A(_2107_),
    .B(_2109_));
 sg13g2_nand2b_1 _6434_ (.Y(_2156_),
    .B(_2155_),
    .A_N(_2154_));
 sg13g2_xor2_1 _6435_ (.B(_2155_),
    .A(_2154_),
    .X(_2157_));
 sg13g2_xor2_1 _6436_ (.B(_2157_),
    .A(_2118_),
    .X(_2158_));
 sg13g2_nand2b_1 _6437_ (.Y(_2159_),
    .B(_2158_),
    .A_N(_2082_));
 sg13g2_xnor2_1 _6438_ (.Y(_2160_),
    .A(_2082_),
    .B(_2158_));
 sg13g2_nand2b_1 _6439_ (.Y(_2161_),
    .B(_2160_),
    .A_N(_2134_));
 sg13g2_xnor2_1 _6440_ (.Y(_2162_),
    .A(_2134_),
    .B(_2160_));
 sg13g2_nand2b_1 _6441_ (.Y(_2163_),
    .B(_2162_),
    .A_N(_2133_));
 sg13g2_xnor2_1 _6442_ (.Y(_2164_),
    .A(_2133_),
    .B(_2162_));
 sg13g2_xor2_1 _6443_ (.B(_2164_),
    .A(_0026_),
    .X(_2165_));
 sg13g2_nand2_1 _6444_ (.Y(_2166_),
    .A(net839),
    .B(_1743_));
 sg13g2_o21ai_1 _6445_ (.B1(_2166_),
    .Y(_2167_),
    .A1(net839),
    .A2(_2165_));
 sg13g2_mux2_1 _6446_ (.A0(_2167_),
    .A1(net200),
    .S(net734),
    .X(_0150_));
 sg13g2_and2_1 _6447_ (.A(\i_coord.y0[-13] ),
    .B(_2164_),
    .X(_2168_));
 sg13g2_nand2_1 _6448_ (.Y(_2169_),
    .A(_2161_),
    .B(_2163_));
 sg13g2_o21ai_1 _6449_ (.B1(_2159_),
    .Y(_2170_),
    .A1(_2118_),
    .A2(_2157_));
 sg13g2_nand2_1 _6450_ (.Y(_2171_),
    .A(net902),
    .B(net930));
 sg13g2_nand2_1 _6451_ (.Y(_2172_),
    .A(net933),
    .B(net894));
 sg13g2_nand2_1 _6452_ (.Y(_2173_),
    .A(net935),
    .B(net896));
 sg13g2_or2_1 _6453_ (.X(_2174_),
    .B(_2173_),
    .A(_2135_));
 sg13g2_xor2_1 _6454_ (.B(_2173_),
    .A(_2135_),
    .X(_2175_));
 sg13g2_nand2b_1 _6455_ (.Y(_2176_),
    .B(_2175_),
    .A_N(_2171_));
 sg13g2_xnor2_1 _6456_ (.Y(_2177_),
    .A(_2171_),
    .B(_2175_));
 sg13g2_nand2_1 _6457_ (.Y(_2178_),
    .A(_2136_),
    .B(_2177_));
 sg13g2_xor2_1 _6458_ (.B(_2177_),
    .A(_2136_),
    .X(_2179_));
 sg13g2_o21ai_1 _6459_ (.B1(_2144_),
    .Y(_2180_),
    .A1(_2091_),
    .A2(_2142_));
 sg13g2_nand2_1 _6460_ (.Y(_2181_),
    .A(net907),
    .B(net923));
 sg13g2_nand2_1 _6461_ (.Y(_2182_),
    .A(net903),
    .B(net926));
 sg13g2_nand2_1 _6462_ (.Y(_2183_),
    .A(net906),
    .B(net927));
 sg13g2_xor2_1 _6463_ (.B(_2183_),
    .A(_2141_),
    .X(_2184_));
 sg13g2_nand2b_1 _6464_ (.Y(_2185_),
    .B(_2184_),
    .A_N(_2181_));
 sg13g2_xnor2_1 _6465_ (.Y(_2186_),
    .A(_2181_),
    .B(_2184_));
 sg13g2_xnor2_1 _6466_ (.Y(_2187_),
    .A(_2180_),
    .B(_2186_));
 sg13g2_nand2_1 _6467_ (.Y(_2188_),
    .A(\i_mandel.i_xy.hc.genblk2[5].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[5].state.D ));
 sg13g2_xnor2_1 _6468_ (.Y(_2189_),
    .A(\i_mandel.i_xy.hc.genblk2[5].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[5].state.D ));
 sg13g2_nor2_1 _6469_ (.A(_2187_),
    .B(_2189_),
    .Y(_2190_));
 sg13g2_xor2_1 _6470_ (.B(_2189_),
    .A(_2187_),
    .X(_2191_));
 sg13g2_a21oi_1 _6471_ (.A1(_2139_),
    .A2(_2145_),
    .Y(_2192_),
    .B1(_2149_));
 sg13g2_nand2b_1 _6472_ (.Y(_2193_),
    .B(_2191_),
    .A_N(_2192_));
 sg13g2_xnor2_1 _6473_ (.Y(_2194_),
    .A(_2191_),
    .B(_2192_));
 sg13g2_nand2_1 _6474_ (.Y(_2195_),
    .A(_2179_),
    .B(_2194_));
 sg13g2_xnor2_1 _6475_ (.Y(_2196_),
    .A(_2179_),
    .B(_2194_));
 sg13g2_a21oi_1 _6476_ (.A1(_2138_),
    .A2(_2153_),
    .Y(_2197_),
    .B1(_2152_));
 sg13g2_nor2_1 _6477_ (.A(_2196_),
    .B(_2197_),
    .Y(_2198_));
 sg13g2_xnor2_1 _6478_ (.Y(_2199_),
    .A(_2196_),
    .B(_2197_));
 sg13g2_xor2_1 _6479_ (.B(_2199_),
    .A(_2156_),
    .X(_2200_));
 sg13g2_nand2b_1 _6480_ (.Y(_2201_),
    .B(_2200_),
    .A_N(_2147_));
 sg13g2_xnor2_1 _6481_ (.Y(_2202_),
    .A(_2147_),
    .B(_2200_));
 sg13g2_xnor2_1 _6482_ (.Y(_2203_),
    .A(_2170_),
    .B(_2202_));
 sg13g2_a21oi_1 _6483_ (.A1(_2161_),
    .A2(_2163_),
    .Y(_2204_),
    .B1(_2203_));
 sg13g2_xnor2_1 _6484_ (.Y(_2205_),
    .A(_2169_),
    .B(_2203_));
 sg13g2_xnor2_1 _6485_ (.Y(_2206_),
    .A(_0025_),
    .B(_2205_));
 sg13g2_xnor2_1 _6486_ (.Y(_2207_),
    .A(_2168_),
    .B(_2206_));
 sg13g2_nand2_1 _6487_ (.Y(_2208_),
    .A(net836),
    .B(_2207_));
 sg13g2_o21ai_1 _6488_ (.B1(_2208_),
    .Y(_2209_),
    .A1(net836),
    .A2(_1754_));
 sg13g2_nand2_1 _6489_ (.Y(_2210_),
    .A(net187),
    .B(net737));
 sg13g2_o21ai_1 _6490_ (.B1(_2210_),
    .Y(_0151_),
    .A1(net737),
    .A2(_2209_));
 sg13g2_a22oi_1 _6491_ (.Y(_2211_),
    .B1(_2206_),
    .B2(_2168_),
    .A2(_2205_),
    .A1(\i_coord.y0[-12] ));
 sg13g2_a21oi_1 _6492_ (.A1(_2170_),
    .A2(_2202_),
    .Y(_2212_),
    .B1(_2204_));
 sg13g2_o21ai_1 _6493_ (.B1(_2201_),
    .Y(_2213_),
    .A1(_2156_),
    .A2(_2199_));
 sg13g2_nand2_2 _6494_ (.Y(_2214_),
    .A(net936),
    .B(net892));
 sg13g2_and2_1 _6495_ (.A(net901),
    .B(net928),
    .X(_2215_));
 sg13g2_nand2_1 _6496_ (.Y(_2216_),
    .A(net897),
    .B(net930));
 sg13g2_nor2_1 _6497_ (.A(_2172_),
    .B(_2216_),
    .Y(_2217_));
 sg13g2_xor2_1 _6498_ (.B(_2216_),
    .A(_2172_),
    .X(_2218_));
 sg13g2_xor2_1 _6499_ (.B(_2218_),
    .A(_2215_),
    .X(_2219_));
 sg13g2_and2_1 _6500_ (.A(_2174_),
    .B(_2176_),
    .X(_2220_));
 sg13g2_nand2b_1 _6501_ (.Y(_2221_),
    .B(_2219_),
    .A_N(_2220_));
 sg13g2_xnor2_1 _6502_ (.Y(_2222_),
    .A(_2219_),
    .B(_2220_));
 sg13g2_nor2b_1 _6503_ (.A(_2214_),
    .B_N(_2222_),
    .Y(_2223_));
 sg13g2_inv_1 _6504_ (.Y(_2224_),
    .A(_2223_));
 sg13g2_xor2_1 _6505_ (.B(_2222_),
    .A(_2214_),
    .X(_2225_));
 sg13g2_a21oi_1 _6506_ (.A1(_2180_),
    .A2(_2186_),
    .Y(_2226_),
    .B1(_2190_));
 sg13g2_nand2_1 _6507_ (.Y(_2227_),
    .A(\i_mandel.i_xy.hc.genblk2[6].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[6].state.D ));
 sg13g2_xnor2_1 _6508_ (.Y(_2228_),
    .A(\i_mandel.i_xy.hc.genblk2[6].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[6].state.D ));
 sg13g2_o21ai_1 _6509_ (.B1(_2185_),
    .Y(_2229_),
    .A1(_2141_),
    .A2(_2183_));
 sg13g2_nand2_1 _6510_ (.Y(_2230_),
    .A(net908),
    .B(net920));
 sg13g2_nand2_1 _6511_ (.Y(_2231_),
    .A(net903),
    .B(net923));
 sg13g2_nand2_1 _6512_ (.Y(_2232_),
    .A(\i_mandel.i_xy.y[-8] ),
    .B(net923));
 sg13g2_xor2_1 _6513_ (.B(_2232_),
    .A(_2182_),
    .X(_2233_));
 sg13g2_nand2b_1 _6514_ (.Y(_2234_),
    .B(_2233_),
    .A_N(_2230_));
 sg13g2_xnor2_1 _6515_ (.Y(_2235_),
    .A(_2230_),
    .B(_2233_));
 sg13g2_nand2_1 _6516_ (.Y(_2236_),
    .A(_2229_),
    .B(_2235_));
 sg13g2_xnor2_1 _6517_ (.Y(_2237_),
    .A(_2229_),
    .B(_2235_));
 sg13g2_xor2_1 _6518_ (.B(_2237_),
    .A(_2228_),
    .X(_2238_));
 sg13g2_nand2b_1 _6519_ (.Y(_2239_),
    .B(_2238_),
    .A_N(_2178_));
 sg13g2_xnor2_1 _6520_ (.Y(_2240_),
    .A(_2178_),
    .B(_2238_));
 sg13g2_nand2b_1 _6521_ (.Y(_2241_),
    .B(_2240_),
    .A_N(_2226_));
 sg13g2_xor2_1 _6522_ (.B(_2240_),
    .A(_2226_),
    .X(_2242_));
 sg13g2_nor2_1 _6523_ (.A(_2225_),
    .B(_2242_),
    .Y(_2243_));
 sg13g2_xnor2_1 _6524_ (.Y(_2244_),
    .A(_2225_),
    .B(_2242_));
 sg13g2_xor2_1 _6525_ (.B(_2244_),
    .A(_2195_),
    .X(_2245_));
 sg13g2_xnor2_1 _6526_ (.Y(_2246_),
    .A(_2193_),
    .B(_2245_));
 sg13g2_nand2_1 _6527_ (.Y(_2247_),
    .A(_2198_),
    .B(_2246_));
 sg13g2_xnor2_1 _6528_ (.Y(_2248_),
    .A(_2198_),
    .B(_2246_));
 sg13g2_xor2_1 _6529_ (.B(_2248_),
    .A(_2188_),
    .X(_2249_));
 sg13g2_nand2_1 _6530_ (.Y(_2250_),
    .A(_2213_),
    .B(_2249_));
 sg13g2_xnor2_1 _6531_ (.Y(_2251_),
    .A(_2213_),
    .B(_2249_));
 sg13g2_xor2_1 _6532_ (.B(_2251_),
    .A(_2212_),
    .X(_2252_));
 sg13g2_nand2_1 _6533_ (.Y(_2253_),
    .A(\i_coord.y0[-11] ),
    .B(_2252_));
 sg13g2_xnor2_1 _6534_ (.Y(_2254_),
    .A(\i_coord.y0[-11] ),
    .B(_2252_));
 sg13g2_nand2_1 _6535_ (.Y(_2255_),
    .A(_2211_),
    .B(_2254_));
 sg13g2_or2_1 _6536_ (.X(_2256_),
    .B(_2254_),
    .A(_2211_));
 sg13g2_a21oi_1 _6537_ (.A1(_2255_),
    .A2(_2256_),
    .Y(_2257_),
    .B1(net839));
 sg13g2_a21oi_1 _6538_ (.A1(net839),
    .A2(_1766_),
    .Y(_2258_),
    .B1(_2257_));
 sg13g2_mux2_1 _6539_ (.A0(_2258_),
    .A1(net202),
    .S(net733),
    .X(_0152_));
 sg13g2_o21ai_1 _6540_ (.B1(_2250_),
    .Y(_2259_),
    .A1(_2212_),
    .A2(_2251_));
 sg13g2_o21ai_1 _6541_ (.B1(_2247_),
    .Y(_2260_),
    .A1(_2188_),
    .A2(_2248_));
 sg13g2_a21oi_2 _6542_ (.B1(_2244_),
    .Y(_2261_),
    .A2(_2195_),
    .A1(_2193_));
 sg13g2_and2_1 _6543_ (.A(_2239_),
    .B(_2241_),
    .X(_2262_));
 sg13g2_nand2_2 _6544_ (.Y(_2263_),
    .A(net933),
    .B(net891));
 sg13g2_nor2_2 _6545_ (.A(_2214_),
    .B(_2263_),
    .Y(_2264_));
 sg13g2_a22oi_1 _6546_ (.Y(_2265_),
    .B1(net891),
    .B2(net936),
    .A2(net892),
    .A1(net933));
 sg13g2_nor2_1 _6547_ (.A(_2264_),
    .B(_2265_),
    .Y(_2266_));
 sg13g2_nand2_1 _6548_ (.Y(_2267_),
    .A(net900),
    .B(net926));
 sg13g2_nand2_2 _6549_ (.Y(_2268_),
    .A(net928),
    .B(net894));
 sg13g2_nor2_1 _6550_ (.A(_2216_),
    .B(_2268_),
    .Y(_2269_));
 sg13g2_a22oi_1 _6551_ (.Y(_2270_),
    .B1(net894),
    .B2(net930),
    .A2(net928),
    .A1(net897));
 sg13g2_nor2_1 _6552_ (.A(_2269_),
    .B(_2270_),
    .Y(_2271_));
 sg13g2_nor3_1 _6553_ (.A(_2267_),
    .B(_2269_),
    .C(_2270_),
    .Y(_2272_));
 sg13g2_xnor2_1 _6554_ (.Y(_2273_),
    .A(_2267_),
    .B(_2271_));
 sg13g2_a21oi_1 _6555_ (.A1(_2215_),
    .A2(_2218_),
    .Y(_2274_),
    .B1(_2217_));
 sg13g2_nand2b_1 _6556_ (.Y(_2275_),
    .B(_2273_),
    .A_N(_2274_));
 sg13g2_xnor2_1 _6557_ (.Y(_2276_),
    .A(_2273_),
    .B(_2274_));
 sg13g2_and2_1 _6558_ (.A(_2266_),
    .B(_2276_),
    .X(_2277_));
 sg13g2_xnor2_1 _6559_ (.Y(_2278_),
    .A(_2266_),
    .B(_2276_));
 sg13g2_nor2_1 _6560_ (.A(_2224_),
    .B(_2278_),
    .Y(_2279_));
 sg13g2_nand2_1 _6561_ (.Y(_2280_),
    .A(_2224_),
    .B(_2278_));
 sg13g2_nand2b_1 _6562_ (.Y(_2281_),
    .B(_2280_),
    .A_N(_2279_));
 sg13g2_o21ai_1 _6563_ (.B1(_2236_),
    .Y(_2282_),
    .A1(_2228_),
    .A2(_2237_));
 sg13g2_nand2_1 _6564_ (.Y(_2283_),
    .A(\i_mandel.i_xy.hc.genblk2[7].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[7].state.D ));
 sg13g2_xnor2_1 _6565_ (.Y(_2284_),
    .A(\i_mandel.i_xy.hc.genblk2[7].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[7].state.D ));
 sg13g2_o21ai_1 _6566_ (.B1(_2234_),
    .Y(_2285_),
    .A1(_2182_),
    .A2(_2232_));
 sg13g2_nand2_1 _6567_ (.Y(_2286_),
    .A(net908),
    .B(net918));
 sg13g2_nand2_1 _6568_ (.Y(_2287_),
    .A(net903),
    .B(net920));
 sg13g2_nand2_1 _6569_ (.Y(_2288_),
    .A(net905),
    .B(net920));
 sg13g2_xor2_1 _6570_ (.B(_2288_),
    .A(_2231_),
    .X(_2289_));
 sg13g2_nand2b_1 _6571_ (.Y(_2290_),
    .B(_2289_),
    .A_N(_2286_));
 sg13g2_xnor2_1 _6572_ (.Y(_2291_),
    .A(_2286_),
    .B(_2289_));
 sg13g2_nand2_1 _6573_ (.Y(_2292_),
    .A(_2285_),
    .B(_2291_));
 sg13g2_xnor2_1 _6574_ (.Y(_2293_),
    .A(_2285_),
    .B(_2291_));
 sg13g2_xnor2_1 _6575_ (.Y(_2294_),
    .A(_2284_),
    .B(_2293_));
 sg13g2_nor2_1 _6576_ (.A(_2221_),
    .B(_2294_),
    .Y(_2295_));
 sg13g2_xor2_1 _6577_ (.B(_2294_),
    .A(_2221_),
    .X(_2296_));
 sg13g2_xor2_1 _6578_ (.B(_2296_),
    .A(_2282_),
    .X(_2297_));
 sg13g2_xnor2_1 _6579_ (.Y(_2298_),
    .A(_2281_),
    .B(_2297_));
 sg13g2_nand2_1 _6580_ (.Y(_2299_),
    .A(_2243_),
    .B(_2298_));
 sg13g2_xnor2_1 _6581_ (.Y(_2300_),
    .A(_2243_),
    .B(_2298_));
 sg13g2_xor2_1 _6582_ (.B(_2300_),
    .A(_2262_),
    .X(_2301_));
 sg13g2_nand2_1 _6583_ (.Y(_2302_),
    .A(_2261_),
    .B(_2301_));
 sg13g2_nor2_1 _6584_ (.A(_2261_),
    .B(_2301_),
    .Y(_2303_));
 sg13g2_xor2_1 _6585_ (.B(_2301_),
    .A(_2261_),
    .X(_2304_));
 sg13g2_xnor2_1 _6586_ (.Y(_2305_),
    .A(_2227_),
    .B(_2304_));
 sg13g2_and2_1 _6587_ (.A(_2260_),
    .B(_2305_),
    .X(_2306_));
 sg13g2_or2_1 _6588_ (.X(_2307_),
    .B(_2305_),
    .A(_2260_));
 sg13g2_xnor2_1 _6589_ (.Y(_2308_),
    .A(_2260_),
    .B(_2305_));
 sg13g2_xnor2_1 _6590_ (.Y(_2309_),
    .A(_2259_),
    .B(_2308_));
 sg13g2_nand2_1 _6591_ (.Y(_2310_),
    .A(\i_coord.y0[-10] ),
    .B(_2309_));
 sg13g2_xnor2_1 _6592_ (.Y(_2311_),
    .A(\i_coord.y0[-10] ),
    .B(_2309_));
 sg13g2_a21o_1 _6593_ (.A2(_2256_),
    .A1(_2253_),
    .B1(_2311_),
    .X(_2312_));
 sg13g2_nand3_1 _6594_ (.B(_2256_),
    .C(_2311_),
    .A(_2253_),
    .Y(_2313_));
 sg13g2_and2_1 _6595_ (.A(net836),
    .B(_2313_),
    .X(_2314_));
 sg13g2_a22oi_1 _6596_ (.Y(_2315_),
    .B1(_2312_),
    .B2(_2314_),
    .A2(_1779_),
    .A1(net839));
 sg13g2_nand2_1 _6597_ (.Y(_2316_),
    .A(net188),
    .B(net734));
 sg13g2_o21ai_1 _6598_ (.B1(_2316_),
    .Y(_0153_),
    .A1(net734),
    .A2(_2315_));
 sg13g2_nor2_1 _6599_ (.A(net836),
    .B(_1790_),
    .Y(_2317_));
 sg13g2_a21oi_1 _6600_ (.A1(_2259_),
    .A2(_2307_),
    .Y(_2318_),
    .B1(_2306_));
 sg13g2_o21ai_1 _6601_ (.B1(_2302_),
    .Y(_2319_),
    .A1(_2227_),
    .A2(_2303_));
 sg13g2_o21ai_1 _6602_ (.B1(_2299_),
    .Y(_2320_),
    .A1(_2262_),
    .A2(_2300_));
 sg13g2_a21oi_1 _6603_ (.A1(_2282_),
    .A2(_2296_),
    .Y(_2321_),
    .B1(_2295_));
 sg13g2_a21o_1 _6604_ (.A2(_2297_),
    .A1(_2280_),
    .B1(_2279_),
    .X(_2322_));
 sg13g2_nand2_1 _6605_ (.Y(_2323_),
    .A(net930),
    .B(net892));
 sg13g2_nand2_1 _6606_ (.Y(_2324_),
    .A(net932),
    .B(net887));
 sg13g2_nand2_1 _6607_ (.Y(_2325_),
    .A(net935),
    .B(net887));
 sg13g2_or2_1 _6608_ (.X(_2326_),
    .B(_2325_),
    .A(_2263_));
 sg13g2_xor2_1 _6609_ (.B(_2325_),
    .A(_2263_),
    .X(_2327_));
 sg13g2_nand2b_1 _6610_ (.Y(_2328_),
    .B(_2327_),
    .A_N(_2323_));
 sg13g2_xnor2_1 _6611_ (.Y(_2329_),
    .A(_2323_),
    .B(_2327_));
 sg13g2_nand2_1 _6612_ (.Y(_2330_),
    .A(net900),
    .B(net924));
 sg13g2_nand2_2 _6613_ (.Y(_2331_),
    .A(net897),
    .B(net926));
 sg13g2_xor2_1 _6614_ (.B(_2331_),
    .A(_2268_),
    .X(_2332_));
 sg13g2_nand2b_1 _6615_ (.Y(_2333_),
    .B(_2332_),
    .A_N(_2330_));
 sg13g2_xnor2_1 _6616_ (.Y(_2334_),
    .A(_2330_),
    .B(_2332_));
 sg13g2_nand2_1 _6617_ (.Y(_2335_),
    .A(_2264_),
    .B(_2334_));
 sg13g2_xor2_1 _6618_ (.B(_2334_),
    .A(_2264_),
    .X(_2336_));
 sg13g2_nor3_1 _6619_ (.A(_2269_),
    .B(_2272_),
    .C(_2336_),
    .Y(_2337_));
 sg13g2_o21ai_1 _6620_ (.B1(_2336_),
    .Y(_2338_),
    .A1(_2269_),
    .A2(_2272_));
 sg13g2_nor2b_1 _6621_ (.A(_2337_),
    .B_N(_2338_),
    .Y(_2339_));
 sg13g2_nand2_1 _6622_ (.Y(_2340_),
    .A(_2329_),
    .B(_2339_));
 sg13g2_inv_1 _6623_ (.Y(_2341_),
    .A(_2340_));
 sg13g2_xor2_1 _6624_ (.B(_2339_),
    .A(_2329_),
    .X(_2342_));
 sg13g2_and2_1 _6625_ (.A(_2277_),
    .B(_2342_),
    .X(_2343_));
 sg13g2_or2_1 _6626_ (.X(_2344_),
    .B(_2342_),
    .A(_2277_));
 sg13g2_nand2b_1 _6627_ (.Y(_2345_),
    .B(_2344_),
    .A_N(_2343_));
 sg13g2_o21ai_1 _6628_ (.B1(_2292_),
    .Y(_2346_),
    .A1(_2284_),
    .A2(_2293_));
 sg13g2_nand2_1 _6629_ (.Y(_2347_),
    .A(\i_mandel.i_xy.hc.genblk2[8].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[8].state.D ));
 sg13g2_xnor2_1 _6630_ (.Y(_2348_),
    .A(\i_mandel.i_xy.hc.genblk2[8].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[8].state.D ));
 sg13g2_o21ai_1 _6631_ (.B1(_2290_),
    .Y(_2349_),
    .A1(_2231_),
    .A2(_2288_));
 sg13g2_nand2_1 _6632_ (.Y(_2350_),
    .A(net908),
    .B(net917));
 sg13g2_nand2_1 _6633_ (.Y(_2351_),
    .A(net903),
    .B(net919));
 sg13g2_nand2_2 _6634_ (.Y(_2352_),
    .A(net905),
    .B(net918));
 sg13g2_xor2_1 _6635_ (.B(_2352_),
    .A(_2287_),
    .X(_2353_));
 sg13g2_nand2b_1 _6636_ (.Y(_2354_),
    .B(_2353_),
    .A_N(_2350_));
 sg13g2_xnor2_1 _6637_ (.Y(_2355_),
    .A(_2350_),
    .B(_2353_));
 sg13g2_nand2_1 _6638_ (.Y(_2356_),
    .A(_2349_),
    .B(_2355_));
 sg13g2_xnor2_1 _6639_ (.Y(_2357_),
    .A(_2349_),
    .B(_2355_));
 sg13g2_xor2_1 _6640_ (.B(_2357_),
    .A(_2348_),
    .X(_2358_));
 sg13g2_nor2b_1 _6641_ (.A(_2275_),
    .B_N(_2358_),
    .Y(_2359_));
 sg13g2_xnor2_1 _6642_ (.Y(_2360_),
    .A(_2275_),
    .B(_2358_));
 sg13g2_xor2_1 _6643_ (.B(_2360_),
    .A(_2346_),
    .X(_2361_));
 sg13g2_xnor2_1 _6644_ (.Y(_2362_),
    .A(_2345_),
    .B(_2361_));
 sg13g2_nand2_1 _6645_ (.Y(_2363_),
    .A(_2322_),
    .B(_2362_));
 sg13g2_xnor2_1 _6646_ (.Y(_2364_),
    .A(_2322_),
    .B(_2362_));
 sg13g2_xor2_1 _6647_ (.B(_2364_),
    .A(_2321_),
    .X(_2365_));
 sg13g2_nand2_1 _6648_ (.Y(_2366_),
    .A(_2320_),
    .B(_2365_));
 sg13g2_xnor2_1 _6649_ (.Y(_2367_),
    .A(_2320_),
    .B(_2365_));
 sg13g2_xor2_1 _6650_ (.B(_2367_),
    .A(_2283_),
    .X(_2368_));
 sg13g2_nand2_1 _6651_ (.Y(_2369_),
    .A(_2319_),
    .B(_2368_));
 sg13g2_xnor2_1 _6652_ (.Y(_2370_),
    .A(_2319_),
    .B(_2368_));
 sg13g2_xor2_1 _6653_ (.B(_2370_),
    .A(_2318_),
    .X(_2371_));
 sg13g2_nand2_1 _6654_ (.Y(_2372_),
    .A(\i_coord.y0[-9] ),
    .B(_2371_));
 sg13g2_xnor2_1 _6655_ (.Y(_2373_),
    .A(\i_coord.y0[-9] ),
    .B(_2371_));
 sg13g2_nand3_1 _6656_ (.B(_2312_),
    .C(_2373_),
    .A(_2310_),
    .Y(_2374_));
 sg13g2_a21o_1 _6657_ (.A2(_2312_),
    .A1(_2310_),
    .B1(_2373_),
    .X(_2375_));
 sg13g2_a21oi_1 _6658_ (.A1(_2374_),
    .A2(_2375_),
    .Y(_2376_),
    .B1(net840));
 sg13g2_nor2_1 _6659_ (.A(_2317_),
    .B(_2376_),
    .Y(_2377_));
 sg13g2_mux2_1 _6660_ (.A0(_2377_),
    .A1(net907),
    .S(net733),
    .X(_0154_));
 sg13g2_nor2_1 _6661_ (.A(net836),
    .B(_1802_),
    .Y(_2378_));
 sg13g2_o21ai_1 _6662_ (.B1(_2369_),
    .Y(_2379_),
    .A1(_2318_),
    .A2(_2370_));
 sg13g2_o21ai_1 _6663_ (.B1(_2366_),
    .Y(_2380_),
    .A1(_2283_),
    .A2(_2367_));
 sg13g2_o21ai_1 _6664_ (.B1(_2363_),
    .Y(_2381_),
    .A1(_2321_),
    .A2(_2364_));
 sg13g2_a21oi_1 _6665_ (.A1(_2346_),
    .A2(_2360_),
    .Y(_2382_),
    .B1(_2359_));
 sg13g2_a21o_1 _6666_ (.A2(_2361_),
    .A1(_2344_),
    .B1(_2343_),
    .X(_2383_));
 sg13g2_nand2_2 _6667_ (.Y(_2384_),
    .A(net935),
    .B(net885));
 sg13g2_nand2_1 _6668_ (.Y(_2385_),
    .A(net928),
    .B(net892));
 sg13g2_nand2_2 _6669_ (.Y(_2386_),
    .A(net930),
    .B(net888));
 sg13g2_nand2_1 _6670_ (.Y(_2387_),
    .A(net930),
    .B(net891));
 sg13g2_or2_1 _6671_ (.X(_2388_),
    .B(_2386_),
    .A(_2263_));
 sg13g2_xor2_1 _6672_ (.B(_2387_),
    .A(_2324_),
    .X(_2389_));
 sg13g2_nand2b_1 _6673_ (.Y(_2390_),
    .B(_2389_),
    .A_N(_2385_));
 sg13g2_xnor2_1 _6674_ (.Y(_2391_),
    .A(_2385_),
    .B(_2389_));
 sg13g2_nand2b_1 _6675_ (.Y(_2392_),
    .B(_2391_),
    .A_N(_2384_));
 sg13g2_xnor2_1 _6676_ (.Y(_2393_),
    .A(_2384_),
    .B(_2391_));
 sg13g2_o21ai_1 _6677_ (.B1(_2333_),
    .Y(_2394_),
    .A1(_2268_),
    .A2(_2331_));
 sg13g2_and2_1 _6678_ (.A(_2326_),
    .B(_2328_),
    .X(_2395_));
 sg13g2_nand2_1 _6679_ (.Y(_2396_),
    .A(net900),
    .B(net921));
 sg13g2_nand2_2 _6680_ (.Y(_2397_),
    .A(net894),
    .B(net924));
 sg13g2_nor2_1 _6681_ (.A(_2331_),
    .B(_2397_),
    .Y(_2398_));
 sg13g2_a22oi_1 _6682_ (.Y(_2399_),
    .B1(net924),
    .B2(net897),
    .A2(net894),
    .A1(net926));
 sg13g2_nor2_1 _6683_ (.A(_2398_),
    .B(_2399_),
    .Y(_2400_));
 sg13g2_nand2b_1 _6684_ (.Y(_2401_),
    .B(_2400_),
    .A_N(_2396_));
 sg13g2_xnor2_1 _6685_ (.Y(_2402_),
    .A(_2396_),
    .B(_2400_));
 sg13g2_nor2b_1 _6686_ (.A(_2395_),
    .B_N(_2402_),
    .Y(_2403_));
 sg13g2_xnor2_1 _6687_ (.Y(_2404_),
    .A(_2395_),
    .B(_2402_));
 sg13g2_xnor2_1 _6688_ (.Y(_2405_),
    .A(_2394_),
    .B(_2404_));
 sg13g2_inv_1 _6689_ (.Y(_2406_),
    .A(_2405_));
 sg13g2_nand2_1 _6690_ (.Y(_2407_),
    .A(_2393_),
    .B(_2406_));
 sg13g2_xnor2_1 _6691_ (.Y(_2408_),
    .A(_2393_),
    .B(_2405_));
 sg13g2_xnor2_1 _6692_ (.Y(_2409_),
    .A(_2340_),
    .B(_2408_));
 sg13g2_inv_1 _6693_ (.Y(_2410_),
    .A(_2409_));
 sg13g2_o21ai_1 _6694_ (.B1(_2356_),
    .Y(_2411_),
    .A1(_2348_),
    .A2(_2357_));
 sg13g2_nand2_1 _6695_ (.Y(_2412_),
    .A(_2335_),
    .B(_2338_));
 sg13g2_nand2_1 _6696_ (.Y(_2413_),
    .A(\i_mandel.i_xy.hc.genblk2[9].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[9].state.D ));
 sg13g2_xnor2_1 _6697_ (.Y(_2414_),
    .A(\i_mandel.i_xy.hc.genblk2[9].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[9].state.D ));
 sg13g2_o21ai_1 _6698_ (.B1(_2354_),
    .Y(_2415_),
    .A1(_2287_),
    .A2(_2352_));
 sg13g2_nand2_1 _6699_ (.Y(_2416_),
    .A(net908),
    .B(net914));
 sg13g2_nand2_2 _6700_ (.Y(_2417_),
    .A(net903),
    .B(net917));
 sg13g2_nand2_1 _6701_ (.Y(_2418_),
    .A(net905),
    .B(net917));
 sg13g2_xor2_1 _6702_ (.B(_2418_),
    .A(_2351_),
    .X(_2419_));
 sg13g2_nand2b_1 _6703_ (.Y(_2420_),
    .B(_2419_),
    .A_N(_2416_));
 sg13g2_xnor2_1 _6704_ (.Y(_2421_),
    .A(_2416_),
    .B(_2419_));
 sg13g2_nand2_1 _6705_ (.Y(_2422_),
    .A(_2415_),
    .B(_2421_));
 sg13g2_xnor2_1 _6706_ (.Y(_2423_),
    .A(_2415_),
    .B(_2421_));
 sg13g2_xor2_1 _6707_ (.B(_2423_),
    .A(_2414_),
    .X(_2424_));
 sg13g2_xnor2_1 _6708_ (.Y(_2425_),
    .A(_2412_),
    .B(_2424_));
 sg13g2_nor2b_1 _6709_ (.A(_2425_),
    .B_N(_2411_),
    .Y(_2426_));
 sg13g2_xor2_1 _6710_ (.B(_2425_),
    .A(_2411_),
    .X(_2427_));
 sg13g2_nor2_1 _6711_ (.A(_2410_),
    .B(_2427_),
    .Y(_2428_));
 sg13g2_xnor2_1 _6712_ (.Y(_2429_),
    .A(_2410_),
    .B(_2427_));
 sg13g2_nand2b_1 _6713_ (.Y(_2430_),
    .B(_2383_),
    .A_N(_2429_));
 sg13g2_xor2_1 _6714_ (.B(_2429_),
    .A(_2383_),
    .X(_2431_));
 sg13g2_xor2_1 _6715_ (.B(_2431_),
    .A(_2382_),
    .X(_2432_));
 sg13g2_nand2_1 _6716_ (.Y(_2433_),
    .A(_2381_),
    .B(_2432_));
 sg13g2_xnor2_1 _6717_ (.Y(_2434_),
    .A(_2381_),
    .B(_2432_));
 sg13g2_xor2_1 _6718_ (.B(_2434_),
    .A(_2347_),
    .X(_2435_));
 sg13g2_and2_1 _6719_ (.A(_2380_),
    .B(_2435_),
    .X(_2436_));
 sg13g2_or2_1 _6720_ (.X(_2437_),
    .B(_2435_),
    .A(_2380_));
 sg13g2_xnor2_1 _6721_ (.Y(_2438_),
    .A(_2380_),
    .B(_2435_));
 sg13g2_xnor2_1 _6722_ (.Y(_2439_),
    .A(_2379_),
    .B(_2438_));
 sg13g2_nand2_1 _6723_ (.Y(_2440_),
    .A(net937),
    .B(_2439_));
 sg13g2_xnor2_1 _6724_ (.Y(_2441_),
    .A(net937),
    .B(_2439_));
 sg13g2_nand3_1 _6725_ (.B(_2375_),
    .C(_2441_),
    .A(_2372_),
    .Y(_2442_));
 sg13g2_a21o_1 _6726_ (.A2(_2375_),
    .A1(_2372_),
    .B1(_2441_),
    .X(_2443_));
 sg13g2_a21oi_1 _6727_ (.A1(_2442_),
    .A2(_2443_),
    .Y(_2444_),
    .B1(net840));
 sg13g2_nor2_1 _6728_ (.A(_2378_),
    .B(_2444_),
    .Y(_2445_));
 sg13g2_mux2_1 _6729_ (.A0(_2445_),
    .A1(net906),
    .S(net735),
    .X(_0155_));
 sg13g2_a21o_1 _6730_ (.A2(_2437_),
    .A1(_2379_),
    .B1(_2436_),
    .X(_2446_));
 sg13g2_o21ai_1 _6731_ (.B1(_2433_),
    .Y(_2447_),
    .A1(_2347_),
    .A2(_2434_));
 sg13g2_o21ai_1 _6732_ (.B1(_2430_),
    .Y(_2448_),
    .A1(_2382_),
    .A2(_2431_));
 sg13g2_a21o_1 _6733_ (.A2(_2424_),
    .A1(_2412_),
    .B1(_2426_),
    .X(_2449_));
 sg13g2_a21oi_1 _6734_ (.A1(_2341_),
    .A2(_2408_),
    .Y(_2450_),
    .B1(_2428_));
 sg13g2_nand2_1 _6735_ (.Y(_2451_),
    .A(net932),
    .B(\i_mandel.i_xy.y[1] ));
 sg13g2_nor2_1 _6736_ (.A(_2384_),
    .B(_2451_),
    .Y(_2452_));
 sg13g2_a22oi_1 _6737_ (.Y(_2453_),
    .B1(net883),
    .B2(net935),
    .A2(net885),
    .A1(net932));
 sg13g2_nor2_1 _6738_ (.A(_2452_),
    .B(_2453_),
    .Y(_2454_));
 sg13g2_nand2_1 _6739_ (.Y(_2455_),
    .A(net926),
    .B(net892));
 sg13g2_nand2_1 _6740_ (.Y(_2456_),
    .A(net928),
    .B(net891));
 sg13g2_or2_1 _6741_ (.X(_2457_),
    .B(_2456_),
    .A(_2386_));
 sg13g2_xor2_1 _6742_ (.B(_2456_),
    .A(_2386_),
    .X(_2458_));
 sg13g2_nand2b_1 _6743_ (.Y(_2459_),
    .B(_2458_),
    .A_N(_2455_));
 sg13g2_xnor2_1 _6744_ (.Y(_2460_),
    .A(_2455_),
    .B(_2458_));
 sg13g2_nand2_1 _6745_ (.Y(_2461_),
    .A(_2454_),
    .B(_2460_));
 sg13g2_xor2_1 _6746_ (.B(_2460_),
    .A(_2454_),
    .X(_2462_));
 sg13g2_nand2b_1 _6747_ (.Y(_2463_),
    .B(_2462_),
    .A_N(_2392_));
 sg13g2_xnor2_1 _6748_ (.Y(_2464_),
    .A(_2392_),
    .B(_2462_));
 sg13g2_inv_1 _6749_ (.Y(_2465_),
    .A(_2464_));
 sg13g2_o21ai_1 _6750_ (.B1(_2401_),
    .Y(_2466_),
    .A1(_2331_),
    .A2(_2397_));
 sg13g2_and2_1 _6751_ (.A(_2388_),
    .B(_2390_),
    .X(_2467_));
 sg13g2_nand2_1 _6752_ (.Y(_2468_),
    .A(net897),
    .B(net920));
 sg13g2_xor2_1 _6753_ (.B(_2468_),
    .A(_2397_),
    .X(_2469_));
 sg13g2_nand3_1 _6754_ (.B(net918),
    .C(_2469_),
    .A(net900),
    .Y(_2470_));
 sg13g2_a21o_1 _6755_ (.A2(net918),
    .A1(net900),
    .B1(_2469_),
    .X(_2471_));
 sg13g2_and2_1 _6756_ (.A(_2470_),
    .B(_2471_),
    .X(_2472_));
 sg13g2_nor2b_1 _6757_ (.A(_2467_),
    .B_N(_2472_),
    .Y(_2473_));
 sg13g2_xnor2_1 _6758_ (.Y(_2474_),
    .A(_2467_),
    .B(_2472_));
 sg13g2_xnor2_1 _6759_ (.Y(_2475_),
    .A(_2466_),
    .B(_2474_));
 sg13g2_xnor2_1 _6760_ (.Y(_2476_),
    .A(_2465_),
    .B(_2475_));
 sg13g2_nor2_1 _6761_ (.A(_2407_),
    .B(_2476_),
    .Y(_2477_));
 sg13g2_xor2_1 _6762_ (.B(_2476_),
    .A(_2407_),
    .X(_2478_));
 sg13g2_inv_1 _6763_ (.Y(_2479_),
    .A(_2478_));
 sg13g2_o21ai_1 _6764_ (.B1(_2422_),
    .Y(_2480_),
    .A1(_2414_),
    .A2(_2423_));
 sg13g2_a21o_1 _6765_ (.A2(_2404_),
    .A1(_2394_),
    .B1(_2403_),
    .X(_2481_));
 sg13g2_o21ai_1 _6766_ (.B1(_2420_),
    .Y(_2482_),
    .A1(_2352_),
    .A2(_2417_));
 sg13g2_nand2_1 _6767_ (.Y(_2483_),
    .A(net908),
    .B(net912));
 sg13g2_nand2_1 _6768_ (.Y(_2484_),
    .A(net903),
    .B(net914));
 sg13g2_nand2_1 _6769_ (.Y(_2485_),
    .A(net905),
    .B(net914));
 sg13g2_xor2_1 _6770_ (.B(_2485_),
    .A(_2417_),
    .X(_2486_));
 sg13g2_nand2b_1 _6771_ (.Y(_2487_),
    .B(_2486_),
    .A_N(_2483_));
 sg13g2_xnor2_1 _6772_ (.Y(_2488_),
    .A(_2483_),
    .B(_2486_));
 sg13g2_nand2_1 _6773_ (.Y(_2489_),
    .A(_2482_),
    .B(_2488_));
 sg13g2_xnor2_1 _6774_ (.Y(_2490_),
    .A(_2482_),
    .B(_2488_));
 sg13g2_nand2_1 _6775_ (.Y(_2491_),
    .A(\i_mandel.i_xy.hc.genblk2[10].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[10].state.D ));
 sg13g2_xnor2_1 _6776_ (.Y(_2492_),
    .A(\i_mandel.i_xy.hc.genblk2[10].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[10].state.D ));
 sg13g2_xor2_1 _6777_ (.B(_2492_),
    .A(_2490_),
    .X(_2493_));
 sg13g2_and2_1 _6778_ (.A(_2481_),
    .B(_2493_),
    .X(_2494_));
 sg13g2_xor2_1 _6779_ (.B(_2493_),
    .A(_2481_),
    .X(_2495_));
 sg13g2_xnor2_1 _6780_ (.Y(_2496_),
    .A(_2480_),
    .B(_2495_));
 sg13g2_nor2_1 _6781_ (.A(_2479_),
    .B(_2496_),
    .Y(_2497_));
 sg13g2_xnor2_1 _6782_ (.Y(_2498_),
    .A(_2479_),
    .B(_2496_));
 sg13g2_nor2_1 _6783_ (.A(_2450_),
    .B(_2498_),
    .Y(_2499_));
 sg13g2_xor2_1 _6784_ (.B(_2498_),
    .A(_2450_),
    .X(_2500_));
 sg13g2_xor2_1 _6785_ (.B(_2500_),
    .A(_2449_),
    .X(_2501_));
 sg13g2_nand2_1 _6786_ (.Y(_2502_),
    .A(_2448_),
    .B(_2501_));
 sg13g2_xnor2_1 _6787_ (.Y(_2503_),
    .A(_2448_),
    .B(_2501_));
 sg13g2_xor2_1 _6788_ (.B(_2503_),
    .A(_2413_),
    .X(_2504_));
 sg13g2_and2_1 _6789_ (.A(_2447_),
    .B(_2504_),
    .X(_2505_));
 sg13g2_or2_1 _6790_ (.X(_2506_),
    .B(_2504_),
    .A(_2447_));
 sg13g2_xor2_1 _6791_ (.B(_2504_),
    .A(_2447_),
    .X(_2507_));
 sg13g2_xnor2_1 _6792_ (.Y(_2508_),
    .A(_2446_),
    .B(_2507_));
 sg13g2_xnor2_1 _6793_ (.Y(_2509_),
    .A(_3121_),
    .B(_2508_));
 sg13g2_a21o_1 _6794_ (.A2(_2443_),
    .A1(_2440_),
    .B1(_2509_),
    .X(_2510_));
 sg13g2_nand3_1 _6795_ (.B(_2443_),
    .C(_2509_),
    .A(_2440_),
    .Y(_2511_));
 sg13g2_a21oi_1 _6796_ (.A1(_2510_),
    .A2(_2511_),
    .Y(_2512_),
    .B1(net840));
 sg13g2_a21oi_1 _6797_ (.A1(net840),
    .A2(_1815_),
    .Y(_2513_),
    .B1(_2512_));
 sg13g2_mux2_1 _6798_ (.A0(_2513_),
    .A1(net904),
    .S(net735),
    .X(_0156_));
 sg13g2_nor2_1 _6799_ (.A(net834),
    .B(_1827_),
    .Y(_2514_));
 sg13g2_or2_1 _6800_ (.X(_2515_),
    .B(_2508_),
    .A(_0024_));
 sg13g2_a21oi_2 _6801_ (.B1(_2505_),
    .Y(_2516_),
    .A2(_2506_),
    .A1(_2446_));
 sg13g2_o21ai_1 _6802_ (.B1(_2502_),
    .Y(_2517_),
    .A1(_2413_),
    .A2(_2503_));
 sg13g2_a21oi_1 _6803_ (.A1(_2449_),
    .A2(_2500_),
    .Y(_2518_),
    .B1(_2499_));
 sg13g2_a21oi_1 _6804_ (.A1(_2480_),
    .A2(_2495_),
    .Y(_2519_),
    .B1(_2494_));
 sg13g2_nor2_1 _6805_ (.A(_2477_),
    .B(_2497_),
    .Y(_2520_));
 sg13g2_o21ai_1 _6806_ (.B1(_2463_),
    .Y(_2521_),
    .A1(_2465_),
    .A2(_2475_));
 sg13g2_nand2_1 _6807_ (.Y(_2522_),
    .A(net927),
    .B(net891));
 sg13g2_nand2_1 _6808_ (.Y(_2523_),
    .A(net928),
    .B(net885));
 sg13g2_nor2_1 _6809_ (.A(_2386_),
    .B(_2523_),
    .Y(_2524_));
 sg13g2_a22oi_1 _6810_ (.Y(_2525_),
    .B1(net885),
    .B2(net931),
    .A2(net887),
    .A1(net928));
 sg13g2_nor3_1 _6811_ (.A(_2522_),
    .B(_2524_),
    .C(_2525_),
    .Y(_2526_));
 sg13g2_o21ai_1 _6812_ (.B1(_2522_),
    .Y(_2527_),
    .A1(_2524_),
    .A2(_2525_));
 sg13g2_nor2b_1 _6813_ (.A(_2526_),
    .B_N(_2527_),
    .Y(_2528_));
 sg13g2_nand2_1 _6814_ (.Y(_2529_),
    .A(net935),
    .B(\i_mandel.i_xy.y[2] ));
 sg13g2_nor2b_1 _6815_ (.A(_2451_),
    .B_N(_2384_),
    .Y(_2530_));
 sg13g2_xnor2_1 _6816_ (.Y(_2531_),
    .A(_2529_),
    .B(_2530_));
 sg13g2_xnor2_1 _6817_ (.Y(_2532_),
    .A(_2528_),
    .B(_2531_));
 sg13g2_nor2_1 _6818_ (.A(_2461_),
    .B(_2532_),
    .Y(_2533_));
 sg13g2_xor2_1 _6819_ (.B(_2532_),
    .A(_2461_),
    .X(_2534_));
 sg13g2_o21ai_1 _6820_ (.B1(_2470_),
    .Y(_2535_),
    .A1(_2397_),
    .A2(_2468_));
 sg13g2_and2_1 _6821_ (.A(_2457_),
    .B(_2459_),
    .X(_2536_));
 sg13g2_nand2_2 _6822_ (.Y(_2537_),
    .A(net897),
    .B(net918));
 sg13g2_nand2_1 _6823_ (.Y(_2538_),
    .A(net892),
    .B(net921));
 sg13g2_nor2_1 _6824_ (.A(_2397_),
    .B(_2538_),
    .Y(_2539_));
 sg13g2_or2_1 _6825_ (.X(_2540_),
    .B(_2538_),
    .A(_2397_));
 sg13g2_a22oi_1 _6826_ (.Y(_2541_),
    .B1(net920),
    .B2(net895),
    .A2(net892),
    .A1(net923));
 sg13g2_nor2_1 _6827_ (.A(_2539_),
    .B(_2541_),
    .Y(_2542_));
 sg13g2_xnor2_1 _6828_ (.Y(_2543_),
    .A(_2537_),
    .B(_2542_));
 sg13g2_nor2b_1 _6829_ (.A(_2536_),
    .B_N(_2543_),
    .Y(_2544_));
 sg13g2_xnor2_1 _6830_ (.Y(_2545_),
    .A(_2536_),
    .B(_2543_));
 sg13g2_xnor2_1 _6831_ (.Y(_2546_),
    .A(_2535_),
    .B(_2545_));
 sg13g2_inv_1 _6832_ (.Y(_2547_),
    .A(_2546_));
 sg13g2_xnor2_1 _6833_ (.Y(_2548_),
    .A(_2534_),
    .B(_2546_));
 sg13g2_and2_1 _6834_ (.A(_2521_),
    .B(_2548_),
    .X(_2549_));
 sg13g2_xor2_1 _6835_ (.B(_2548_),
    .A(_2521_),
    .X(_2550_));
 sg13g2_o21ai_1 _6836_ (.B1(_2489_),
    .Y(_2551_),
    .A1(_2490_),
    .A2(_2492_));
 sg13g2_a21o_1 _6837_ (.A2(_2474_),
    .A1(_2466_),
    .B1(_2473_),
    .X(_2552_));
 sg13g2_nand2_2 _6838_ (.Y(_2553_),
    .A(net908),
    .B(net909));
 sg13g2_xor2_1 _6839_ (.B(_2553_),
    .A(_1304_),
    .X(_2554_));
 sg13g2_nand2_1 _6840_ (.Y(_2555_),
    .A(\i_mandel.i_xy.hc.genblk2[11].state.Q ),
    .B(_2554_));
 sg13g2_xnor2_1 _6841_ (.Y(_2556_),
    .A(\i_mandel.i_xy.hc.genblk2[11].state.Q ),
    .B(_2554_));
 sg13g2_o21ai_1 _6842_ (.B1(_2487_),
    .Y(_2557_),
    .A1(_2418_),
    .A2(_2484_));
 sg13g2_nand2_1 _6843_ (.Y(_2558_),
    .A(net906),
    .B(net912));
 sg13g2_nand2_1 _6844_ (.Y(_2559_),
    .A(net901),
    .B(net914));
 sg13g2_nand2_1 _6845_ (.Y(_2560_),
    .A(net900),
    .B(net917));
 sg13g2_xor2_1 _6846_ (.B(_2560_),
    .A(_2484_),
    .X(_2561_));
 sg13g2_nand2b_1 _6847_ (.Y(_2562_),
    .B(_2561_),
    .A_N(_2558_));
 sg13g2_xnor2_1 _6848_ (.Y(_2563_),
    .A(_2558_),
    .B(_2561_));
 sg13g2_nand2_1 _6849_ (.Y(_2564_),
    .A(_2557_),
    .B(_2563_));
 sg13g2_xnor2_1 _6850_ (.Y(_2565_),
    .A(_2557_),
    .B(_2563_));
 sg13g2_xor2_1 _6851_ (.B(_2565_),
    .A(_2556_),
    .X(_2566_));
 sg13g2_xnor2_1 _6852_ (.Y(_2567_),
    .A(_2552_),
    .B(_2566_));
 sg13g2_nor2b_1 _6853_ (.A(_2567_),
    .B_N(_2551_),
    .Y(_2568_));
 sg13g2_xnor2_1 _6854_ (.Y(_2569_),
    .A(_2551_),
    .B(_2567_));
 sg13g2_xnor2_1 _6855_ (.Y(_2570_),
    .A(_2550_),
    .B(_2569_));
 sg13g2_nor2_1 _6856_ (.A(_2520_),
    .B(_2570_),
    .Y(_2571_));
 sg13g2_xor2_1 _6857_ (.B(_2570_),
    .A(_2520_),
    .X(_2572_));
 sg13g2_nor2b_1 _6858_ (.A(_2519_),
    .B_N(_2572_),
    .Y(_2573_));
 sg13g2_xnor2_1 _6859_ (.Y(_2574_),
    .A(_2519_),
    .B(_2572_));
 sg13g2_nand2b_1 _6860_ (.Y(_2575_),
    .B(_2574_),
    .A_N(_2518_));
 sg13g2_xnor2_1 _6861_ (.Y(_2576_),
    .A(_2518_),
    .B(_2574_));
 sg13g2_nand2b_1 _6862_ (.Y(_2577_),
    .B(_2576_),
    .A_N(_2491_));
 sg13g2_xnor2_1 _6863_ (.Y(_2578_),
    .A(_2491_),
    .B(_2576_));
 sg13g2_nand2_1 _6864_ (.Y(_2579_),
    .A(_2517_),
    .B(_2578_));
 sg13g2_xnor2_1 _6865_ (.Y(_2580_),
    .A(_2517_),
    .B(_2578_));
 sg13g2_xor2_1 _6866_ (.B(_2580_),
    .A(_2516_),
    .X(_2581_));
 sg13g2_and2_1 _6867_ (.A(\i_coord.y0[-6] ),
    .B(_2581_),
    .X(_2582_));
 sg13g2_xnor2_1 _6868_ (.Y(_2583_),
    .A(\i_coord.y0[-6] ),
    .B(_2581_));
 sg13g2_and3_1 _6869_ (.X(_2584_),
    .A(_2510_),
    .B(_2515_),
    .C(_2583_));
 sg13g2_a21oi_1 _6870_ (.A1(_2510_),
    .A2(_2515_),
    .Y(_2585_),
    .B1(_2583_));
 sg13g2_or2_1 _6871_ (.X(_2586_),
    .B(_2585_),
    .A(_2584_));
 sg13g2_a21oi_1 _6872_ (.A1(net834),
    .A2(_2586_),
    .Y(_2587_),
    .B1(_2514_));
 sg13g2_mux2_1 _6873_ (.A0(_2587_),
    .A1(net319),
    .S(net736),
    .X(_0157_));
 sg13g2_o21ai_1 _6874_ (.B1(_2579_),
    .Y(_2588_),
    .A1(_2516_),
    .A2(_2580_));
 sg13g2_nand2_2 _6875_ (.Y(_2589_),
    .A(_2575_),
    .B(_2577_));
 sg13g2_o21ai_1 _6876_ (.B1(_2555_),
    .Y(_2590_),
    .A1(_1304_),
    .A2(_2553_));
 sg13g2_nor2_2 _6877_ (.A(_2571_),
    .B(_2573_),
    .Y(_2591_));
 sg13g2_a21o_1 _6878_ (.A2(_2566_),
    .A1(_2552_),
    .B1(_2568_),
    .X(_2592_));
 sg13g2_a21o_1 _6879_ (.A2(_2569_),
    .A1(_2550_),
    .B1(_2549_),
    .X(_2593_));
 sg13g2_a21oi_1 _6880_ (.A1(_2534_),
    .A2(_2547_),
    .Y(_2594_),
    .B1(_2533_));
 sg13g2_a22oi_1 _6881_ (.Y(_2595_),
    .B1(_2528_),
    .B2(_2531_),
    .A2(_2452_),
    .A1(_3135_));
 sg13g2_a21oi_1 _6882_ (.A1(net935),
    .A2(_2451_),
    .Y(_2596_),
    .B1(_3135_));
 sg13g2_nor2_1 _6883_ (.A(net932),
    .B(_3135_),
    .Y(_2597_));
 sg13g2_nand3_1 _6884_ (.B(net883),
    .C(_2597_),
    .A(net931),
    .Y(_2598_));
 sg13g2_a21o_1 _6885_ (.A2(net883),
    .A1(net930),
    .B1(_2597_),
    .X(_2599_));
 sg13g2_and2_1 _6886_ (.A(_2598_),
    .B(_2599_),
    .X(_2600_));
 sg13g2_nand2b_1 _6887_ (.Y(_2601_),
    .B(_2600_),
    .A_N(_2523_));
 sg13g2_xnor2_1 _6888_ (.Y(_2602_),
    .A(_2523_),
    .B(_2600_));
 sg13g2_xnor2_1 _6889_ (.Y(_2603_),
    .A(_2596_),
    .B(_2602_));
 sg13g2_nand2_1 _6890_ (.Y(_2604_),
    .A(net924),
    .B(net887));
 sg13g2_nor2_1 _6891_ (.A(_2522_),
    .B(_2604_),
    .Y(_2605_));
 sg13g2_a22oi_1 _6892_ (.Y(_2606_),
    .B1(net887),
    .B2(net927),
    .A2(net891),
    .A1(net924));
 sg13g2_nor3_1 _6893_ (.A(_2538_),
    .B(_2605_),
    .C(_2606_),
    .Y(_2607_));
 sg13g2_o21ai_1 _6894_ (.B1(_2538_),
    .Y(_2608_),
    .A1(_2605_),
    .A2(_2606_));
 sg13g2_nor2b_1 _6895_ (.A(_2607_),
    .B_N(_2608_),
    .Y(_2609_));
 sg13g2_nor2b_1 _6896_ (.A(_2603_),
    .B_N(_2609_),
    .Y(_2610_));
 sg13g2_xnor2_1 _6897_ (.Y(_2611_),
    .A(_2603_),
    .B(_2609_));
 sg13g2_nor2b_1 _6898_ (.A(_2595_),
    .B_N(_2611_),
    .Y(_2612_));
 sg13g2_xnor2_1 _6899_ (.Y(_2613_),
    .A(_2595_),
    .B(_2611_));
 sg13g2_o21ai_1 _6900_ (.B1(_2540_),
    .Y(_2614_),
    .A1(_2537_),
    .A2(_2541_));
 sg13g2_or2_1 _6901_ (.X(_2615_),
    .B(_2526_),
    .A(_2524_));
 sg13g2_nand2_1 _6902_ (.Y(_2616_),
    .A(net895),
    .B(net917));
 sg13g2_nor2_1 _6903_ (.A(_2537_),
    .B(_2616_),
    .Y(_2617_));
 sg13g2_a22oi_1 _6904_ (.Y(_2618_),
    .B1(net917),
    .B2(net898),
    .A2(net918),
    .A1(net895));
 sg13g2_nor3_1 _6905_ (.A(_2559_),
    .B(_2617_),
    .C(_2618_),
    .Y(_2619_));
 sg13g2_o21ai_1 _6906_ (.B1(_2559_),
    .Y(_2620_),
    .A1(_2617_),
    .A2(_2618_));
 sg13g2_nor2b_1 _6907_ (.A(_2619_),
    .B_N(_2620_),
    .Y(_2621_));
 sg13g2_xnor2_1 _6908_ (.Y(_2622_),
    .A(_2615_),
    .B(_2621_));
 sg13g2_nor2b_1 _6909_ (.A(_2622_),
    .B_N(_2614_),
    .Y(_2623_));
 sg13g2_xor2_1 _6910_ (.B(_2622_),
    .A(_2614_),
    .X(_2624_));
 sg13g2_inv_1 _6911_ (.Y(_2625_),
    .A(_2624_));
 sg13g2_xnor2_1 _6912_ (.Y(_2626_),
    .A(_2613_),
    .B(_2625_));
 sg13g2_nor2_1 _6913_ (.A(_2594_),
    .B(_2626_),
    .Y(_2627_));
 sg13g2_xor2_1 _6914_ (.B(_2626_),
    .A(_2594_),
    .X(_2628_));
 sg13g2_o21ai_1 _6915_ (.B1(_2564_),
    .Y(_2629_),
    .A1(_2556_),
    .A2(_2565_));
 sg13g2_a21o_1 _6916_ (.A2(_2545_),
    .A1(_2535_),
    .B1(_2544_),
    .X(_2630_));
 sg13g2_inv_1 _6917_ (.Y(_2631_),
    .A(_2630_));
 sg13g2_nand2_1 _6918_ (.Y(_2632_),
    .A(\i_mandel.i_xy.hc.genblk2[11].state.Q ),
    .B(\i_mandel.i_xy.hc.genblk2[11].state.D ));
 sg13g2_xnor2_1 _6919_ (.Y(_2633_),
    .A(\i_mandel.i_xy.hc.genblk2[11].state.Q ),
    .B(_1304_));
 sg13g2_inv_1 _6920_ (.Y(_2634_),
    .A(_2633_));
 sg13g2_o21ai_1 _6921_ (.B1(_2562_),
    .Y(_2635_),
    .A1(_2417_),
    .A2(_2559_));
 sg13g2_and4_1 _6922_ (.A(net904),
    .B(net905),
    .C(net912),
    .D(net910),
    .X(_2636_));
 sg13g2_a22oi_1 _6923_ (.Y(_2637_),
    .B1(net910),
    .B2(net905),
    .A2(net912),
    .A1(\i_mandel.i_xy.y[-7] ));
 sg13g2_nor3_1 _6924_ (.A(_2553_),
    .B(_2636_),
    .C(_2637_),
    .Y(_2638_));
 sg13g2_o21ai_1 _6925_ (.B1(_2553_),
    .Y(_2639_),
    .A1(_2636_),
    .A2(_2637_));
 sg13g2_nor2b_1 _6926_ (.A(_2638_),
    .B_N(_2639_),
    .Y(_2640_));
 sg13g2_xnor2_1 _6927_ (.Y(_2641_),
    .A(_2635_),
    .B(_2640_));
 sg13g2_nor2_1 _6928_ (.A(_2634_),
    .B(_2641_),
    .Y(_2642_));
 sg13g2_xor2_1 _6929_ (.B(_2641_),
    .A(_2633_),
    .X(_2643_));
 sg13g2_xnor2_1 _6930_ (.Y(_2644_),
    .A(_2631_),
    .B(_2643_));
 sg13g2_nand2b_1 _6931_ (.Y(_2645_),
    .B(_2629_),
    .A_N(_2644_));
 sg13g2_xor2_1 _6932_ (.B(_2644_),
    .A(_2629_),
    .X(_2646_));
 sg13g2_inv_1 _6933_ (.Y(_2647_),
    .A(_2646_));
 sg13g2_xnor2_1 _6934_ (.Y(_2648_),
    .A(_2628_),
    .B(_2646_));
 sg13g2_xnor2_1 _6935_ (.Y(_2649_),
    .A(_2593_),
    .B(_2648_));
 sg13g2_nor2b_1 _6936_ (.A(_2649_),
    .B_N(_2592_),
    .Y(_2650_));
 sg13g2_xor2_1 _6937_ (.B(_2649_),
    .A(_2592_),
    .X(_2651_));
 sg13g2_nor2_1 _6938_ (.A(_2591_),
    .B(_2651_),
    .Y(_2652_));
 sg13g2_xor2_1 _6939_ (.B(_2651_),
    .A(_2591_),
    .X(_2653_));
 sg13g2_xnor2_1 _6940_ (.Y(_2654_),
    .A(_2590_),
    .B(_2653_));
 sg13g2_nor2b_1 _6941_ (.A(_2654_),
    .B_N(_2589_),
    .Y(_2655_));
 sg13g2_nand2b_1 _6942_ (.Y(_2656_),
    .B(_2654_),
    .A_N(_2589_));
 sg13g2_xor2_1 _6943_ (.B(_2654_),
    .A(_2589_),
    .X(_2657_));
 sg13g2_xnor2_1 _6944_ (.Y(_2658_),
    .A(_2588_),
    .B(_2657_));
 sg13g2_nand2_1 _6945_ (.Y(_2659_),
    .A(\i_coord.y0[-5] ),
    .B(_2658_));
 sg13g2_xnor2_1 _6946_ (.Y(_2660_),
    .A(_3123_),
    .B(_2658_));
 sg13g2_nor3_1 _6947_ (.A(_2582_),
    .B(_2585_),
    .C(_2660_),
    .Y(_2661_));
 sg13g2_o21ai_1 _6948_ (.B1(_2660_),
    .Y(_2662_),
    .A1(_2582_),
    .A2(_2585_));
 sg13g2_nor2b_1 _6949_ (.A(_2661_),
    .B_N(_2662_),
    .Y(_2663_));
 sg13g2_mux2_1 _6950_ (.A0(_1838_),
    .A1(_2663_),
    .S(net834),
    .X(_2664_));
 sg13g2_mux2_1 _6951_ (.A0(_2664_),
    .A1(net338),
    .S(net736),
    .X(_0158_));
 sg13g2_a21o_1 _6952_ (.A2(_2656_),
    .A1(_2588_),
    .B1(_2655_),
    .X(_2665_));
 sg13g2_a21oi_2 _6953_ (.B1(_2652_),
    .Y(_2666_),
    .A2(_2653_),
    .A1(_2590_));
 sg13g2_a21o_1 _6954_ (.A2(_2648_),
    .A1(_2593_),
    .B1(_2650_),
    .X(_2667_));
 sg13g2_o21ai_1 _6955_ (.B1(_2645_),
    .Y(_2668_),
    .A1(_2631_),
    .A2(_2643_));
 sg13g2_a21oi_2 _6956_ (.B1(_2627_),
    .Y(_2669_),
    .A2(_2647_),
    .A1(_2628_));
 sg13g2_a21oi_2 _6957_ (.B1(_2612_),
    .Y(_2670_),
    .A2(_2625_),
    .A1(_2613_));
 sg13g2_a21o_1 _6958_ (.A2(_2602_),
    .A1(_2596_),
    .B1(_2610_),
    .X(_2671_));
 sg13g2_nand2_1 _6959_ (.Y(_2672_),
    .A(_2598_),
    .B(_2601_));
 sg13g2_nand2_1 _6960_ (.Y(_2673_),
    .A(net926),
    .B(net885));
 sg13g2_nor2_1 _6961_ (.A(net930),
    .B(net879),
    .Y(_2674_));
 sg13g2_nand3_1 _6962_ (.B(net883),
    .C(_2674_),
    .A(net929),
    .Y(_2675_));
 sg13g2_a21o_1 _6963_ (.A2(\i_mandel.i_xy.y[1] ),
    .A1(net929),
    .B1(_2674_),
    .X(_2676_));
 sg13g2_and2_1 _6964_ (.A(_2675_),
    .B(_2676_),
    .X(_2677_));
 sg13g2_nand2b_1 _6965_ (.Y(_2678_),
    .B(_2677_),
    .A_N(_2673_));
 sg13g2_xnor2_1 _6966_ (.Y(_2679_),
    .A(_2673_),
    .B(_2677_));
 sg13g2_xnor2_1 _6967_ (.Y(_2680_),
    .A(_2672_),
    .B(_2679_));
 sg13g2_nand2_1 _6968_ (.Y(_2681_),
    .A(net893),
    .B(net918));
 sg13g2_nand2_1 _6969_ (.Y(_2682_),
    .A(net921),
    .B(net888));
 sg13g2_nand2_1 _6970_ (.Y(_2683_),
    .A(net921),
    .B(net890));
 sg13g2_xor2_1 _6971_ (.B(_2683_),
    .A(_2604_),
    .X(_2684_));
 sg13g2_nand2b_1 _6972_ (.Y(_2685_),
    .B(_2684_),
    .A_N(_2681_));
 sg13g2_xnor2_1 _6973_ (.Y(_2686_),
    .A(_2681_),
    .B(_2684_));
 sg13g2_nor2b_1 _6974_ (.A(_2680_),
    .B_N(_2686_),
    .Y(_2687_));
 sg13g2_xnor2_1 _6975_ (.Y(_2688_),
    .A(_2680_),
    .B(_2686_));
 sg13g2_nand2_1 _6976_ (.Y(_2689_),
    .A(_2671_),
    .B(_2688_));
 sg13g2_xnor2_1 _6977_ (.Y(_2690_),
    .A(_2671_),
    .B(_2688_));
 sg13g2_or2_1 _6978_ (.X(_2691_),
    .B(_2619_),
    .A(_2617_));
 sg13g2_or2_1 _6979_ (.X(_2692_),
    .B(_2607_),
    .A(_2605_));
 sg13g2_nand2_1 _6980_ (.Y(_2693_),
    .A(net897),
    .B(net915));
 sg13g2_xor2_1 _6981_ (.B(_2693_),
    .A(_2616_),
    .X(_2694_));
 sg13g2_nand3_1 _6982_ (.B(net912),
    .C(_2694_),
    .A(net900),
    .Y(_2695_));
 sg13g2_a21o_1 _6983_ (.A2(net911),
    .A1(net900),
    .B1(_2694_),
    .X(_2696_));
 sg13g2_and2_1 _6984_ (.A(_2695_),
    .B(_2696_),
    .X(_2697_));
 sg13g2_xnor2_1 _6985_ (.Y(_2698_),
    .A(_2692_),
    .B(_2697_));
 sg13g2_nor2b_1 _6986_ (.A(_2698_),
    .B_N(_2691_),
    .Y(_2699_));
 sg13g2_xor2_1 _6987_ (.B(_2698_),
    .A(_2691_),
    .X(_2700_));
 sg13g2_xor2_1 _6988_ (.B(_2700_),
    .A(_2690_),
    .X(_2701_));
 sg13g2_nor2b_1 _6989_ (.A(_2670_),
    .B_N(_2701_),
    .Y(_2702_));
 sg13g2_xnor2_1 _6990_ (.Y(_2703_),
    .A(_2670_),
    .B(_2701_));
 sg13g2_a21oi_1 _6991_ (.A1(_2635_),
    .A2(_2640_),
    .Y(_2704_),
    .B1(_2642_));
 sg13g2_a21o_1 _6992_ (.A2(_2621_),
    .A1(_2615_),
    .B1(_2623_),
    .X(_2705_));
 sg13g2_or2_1 _6993_ (.X(_2706_),
    .B(_2638_),
    .A(_2636_));
 sg13g2_o21ai_1 _6994_ (.B1(net909),
    .Y(_2707_),
    .A1(net903),
    .A2(net905));
 sg13g2_nand3_1 _6995_ (.B(net905),
    .C(net909),
    .A(net903),
    .Y(_2708_));
 sg13g2_nand2b_1 _6996_ (.Y(_2709_),
    .B(_2708_),
    .A_N(_2707_));
 sg13g2_xnor2_1 _6997_ (.Y(_2710_),
    .A(_2553_),
    .B(_2709_));
 sg13g2_nor2b_1 _6998_ (.A(_2710_),
    .B_N(_2706_),
    .Y(_2711_));
 sg13g2_nand2b_1 _6999_ (.Y(_2712_),
    .B(_2706_),
    .A_N(_2710_));
 sg13g2_xnor2_1 _7000_ (.Y(_2713_),
    .A(_2706_),
    .B(_2710_));
 sg13g2_xor2_1 _7001_ (.B(_2713_),
    .A(_2633_),
    .X(_2714_));
 sg13g2_nand2_1 _7002_ (.Y(_2715_),
    .A(_2705_),
    .B(_2714_));
 sg13g2_xnor2_1 _7003_ (.Y(_2716_),
    .A(_2705_),
    .B(_2714_));
 sg13g2_xor2_1 _7004_ (.B(_2716_),
    .A(_2704_),
    .X(_2717_));
 sg13g2_xnor2_1 _7005_ (.Y(_2718_),
    .A(_2703_),
    .B(_2717_));
 sg13g2_nor2_1 _7006_ (.A(_2669_),
    .B(_2718_),
    .Y(_2719_));
 sg13g2_xor2_1 _7007_ (.B(_2718_),
    .A(_2669_),
    .X(_2720_));
 sg13g2_xor2_1 _7008_ (.B(_2720_),
    .A(_2668_),
    .X(_2721_));
 sg13g2_nand2_1 _7009_ (.Y(_2722_),
    .A(_2667_),
    .B(_2721_));
 sg13g2_xnor2_1 _7010_ (.Y(_2723_),
    .A(_2667_),
    .B(_2721_));
 sg13g2_xor2_1 _7011_ (.B(_2723_),
    .A(net743),
    .X(_2724_));
 sg13g2_nor2b_1 _7012_ (.A(_2666_),
    .B_N(_2724_),
    .Y(_2725_));
 sg13g2_xnor2_1 _7013_ (.Y(_2726_),
    .A(_2666_),
    .B(_2724_));
 sg13g2_xor2_1 _7014_ (.B(_2726_),
    .A(_2665_),
    .X(_2727_));
 sg13g2_and2_1 _7015_ (.A(\i_coord.y0[-4] ),
    .B(_2727_),
    .X(_2728_));
 sg13g2_xnor2_1 _7016_ (.Y(_2729_),
    .A(\i_coord.y0[-4] ),
    .B(_2727_));
 sg13g2_and3_1 _7017_ (.X(_2730_),
    .A(_2659_),
    .B(_2662_),
    .C(_2729_));
 sg13g2_a21oi_2 _7018_ (.B1(_2729_),
    .Y(_2731_),
    .A2(_2662_),
    .A1(_2659_));
 sg13g2_o21ai_1 _7019_ (.B1(net834),
    .Y(_2732_),
    .A1(_2730_),
    .A2(_2731_));
 sg13g2_o21ai_1 _7020_ (.B1(_2732_),
    .Y(_2733_),
    .A1(net834),
    .A2(_1848_));
 sg13g2_nand2_1 _7021_ (.Y(_2734_),
    .A(net896),
    .B(net735));
 sg13g2_o21ai_1 _7022_ (.B1(_2734_),
    .Y(_0159_),
    .A1(net735),
    .A2(_2733_));
 sg13g2_nor2_1 _7023_ (.A(net834),
    .B(_1859_),
    .Y(_2735_));
 sg13g2_a21oi_1 _7024_ (.A1(_2665_),
    .A2(_2726_),
    .Y(_2736_),
    .B1(_2725_));
 sg13g2_o21ai_1 _7025_ (.B1(_2722_),
    .Y(_2737_),
    .A1(net743),
    .A2(_2723_));
 sg13g2_a21oi_2 _7026_ (.B1(_2719_),
    .Y(_2738_),
    .A2(_2720_),
    .A1(_2668_));
 sg13g2_o21ai_1 _7027_ (.B1(_2715_),
    .Y(_2739_),
    .A1(_2704_),
    .A2(_2716_));
 sg13g2_a21o_1 _7028_ (.A2(_2717_),
    .A1(_2703_),
    .B1(_2702_),
    .X(_2740_));
 sg13g2_o21ai_1 _7029_ (.B1(_2689_),
    .Y(_2741_),
    .A1(_2690_),
    .A2(_2700_));
 sg13g2_a21oi_2 _7030_ (.B1(_2687_),
    .Y(_2742_),
    .A2(_2679_),
    .A1(_2672_));
 sg13g2_nand2_1 _7031_ (.Y(_2743_),
    .A(_2675_),
    .B(_2678_));
 sg13g2_nand2_1 _7032_ (.Y(_2744_),
    .A(net923),
    .B(net885));
 sg13g2_nor2_1 _7033_ (.A(net928),
    .B(net879),
    .Y(_2745_));
 sg13g2_nand3_1 _7034_ (.B(net883),
    .C(_2745_),
    .A(net926),
    .Y(_2746_));
 sg13g2_a21o_1 _7035_ (.A2(net883),
    .A1(net926),
    .B1(_2745_),
    .X(_2747_));
 sg13g2_and2_1 _7036_ (.A(_2746_),
    .B(_2747_),
    .X(_2748_));
 sg13g2_nand2b_1 _7037_ (.Y(_2749_),
    .B(_2748_),
    .A_N(_2744_));
 sg13g2_xnor2_1 _7038_ (.Y(_2750_),
    .A(_2744_),
    .B(_2748_));
 sg13g2_xnor2_1 _7039_ (.Y(_2751_),
    .A(_2743_),
    .B(_2750_));
 sg13g2_nand2_1 _7040_ (.Y(_2752_),
    .A(net893),
    .B(net917));
 sg13g2_nand2_1 _7041_ (.Y(_2753_),
    .A(net919),
    .B(net887));
 sg13g2_nand2_1 _7042_ (.Y(_2754_),
    .A(net891),
    .B(net918));
 sg13g2_xor2_1 _7043_ (.B(_2754_),
    .A(_2682_),
    .X(_2755_));
 sg13g2_nand2b_1 _7044_ (.Y(_2756_),
    .B(_2755_),
    .A_N(_2752_));
 sg13g2_xnor2_1 _7045_ (.Y(_2757_),
    .A(_2752_),
    .B(_2755_));
 sg13g2_nor2b_1 _7046_ (.A(_2751_),
    .B_N(_2757_),
    .Y(_2758_));
 sg13g2_xnor2_1 _7047_ (.Y(_2759_),
    .A(_2751_),
    .B(_2757_));
 sg13g2_nand2b_1 _7048_ (.Y(_2760_),
    .B(_2759_),
    .A_N(_2742_));
 sg13g2_xnor2_1 _7049_ (.Y(_2761_),
    .A(_2742_),
    .B(_2759_));
 sg13g2_inv_1 _7050_ (.Y(_2762_),
    .A(_2761_));
 sg13g2_o21ai_1 _7051_ (.B1(_2695_),
    .Y(_2763_),
    .A1(_2616_),
    .A2(_2693_));
 sg13g2_o21ai_1 _7052_ (.B1(_2685_),
    .Y(_2764_),
    .A1(_2604_),
    .A2(_2683_));
 sg13g2_nand2_2 _7053_ (.Y(_2765_),
    .A(net901),
    .B(net909));
 sg13g2_inv_1 _7054_ (.Y(_2766_),
    .A(_2765_));
 sg13g2_nor3_1 _7055_ (.A(_3131_),
    .B(_3133_),
    .C(_2693_),
    .Y(_2767_));
 sg13g2_a22oi_1 _7056_ (.Y(_2768_),
    .B1(net911),
    .B2(net897),
    .A2(net914),
    .A1(net895));
 sg13g2_nor2_1 _7057_ (.A(_2767_),
    .B(_2768_),
    .Y(_2769_));
 sg13g2_xnor2_1 _7058_ (.Y(_2770_),
    .A(_2765_),
    .B(_2769_));
 sg13g2_xnor2_1 _7059_ (.Y(_2771_),
    .A(_2764_),
    .B(_2770_));
 sg13g2_nor2b_1 _7060_ (.A(_2771_),
    .B_N(_2763_),
    .Y(_2772_));
 sg13g2_xor2_1 _7061_ (.B(_2771_),
    .A(_2763_),
    .X(_2773_));
 sg13g2_xor2_1 _7062_ (.B(_2773_),
    .A(_2761_),
    .X(_2774_));
 sg13g2_nand2b_1 _7063_ (.Y(_2775_),
    .B(_2741_),
    .A_N(_2774_));
 sg13g2_xor2_1 _7064_ (.B(_2774_),
    .A(_2741_),
    .X(_2776_));
 sg13g2_a21oi_1 _7065_ (.A1(_2633_),
    .A2(_2713_),
    .Y(_2777_),
    .B1(_2711_));
 sg13g2_nand2_1 _7066_ (.Y(_2778_),
    .A(_2553_),
    .B(_2707_));
 sg13g2_nand2_1 _7067_ (.Y(_2779_),
    .A(_2712_),
    .B(_2778_));
 sg13g2_xnor2_1 _7068_ (.Y(_2780_),
    .A(_2633_),
    .B(_2779_));
 sg13g2_a21o_1 _7069_ (.A2(_2697_),
    .A1(_2692_),
    .B1(_2699_),
    .X(_2781_));
 sg13g2_xor2_1 _7070_ (.B(_2781_),
    .A(net741),
    .X(_2782_));
 sg13g2_nor2b_1 _7071_ (.A(_2777_),
    .B_N(_2782_),
    .Y(_2783_));
 sg13g2_xnor2_1 _7072_ (.Y(_2784_),
    .A(_2777_),
    .B(_2782_));
 sg13g2_inv_1 _7073_ (.Y(_2785_),
    .A(_2784_));
 sg13g2_xnor2_1 _7074_ (.Y(_2786_),
    .A(_2776_),
    .B(_2784_));
 sg13g2_and2_1 _7075_ (.A(_2740_),
    .B(_2786_),
    .X(_2787_));
 sg13g2_xor2_1 _7076_ (.B(_2786_),
    .A(_2740_),
    .X(_2788_));
 sg13g2_xnor2_1 _7077_ (.Y(_2789_),
    .A(_2739_),
    .B(_2788_));
 sg13g2_xor2_1 _7078_ (.B(_2789_),
    .A(_2738_),
    .X(_2790_));
 sg13g2_nand2b_1 _7079_ (.Y(_2791_),
    .B(_2790_),
    .A_N(net743));
 sg13g2_xnor2_1 _7080_ (.Y(_2792_),
    .A(net743),
    .B(_2790_));
 sg13g2_nand2_1 _7081_ (.Y(_2793_),
    .A(_2737_),
    .B(_2792_));
 sg13g2_xnor2_1 _7082_ (.Y(_2794_),
    .A(_2737_),
    .B(_2792_));
 sg13g2_xor2_1 _7083_ (.B(_2794_),
    .A(_2736_),
    .X(_2795_));
 sg13g2_xor2_1 _7084_ (.B(_2795_),
    .A(\i_coord.y0[-3] ),
    .X(_2796_));
 sg13g2_nor3_1 _7085_ (.A(_2728_),
    .B(_2731_),
    .C(_2796_),
    .Y(_2797_));
 sg13g2_o21ai_1 _7086_ (.B1(_2796_),
    .Y(_2798_),
    .A1(_2728_),
    .A2(_2731_));
 sg13g2_nand2b_1 _7087_ (.Y(_2799_),
    .B(_2798_),
    .A_N(_2797_));
 sg13g2_a21oi_2 _7088_ (.B1(_2735_),
    .Y(_2800_),
    .A2(_2799_),
    .A1(net835));
 sg13g2_mux2_1 _7089_ (.A0(_2800_),
    .A1(net893),
    .S(net735),
    .X(_0160_));
 sg13g2_nand2b_1 _7090_ (.Y(_2801_),
    .B(_2795_),
    .A_N(_0023_));
 sg13g2_o21ai_1 _7091_ (.B1(_2793_),
    .Y(_2802_),
    .A1(_2736_),
    .A2(_2794_));
 sg13g2_o21ai_1 _7092_ (.B1(_2791_),
    .Y(_2803_),
    .A1(_2738_),
    .A2(_2789_));
 sg13g2_a21oi_1 _7093_ (.A1(_2739_),
    .A2(_2788_),
    .Y(_2804_),
    .B1(_2787_));
 sg13g2_a21o_1 _7094_ (.A2(_2781_),
    .A1(net741),
    .B1(_2783_),
    .X(_2805_));
 sg13g2_o21ai_1 _7095_ (.B1(_2775_),
    .Y(_2806_),
    .A1(_2776_),
    .A2(_2785_));
 sg13g2_o21ai_1 _7096_ (.B1(_2760_),
    .Y(_2807_),
    .A1(_2762_),
    .A2(_2773_));
 sg13g2_a21o_1 _7097_ (.A2(_2750_),
    .A1(_2743_),
    .B1(_2758_),
    .X(_2808_));
 sg13g2_nand2_1 _7098_ (.Y(_2809_),
    .A(_2746_),
    .B(_2749_));
 sg13g2_nand2_1 _7099_ (.Y(_2810_),
    .A(net920),
    .B(net885));
 sg13g2_nor2_1 _7100_ (.A(net927),
    .B(net879),
    .Y(_2811_));
 sg13g2_nand3_1 _7101_ (.B(net883),
    .C(_2811_),
    .A(net923),
    .Y(_2812_));
 sg13g2_a21o_1 _7102_ (.A2(net883),
    .A1(net923),
    .B1(_2811_),
    .X(_2813_));
 sg13g2_and2_1 _7103_ (.A(_2812_),
    .B(_2813_),
    .X(_2814_));
 sg13g2_nand2b_1 _7104_ (.Y(_2815_),
    .B(_2814_),
    .A_N(_2810_));
 sg13g2_xnor2_1 _7105_ (.Y(_2816_),
    .A(_2810_),
    .B(_2814_));
 sg13g2_xnor2_1 _7106_ (.Y(_2817_),
    .A(_2809_),
    .B(_2816_));
 sg13g2_nand2_1 _7107_ (.Y(_2818_),
    .A(net890),
    .B(net916));
 sg13g2_xor2_1 _7108_ (.B(_2818_),
    .A(_2753_),
    .X(_2819_));
 sg13g2_nand3_1 _7109_ (.B(net914),
    .C(_2819_),
    .A(net893),
    .Y(_2820_));
 sg13g2_a21o_1 _7110_ (.A2(net914),
    .A1(net892),
    .B1(_2819_),
    .X(_2821_));
 sg13g2_and2_1 _7111_ (.A(_2820_),
    .B(_2821_),
    .X(_2822_));
 sg13g2_nor2b_1 _7112_ (.A(_2817_),
    .B_N(_2822_),
    .Y(_2823_));
 sg13g2_xnor2_1 _7113_ (.Y(_2824_),
    .A(_2817_),
    .B(_2822_));
 sg13g2_nand2_1 _7114_ (.Y(_2825_),
    .A(_2808_),
    .B(_2824_));
 sg13g2_nor2_1 _7115_ (.A(_2808_),
    .B(_2824_),
    .Y(_2826_));
 sg13g2_xor2_1 _7116_ (.B(_2824_),
    .A(_2808_),
    .X(_2827_));
 sg13g2_a21o_1 _7117_ (.A2(_2769_),
    .A1(_2766_),
    .B1(_2767_),
    .X(_2828_));
 sg13g2_o21ai_1 _7118_ (.B1(_2756_),
    .Y(_2829_),
    .A1(_2682_),
    .A2(_2754_));
 sg13g2_a22oi_1 _7119_ (.Y(_2830_),
    .B1(net909),
    .B2(net898),
    .A2(net911),
    .A1(net895));
 sg13g2_and3_1 _7120_ (.X(_2831_),
    .A(net898),
    .B(net894),
    .C(net909));
 sg13g2_a21oi_1 _7121_ (.A1(net911),
    .A2(_2831_),
    .Y(_2832_),
    .B1(_2830_));
 sg13g2_xnor2_1 _7122_ (.Y(_2833_),
    .A(_2765_),
    .B(_2832_));
 sg13g2_xnor2_1 _7123_ (.Y(_2834_),
    .A(_2829_),
    .B(_2833_));
 sg13g2_nor2b_1 _7124_ (.A(_2834_),
    .B_N(_2828_),
    .Y(_2835_));
 sg13g2_xor2_1 _7125_ (.B(_2834_),
    .A(_2828_),
    .X(_2836_));
 sg13g2_xnor2_1 _7126_ (.Y(_2837_),
    .A(_2827_),
    .B(_2836_));
 sg13g2_nand2_1 _7127_ (.Y(_2838_),
    .A(_2807_),
    .B(_2837_));
 sg13g2_xnor2_1 _7128_ (.Y(_2839_),
    .A(_2807_),
    .B(_2837_));
 sg13g2_a21oi_2 _7129_ (.B1(_2711_),
    .Y(_2840_),
    .A2(_2778_),
    .A1(_2633_));
 sg13g2_a21o_1 _7130_ (.A2(_2770_),
    .A1(_2764_),
    .B1(_2772_),
    .X(_2841_));
 sg13g2_nand2_1 _7131_ (.Y(_2842_),
    .A(_2780_),
    .B(_2841_));
 sg13g2_xor2_1 _7132_ (.B(_2841_),
    .A(_2780_),
    .X(_2843_));
 sg13g2_inv_1 _7133_ (.Y(_2844_),
    .A(_2843_));
 sg13g2_xnor2_1 _7134_ (.Y(_2845_),
    .A(_2840_),
    .B(_2843_));
 sg13g2_inv_1 _7135_ (.Y(_2846_),
    .A(_2845_));
 sg13g2_xnor2_1 _7136_ (.Y(_2847_),
    .A(_2839_),
    .B(_2845_));
 sg13g2_and2_1 _7137_ (.A(_2806_),
    .B(_2847_),
    .X(_2848_));
 sg13g2_xor2_1 _7138_ (.B(_2847_),
    .A(_2806_),
    .X(_2849_));
 sg13g2_xnor2_1 _7139_ (.Y(_2850_),
    .A(_2805_),
    .B(_2849_));
 sg13g2_xor2_1 _7140_ (.B(_2850_),
    .A(_2804_),
    .X(_2851_));
 sg13g2_nand2b_1 _7141_ (.Y(_2852_),
    .B(_2851_),
    .A_N(net743));
 sg13g2_xnor2_1 _7142_ (.Y(_2853_),
    .A(net742),
    .B(_2851_));
 sg13g2_and2_1 _7143_ (.A(_2803_),
    .B(_2853_),
    .X(_2854_));
 sg13g2_xor2_1 _7144_ (.B(_2853_),
    .A(_2803_),
    .X(_2855_));
 sg13g2_xnor2_1 _7145_ (.Y(_2856_),
    .A(_2802_),
    .B(_2855_));
 sg13g2_xor2_1 _7146_ (.B(_2856_),
    .A(\i_coord.y0[-2] ),
    .X(_2857_));
 sg13g2_a21o_1 _7147_ (.A2(_2801_),
    .A1(_2798_),
    .B1(_2857_),
    .X(_2858_));
 sg13g2_nand3_1 _7148_ (.B(_2801_),
    .C(_2857_),
    .A(_2798_),
    .Y(_2859_));
 sg13g2_a21oi_1 _7149_ (.A1(_2858_),
    .A2(_2859_),
    .Y(_2860_),
    .B1(net840));
 sg13g2_nor2_1 _7150_ (.A(net835),
    .B(_1872_),
    .Y(_2861_));
 sg13g2_nor2_1 _7151_ (.A(_2860_),
    .B(_2861_),
    .Y(_2862_));
 sg13g2_mux2_1 _7152_ (.A0(_2862_),
    .A1(net890),
    .S(net736),
    .X(_0161_));
 sg13g2_nor2_1 _7153_ (.A(_0022_),
    .B(_2856_),
    .Y(_2863_));
 sg13g2_inv_1 _7154_ (.Y(_2864_),
    .A(_2863_));
 sg13g2_nand2_1 _7155_ (.Y(_2865_),
    .A(_2858_),
    .B(_2864_));
 sg13g2_a21o_1 _7156_ (.A2(_2855_),
    .A1(_2802_),
    .B1(_2854_),
    .X(_2866_));
 sg13g2_o21ai_1 _7157_ (.B1(_2852_),
    .Y(_2867_),
    .A1(_2804_),
    .A2(_2850_));
 sg13g2_a21oi_1 _7158_ (.A1(_2805_),
    .A2(_2849_),
    .Y(_2868_),
    .B1(_2848_));
 sg13g2_o21ai_1 _7159_ (.B1(_2842_),
    .Y(_2869_),
    .A1(_2840_),
    .A2(_2844_));
 sg13g2_o21ai_1 _7160_ (.B1(_2838_),
    .Y(_2870_),
    .A1(_2839_),
    .A2(_2846_));
 sg13g2_o21ai_1 _7161_ (.B1(_2825_),
    .Y(_2871_),
    .A1(_2826_),
    .A2(_2836_));
 sg13g2_a21o_1 _7162_ (.A2(_2816_),
    .A1(_2809_),
    .B1(_2823_),
    .X(_2872_));
 sg13g2_nand2_1 _7163_ (.Y(_2873_),
    .A(_2812_),
    .B(_2815_));
 sg13g2_nand2_1 _7164_ (.Y(_2874_),
    .A(net919),
    .B(net885));
 sg13g2_nor2_1 _7165_ (.A(net923),
    .B(net879),
    .Y(_2875_));
 sg13g2_nand3_1 _7166_ (.B(net884),
    .C(_2875_),
    .A(net920),
    .Y(_2876_));
 sg13g2_a21o_1 _7167_ (.A2(net884),
    .A1(net920),
    .B1(_2875_),
    .X(_2877_));
 sg13g2_and2_1 _7168_ (.A(_2876_),
    .B(_2877_),
    .X(_2878_));
 sg13g2_nand2b_1 _7169_ (.Y(_2879_),
    .B(_2878_),
    .A_N(_2874_));
 sg13g2_xnor2_1 _7170_ (.Y(_2880_),
    .A(_2874_),
    .B(_2878_));
 sg13g2_xnor2_1 _7171_ (.Y(_2881_),
    .A(_2873_),
    .B(_2880_));
 sg13g2_nand2_1 _7172_ (.Y(_2882_),
    .A(net893),
    .B(net911));
 sg13g2_nand2_1 _7173_ (.Y(_2883_),
    .A(net888),
    .B(net915));
 sg13g2_nor2_1 _7174_ (.A(_2818_),
    .B(_2883_),
    .Y(_2884_));
 sg13g2_a22oi_1 _7175_ (.Y(_2885_),
    .B1(net914),
    .B2(net890),
    .A2(net916),
    .A1(net887));
 sg13g2_nor3_1 _7176_ (.A(_2882_),
    .B(_2884_),
    .C(_2885_),
    .Y(_2886_));
 sg13g2_o21ai_1 _7177_ (.B1(_2882_),
    .Y(_2887_),
    .A1(_2884_),
    .A2(_2885_));
 sg13g2_nor2b_1 _7178_ (.A(_2886_),
    .B_N(_2887_),
    .Y(_2888_));
 sg13g2_nor2b_1 _7179_ (.A(_2881_),
    .B_N(_2888_),
    .Y(_2889_));
 sg13g2_xnor2_1 _7180_ (.Y(_2890_),
    .A(_2881_),
    .B(_2888_));
 sg13g2_nand2_1 _7181_ (.Y(_2891_),
    .A(_2872_),
    .B(_2890_));
 sg13g2_nor2_1 _7182_ (.A(_2872_),
    .B(_2890_),
    .Y(_2892_));
 sg13g2_xor2_1 _7183_ (.B(_2890_),
    .A(_2872_),
    .X(_2893_));
 sg13g2_a22oi_1 _7184_ (.Y(_2894_),
    .B1(_2832_),
    .B2(_2766_),
    .A2(_2831_),
    .A1(net911));
 sg13g2_o21ai_1 _7185_ (.B1(_2820_),
    .Y(_2895_),
    .A1(_2753_),
    .A2(_2818_));
 sg13g2_o21ai_1 _7186_ (.B1(net909),
    .Y(_2896_),
    .A1(net898),
    .A2(net894));
 sg13g2_nor2_1 _7187_ (.A(_2831_),
    .B(_2896_),
    .Y(_2897_));
 sg13g2_xnor2_1 _7188_ (.Y(_2898_),
    .A(_2765_),
    .B(_2897_));
 sg13g2_nand2_1 _7189_ (.Y(_2899_),
    .A(_2895_),
    .B(_2898_));
 sg13g2_xnor2_1 _7190_ (.Y(_2900_),
    .A(_2895_),
    .B(_2898_));
 sg13g2_xnor2_1 _7191_ (.Y(_2901_),
    .A(_2894_),
    .B(_2900_));
 sg13g2_xnor2_1 _7192_ (.Y(_2902_),
    .A(_2893_),
    .B(_2901_));
 sg13g2_nand2_1 _7193_ (.Y(_2903_),
    .A(_2871_),
    .B(_2902_));
 sg13g2_xnor2_1 _7194_ (.Y(_2904_),
    .A(_2871_),
    .B(_2902_));
 sg13g2_a21o_1 _7195_ (.A2(_2833_),
    .A1(_2829_),
    .B1(_2835_),
    .X(_2905_));
 sg13g2_nand2_1 _7196_ (.Y(_2906_),
    .A(net741),
    .B(_2905_));
 sg13g2_xor2_1 _7197_ (.B(_2905_),
    .A(net741),
    .X(_2907_));
 sg13g2_inv_1 _7198_ (.Y(_2908_),
    .A(_2907_));
 sg13g2_xnor2_1 _7199_ (.Y(_2909_),
    .A(_2840_),
    .B(_2907_));
 sg13g2_inv_1 _7200_ (.Y(_2910_),
    .A(_2909_));
 sg13g2_xnor2_1 _7201_ (.Y(_2911_),
    .A(_2904_),
    .B(_2909_));
 sg13g2_and2_1 _7202_ (.A(_2870_),
    .B(_2911_),
    .X(_2912_));
 sg13g2_xor2_1 _7203_ (.B(_2911_),
    .A(_2870_),
    .X(_2913_));
 sg13g2_xnor2_1 _7204_ (.Y(_2914_),
    .A(_2869_),
    .B(_2913_));
 sg13g2_xor2_1 _7205_ (.B(_2914_),
    .A(_2868_),
    .X(_2915_));
 sg13g2_nand2b_1 _7206_ (.Y(_2916_),
    .B(_2915_),
    .A_N(net742));
 sg13g2_xnor2_1 _7207_ (.Y(_2917_),
    .A(net742),
    .B(_2915_));
 sg13g2_and2_1 _7208_ (.A(_2867_),
    .B(_2917_),
    .X(_2918_));
 sg13g2_xnor2_1 _7209_ (.Y(_2919_),
    .A(_2867_),
    .B(_2917_));
 sg13g2_inv_1 _7210_ (.Y(_2920_),
    .A(_2919_));
 sg13g2_xnor2_1 _7211_ (.Y(_2921_),
    .A(_2866_),
    .B(_2920_));
 sg13g2_xnor2_1 _7212_ (.Y(_2922_),
    .A(_3125_),
    .B(_2921_));
 sg13g2_a21oi_1 _7213_ (.A1(_2858_),
    .A2(_2864_),
    .Y(_2923_),
    .B1(_2922_));
 sg13g2_xnor2_1 _7214_ (.Y(_2924_),
    .A(_2865_),
    .B(_2922_));
 sg13g2_mux2_1 _7215_ (.A0(_1883_),
    .A1(_2924_),
    .S(net834),
    .X(_2925_));
 sg13g2_mux2_1 _7216_ (.A0(_2925_),
    .A1(net888),
    .S(net735),
    .X(_0162_));
 sg13g2_nor2_1 _7217_ (.A(_0021_),
    .B(_2921_),
    .Y(_2926_));
 sg13g2_nor2_1 _7218_ (.A(_2923_),
    .B(_2926_),
    .Y(_2927_));
 sg13g2_a21oi_1 _7219_ (.A1(_2866_),
    .A2(_2920_),
    .Y(_2928_),
    .B1(_2918_));
 sg13g2_o21ai_1 _7220_ (.B1(_2916_),
    .Y(_2929_),
    .A1(_2868_),
    .A2(_2914_));
 sg13g2_a21oi_1 _7221_ (.A1(_2869_),
    .A2(_2913_),
    .Y(_2930_),
    .B1(_2912_));
 sg13g2_o21ai_1 _7222_ (.B1(_2906_),
    .Y(_2931_),
    .A1(_2840_),
    .A2(_2908_));
 sg13g2_o21ai_1 _7223_ (.B1(_2903_),
    .Y(_2932_),
    .A1(_2904_),
    .A2(_2910_));
 sg13g2_o21ai_1 _7224_ (.B1(_2891_),
    .Y(_2933_),
    .A1(_2892_),
    .A2(_2901_));
 sg13g2_a21o_1 _7225_ (.A2(_2880_),
    .A1(_2873_),
    .B1(_2889_),
    .X(_2934_));
 sg13g2_nand2_1 _7226_ (.Y(_2935_),
    .A(_2876_),
    .B(_2879_));
 sg13g2_nand2_1 _7227_ (.Y(_2936_),
    .A(net916),
    .B(net886));
 sg13g2_nor2_1 _7228_ (.A(net922),
    .B(net879),
    .Y(_2937_));
 sg13g2_nand3_1 _7229_ (.B(net884),
    .C(_2937_),
    .A(net919),
    .Y(_2938_));
 sg13g2_a21o_1 _7230_ (.A2(net884),
    .A1(net919),
    .B1(_2937_),
    .X(_2939_));
 sg13g2_and2_1 _7231_ (.A(_2938_),
    .B(_2939_),
    .X(_2940_));
 sg13g2_nand2b_1 _7232_ (.Y(_2941_),
    .B(_2940_),
    .A_N(_2936_));
 sg13g2_xnor2_1 _7233_ (.Y(_2942_),
    .A(_2936_),
    .B(_2940_));
 sg13g2_nand2_1 _7234_ (.Y(_2943_),
    .A(_2935_),
    .B(_2942_));
 sg13g2_xnor2_1 _7235_ (.Y(_2944_),
    .A(_2935_),
    .B(_2942_));
 sg13g2_nand2_2 _7236_ (.Y(_2945_),
    .A(net893),
    .B(net910));
 sg13g2_nand2_1 _7237_ (.Y(_2946_),
    .A(net890),
    .B(net913));
 sg13g2_or2_1 _7238_ (.X(_2947_),
    .B(_2946_),
    .A(_2883_));
 sg13g2_xnor2_1 _7239_ (.Y(_2948_),
    .A(_2883_),
    .B(_2946_));
 sg13g2_xor2_1 _7240_ (.B(_2948_),
    .A(_2945_),
    .X(_2949_));
 sg13g2_inv_1 _7241_ (.Y(_2950_),
    .A(_2949_));
 sg13g2_xnor2_1 _7242_ (.Y(_2951_),
    .A(_2944_),
    .B(_2949_));
 sg13g2_nand2_1 _7243_ (.Y(_2952_),
    .A(_2934_),
    .B(_2951_));
 sg13g2_xor2_1 _7244_ (.B(_2951_),
    .A(_2934_),
    .X(_2953_));
 sg13g2_inv_1 _7245_ (.Y(_2954_),
    .A(_2953_));
 sg13g2_a21o_2 _7246_ (.A2(_2897_),
    .A1(_2766_),
    .B1(_2831_),
    .X(_2955_));
 sg13g2_or2_1 _7247_ (.X(_2956_),
    .B(_2886_),
    .A(_2884_));
 sg13g2_and2_1 _7248_ (.A(_2898_),
    .B(_2956_),
    .X(_2957_));
 sg13g2_xor2_1 _7249_ (.B(_2956_),
    .A(_2898_),
    .X(_2958_));
 sg13g2_xnor2_1 _7250_ (.Y(_2959_),
    .A(_2955_),
    .B(_2958_));
 sg13g2_xnor2_1 _7251_ (.Y(_2960_),
    .A(_2953_),
    .B(_2959_));
 sg13g2_nand2_1 _7252_ (.Y(_2961_),
    .A(_2933_),
    .B(_2960_));
 sg13g2_xnor2_1 _7253_ (.Y(_2962_),
    .A(_2933_),
    .B(_2960_));
 sg13g2_o21ai_1 _7254_ (.B1(_2899_),
    .Y(_2963_),
    .A1(_2894_),
    .A2(_2900_));
 sg13g2_nand2_1 _7255_ (.Y(_2964_),
    .A(net741),
    .B(_2963_));
 sg13g2_xor2_1 _7256_ (.B(_2963_),
    .A(net741),
    .X(_2965_));
 sg13g2_inv_1 _7257_ (.Y(_2966_),
    .A(_2965_));
 sg13g2_xnor2_1 _7258_ (.Y(_2967_),
    .A(_2840_),
    .B(_2965_));
 sg13g2_inv_1 _7259_ (.Y(_2968_),
    .A(_2967_));
 sg13g2_xnor2_1 _7260_ (.Y(_2969_),
    .A(_2962_),
    .B(_2967_));
 sg13g2_and2_1 _7261_ (.A(_2932_),
    .B(_2969_),
    .X(_2970_));
 sg13g2_xor2_1 _7262_ (.B(_2969_),
    .A(_2932_),
    .X(_2971_));
 sg13g2_xnor2_1 _7263_ (.Y(_2972_),
    .A(_2931_),
    .B(_2971_));
 sg13g2_xor2_1 _7264_ (.B(_2972_),
    .A(_2930_),
    .X(_2973_));
 sg13g2_nand2b_1 _7265_ (.Y(_2974_),
    .B(_2973_),
    .A_N(net742));
 sg13g2_xnor2_1 _7266_ (.Y(_2975_),
    .A(net742),
    .B(_2973_));
 sg13g2_nand2_1 _7267_ (.Y(_2976_),
    .A(_2929_),
    .B(_2975_));
 sg13g2_xnor2_1 _7268_ (.Y(_2977_),
    .A(_2929_),
    .B(_2975_));
 sg13g2_xnor2_1 _7269_ (.Y(_2978_),
    .A(_2928_),
    .B(_2977_));
 sg13g2_or2_1 _7270_ (.X(_2979_),
    .B(_2978_),
    .A(_3127_));
 sg13g2_xnor2_1 _7271_ (.Y(_2980_),
    .A(_3127_),
    .B(_2978_));
 sg13g2_xnor2_1 _7272_ (.Y(_2981_),
    .A(_2927_),
    .B(_2980_));
 sg13g2_nand2_1 _7273_ (.Y(_2982_),
    .A(net835),
    .B(_2981_));
 sg13g2_o21ai_1 _7274_ (.B1(_2982_),
    .Y(_2983_),
    .A1(net834),
    .A2(_1893_));
 sg13g2_nand2_1 _7275_ (.Y(_2984_),
    .A(net886),
    .B(net736));
 sg13g2_o21ai_1 _7276_ (.B1(_2984_),
    .Y(_0163_),
    .A1(net735),
    .A2(_2983_));
 sg13g2_a21oi_2 _7277_ (.B1(net735),
    .Y(_2985_),
    .A2(_1905_),
    .A1(net840));
 sg13g2_o21ai_1 _7278_ (.B1(_2979_),
    .Y(_2986_),
    .A1(_2927_),
    .A2(_2980_));
 sg13g2_o21ai_1 _7279_ (.B1(_2976_),
    .Y(_2987_),
    .A1(_2928_),
    .A2(_2977_));
 sg13g2_o21ai_1 _7280_ (.B1(_2974_),
    .Y(_2988_),
    .A1(_2930_),
    .A2(_2972_));
 sg13g2_a21oi_1 _7281_ (.A1(_2931_),
    .A2(_2971_),
    .Y(_2989_),
    .B1(_2970_));
 sg13g2_o21ai_1 _7282_ (.B1(_2964_),
    .Y(_2990_),
    .A1(_2840_),
    .A2(_2966_));
 sg13g2_o21ai_1 _7283_ (.B1(_2961_),
    .Y(_2991_),
    .A1(_2962_),
    .A2(_2968_));
 sg13g2_o21ai_1 _7284_ (.B1(_2952_),
    .Y(_2992_),
    .A1(_2954_),
    .A2(_2959_));
 sg13g2_o21ai_1 _7285_ (.B1(_2943_),
    .Y(_2993_),
    .A1(_2944_),
    .A2(_2950_));
 sg13g2_nand2_1 _7286_ (.Y(_2994_),
    .A(_2938_),
    .B(_2941_));
 sg13g2_nand2_1 _7287_ (.Y(_2995_),
    .A(net886),
    .B(net915));
 sg13g2_nor2_1 _7288_ (.A(net919),
    .B(net879),
    .Y(_2996_));
 sg13g2_nand3_1 _7289_ (.B(net884),
    .C(_2996_),
    .A(net916),
    .Y(_2997_));
 sg13g2_a21o_1 _7290_ (.A2(net884),
    .A1(net916),
    .B1(_2996_),
    .X(_2998_));
 sg13g2_and2_1 _7291_ (.A(_2997_),
    .B(_2998_),
    .X(_2999_));
 sg13g2_nand2b_1 _7292_ (.Y(_3000_),
    .B(_2999_),
    .A_N(_2995_));
 sg13g2_xnor2_1 _7293_ (.Y(_3001_),
    .A(_2995_),
    .B(_2999_));
 sg13g2_and2_1 _7294_ (.A(_2994_),
    .B(_3001_),
    .X(_3002_));
 sg13g2_or2_1 _7295_ (.X(_3003_),
    .B(_3001_),
    .A(_2994_));
 sg13g2_nand2b_1 _7296_ (.Y(_3004_),
    .B(_3003_),
    .A_N(_3002_));
 sg13g2_and4_1 _7297_ (.A(net890),
    .B(net889),
    .C(net913),
    .D(net910),
    .X(_3005_));
 sg13g2_a22oi_1 _7298_ (.Y(_3006_),
    .B1(net910),
    .B2(net890),
    .A2(net913),
    .A1(net889));
 sg13g2_nor3_1 _7299_ (.A(_2945_),
    .B(_3005_),
    .C(_3006_),
    .Y(_3007_));
 sg13g2_o21ai_1 _7300_ (.B1(_2945_),
    .Y(_3008_),
    .A1(_3005_),
    .A2(_3006_));
 sg13g2_nor2b_1 _7301_ (.A(_3007_),
    .B_N(_3008_),
    .Y(_3009_));
 sg13g2_xnor2_1 _7302_ (.Y(_3010_),
    .A(_3004_),
    .B(_3009_));
 sg13g2_and2_1 _7303_ (.A(_2993_),
    .B(_3010_),
    .X(_3011_));
 sg13g2_or2_1 _7304_ (.X(_3012_),
    .B(_3010_),
    .A(_2993_));
 sg13g2_nand2b_1 _7305_ (.Y(_3013_),
    .B(_3012_),
    .A_N(_3011_));
 sg13g2_o21ai_1 _7306_ (.B1(_2947_),
    .Y(_3014_),
    .A1(_2945_),
    .A2(_2948_));
 sg13g2_and2_1 _7307_ (.A(_2898_),
    .B(_3014_),
    .X(_3015_));
 sg13g2_xor2_1 _7308_ (.B(_3014_),
    .A(_2898_),
    .X(_3016_));
 sg13g2_xor2_1 _7309_ (.B(_3016_),
    .A(_2955_),
    .X(_3017_));
 sg13g2_xnor2_1 _7310_ (.Y(_3018_),
    .A(_3013_),
    .B(_3017_));
 sg13g2_xnor2_1 _7311_ (.Y(_3019_),
    .A(_2992_),
    .B(_3018_));
 sg13g2_a21o_1 _7312_ (.A2(_2958_),
    .A1(_2955_),
    .B1(_2957_),
    .X(_3020_));
 sg13g2_xor2_1 _7313_ (.B(_3020_),
    .A(net741),
    .X(_3021_));
 sg13g2_nor2b_1 _7314_ (.A(_2840_),
    .B_N(_3021_),
    .Y(_3022_));
 sg13g2_xnor2_1 _7315_ (.Y(_3023_),
    .A(_2840_),
    .B(_3021_));
 sg13g2_nor2b_1 _7316_ (.A(_3019_),
    .B_N(_3023_),
    .Y(_3024_));
 sg13g2_xnor2_1 _7317_ (.Y(_3025_),
    .A(_3019_),
    .B(_3023_));
 sg13g2_and2_1 _7318_ (.A(_2991_),
    .B(_3025_),
    .X(_3026_));
 sg13g2_xor2_1 _7319_ (.B(_3025_),
    .A(_2991_),
    .X(_3027_));
 sg13g2_xnor2_1 _7320_ (.Y(_3028_),
    .A(_2990_),
    .B(_3027_));
 sg13g2_xor2_1 _7321_ (.B(_3028_),
    .A(_2989_),
    .X(_3029_));
 sg13g2_nand2b_1 _7322_ (.Y(_3030_),
    .B(_3029_),
    .A_N(net742));
 sg13g2_xnor2_1 _7323_ (.Y(_3031_),
    .A(net742),
    .B(_3029_));
 sg13g2_xnor2_1 _7324_ (.Y(_3032_),
    .A(_2988_),
    .B(_3031_));
 sg13g2_nor2b_1 _7325_ (.A(_3032_),
    .B_N(_2987_),
    .Y(_3033_));
 sg13g2_xor2_1 _7326_ (.B(_3032_),
    .A(_2987_),
    .X(_3034_));
 sg13g2_xnor2_1 _7327_ (.Y(_3035_),
    .A(\i_coord.y0[1] ),
    .B(_3034_));
 sg13g2_o21ai_1 _7328_ (.B1(net835),
    .Y(_3036_),
    .A1(_2986_),
    .A2(_3035_));
 sg13g2_a21o_1 _7329_ (.A2(_3035_),
    .A1(_2986_),
    .B1(_3036_),
    .X(_3037_));
 sg13g2_a22oi_1 _7330_ (.Y(_0164_),
    .B1(_2985_),
    .B2(_3037_),
    .A2(net736),
    .A1(_3132_));
 sg13g2_nor2_1 _7331_ (.A(_0020_),
    .B(_3034_),
    .Y(_3038_));
 sg13g2_a21oi_1 _7332_ (.A1(_2986_),
    .A2(_3035_),
    .Y(_3039_),
    .B1(_3038_));
 sg13g2_a21oi_1 _7333_ (.A1(_2988_),
    .A2(_3031_),
    .Y(_3040_),
    .B1(_3033_));
 sg13g2_o21ai_1 _7334_ (.B1(_3030_),
    .Y(_3041_),
    .A1(_2989_),
    .A2(_3028_));
 sg13g2_a21oi_1 _7335_ (.A1(_2990_),
    .A2(_3027_),
    .Y(_3042_),
    .B1(_3026_));
 sg13g2_a21oi_1 _7336_ (.A1(net741),
    .A2(_3020_),
    .Y(_3043_),
    .B1(_3022_));
 sg13g2_o21ai_1 _7337_ (.B1(_2712_),
    .Y(_3044_),
    .A1(_2633_),
    .A2(_2778_));
 sg13g2_o21ai_1 _7338_ (.B1(_3044_),
    .Y(_3045_),
    .A1(_2633_),
    .A2(_2712_));
 sg13g2_a21oi_1 _7339_ (.A1(_2955_),
    .A2(_3016_),
    .Y(_3046_),
    .B1(_3015_));
 sg13g2_a21oi_1 _7340_ (.A1(_3012_),
    .A2(_3017_),
    .Y(_3047_),
    .B1(_3011_));
 sg13g2_nor2_1 _7341_ (.A(net916),
    .B(net879),
    .Y(_3048_));
 sg13g2_nand2_1 _7342_ (.Y(_3049_),
    .A(net915),
    .B(net884));
 sg13g2_xnor2_1 _7343_ (.Y(_3050_),
    .A(_3048_),
    .B(_3049_));
 sg13g2_a22oi_1 _7344_ (.Y(_3051_),
    .B1(_2896_),
    .B2(_2765_),
    .A2(_2831_),
    .A1(net901));
 sg13g2_nand2_1 _7345_ (.Y(_3052_),
    .A(net886),
    .B(net911));
 sg13g2_xnor2_1 _7346_ (.Y(_3053_),
    .A(_3051_),
    .B(_3052_));
 sg13g2_nor2_1 _7347_ (.A(_3005_),
    .B(_3007_),
    .Y(_3054_));
 sg13g2_nand2_1 _7348_ (.Y(_3055_),
    .A(_2997_),
    .B(_3000_));
 sg13g2_a21oi_1 _7349_ (.A1(_3003_),
    .A2(_3009_),
    .Y(_3056_),
    .B1(_3002_));
 sg13g2_xnor2_1 _7350_ (.Y(_3057_),
    .A(net893),
    .B(net890));
 sg13g2_xnor2_1 _7351_ (.Y(_3058_),
    .A(net887),
    .B(_3057_));
 sg13g2_nand2_1 _7352_ (.Y(_3059_),
    .A(net909),
    .B(_3058_));
 sg13g2_xor2_1 _7353_ (.B(_3055_),
    .A(_3050_),
    .X(_3060_));
 sg13g2_xnor2_1 _7354_ (.Y(_3061_),
    .A(_3054_),
    .B(_3060_));
 sg13g2_xnor2_1 _7355_ (.Y(_3062_),
    .A(_3056_),
    .B(_3061_));
 sg13g2_xnor2_1 _7356_ (.Y(_3063_),
    .A(_3053_),
    .B(_3059_));
 sg13g2_xnor2_1 _7357_ (.Y(_3064_),
    .A(_3062_),
    .B(_3063_));
 sg13g2_xnor2_1 _7358_ (.Y(_3065_),
    .A(_3047_),
    .B(_3064_));
 sg13g2_xnor2_1 _7359_ (.Y(_3066_),
    .A(_3046_),
    .B(_3065_));
 sg13g2_xnor2_1 _7360_ (.Y(_3067_),
    .A(_3045_),
    .B(_3066_));
 sg13g2_xnor2_1 _7361_ (.Y(_3068_),
    .A(_3043_),
    .B(_3067_));
 sg13g2_xnor2_1 _7362_ (.Y(_3069_),
    .A(\i_coord.y0[1] ),
    .B(net742));
 sg13g2_a21oi_1 _7363_ (.A1(_2992_),
    .A2(_3018_),
    .Y(_3070_),
    .B1(_3024_));
 sg13g2_xnor2_1 _7364_ (.Y(_3071_),
    .A(_3069_),
    .B(_3070_));
 sg13g2_xnor2_1 _7365_ (.Y(_3072_),
    .A(_3068_),
    .B(_3071_));
 sg13g2_xnor2_1 _7366_ (.Y(_3073_),
    .A(_3042_),
    .B(_3072_));
 sg13g2_xnor2_1 _7367_ (.Y(_3074_),
    .A(_3041_),
    .B(_3073_));
 sg13g2_xnor2_1 _7368_ (.Y(_3075_),
    .A(_3040_),
    .B(_3074_));
 sg13g2_xnor2_1 _7369_ (.Y(_3076_),
    .A(_3039_),
    .B(_3075_));
 sg13g2_nand2_1 _7370_ (.Y(_3077_),
    .A(net835),
    .B(_3076_));
 sg13g2_a22oi_1 _7371_ (.Y(_0165_),
    .B1(_2985_),
    .B2(_3077_),
    .A2(net736),
    .A1(net879));
 sg13g2_a21oi_1 _7372_ (.A1(\i_coord.l_xir.genblk2[0].state.Q ),
    .A2(net798),
    .Y(_3078_),
    .B1(net206));
 sg13g2_nor2_1 _7373_ (.A(net795),
    .B(_1314_),
    .Y(_3079_));
 sg13g2_nor3_1 _7374_ (.A(net782),
    .B(_3078_),
    .C(_3079_),
    .Y(_0170_));
 sg13g2_xor2_1 _7375_ (.B(_1315_),
    .A(_1314_),
    .X(_3080_));
 sg13g2_o21ai_1 _7376_ (.B1(net771),
    .Y(_3081_),
    .A1(net271),
    .A2(net798));
 sg13g2_a21oi_1 _7377_ (.A1(net798),
    .A2(_3080_),
    .Y(_0171_),
    .B1(_3081_));
 sg13g2_xor2_1 _7378_ (.B(_1317_),
    .A(_1313_),
    .X(_3082_));
 sg13g2_o21ai_1 _7379_ (.B1(net771),
    .Y(_3083_),
    .A1(net247),
    .A2(net798));
 sg13g2_a21oi_1 _7380_ (.A1(net798),
    .A2(_3082_),
    .Y(_0172_),
    .B1(_3083_));
 sg13g2_buf_1 _7381_ (.A(net204),
    .X(\i_vga.timing_ver.blank ));
 sg13g2_dfrbp_1 _7382_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net51),
    .D(_0033_),
    .Q_N(\i_mandel.i_xy.hc.genblk1.genblk1.CG.GATE ),
    .Q(\i_mandel.i_xy.phase ));
 sg13g2_dfrbp_1 _7383_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net42),
    .D(net215),
    .Q_N(_3643_),
    .Q(\step[1] ));
 sg13g2_dfrbp_1 _7384_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net41),
    .D(_0035_),
    .Q_N(_3642_),
    .Q(\step[2] ));
 sg13g2_dfrbp_1 _7385_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net40),
    .D(net195),
    .Q_N(_3641_),
    .Q(\step[3] ));
 sg13g2_dfrbp_1 _7386_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net39),
    .D(_0037_),
    .Q_N(_3640_),
    .Q(\step[4] ));
 sg13g2_dfrbp_1 _7387_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net38),
    .D(_0038_),
    .Q_N(_3639_),
    .Q(\i_coord.x_row_start[-10] ));
 sg13g2_dfrbp_1 _7388_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0039_),
    .Q_N(_3638_),
    .Q(\i_coord.x_row_start[-9] ));
 sg13g2_dfrbp_1 _7389_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net36),
    .D(_0040_),
    .Q_N(_3637_),
    .Q(\i_coord.x_row_start[-8] ));
 sg13g2_dfrbp_1 _7390_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net35),
    .D(_0041_),
    .Q_N(_3636_),
    .Q(\i_coord.x_row_start[-7] ));
 sg13g2_dfrbp_1 _7391_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net34),
    .D(_0042_),
    .Q_N(_3635_),
    .Q(\i_coord.x_row_start[-6] ));
 sg13g2_dfrbp_1 _7392_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net33),
    .D(_0043_),
    .Q_N(_3634_),
    .Q(\i_coord.x_row_start[-5] ));
 sg13g2_dfrbp_1 _7393_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net179),
    .D(_0044_),
    .Q_N(_3633_),
    .Q(\i_coord.x_row_start[-4] ));
 sg13g2_dfrbp_1 _7394_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net178),
    .D(_0045_),
    .Q_N(_3632_),
    .Q(\i_coord.x_row_start[-3] ));
 sg13g2_dfrbp_1 _7395_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net177),
    .D(_0046_),
    .Q_N(_3631_),
    .Q(\i_coord.x_row_start[-2] ));
 sg13g2_dfrbp_1 _7396_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net176),
    .D(_0047_),
    .Q_N(_3630_),
    .Q(\i_coord.x_row_start[-1] ));
 sg13g2_dfrbp_1 _7397_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net175),
    .D(_0048_),
    .Q_N(_3629_),
    .Q(\i_coord.x_row_start[0] ));
 sg13g2_dfrbp_1 _7398_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net174),
    .D(_0049_),
    .Q_N(_3628_),
    .Q(\i_coord.x_row_start[1] ));
 sg13g2_dfrbp_1 _7399_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net52),
    .D(net226),
    .Q_N(_3644_),
    .Q(\i_coord.x_row_start[2] ));
 sg13g2_dlhq_1 _7400_ (.D(\i_coord.l_xir.genblk2[0].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xir.gated_clk ),
    .Q(\i_coord.l_xir.genblk2[0].state.Q ));
 sg13g2_dlhq_1 _7401_ (.D(\i_coord.l_xir.genblk2[1].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xir.gated_clk ),
    .Q(\i_coord.l_xir.genblk2[1].state.Q ));
 sg13g2_dlhq_1 _7402_ (.D(\i_coord.l_xir.genblk2[2].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xir.gated_clk ),
    .Q(\i_coord.l_xir.genblk2[2].state.Q ));
 sg13g2_dlhq_1 _7403_ (.D(\i_coord.l_xir.genblk2[3].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xir.gated_clk ),
    .Q(\i_coord.l_xir.genblk2[3].state.Q ));
 sg13g2_dlhq_1 _7404_ (.D(\i_coord.l_xir.genblk2[4].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xir.gated_clk ),
    .Q(\i_coord.l_xir.genblk2[4].state.Q ));
 sg13g2_dlhq_1 _7405_ (.D(\i_coord.l_xir.genblk2[5].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xir.gated_clk ),
    .Q(\i_coord.l_xir.genblk2[5].state.Q ));
 sg13g2_dlhq_1 _7406_ (.D(\i_coord.l_xir.genblk2[6].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xir.gated_clk ),
    .Q(\i_coord.l_xir.genblk2[6].state.Q ));
 sg13g2_dlhq_1 _7407_ (.D(\i_coord.l_xir.genblk2[7].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xir.gated_clk ),
    .Q(\i_coord.l_xir.genblk2[7].state.Q ));
 sg13g2_dlhq_1 _7408_ (.D(\i_coord.l_xir.genblk2[0].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[0].state.Q ));
 sg13g2_dlhq_1 _7409_ (.D(\i_coord.l_xir.genblk2[1].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[1].state.Q ));
 sg13g2_dlhq_1 _7410_ (.D(\i_coord.l_xir.genblk2[2].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[2].state.Q ));
 sg13g2_dlhq_1 _7411_ (.D(\i_coord.l_xir.genblk2[3].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[3].state.Q ));
 sg13g2_dlhq_1 _7412_ (.D(\i_coord.l_xir.genblk2[4].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[4].state.Q ));
 sg13g2_dlhq_1 _7413_ (.D(\i_coord.l_xir.genblk2[5].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[5].state.Q ));
 sg13g2_dlhq_1 _7414_ (.D(\i_coord.l_xir.genblk2[6].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[6].state.Q ));
 sg13g2_dlhq_1 _7415_ (.D(\i_coord.l_xir.genblk2[7].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[7].state.Q ));
 sg13g2_dlhq_1 _7416_ (.D(\i_coord.l_xl.genblk2[11].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[8].state.Q ));
 sg13g2_dlhq_1 _7417_ (.D(\i_coord.l_xl.genblk2[12].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_yip.gated_clk ),
    .Q(\i_coord.l_yip.genblk2[9].state.Q ));
 sg13g2_dlhq_1 _7418_ (.D(\i_coord.l_xip.genblk2[0].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[0].state.Q ));
 sg13g2_dlhq_1 _7419_ (.D(\i_coord.l_xip.genblk2[1].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[1].state.Q ));
 sg13g2_dlhq_1 _7420_ (.D(\i_coord.l_xip.genblk2[2].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[2].state.Q ));
 sg13g2_dlhq_1 _7421_ (.D(\i_coord.l_xip.genblk2[3].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[3].state.Q ));
 sg13g2_dlhq_1 _7422_ (.D(\i_coord.l_xip.genblk2[4].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[4].state.Q ));
 sg13g2_dlhq_1 _7423_ (.D(\i_coord.l_xip.genblk2[5].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[5].state.Q ));
 sg13g2_dlhq_1 _7424_ (.D(\i_coord.l_xip.genblk2[6].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[6].state.Q ));
 sg13g2_dlhq_1 _7425_ (.D(\i_coord.l_xip.genblk2[7].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[7].state.Q ));
 sg13g2_dlhq_1 _7426_ (.D(\i_coord.l_xip.genblk2[8].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[8].state.Q ));
 sg13g2_dlhq_1 _7427_ (.D(\i_coord.l_xip.genblk2[9].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xip.gated_clk ),
    .Q(\i_coord.l_xip.genblk2[9].state.Q ));
 sg13g2_dlhq_1 _7428_ (.D(net334),
    .GATE(\clknet_2_0__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[0].state.Q ));
 sg13g2_dlhq_1 _7429_ (.D(net336),
    .GATE(\clknet_2_0__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[1].state.Q ));
 sg13g2_dlhq_1 _7430_ (.D(\i_coord.l_yt.genblk2[2].state.D ),
    .GATE(\clknet_2_0__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[2].state.Q ));
 sg13g2_dlhq_1 _7431_ (.D(\i_coord.l_yt.genblk2[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[3].state.Q ));
 sg13g2_dlhq_1 _7432_ (.D(\i_coord.l_yt.genblk2[4].state.D ),
    .GATE(\clknet_2_1__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[4].state.Q ));
 sg13g2_dlhq_1 _7433_ (.D(\i_coord.l_yt.genblk2[5].state.D ),
    .GATE(\clknet_2_1__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[5].state.Q ));
 sg13g2_dlhq_1 _7434_ (.D(\i_coord.l_yt.genblk2[6].state.D ),
    .GATE(\clknet_2_1__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[6].state.Q ));
 sg13g2_dlhq_1 _7435_ (.D(\i_coord.l_yt.genblk2[7].state.D ),
    .GATE(\clknet_2_1__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[7].state.Q ));
 sg13g2_dlhq_1 _7436_ (.D(\i_coord.l_yt.genblk2[8].state.D ),
    .GATE(\clknet_2_3__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[8].state.Q ));
 sg13g2_dlhq_1 _7437_ (.D(\i_coord.l_yt.genblk2[9].state.D ),
    .GATE(\clknet_2_3__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[9].state.Q ));
 sg13g2_dlhq_1 _7438_ (.D(\i_coord.l_yt.genblk2[10].state.D ),
    .GATE(\clknet_2_3__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[10].state.Q ));
 sg13g2_dlhq_1 _7439_ (.D(\i_coord.l_yt.genblk2[11].state.D ),
    .GATE(\clknet_2_2__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[11].state.Q ));
 sg13g2_dlhq_1 _7440_ (.D(\i_coord.l_yt.genblk2[12].state.D ),
    .GATE(\clknet_2_2__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[12].state.Q ));
 sg13g2_dlhq_1 _7441_ (.D(\i_coord.l_yt.genblk2[13].state.D ),
    .GATE(\clknet_2_2__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[13].state.Q ));
 sg13g2_dlhq_1 _7442_ (.D(\i_coord.l_yt.genblk2[14].state.D ),
    .GATE(\clknet_2_2__leaf_i_coord.l_yt.gated_clk ),
    .Q(\i_coord.l_yt.genblk2[14].state.Q ));
 sg13g2_dfrbp_1 _7443_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net53),
    .D(net351),
    .Q_N(_3645_),
    .Q(\video_colour[0] ));
 sg13g2_dfrbp_1 _7444_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net54),
    .D(_0001_),
    .Q_N(_3646_),
    .Q(\video_colour[1] ));
 sg13g2_dfrbp_1 _7445_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net91),
    .D(_0002_),
    .Q_N(_3647_),
    .Q(\video_colour[2] ));
 sg13g2_dfrbp_1 _7446_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net173),
    .D(_0003_),
    .Q_N(_3627_),
    .Q(\video_colour[3] ));
 sg13g2_dlhq_1 _7447_ (.D(\i_coord.l_xir.genblk2[0].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[3].state.Q ));
 sg13g2_dlhq_1 _7448_ (.D(\i_coord.l_xir.genblk2[1].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[4].state.Q ));
 sg13g2_dlhq_1 _7449_ (.D(\i_coord.l_xir.genblk2[2].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[5].state.Q ));
 sg13g2_dlhq_1 _7450_ (.D(\i_coord.l_xir.genblk2[3].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[6].state.Q ));
 sg13g2_dlhq_1 _7451_ (.D(\i_coord.l_xir.genblk2[4].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[7].state.Q ));
 sg13g2_dlhq_1 _7452_ (.D(\i_coord.l_xir.genblk2[5].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[8].state.Q ));
 sg13g2_dlhq_1 _7453_ (.D(\i_coord.l_xir.genblk2[6].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[9].state.Q ));
 sg13g2_dlhq_1 _7454_ (.D(\i_coord.l_xir.genblk2[7].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[10].state.Q ));
 sg13g2_dlhq_1 _7455_ (.D(\i_coord.l_xl.genblk2[11].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[11].state.Q ));
 sg13g2_dlhq_1 _7456_ (.D(\i_coord.l_xl.genblk2[12].state.D ),
    .GATE(\clknet_1_1__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[12].state.Q ));
 sg13g2_dlhq_1 _7457_ (.D(\i_coord.l_xl.genblk2[13].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[13].state.Q ));
 sg13g2_dlhq_1 _7458_ (.D(\i_coord.l_xl.genblk2[14].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[14].state.Q ));
 sg13g2_dlhq_1 _7459_ (.D(\i_coord.l_xl.genblk2[15].state.D ),
    .GATE(\clknet_1_0__leaf_i_coord.l_xl.gated_clk ),
    .Q(\i_coord.l_xl.genblk2[15].state.Q ));
 sg13g2_dfrbp_1 _7460_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net172),
    .D(_0051_),
    .Q_N(_3626_),
    .Q(\i_coord.y_inc_row[-13] ));
 sg13g2_dfrbp_1 _7461_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net170),
    .D(_0052_),
    .Q_N(_3625_),
    .Q(\i_coord.y_inc_row[-12] ));
 sg13g2_dfrbp_1 _7462_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net168),
    .D(_0053_),
    .Q_N(_3624_),
    .Q(\i_coord.y_inc_row[-11] ));
 sg13g2_dfrbp_1 _7463_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net166),
    .D(_0054_),
    .Q_N(_3623_),
    .Q(\i_coord.y_inc_row[-10] ));
 sg13g2_dfrbp_1 _7464_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net164),
    .D(_0055_),
    .Q_N(_3622_),
    .Q(\i_coord.y_inc_row[-9] ));
 sg13g2_dfrbp_1 _7465_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net162),
    .D(_0056_),
    .Q_N(_3621_),
    .Q(\i_coord.y_inc_row[-8] ));
 sg13g2_dfrbp_1 _7466_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net160),
    .D(_0057_),
    .Q_N(_3620_),
    .Q(\i_coord.y_inc_row[-7] ));
 sg13g2_dfrbp_1 _7467_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net158),
    .D(_0058_),
    .Q_N(_3619_),
    .Q(\i_coord.y_inc_row[-6] ));
 sg13g2_dfrbp_1 _7468_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net156),
    .D(_0059_),
    .Q_N(_3618_),
    .Q(\i_coord.y_row_start[-13] ));
 sg13g2_dfrbp_1 _7469_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net155),
    .D(net234),
    .Q_N(_3617_),
    .Q(\i_coord.y_row_start[-12] ));
 sg13g2_dfrbp_1 _7470_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net154),
    .D(net293),
    .Q_N(_3616_),
    .Q(\i_coord.y_row_start[-11] ));
 sg13g2_dfrbp_1 _7471_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net153),
    .D(_0062_),
    .Q_N(_3615_),
    .Q(\i_coord.y_row_start[-10] ));
 sg13g2_dfrbp_1 _7472_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net152),
    .D(net283),
    .Q_N(_3614_),
    .Q(\i_coord.y_row_start[-9] ));
 sg13g2_dfrbp_1 _7473_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net151),
    .D(_0064_),
    .Q_N(_3613_),
    .Q(\i_coord.y_row_start[-8] ));
 sg13g2_dfrbp_1 _7474_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net150),
    .D(_0065_),
    .Q_N(_3612_),
    .Q(\i_coord.y_row_start[-7] ));
 sg13g2_dfrbp_1 _7475_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net149),
    .D(net253),
    .Q_N(_3611_),
    .Q(\i_coord.y_row_start[-6] ));
 sg13g2_dfrbp_1 _7476_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net148),
    .D(_0067_),
    .Q_N(_3610_),
    .Q(\i_coord.y_row_start[-5] ));
 sg13g2_dfrbp_1 _7477_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net147),
    .D(_0068_),
    .Q_N(_3609_),
    .Q(\i_coord.y_row_start[-4] ));
 sg13g2_dfrbp_1 _7478_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net146),
    .D(_0069_),
    .Q_N(_3608_),
    .Q(\i_coord.y_row_start[-3] ));
 sg13g2_dfrbp_1 _7479_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net145),
    .D(_0070_),
    .Q_N(_3607_),
    .Q(\i_coord.y_row_start[-2] ));
 sg13g2_dfrbp_1 _7480_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net144),
    .D(_0071_),
    .Q_N(_3606_),
    .Q(\i_coord.y_row_start[-1] ));
 sg13g2_dfrbp_1 _7481_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net143),
    .D(_0072_),
    .Q_N(_3605_),
    .Q(\i_coord.y_row_start[0] ));
 sg13g2_dfrbp_1 _7482_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net142),
    .D(_0073_),
    .Q_N(_3604_),
    .Q(\i_coord.y_row_start[1] ));
 sg13g2_dfrbp_1 _7483_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net141),
    .D(net183),
    .Q_N(_0030_),
    .Q(\i_coord.demo_update_delay ));
 sg13g2_dfrbp_1 _7484_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net139),
    .D(_0075_),
    .Q_N(_3603_),
    .Q(\video_colour[4] ));
 sg13g2_dfrbp_1 _7485_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net138),
    .D(_0076_),
    .Q_N(_3602_),
    .Q(\video_colour[5] ));
 sg13g2_dlhq_1 _7486_ (.D(\i_mandel.i_xy.hc.genblk2[11].state.D ),
    .GATE(\clknet_3_7__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[11].state.Q ));
 sg13g2_dlhq_1 _7487_ (.D(\i_mandel.i_xy.hc.genblk2[10].state.D ),
    .GATE(\clknet_3_5__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[10].state.Q ));
 sg13g2_dlhq_1 _7488_ (.D(\i_mandel.i_xy.hc.genblk2[9].state.D ),
    .GATE(\clknet_3_5__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[9].state.Q ));
 sg13g2_dlhq_1 _7489_ (.D(\i_mandel.i_xy.hc.genblk2[8].state.D ),
    .GATE(\clknet_3_5__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[8].state.Q ));
 sg13g2_dlhq_1 _7490_ (.D(\i_mandel.i_xy.hc.genblk2[7].state.D ),
    .GATE(\clknet_3_5__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[7].state.Q ));
 sg13g2_dlhq_1 _7491_ (.D(\i_mandel.i_xy.hc.genblk2[6].state.D ),
    .GATE(\clknet_3_4__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[6].state.Q ));
 sg13g2_dlhq_1 _7492_ (.D(\i_mandel.i_xy.hc.genblk2[5].state.D ),
    .GATE(\clknet_3_4__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[5].state.Q ));
 sg13g2_dlhq_1 _7493_ (.D(\i_mandel.i_xy.hc.genblk2[4].state.D ),
    .GATE(\clknet_3_7__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[4].state.Q ));
 sg13g2_dlhq_1 _7494_ (.D(\i_mandel.i_xy.hc.genblk2[3].state.D ),
    .GATE(\clknet_3_7__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[3].state.Q ));
 sg13g2_dlhq_1 _7495_ (.D(\i_mandel.i_xy.hc.genblk2[2].state.D ),
    .GATE(\clknet_3_6__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[2].state.Q ));
 sg13g2_dlhq_1 _7496_ (.D(\i_mandel.i_xy.hc.genblk2[1].state.D ),
    .GATE(\clknet_3_4__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[1].state.Q ));
 sg13g2_dlhq_1 _7497_ (.D(\i_mandel.i_xy.hc.genblk2[0].state.D ),
    .GATE(\clknet_3_4__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.i_xy.hc.genblk2[0].state.Q ));
 sg13g2_dlhq_1 _7498_ (.D(\i_mandel.l_sq.genblk2[0].state.D ),
    .GATE(\clknet_3_6__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[0].state.Q ));
 sg13g2_dlhq_1 _7499_ (.D(\i_mandel.l_sq.genblk2[1].state.D ),
    .GATE(\clknet_3_6__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[1].state.Q ));
 sg13g2_dlhq_1 _7500_ (.D(\i_mandel.l_sq.genblk2[2].state.D ),
    .GATE(\clknet_3_6__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[2].state.Q ));
 sg13g2_dlhq_1 _7501_ (.D(\i_mandel.l_sq.genblk2[3].state.D ),
    .GATE(\clknet_3_1__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[3].state.Q ));
 sg13g2_dlhq_1 _7502_ (.D(\i_mandel.l_sq.genblk2[4].state.D ),
    .GATE(\clknet_3_1__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[4].state.Q ));
 sg13g2_dlhq_1 _7503_ (.D(\i_mandel.l_sq.genblk2[5].state.D ),
    .GATE(\clknet_3_1__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[5].state.Q ));
 sg13g2_dlhq_1 _7504_ (.D(\i_mandel.l_sq.genblk2[6].state.D ),
    .GATE(\clknet_3_1__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[6].state.Q ));
 sg13g2_dlhq_1 _7505_ (.D(\i_mandel.l_sq.genblk2[7].state.D ),
    .GATE(\clknet_3_3__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[7].state.Q ));
 sg13g2_dlhq_1 _7506_ (.D(\i_mandel.l_sq.genblk2[8].state.D ),
    .GATE(\clknet_3_0__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[8].state.Q ));
 sg13g2_dlhq_1 _7507_ (.D(\i_mandel.l_sq.genblk2[9].state.D ),
    .GATE(\clknet_3_0__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[9].state.Q ));
 sg13g2_dlhq_1 _7508_ (.D(\i_mandel.l_sq.genblk2[10].state.D ),
    .GATE(\clknet_3_3__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[10].state.Q ));
 sg13g2_dlhq_1 _7509_ (.D(\i_mandel.l_sq.genblk2[11].state.D ),
    .GATE(\clknet_3_3__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[11].state.Q ));
 sg13g2_dlhq_1 _7510_ (.D(\i_mandel.l_sq.genblk2[12].state.D ),
    .GATE(\clknet_3_2__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[12].state.Q ));
 sg13g2_dlhq_1 _7511_ (.D(\i_mandel.l_sq.genblk2[13].state.D ),
    .GATE(\clknet_3_0__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[13].state.Q ));
 sg13g2_dlhq_1 _7512_ (.D(\i_mandel.l_sq.genblk2[14].state.D ),
    .GATE(\clknet_3_2__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[14].state.Q ));
 sg13g2_dlhq_1 _7513_ (.D(\i_mandel.l_sq.genblk2[15].state.D ),
    .GATE(\clknet_3_0__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[15].state.Q ));
 sg13g2_dlhq_1 _7514_ (.D(\i_mandel.l_sq.genblk2[16].state.D ),
    .GATE(\clknet_3_3__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[16].state.Q ));
 sg13g2_dlhq_1 _7515_ (.D(\i_mandel.l_sq.genblk2[17].state.D ),
    .GATE(\clknet_3_2__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[17].state.Q ));
 sg13g2_dlhq_1 _7516_ (.D(\i_mandel.l_sq.genblk2[18].state.D ),
    .GATE(\clknet_3_2__leaf_i_mandel.i_xy.hc.gated_clk ),
    .Q(\i_mandel.l_sq.genblk2[18].state.Q ));
 sg13g2_dfrbp_1 _7517_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net137),
    .D(net317),
    .Q_N(_3601_),
    .Q(\i_vga.timing_ver.counter[0] ));
 sg13g2_dfrbp_1 _7518_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net135),
    .D(_0078_),
    .Q_N(_3600_),
    .Q(\i_vga.timing_ver.counter[1] ));
 sg13g2_dfrbp_1 _7519_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net133),
    .D(net323),
    .Q_N(_3599_),
    .Q(\i_vga.timing_ver.counter[2] ));
 sg13g2_dfrbp_1 _7520_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net131),
    .D(_0080_),
    .Q_N(_3598_),
    .Q(\i_vga.timing_ver.counter[3] ));
 sg13g2_dfrbp_1 _7521_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net129),
    .D(_0081_),
    .Q_N(_3597_),
    .Q(\i_vga.timing_ver.counter[4] ));
 sg13g2_dfrbp_1 _7522_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net127),
    .D(_0082_),
    .Q_N(_3596_),
    .Q(\i_vga.timing_ver.counter[5] ));
 sg13g2_dfrbp_1 _7523_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net125),
    .D(_0083_),
    .Q_N(_3595_),
    .Q(\i_vga.timing_ver.counter[6] ));
 sg13g2_dfrbp_1 _7524_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net123),
    .D(net223),
    .Q_N(_3594_),
    .Q(\i_vga.timing_ver.counter[7] ));
 sg13g2_dfrbp_1 _7525_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net121),
    .D(_0085_),
    .Q_N(_0029_),
    .Q(\i_vga.timing_ver.counter[8] ));
 sg13g2_dfrbp_1 _7526_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net103),
    .D(_0086_),
    .Q_N(_0031_),
    .Q(\i_vga.timing_ver.counter[9] ));
 sg13g2_dfrbp_1 _7527_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net119),
    .D(net181),
    .Q_N(_3593_),
    .Q(\i_vga.timing_ver.sync ));
 sg13g2_dfrbp_1 _7528_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net117),
    .D(_0087_),
    .Q_N(_3592_),
    .Q(\i_vga.timing_hor.counter[0] ));
 sg13g2_dfrbp_1 _7529_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net115),
    .D(_0088_),
    .Q_N(_3591_),
    .Q(\i_vga.timing_hor.counter[1] ));
 sg13g2_dfrbp_1 _7530_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net113),
    .D(net198),
    .Q_N(_3590_),
    .Q(\i_vga.timing_hor.counter[2] ));
 sg13g2_dfrbp_1 _7531_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net111),
    .D(net236),
    .Q_N(_3589_),
    .Q(\i_vga.timing_hor.counter[3] ));
 sg13g2_dfrbp_1 _7532_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net109),
    .D(_0091_),
    .Q_N(_3588_),
    .Q(\i_vga.timing_hor.counter[4] ));
 sg13g2_dfrbp_1 _7533_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net107),
    .D(_0092_),
    .Q_N(_0028_),
    .Q(\i_vga.timing_hor.counter[5] ));
 sg13g2_dfrbp_1 _7534_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net105),
    .D(net329),
    .Q_N(_3587_),
    .Q(\i_vga.timing_hor.counter[6] ));
 sg13g2_dfrbp_1 _7535_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net101),
    .D(net256),
    .Q_N(_3586_),
    .Q(\i_vga.timing_hor.counter[7] ));
 sg13g2_dfrbp_1 _7536_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net99),
    .D(_0095_),
    .Q_N(_3585_),
    .Q(\i_vga.timing_hor.counter[8] ));
 sg13g2_dfrbp_1 _7537_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net97),
    .D(_0096_),
    .Q_N(_3584_),
    .Q(\i_vga.timing_hor.counter[9] ));
 sg13g2_dfrbp_1 _7538_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net104),
    .D(_0097_),
    .Q_N(_0032_),
    .Q(\i_vga.timing_hor.counter[10] ));
 sg13g2_dfrbp_1 _7539_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net136),
    .D(_0004_),
    .Q_N(_3648_),
    .Q(\i_vga.hsync ));
 sg13g2_dfrbp_1 _7540_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net95),
    .D(\i_vga.timing_ver.blank ),
    .Q_N(_3583_),
    .Q(\i_vga.vblank ));
 sg13g2_dfrbp_1 _7541_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net93),
    .D(_0098_),
    .Q_N(_0027_),
    .Q(\i_coord.demo_update ));
 sg13g2_dfrbp_1 _7542_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net92),
    .D(_0099_),
    .Q_N(_3582_),
    .Q(\i_coord.x0[-13] ));
 sg13g2_dfrbp_1 _7543_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net90),
    .D(_0100_),
    .Q_N(_3581_),
    .Q(\i_coord.x0[-12] ));
 sg13g2_dfrbp_1 _7544_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net89),
    .D(_0101_),
    .Q_N(_3580_),
    .Q(\i_coord.x0[-11] ));
 sg13g2_dfrbp_1 _7545_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net88),
    .D(_0102_),
    .Q_N(_3579_),
    .Q(\i_coord.x0[-10] ));
 sg13g2_dfrbp_1 _7546_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net87),
    .D(_0103_),
    .Q_N(_3578_),
    .Q(\i_coord.x0[-9] ));
 sg13g2_dfrbp_1 _7547_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net86),
    .D(_0104_),
    .Q_N(_3577_),
    .Q(\i_coord.x0[-8] ));
 sg13g2_dfrbp_1 _7548_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net85),
    .D(_0105_),
    .Q_N(_3576_),
    .Q(\i_coord.x0[-7] ));
 sg13g2_dfrbp_1 _7549_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net84),
    .D(_0106_),
    .Q_N(_3575_),
    .Q(\i_coord.x0[-6] ));
 sg13g2_dfrbp_1 _7550_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net83),
    .D(_0107_),
    .Q_N(_3574_),
    .Q(\i_coord.x0[-5] ));
 sg13g2_dfrbp_1 _7551_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net82),
    .D(_0108_),
    .Q_N(_3573_),
    .Q(\i_coord.x0[-4] ));
 sg13g2_dfrbp_1 _7552_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net81),
    .D(_0109_),
    .Q_N(_3572_),
    .Q(\i_coord.x0[-3] ));
 sg13g2_dfrbp_1 _7553_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net80),
    .D(_0110_),
    .Q_N(_3571_),
    .Q(\i_coord.x0[-2] ));
 sg13g2_dfrbp_1 _7554_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net79),
    .D(_0111_),
    .Q_N(_3570_),
    .Q(\i_coord.x0[-1] ));
 sg13g2_dfrbp_1 _7555_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net78),
    .D(_0112_),
    .Q_N(_3569_),
    .Q(\i_coord.x0[0] ));
 sg13g2_dfrbp_1 _7556_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net77),
    .D(_0113_),
    .Q_N(_3568_),
    .Q(\i_coord.x0[1] ));
 sg13g2_dfrbp_1 _7557_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net76),
    .D(_0114_),
    .Q_N(_3567_),
    .Q(\i_coord.x0[2] ));
 sg13g2_dfrbp_1 _7558_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net75),
    .D(_0115_),
    .Q_N(_0026_),
    .Q(\i_coord.y0[-13] ));
 sg13g2_dfrbp_1 _7559_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net74),
    .D(_0116_),
    .Q_N(_0025_),
    .Q(\i_coord.y0[-12] ));
 sg13g2_dfrbp_1 _7560_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net73),
    .D(_0117_),
    .Q_N(_3566_),
    .Q(\i_coord.y0[-11] ));
 sg13g2_dfrbp_1 _7561_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net72),
    .D(_0118_),
    .Q_N(_3565_),
    .Q(\i_coord.y0[-10] ));
 sg13g2_dfrbp_1 _7562_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net71),
    .D(_0119_),
    .Q_N(_3564_),
    .Q(\i_coord.y0[-9] ));
 sg13g2_dfrbp_1 _7563_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net70),
    .D(_0120_),
    .Q_N(_3563_),
    .Q(\i_coord.y0[-8] ));
 sg13g2_dfrbp_1 _7564_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net69),
    .D(_0121_),
    .Q_N(_0024_),
    .Q(\i_coord.y0[-7] ));
 sg13g2_dfrbp_1 _7565_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net68),
    .D(_0122_),
    .Q_N(_3562_),
    .Q(\i_coord.y0[-6] ));
 sg13g2_dfrbp_1 _7566_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net67),
    .D(_0123_),
    .Q_N(_3561_),
    .Q(\i_coord.y0[-5] ));
 sg13g2_dfrbp_1 _7567_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net66),
    .D(_0124_),
    .Q_N(_3560_),
    .Q(\i_coord.y0[-4] ));
 sg13g2_dfrbp_1 _7568_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net65),
    .D(_0125_),
    .Q_N(_0023_),
    .Q(\i_coord.y0[-3] ));
 sg13g2_dfrbp_1 _7569_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net64),
    .D(_0126_),
    .Q_N(_0022_),
    .Q(\i_coord.y0[-2] ));
 sg13g2_dfrbp_1 _7570_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net63),
    .D(_0127_),
    .Q_N(_0021_),
    .Q(\i_coord.y0[-1] ));
 sg13g2_dfrbp_1 _7571_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net62),
    .D(_0128_),
    .Q_N(_3559_),
    .Q(\i_coord.y0[0] ));
 sg13g2_dfrbp_1 _7572_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net61),
    .D(_0129_),
    .Q_N(_0020_),
    .Q(\i_coord.y0[1] ));
 sg13g2_dfrbp_1 _7573_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net60),
    .D(_0130_),
    .Q_N(_0019_),
    .Q(\i_mandel.i_xy.x[-13] ));
 sg13g2_dfrbp_1 _7574_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0131_),
    .Q_N(_0018_),
    .Q(\i_mandel.i_xy.x[-12] ));
 sg13g2_dfrbp_1 _7575_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net58),
    .D(_0132_),
    .Q_N(_0017_),
    .Q(\i_mandel.i_xy.x[-11] ));
 sg13g2_dfrbp_1 _7576_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net57),
    .D(_0133_),
    .Q_N(_0016_),
    .Q(\i_mandel.i_xy.x[-10] ));
 sg13g2_dfrbp_1 _7577_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net56),
    .D(_0134_),
    .Q_N(_3558_),
    .Q(\i_mandel.i_xy.x[-9] ));
 sg13g2_dfrbp_1 _7578_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net55),
    .D(_0135_),
    .Q_N(_3557_),
    .Q(\i_mandel.i_xy.x[-8] ));
 sg13g2_dfrbp_1 _7579_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net50),
    .D(_0136_),
    .Q_N(_3556_),
    .Q(\i_mandel.i_xy.x[-7] ));
 sg13g2_dfrbp_1 _7580_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net49),
    .D(_0137_),
    .Q_N(_3555_),
    .Q(\i_mandel.i_xy.x[-6] ));
 sg13g2_dfrbp_1 _7581_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net48),
    .D(_0138_),
    .Q_N(_3554_),
    .Q(\i_mandel.i_xy.x[-5] ));
 sg13g2_dfrbp_1 _7582_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net47),
    .D(_0139_),
    .Q_N(_3553_),
    .Q(\i_mandel.i_xy.x[-4] ));
 sg13g2_dfrbp_1 _7583_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0140_),
    .Q_N(_3552_),
    .Q(\i_mandel.i_xy.x[-3] ));
 sg13g2_dfrbp_1 _7584_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net45),
    .D(_0141_),
    .Q_N(_0015_),
    .Q(\i_mandel.i_xy.x[-2] ));
 sg13g2_dfrbp_1 _7585_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0142_),
    .Q_N(_3551_),
    .Q(\i_mandel.i_xy.x[-1] ));
 sg13g2_dfrbp_1 _7586_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net43),
    .D(_0143_),
    .Q_N(_3550_),
    .Q(\i_mandel.i_xy.x[0] ));
 sg13g2_dfrbp_1 _7587_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net171),
    .D(_0144_),
    .Q_N(_3549_),
    .Q(\i_mandel.i_xy.x[1] ));
 sg13g2_dfrbp_1 _7588_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net169),
    .D(_0145_),
    .Q_N(_0014_),
    .Q(\i_mandel.i_xy.x[2] ));
 sg13g2_dfrbp_1 _7589_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net167),
    .D(_0146_),
    .Q_N(_3548_),
    .Q(\iter[0] ));
 sg13g2_dfrbp_1 _7590_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net163),
    .D(_0147_),
    .Q_N(_0013_),
    .Q(\iter[1] ));
 sg13g2_dfrbp_1 _7591_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net159),
    .D(net213),
    .Q_N(_3547_),
    .Q(\iter[2] ));
 sg13g2_dfrbp_1 _7592_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net140),
    .D(net190),
    .Q_N(_3546_),
    .Q(\iter[3] ));
 sg13g2_dfrbp_1 _7593_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net134),
    .D(net201),
    .Q_N(_0012_),
    .Q(\i_mandel.i_xy.y[-13] ));
 sg13g2_dfrbp_1 _7594_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net132),
    .D(_0151_),
    .Q_N(_0011_),
    .Q(\i_mandel.i_xy.y[-12] ));
 sg13g2_dfrbp_1 _7595_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net130),
    .D(_0152_),
    .Q_N(_0010_),
    .Q(\i_mandel.i_xy.y[-11] ));
 sg13g2_dfrbp_1 _7596_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net128),
    .D(_0153_),
    .Q_N(_0009_),
    .Q(\i_mandel.i_xy.y[-10] ));
 sg13g2_dfrbp_1 _7597_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net126),
    .D(_0154_),
    .Q_N(_3545_),
    .Q(\i_mandel.i_xy.y[-9] ));
 sg13g2_dfrbp_1 _7598_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net124),
    .D(_0155_),
    .Q_N(_3544_),
    .Q(\i_mandel.i_xy.y[-8] ));
 sg13g2_dfrbp_1 _7599_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net122),
    .D(_0156_),
    .Q_N(_3543_),
    .Q(\i_mandel.i_xy.y[-7] ));
 sg13g2_dfrbp_1 _7600_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net120),
    .D(_0157_),
    .Q_N(_3542_),
    .Q(\i_mandel.i_xy.y[-6] ));
 sg13g2_dfrbp_1 _7601_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net118),
    .D(_0158_),
    .Q_N(_3541_),
    .Q(\i_mandel.i_xy.y[-5] ));
 sg13g2_dfrbp_1 _7602_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net116),
    .D(_0159_),
    .Q_N(_3540_),
    .Q(\i_mandel.i_xy.y[-4] ));
 sg13g2_dfrbp_1 _7603_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net114),
    .D(_0160_),
    .Q_N(_3539_),
    .Q(\i_mandel.i_xy.y[-3] ));
 sg13g2_dfrbp_1 _7604_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net112),
    .D(_0161_),
    .Q_N(_0008_),
    .Q(\i_mandel.i_xy.y[-2] ));
 sg13g2_dfrbp_1 _7605_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net110),
    .D(_0162_),
    .Q_N(_3538_),
    .Q(\i_mandel.i_xy.y[-1] ));
 sg13g2_dfrbp_1 _7606_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net108),
    .D(_0163_),
    .Q_N(_3537_),
    .Q(\i_mandel.i_xy.y[0] ));
 sg13g2_dfrbp_1 _7607_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net106),
    .D(_0164_),
    .Q_N(_3536_),
    .Q(\i_mandel.i_xy.y[1] ));
 sg13g2_dfrbp_1 _7608_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net102),
    .D(_0165_),
    .Q_N(_0007_),
    .Q(\i_mandel.i_xy.y[2] ));
 sg13g2_dfrbp_1 _7609_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net100),
    .D(_0166_),
    .Q_N(_3535_),
    .Q(\last_iter[0] ));
 sg13g2_dfrbp_1 _7610_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net98),
    .D(_0167_),
    .Q_N(_0006_),
    .Q(\last_iter[1] ));
 sg13g2_dfrbp_1 _7611_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net96),
    .D(_0168_),
    .Q_N(_0005_),
    .Q(\last_iter[2] ));
 sg13g2_dfrbp_1 _7612_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net94),
    .D(_0169_),
    .Q_N(_3534_),
    .Q(\last_iter[3] ));
 sg13g2_dfrbp_1 _7613_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net165),
    .D(_0170_),
    .Q_N(_3533_),
    .Q(\i_coord.x_row_start[-13] ));
 sg13g2_dfrbp_1 _7614_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net157),
    .D(_0171_),
    .Q_N(_3532_),
    .Q(\i_coord.x_row_start[-12] ));
 sg13g2_dfrbp_1 _7615_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net161),
    .D(_0172_),
    .Q_N(_3531_),
    .Q(\i_coord.x_row_start[-11] ));
 sg13g2_tiehi _7391__34 (.L_HI(net34));
 sg13g2_tiehi _7390__35 (.L_HI(net35));
 sg13g2_tiehi _7389__36 (.L_HI(net36));
 sg13g2_tiehi _7388__37 (.L_HI(net37));
 sg13g2_tiehi _7387__38 (.L_HI(net38));
 sg13g2_tiehi _7386__39 (.L_HI(net39));
 sg13g2_tiehi _7385__40 (.L_HI(net40));
 sg13g2_tiehi _7384__41 (.L_HI(net41));
 sg13g2_tiehi _7383__42 (.L_HI(net42));
 sg13g2_tiehi _7586__43 (.L_HI(net43));
 sg13g2_tiehi _7585__44 (.L_HI(net44));
 sg13g2_tiehi _7584__45 (.L_HI(net45));
 sg13g2_tiehi _7583__46 (.L_HI(net46));
 sg13g2_tiehi _7582__47 (.L_HI(net47));
 sg13g2_tiehi _7581__48 (.L_HI(net48));
 sg13g2_tiehi _7580__49 (.L_HI(net49));
 sg13g2_tiehi _7579__50 (.L_HI(net50));
 sg13g2_tiehi _7382__51 (.L_HI(net51));
 sg13g2_tiehi _7399__52 (.L_HI(net52));
 sg13g2_tiehi _7443__53 (.L_HI(net53));
 sg13g2_tiehi _7444__54 (.L_HI(net54));
 sg13g2_tiehi _7578__55 (.L_HI(net55));
 sg13g2_tiehi _7577__56 (.L_HI(net56));
 sg13g2_tiehi _7576__57 (.L_HI(net57));
 sg13g2_tiehi _7575__58 (.L_HI(net58));
 sg13g2_tiehi _7574__59 (.L_HI(net59));
 sg13g2_tiehi _7573__60 (.L_HI(net60));
 sg13g2_tiehi _7572__61 (.L_HI(net61));
 sg13g2_tiehi _7571__62 (.L_HI(net62));
 sg13g2_tiehi _7570__63 (.L_HI(net63));
 sg13g2_tiehi _7569__64 (.L_HI(net64));
 sg13g2_tiehi _7568__65 (.L_HI(net65));
 sg13g2_tiehi _7567__66 (.L_HI(net66));
 sg13g2_tiehi _7566__67 (.L_HI(net67));
 sg13g2_tiehi _7565__68 (.L_HI(net68));
 sg13g2_tiehi _7564__69 (.L_HI(net69));
 sg13g2_tiehi _7563__70 (.L_HI(net70));
 sg13g2_tiehi _7562__71 (.L_HI(net71));
 sg13g2_tiehi _7561__72 (.L_HI(net72));
 sg13g2_tiehi _7560__73 (.L_HI(net73));
 sg13g2_tiehi _7559__74 (.L_HI(net74));
 sg13g2_tiehi _7558__75 (.L_HI(net75));
 sg13g2_tiehi _7557__76 (.L_HI(net76));
 sg13g2_tiehi _7556__77 (.L_HI(net77));
 sg13g2_tiehi _7555__78 (.L_HI(net78));
 sg13g2_tiehi _7554__79 (.L_HI(net79));
 sg13g2_tiehi _7553__80 (.L_HI(net80));
 sg13g2_tiehi _7552__81 (.L_HI(net81));
 sg13g2_tiehi _7551__82 (.L_HI(net82));
 sg13g2_tiehi _7550__83 (.L_HI(net83));
 sg13g2_tiehi _7549__84 (.L_HI(net84));
 sg13g2_tiehi _7548__85 (.L_HI(net85));
 sg13g2_tiehi _7547__86 (.L_HI(net86));
 sg13g2_tiehi _7546__87 (.L_HI(net87));
 sg13g2_tiehi _7545__88 (.L_HI(net88));
 sg13g2_tiehi _7544__89 (.L_HI(net89));
 sg13g2_tiehi _7543__90 (.L_HI(net90));
 sg13g2_tiehi _7445__91 (.L_HI(net91));
 sg13g2_tiehi _7542__92 (.L_HI(net92));
 sg13g2_tiehi _7541__93 (.L_HI(net93));
 sg13g2_tiehi _7612__94 (.L_HI(net94));
 sg13g2_tiehi _7540__95 (.L_HI(net95));
 sg13g2_tiehi _7611__96 (.L_HI(net96));
 sg13g2_tiehi _7537__97 (.L_HI(net97));
 sg13g2_tiehi _7610__98 (.L_HI(net98));
 sg13g2_tiehi _7536__99 (.L_HI(net99));
 sg13g2_tiehi _7609__100 (.L_HI(net100));
 sg13g2_tiehi _7535__101 (.L_HI(net101));
 sg13g2_tiehi _7608__102 (.L_HI(net102));
 sg13g2_tiehi _7526__103 (.L_HI(net103));
 sg13g2_tiehi _7538__104 (.L_HI(net104));
 sg13g2_tiehi _7534__105 (.L_HI(net105));
 sg13g2_tiehi _7607__106 (.L_HI(net106));
 sg13g2_tiehi _7533__107 (.L_HI(net107));
 sg13g2_tiehi _7606__108 (.L_HI(net108));
 sg13g2_tiehi _7532__109 (.L_HI(net109));
 sg13g2_tiehi _7605__110 (.L_HI(net110));
 sg13g2_tiehi _7531__111 (.L_HI(net111));
 sg13g2_tiehi _7604__112 (.L_HI(net112));
 sg13g2_tiehi _7530__113 (.L_HI(net113));
 sg13g2_tiehi _7603__114 (.L_HI(net114));
 sg13g2_tiehi _7529__115 (.L_HI(net115));
 sg13g2_tiehi _7602__116 (.L_HI(net116));
 sg13g2_tiehi _7528__117 (.L_HI(net117));
 sg13g2_tiehi _7601__118 (.L_HI(net118));
 sg13g2_tiehi _7527__119 (.L_HI(net119));
 sg13g2_tiehi _7600__120 (.L_HI(net120));
 sg13g2_tiehi _7525__121 (.L_HI(net121));
 sg13g2_tiehi _7599__122 (.L_HI(net122));
 sg13g2_tiehi _7524__123 (.L_HI(net123));
 sg13g2_tiehi _7598__124 (.L_HI(net124));
 sg13g2_tiehi _7523__125 (.L_HI(net125));
 sg13g2_tiehi _7597__126 (.L_HI(net126));
 sg13g2_tiehi _7522__127 (.L_HI(net127));
 sg13g2_tiehi _7596__128 (.L_HI(net128));
 sg13g2_tiehi _7521__129 (.L_HI(net129));
 sg13g2_tiehi _7595__130 (.L_HI(net130));
 sg13g2_tiehi _7520__131 (.L_HI(net131));
 sg13g2_tiehi _7594__132 (.L_HI(net132));
 sg13g2_tiehi _7519__133 (.L_HI(net133));
 sg13g2_tiehi _7593__134 (.L_HI(net134));
 sg13g2_tiehi _7518__135 (.L_HI(net135));
 sg13g2_tiehi _7539__136 (.L_HI(net136));
 sg13g2_tiehi _7517__137 (.L_HI(net137));
 sg13g2_tiehi _7485__138 (.L_HI(net138));
 sg13g2_tiehi _7484__139 (.L_HI(net139));
 sg13g2_tiehi _7592__140 (.L_HI(net140));
 sg13g2_tiehi _7483__141 (.L_HI(net141));
 sg13g2_tiehi _7482__142 (.L_HI(net142));
 sg13g2_tiehi _7481__143 (.L_HI(net143));
 sg13g2_tiehi _7480__144 (.L_HI(net144));
 sg13g2_tiehi _7479__145 (.L_HI(net145));
 sg13g2_tiehi _7478__146 (.L_HI(net146));
 sg13g2_tiehi _7477__147 (.L_HI(net147));
 sg13g2_tiehi _7476__148 (.L_HI(net148));
 sg13g2_tiehi _7475__149 (.L_HI(net149));
 sg13g2_tiehi _7474__150 (.L_HI(net150));
 sg13g2_tiehi _7473__151 (.L_HI(net151));
 sg13g2_tiehi _7472__152 (.L_HI(net152));
 sg13g2_tiehi _7471__153 (.L_HI(net153));
 sg13g2_tiehi _7470__154 (.L_HI(net154));
 sg13g2_tiehi _7469__155 (.L_HI(net155));
 sg13g2_tiehi _7468__156 (.L_HI(net156));
 sg13g2_tiehi _7614__157 (.L_HI(net157));
 sg13g2_tiehi _7467__158 (.L_HI(net158));
 sg13g2_tiehi _7591__159 (.L_HI(net159));
 sg13g2_tiehi _7466__160 (.L_HI(net160));
 sg13g2_tiehi _7615__161 (.L_HI(net161));
 sg13g2_tiehi _7465__162 (.L_HI(net162));
 sg13g2_tiehi _7590__163 (.L_HI(net163));
 sg13g2_tiehi _7464__164 (.L_HI(net164));
 sg13g2_tiehi _7613__165 (.L_HI(net165));
 sg13g2_tiehi _7463__166 (.L_HI(net166));
 sg13g2_tiehi _7589__167 (.L_HI(net167));
 sg13g2_tiehi _7462__168 (.L_HI(net168));
 sg13g2_tiehi _7588__169 (.L_HI(net169));
 sg13g2_tiehi _7461__170 (.L_HI(net170));
 sg13g2_tiehi _7587__171 (.L_HI(net171));
 sg13g2_tiehi _7460__172 (.L_HI(net172));
 sg13g2_tiehi _7446__173 (.L_HI(net173));
 sg13g2_tiehi _7398__174 (.L_HI(net174));
 sg13g2_tiehi _7397__175 (.L_HI(net175));
 sg13g2_tiehi _7396__176 (.L_HI(net176));
 sg13g2_tiehi _7395__177 (.L_HI(net177));
 sg13g2_tiehi _7394__178 (.L_HI(net178));
 sg13g2_tiehi _7393__179 (.L_HI(net179));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_18 (.L_LO(net18));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_19 (.L_LO(net19));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_20 (.L_LO(net20));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_21 (.L_LO(net21));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_22 (.L_LO(net22));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_23 (.L_LO(net23));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_24 (.L_LO(net24));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_25 (.L_LO(net25));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_26 (.L_LO(net26));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_27 (.L_LO(net27));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_28 (.L_LO(net28));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_29 (.L_LO(net29));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_30 (.L_LO(net30));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_31 (.L_LO(net31));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_32 (.L_LO(net32));
 sg13g2_tiehi _7392__33 (.L_HI(net33));
 sg13g2_buf_1 _7779_ (.A(\i_vga.timing_ver.sync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _7780_ (.A(\i_vga.hsync ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(net738));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(net734));
 sg13g2_buf_2 fanout734 (.A(net737),
    .X(net734));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(net736));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(net737));
 sg13g2_buf_2 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_1909_),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(net740));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(_0177_));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(_2780_));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(_2632_));
 sg13g2_buf_2 fanout743 (.A(_2632_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net746),
    .X(net744));
 sg13g2_buf_1 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net749),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(net749),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_1566_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(net751),
    .X(net750));
 sg13g2_buf_4 fanout751 (.X(net751),
    .A(net753));
 sg13g2_buf_2 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(_1565_));
 sg13g2_buf_2 fanout754 (.A(_3269_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_1413_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_1413_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(net760),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(net760),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(net760),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(_3265_));
 sg13g2_buf_4 fanout762 (.X(net762),
    .A(net763));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(_3261_));
 sg13g2_buf_2 fanout764 (.A(net768),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(net768),
    .X(net765));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(net768));
 sg13g2_buf_1 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_3260_),
    .X(net768));
 sg13g2_buf_4 fanout769 (.X(net769),
    .A(net774));
 sg13g2_buf_2 fanout770 (.A(net774),
    .X(net770));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(net772));
 sg13g2_buf_2 fanout772 (.A(net774),
    .X(net772));
 sg13g2_buf_1 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_3251_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(net776),
    .X(net775));
 sg13g2_buf_1 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_1 fanout778 (.A(_3250_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(net781),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(net781),
    .X(net780));
 sg13g2_buf_1 fanout781 (.A(_3250_),
    .X(net781));
 sg13g2_buf_4 fanout782 (.X(net782),
    .A(net785));
 sg13g2_buf_2 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_3250_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_3354_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_3345_),
    .X(net787));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(net789));
 sg13g2_buf_2 fanout789 (.A(\i_coord.l_xip.genblk2[9].state.Q ),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_3331_),
    .X(net790));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(net792));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(_3264_));
 sg13g2_buf_2 fanout793 (.A(_3259_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_3259_),
    .X(net794));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(net797));
 sg13g2_buf_2 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_3259_),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(net799),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(net801),
    .X(net800));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(_3258_));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_3202_));
 sg13g2_buf_2 fanout803 (.A(\i_coord.l_yip.genblk2[9].state.Q ),
    .X(net803));
 sg13g2_buf_1 fanout804 (.A(\i_coord.l_yip.genblk2[9].state.Q ),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(\i_coord.l_xir.genblk2[7].state.Q ),
    .X(net805));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(\i_coord.l_xir.genblk2[7].state.Q ));
 sg13g2_buf_2 fanout807 (.A(_0187_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_0187_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_3420_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_1148_),
    .X(net810));
 sg13g2_buf_1 fanout811 (.A(_1148_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_1137_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_1 fanout814 (.A(_1136_),
    .X(net814));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(_0184_));
 sg13g2_buf_2 fanout816 (.A(net818),
    .X(net816));
 sg13g2_buf_1 fanout817 (.A(net818),
    .X(net817));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(net819));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(_3342_));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(net822));
 sg13g2_buf_1 fanout821 (.A(net822),
    .X(net821));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(_3323_));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(_3301_));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(_3286_));
 sg13g2_buf_1 fanout825 (.A(_3286_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_3284_),
    .X(net826));
 sg13g2_buf_1 fanout827 (.A(_3284_),
    .X(net827));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(_3278_));
 sg13g2_buf_1 fanout829 (.A(_3278_),
    .X(net829));
 sg13g2_buf_4 fanout830 (.X(net830),
    .A(_3272_));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_1 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net837),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(net837),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(net837),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_3238_),
    .X(net837));
 sg13g2_buf_4 fanout838 (.X(net838),
    .A(net841));
 sg13g2_buf_2 fanout839 (.A(net841),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(_3237_));
 sg13g2_buf_2 fanout842 (.A(net843),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(_3300_));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_4 fanout846 (.X(net846),
    .A(_3297_));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(net848));
 sg13g2_buf_4 fanout848 (.X(net848),
    .A(_3292_));
 sg13g2_buf_2 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_4 fanout850 (.X(net850),
    .A(net851));
 sg13g2_buf_2 fanout851 (.A(_3288_),
    .X(net851));
 sg13g2_buf_4 fanout852 (.X(net852),
    .A(_3287_));
 sg13g2_buf_2 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_3277_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_3276_),
    .X(net855));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(_3276_));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(net860));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(net860));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_3274_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(net862),
    .X(net861));
 sg13g2_buf_4 fanout862 (.X(net862),
    .A(net864));
 sg13g2_buf_1 fanout863 (.A(net864),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_4 fanout865 (.X(net865),
    .A(_3273_));
 sg13g2_buf_2 fanout866 (.A(_3239_),
    .X(net866));
 sg13g2_buf_1 fanout867 (.A(_3239_),
    .X(net867));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(_3152_));
 sg13g2_buf_2 fanout869 (.A(_3152_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(net872),
    .X(net870));
 sg13g2_buf_1 fanout871 (.A(net872),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_4 fanout873 (.X(net873),
    .A(net878));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net878),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net878),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_4 fanout878 (.X(net878),
    .A(_3151_));
 sg13g2_buf_2 fanout879 (.A(_3135_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_3095_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(\i_mandel.i_xy.y[1] ),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(\i_mandel.i_xy.y[1] ),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(net886),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(net340),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net889),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(\i_mandel.i_xy.y[-1] ),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net356),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(\i_mandel.i_xy.y[-2] ),
    .X(net891));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(net893));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net362));
 sg13g2_buf_4 fanout894 (.X(net894),
    .A(net896));
 sg13g2_buf_2 fanout895 (.A(net896),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net355),
    .X(net896));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(net898));
 sg13g2_buf_2 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(\i_mandel.i_xy.y[-5] ),
    .X(net899));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(net901));
 sg13g2_buf_2 fanout901 (.A(net902),
    .X(net901));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(\i_mandel.i_xy.y[-6] ));
 sg13g2_buf_4 fanout903 (.X(net903),
    .A(net904));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(net352));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(\i_mandel.i_xy.y[-8] ));
 sg13g2_buf_4 fanout906 (.X(net906),
    .A(net358));
 sg13g2_buf_2 fanout907 (.A(net354),
    .X(net907));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(\i_mandel.i_xy.y[-9] ));
 sg13g2_buf_2 fanout909 (.A(net910),
    .X(net909));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(\i_mandel.i_xy.x[2] ));
 sg13g2_buf_2 fanout911 (.A(net913),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(\i_mandel.i_xy.x[1] ));
 sg13g2_buf_2 fanout914 (.A(net915),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(\i_mandel.i_xy.x[0] ),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(\i_mandel.i_xy.x[-1] ),
    .X(net916));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(\i_mandel.i_xy.x[-1] ));
 sg13g2_buf_4 fanout918 (.X(net918),
    .A(net919));
 sg13g2_buf_4 fanout919 (.X(net919),
    .A(\i_mandel.i_xy.x[-2] ));
 sg13g2_buf_2 fanout920 (.A(net922),
    .X(net920));
 sg13g2_buf_1 fanout921 (.A(net922),
    .X(net921));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(net324));
 sg13g2_buf_2 fanout923 (.A(net925),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(net344),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(\i_mandel.i_xy.x[-5] ),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(net929),
    .X(net928));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(\i_mandel.i_xy.x[-6] ));
 sg13g2_buf_2 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(\i_mandel.i_xy.x[-7] ),
    .X(net931));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(net934));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(net327),
    .X(net934));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(net936));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(net330));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(\i_coord.y0[-8] ));
 sg13g2_buf_2 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(\i_coord.demo_update ));
 sg13g2_buf_2 fanout941 (.A(net328),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(net943),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(net944),
    .X(net943));
 sg13g2_buf_1 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(net359),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(net360),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(net948),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(net273),
    .X(net948));
 sg13g2_buf_4 fanout949 (.X(net949),
    .A(net957));
 sg13g2_buf_2 fanout950 (.A(net957),
    .X(net950));
 sg13g2_buf_1 fanout951 (.A(net957),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(net954),
    .X(net952));
 sg13g2_buf_1 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(net955),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(net957),
    .X(net956));
 sg13g2_buf_4 fanout957 (.X(net957),
    .A(\i_mandel.i_xy.phase ));
 sg13g2_buf_2 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_4 fanout960 (.X(net960),
    .A(_3115_));
 sg13g2_buf_2 fanout961 (.A(net963),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net963),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(rst_n),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(net966),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(rst_n),
    .X(net967));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_2 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_2 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_4 input16 (.X(net16),
    .A(uio_in[7]));
 sg13g2_tielo tt_um_MichaelBell_mandelbrot_17 (.L_LO(net17));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_5_21__leaf_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk_regs));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_inv_1 clkload13 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_2 \clkbuf_0_i_mandel.i_xy.hc.gated_clk  (.A(\i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_0_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_3_0__f_i_mandel.i_xy.hc.gated_clk  (.A(\clknet_0_i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_3_0__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_3_1__f_i_mandel.i_xy.hc.gated_clk  (.A(\clknet_0_i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_3_1__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_3_2__f_i_mandel.i_xy.hc.gated_clk  (.A(\clknet_0_i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_3_2__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_3_3__f_i_mandel.i_xy.hc.gated_clk  (.A(\clknet_0_i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_3_3__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_3_4__f_i_mandel.i_xy.hc.gated_clk  (.A(\clknet_0_i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_3_4__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_3_5__f_i_mandel.i_xy.hc.gated_clk  (.A(\clknet_0_i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_3_5__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_3_6__f_i_mandel.i_xy.hc.gated_clk  (.A(\clknet_0_i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_3_6__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_3_7__f_i_mandel.i_xy.hc.gated_clk  (.A(\clknet_0_i_mandel.i_xy.hc.gated_clk ),
    .X(\clknet_3_7__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_inv_1 clkload14 (.A(\clknet_3_7__leaf_i_mandel.i_xy.hc.gated_clk ));
 sg13g2_buf_2 \clkbuf_0_i_coord.l_xl.gated_clk  (.A(\i_coord.l_xl.gated_clk ),
    .X(\clknet_0_i_coord.l_xl.gated_clk ));
 sg13g2_buf_2 \clkbuf_1_0__f_i_coord.l_xl.gated_clk  (.A(\clknet_0_i_coord.l_xl.gated_clk ),
    .X(\clknet_1_0__leaf_i_coord.l_xl.gated_clk ));
 sg13g2_buf_2 \clkbuf_1_1__f_i_coord.l_xl.gated_clk  (.A(\clknet_0_i_coord.l_xl.gated_clk ),
    .X(\clknet_1_1__leaf_i_coord.l_xl.gated_clk ));
 sg13g2_inv_1 clkload15 (.A(\clknet_1_1__leaf_i_coord.l_xl.gated_clk ));
 sg13g2_buf_2 \clkbuf_0_i_coord.l_yt.gated_clk  (.A(\i_coord.l_yt.gated_clk ),
    .X(\clknet_0_i_coord.l_yt.gated_clk ));
 sg13g2_buf_2 \clkbuf_2_0__f_i_coord.l_yt.gated_clk  (.A(\clknet_0_i_coord.l_yt.gated_clk ),
    .X(\clknet_2_0__leaf_i_coord.l_yt.gated_clk ));
 sg13g2_buf_2 \clkbuf_2_1__f_i_coord.l_yt.gated_clk  (.A(\clknet_0_i_coord.l_yt.gated_clk ),
    .X(\clknet_2_1__leaf_i_coord.l_yt.gated_clk ));
 sg13g2_buf_2 \clkbuf_2_2__f_i_coord.l_yt.gated_clk  (.A(\clknet_0_i_coord.l_yt.gated_clk ),
    .X(\clknet_2_2__leaf_i_coord.l_yt.gated_clk ));
 sg13g2_buf_2 \clkbuf_2_3__f_i_coord.l_yt.gated_clk  (.A(\clknet_0_i_coord.l_yt.gated_clk ),
    .X(\clknet_2_3__leaf_i_coord.l_yt.gated_clk ));
 sg13g2_inv_1 clkload16 (.A(\clknet_2_3__leaf_i_coord.l_yt.gated_clk ));
 sg13g2_buf_2 \clkbuf_0_i_coord.l_xip.gated_clk  (.A(\i_coord.l_xip.gated_clk ),
    .X(\clknet_0_i_coord.l_xip.gated_clk ));
 sg13g2_buf_2 \clkbuf_1_0__f_i_coord.l_xip.gated_clk  (.A(\clknet_0_i_coord.l_xip.gated_clk ),
    .X(\clknet_1_0__leaf_i_coord.l_xip.gated_clk ));
 sg13g2_buf_2 \clkbuf_1_1__f_i_coord.l_xip.gated_clk  (.A(\clknet_0_i_coord.l_xip.gated_clk ),
    .X(\clknet_1_1__leaf_i_coord.l_xip.gated_clk ));
 sg13g2_buf_2 \clkbuf_0_i_coord.l_yip.gated_clk  (.A(\i_coord.l_yip.gated_clk ),
    .X(\clknet_0_i_coord.l_yip.gated_clk ));
 sg13g2_buf_2 \clkbuf_1_0__f_i_coord.l_yip.gated_clk  (.A(\clknet_0_i_coord.l_yip.gated_clk ),
    .X(\clknet_1_0__leaf_i_coord.l_yip.gated_clk ));
 sg13g2_buf_2 \clkbuf_1_1__f_i_coord.l_yip.gated_clk  (.A(\clknet_0_i_coord.l_yip.gated_clk ),
    .X(\clknet_1_1__leaf_i_coord.l_yip.gated_clk ));
 sg13g2_buf_2 \clkbuf_0_i_coord.l_xir.gated_clk  (.A(\i_coord.l_xir.gated_clk ),
    .X(\clknet_0_i_coord.l_xir.gated_clk ));
 sg13g2_buf_2 \clkbuf_1_0__f_i_coord.l_xir.gated_clk  (.A(\clknet_0_i_coord.l_xir.gated_clk ),
    .X(\clknet_1_0__leaf_i_coord.l_xir.gated_clk ));
 sg13g2_buf_2 \clkbuf_1_1__f_i_coord.l_xir.gated_clk  (.A(\clknet_0_i_coord.l_xir.gated_clk ),
    .X(\clknet_1_1__leaf_i_coord.l_xir.gated_clk ));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0031_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold2 (.A(\i_vga.timing_ver.sync_tmp ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0030_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0074_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_mandel.i_xy.hc.genblk1.genblk1.CG.GATE ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_mandel.i_xy.x[-10] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_mandel.i_xy.x[-11] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_mandel.i_xy.y[-12] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_mandel.i_xy.y[-10] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold10 (.A(\iter[3] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0149_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_mandel.i_xy.x[2] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold13 (.A(\iter[1] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold14 (.A(\step[3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold15 (.A(_1309_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0036_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_vga.timing_hor.counter[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold18 (.A(_1538_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0089_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_mandel.i_xy.x[-12] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_mandel.i_xy.y[-13] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0150_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_mandel.i_xy.y[-11] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_mandel.i_xy.x[-13] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_vga.timing_ver.counter[9] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold26 (.A(\iter[0] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_coord.x_row_start[-13] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_coord.y0[-8] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_vga.timing_ver.counter[1] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold30 (.A(_1521_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_coord.y_row_start[1] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_mandel.i_xy.x[-2] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold33 (.A(\iter[2] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0148_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold35 (.A(\step[1] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0034_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0029_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold38 (.A(_1534_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_coord.x_row_start[-6] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold40 (.A(\step[4] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold41 (.A(_1310_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_vga.timing_ver.counter[7] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold43 (.A(_1530_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0084_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_coord.demo_update_delay ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_coord.x_row_start[2] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0050_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold48 (.A(\step[2] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_coord.y0[-2] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0028_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold51 (.A(_1545_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold52 (.A(_1546_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_coord.y_row_start[-3] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_coord.y_row_start[-12] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0060_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_vga.timing_hor.counter[3] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0090_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_coord.x_row_start[-9] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_coord.x_row_start[-2] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_coord.x_row_start[-7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_coord.x0[-6] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_vga.timing_hor.counter[4] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_vga.timing_ver.counter[5] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold64 (.A(_1527_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_coord.y_row_start[-8] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_coord.y_row_start[-2] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold67 (.A(\i_coord.y0[-13] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_coord.x_row_start[-11] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_coord.y0[-3] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_coord.y_row_start[-7] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_coord.y0[-12] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_coord.x_row_start[1] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_coord.y_row_start[-6] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0066_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_vga.timing_hor.counter[7] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold76 (.A(_1553_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0094_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_coord.x_row_start[-3] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_coord.x_row_start[-10] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_coord.x_row_start[-4] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_coord.x0[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_vga.timing_ver.counter[8] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold83 (.A(_1533_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_coord.y_row_start[0] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0032_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_coord.x_row_start[-8] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_vga.timing_ver.counter[6] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_mandel.i_xy.x[-5] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_coord.x_row_start[-5] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_coord.x_row_start[0] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_coord.y_row_start[-4] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_coord.x_row_start[-12] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_coord.y0[-7] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_coord.y_inc_row[-13] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_mandel.i_xy.x[-7] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_coord.y_row_start[-1] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_coord.y_row_start[-13] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_coord.x0[-12] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_vga.timing_hor.counter[0] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold100 (.A(\i_coord.y_row_start[-5] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_vga.timing_hor.counter[1] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold102 (.A(\i_coord.x_row_start[-1] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_coord.y_row_start[-9] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0063_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_vga.timing_ver.counter[4] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold106 (.A(_1526_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_mandel.i_xy.x[0] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_coord.x0[-9] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_coord.y0[1] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_coord.x0[-10] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_vga.timing_hor.counter[10] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold112 (.A(_1562_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_coord.y_row_start[-11] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0061_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_coord.x0[-13] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_vga.timing_hor.counter[9] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold117 (.A(_1559_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_coord.x0[1] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_coord.y_row_start[-10] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0005_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold121 (.A(\i_coord.x0[-11] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_coord.x0[-5] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_coord.x0[0] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_coord.x0[-7] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_coord.y0[-10] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_vga.timing_hor.counter[8] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_coord.x0[-8] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_coord.y0[-1] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_coord.y_inc_row[-8] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_coord.y0[0] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_coord.x0[-3] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_coord.x0[-2] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_coord.x0[-4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_coord.x0[-1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_coord.y0[-5] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_vga.timing_ver.counter[0] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold137 (.A(_1520_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0077_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold140 (.A(net902),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold142 (.A(net929),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_vga.timing_ver.counter[2] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0079_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_mandel.i_xy.x[-3] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_coord.y0[-11] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_coord.y_inc_row[-10] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_mandel.i_xy.x[-8] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_vga.timing_hor.counter[6] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0093_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_mandel.i_xy.x[-9] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_vga.timing_ver.counter[3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold153 (.A(_1525_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0026_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_coord.l_yt.genblk2[0].state.D ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0025_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_coord.l_yt.genblk2[1].state.D ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold159 (.A(net899),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_coord.y_inc_row[-9] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_mandel.i_xy.y[0] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_coord.y0[-6] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold163 (.A(\last_iter[1] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_coord.y_inc_row[-7] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_mandel.i_xy.x[-4] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_coord.y_inc_row[-11] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold168 (.A(net916),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0006_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_coord.y0[-4] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold171 (.A(\last_iter[3] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0000_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_mandel.i_xy.y[-7] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold174 (.A(\last_iter[2] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_mandel.i_xy.y[-9] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_mandel.i_xy.y[-4] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_mandel.i_xy.y[-2] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold178 (.A(\last_iter[0] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_mandel.i_xy.y[-8] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold180 (.A(\i_coord.y_inc_row[-6] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_coord.y_inc_row[-12] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_coord.y0[-9] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_mandel.i_xy.y[-3] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0021_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_vga.timing_ver.counter[4] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_vga.timing_ver.counter[3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_vga.timing_hor.counter[0] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold188 (.A(\iter[0] ),
    .X(net367));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_4 FILLER_23_546 ();
 sg13g2_fill_1 FILLER_23_550 ();
 sg13g2_decap_8 FILLER_23_554 ();
 sg13g2_decap_8 FILLER_23_561 ();
 sg13g2_decap_8 FILLER_23_568 ();
 sg13g2_decap_8 FILLER_23_575 ();
 sg13g2_decap_8 FILLER_23_582 ();
 sg13g2_decap_8 FILLER_23_589 ();
 sg13g2_decap_8 FILLER_23_596 ();
 sg13g2_decap_8 FILLER_23_603 ();
 sg13g2_decap_8 FILLER_23_610 ();
 sg13g2_decap_8 FILLER_23_617 ();
 sg13g2_decap_8 FILLER_23_624 ();
 sg13g2_decap_8 FILLER_23_631 ();
 sg13g2_decap_8 FILLER_23_638 ();
 sg13g2_decap_8 FILLER_23_645 ();
 sg13g2_decap_8 FILLER_23_652 ();
 sg13g2_decap_8 FILLER_23_659 ();
 sg13g2_decap_8 FILLER_23_666 ();
 sg13g2_decap_8 FILLER_23_673 ();
 sg13g2_decap_8 FILLER_23_680 ();
 sg13g2_decap_8 FILLER_23_687 ();
 sg13g2_decap_8 FILLER_23_694 ();
 sg13g2_decap_8 FILLER_23_701 ();
 sg13g2_decap_8 FILLER_23_708 ();
 sg13g2_decap_8 FILLER_23_715 ();
 sg13g2_decap_8 FILLER_23_722 ();
 sg13g2_decap_8 FILLER_23_729 ();
 sg13g2_decap_8 FILLER_23_736 ();
 sg13g2_decap_8 FILLER_23_743 ();
 sg13g2_decap_8 FILLER_23_750 ();
 sg13g2_decap_8 FILLER_23_757 ();
 sg13g2_decap_8 FILLER_23_764 ();
 sg13g2_decap_8 FILLER_23_771 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_decap_8 FILLER_23_785 ();
 sg13g2_decap_8 FILLER_23_792 ();
 sg13g2_decap_8 FILLER_23_799 ();
 sg13g2_decap_8 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_813 ();
 sg13g2_decap_8 FILLER_23_820 ();
 sg13g2_decap_8 FILLER_23_827 ();
 sg13g2_decap_8 FILLER_23_834 ();
 sg13g2_decap_8 FILLER_23_841 ();
 sg13g2_decap_8 FILLER_23_848 ();
 sg13g2_decap_8 FILLER_23_855 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_51 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_4 FILLER_24_66 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_113 ();
 sg13g2_fill_1 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_fill_2 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_fill_2 FILLER_24_323 ();
 sg13g2_fill_1 FILLER_24_325 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_fill_2 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_fill_2 FILLER_24_385 ();
 sg13g2_fill_1 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_8 FILLER_24_425 ();
 sg13g2_decap_8 FILLER_24_432 ();
 sg13g2_decap_8 FILLER_24_439 ();
 sg13g2_decap_8 FILLER_24_446 ();
 sg13g2_fill_2 FILLER_24_453 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_8 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_477 ();
 sg13g2_decap_8 FILLER_24_494 ();
 sg13g2_fill_2 FILLER_24_501 ();
 sg13g2_fill_1 FILLER_24_503 ();
 sg13g2_fill_2 FILLER_24_508 ();
 sg13g2_fill_1 FILLER_24_510 ();
 sg13g2_fill_2 FILLER_24_515 ();
 sg13g2_decap_4 FILLER_24_525 ();
 sg13g2_fill_1 FILLER_24_529 ();
 sg13g2_decap_8 FILLER_24_534 ();
 sg13g2_decap_4 FILLER_24_541 ();
 sg13g2_fill_1 FILLER_24_545 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_decap_8 FILLER_24_571 ();
 sg13g2_decap_4 FILLER_24_578 ();
 sg13g2_fill_2 FILLER_24_582 ();
 sg13g2_decap_8 FILLER_24_594 ();
 sg13g2_decap_8 FILLER_24_601 ();
 sg13g2_decap_8 FILLER_24_608 ();
 sg13g2_decap_8 FILLER_24_615 ();
 sg13g2_decap_8 FILLER_24_622 ();
 sg13g2_decap_8 FILLER_24_629 ();
 sg13g2_decap_8 FILLER_24_636 ();
 sg13g2_decap_8 FILLER_24_643 ();
 sg13g2_decap_8 FILLER_24_650 ();
 sg13g2_decap_8 FILLER_24_657 ();
 sg13g2_decap_8 FILLER_24_664 ();
 sg13g2_decap_8 FILLER_24_671 ();
 sg13g2_decap_8 FILLER_24_678 ();
 sg13g2_decap_8 FILLER_24_685 ();
 sg13g2_decap_8 FILLER_24_692 ();
 sg13g2_decap_8 FILLER_24_699 ();
 sg13g2_decap_8 FILLER_24_706 ();
 sg13g2_decap_8 FILLER_24_713 ();
 sg13g2_decap_8 FILLER_24_720 ();
 sg13g2_decap_8 FILLER_24_727 ();
 sg13g2_decap_8 FILLER_24_734 ();
 sg13g2_decap_8 FILLER_24_741 ();
 sg13g2_decap_8 FILLER_24_748 ();
 sg13g2_decap_8 FILLER_24_755 ();
 sg13g2_decap_8 FILLER_24_762 ();
 sg13g2_decap_8 FILLER_24_769 ();
 sg13g2_decap_8 FILLER_24_776 ();
 sg13g2_decap_8 FILLER_24_783 ();
 sg13g2_decap_8 FILLER_24_790 ();
 sg13g2_decap_8 FILLER_24_797 ();
 sg13g2_decap_8 FILLER_24_804 ();
 sg13g2_decap_8 FILLER_24_811 ();
 sg13g2_decap_8 FILLER_24_818 ();
 sg13g2_decap_8 FILLER_24_825 ();
 sg13g2_decap_8 FILLER_24_832 ();
 sg13g2_decap_8 FILLER_24_839 ();
 sg13g2_decap_8 FILLER_24_846 ();
 sg13g2_decap_8 FILLER_24_853 ();
 sg13g2_fill_2 FILLER_24_860 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_4 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_30 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_decap_8 FILLER_25_80 ();
 sg13g2_fill_2 FILLER_25_104 ();
 sg13g2_decap_4 FILLER_25_122 ();
 sg13g2_fill_2 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_141 ();
 sg13g2_decap_8 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_178 ();
 sg13g2_decap_8 FILLER_25_185 ();
 sg13g2_decap_8 FILLER_25_192 ();
 sg13g2_decap_8 FILLER_25_199 ();
 sg13g2_decap_8 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_decap_8 FILLER_25_220 ();
 sg13g2_decap_8 FILLER_25_227 ();
 sg13g2_decap_8 FILLER_25_234 ();
 sg13g2_decap_8 FILLER_25_241 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_decap_4 FILLER_25_255 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_decap_4 FILLER_25_268 ();
 sg13g2_decap_4 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_decap_4 FILLER_25_309 ();
 sg13g2_decap_4 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_decap_4 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_fill_1 FILLER_25_445 ();
 sg13g2_fill_2 FILLER_25_456 ();
 sg13g2_fill_1 FILLER_25_458 ();
 sg13g2_fill_1 FILLER_25_474 ();
 sg13g2_fill_2 FILLER_25_499 ();
 sg13g2_fill_2 FILLER_25_506 ();
 sg13g2_fill_1 FILLER_25_508 ();
 sg13g2_fill_2 FILLER_25_534 ();
 sg13g2_fill_2 FILLER_25_554 ();
 sg13g2_fill_1 FILLER_25_556 ();
 sg13g2_fill_2 FILLER_25_601 ();
 sg13g2_decap_8 FILLER_25_607 ();
 sg13g2_decap_8 FILLER_25_614 ();
 sg13g2_decap_8 FILLER_25_621 ();
 sg13g2_decap_8 FILLER_25_628 ();
 sg13g2_decap_8 FILLER_25_635 ();
 sg13g2_decap_8 FILLER_25_642 ();
 sg13g2_decap_8 FILLER_25_649 ();
 sg13g2_decap_8 FILLER_25_656 ();
 sg13g2_decap_8 FILLER_25_663 ();
 sg13g2_decap_8 FILLER_25_670 ();
 sg13g2_decap_8 FILLER_25_677 ();
 sg13g2_decap_8 FILLER_25_684 ();
 sg13g2_decap_8 FILLER_25_691 ();
 sg13g2_decap_8 FILLER_25_698 ();
 sg13g2_decap_8 FILLER_25_705 ();
 sg13g2_decap_8 FILLER_25_712 ();
 sg13g2_decap_8 FILLER_25_719 ();
 sg13g2_decap_8 FILLER_25_726 ();
 sg13g2_decap_8 FILLER_25_733 ();
 sg13g2_decap_8 FILLER_25_740 ();
 sg13g2_decap_8 FILLER_25_747 ();
 sg13g2_decap_8 FILLER_25_754 ();
 sg13g2_decap_8 FILLER_25_761 ();
 sg13g2_decap_8 FILLER_25_768 ();
 sg13g2_decap_8 FILLER_25_775 ();
 sg13g2_decap_8 FILLER_25_782 ();
 sg13g2_decap_8 FILLER_25_789 ();
 sg13g2_decap_8 FILLER_25_796 ();
 sg13g2_decap_8 FILLER_25_803 ();
 sg13g2_decap_8 FILLER_25_810 ();
 sg13g2_decap_8 FILLER_25_817 ();
 sg13g2_decap_8 FILLER_25_824 ();
 sg13g2_decap_8 FILLER_25_831 ();
 sg13g2_decap_8 FILLER_25_838 ();
 sg13g2_decap_8 FILLER_25_845 ();
 sg13g2_decap_8 FILLER_25_852 ();
 sg13g2_fill_2 FILLER_25_859 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_11 ();
 sg13g2_decap_4 FILLER_26_29 ();
 sg13g2_decap_4 FILLER_26_52 ();
 sg13g2_fill_2 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_decap_4 FILLER_26_76 ();
 sg13g2_fill_2 FILLER_26_80 ();
 sg13g2_decap_8 FILLER_26_106 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_decap_4 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_183 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_fill_2 FILLER_26_197 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_decap_4 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_decap_4 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_326 ();
 sg13g2_decap_4 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_366 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_fill_2 FILLER_26_400 ();
 sg13g2_decap_4 FILLER_26_428 ();
 sg13g2_fill_1 FILLER_26_432 ();
 sg13g2_decap_8 FILLER_26_438 ();
 sg13g2_decap_4 FILLER_26_445 ();
 sg13g2_fill_1 FILLER_26_449 ();
 sg13g2_fill_2 FILLER_26_464 ();
 sg13g2_decap_4 FILLER_26_476 ();
 sg13g2_fill_1 FILLER_26_480 ();
 sg13g2_decap_4 FILLER_26_491 ();
 sg13g2_fill_2 FILLER_26_495 ();
 sg13g2_fill_1 FILLER_26_501 ();
 sg13g2_fill_2 FILLER_26_519 ();
 sg13g2_fill_1 FILLER_26_521 ();
 sg13g2_fill_2 FILLER_26_536 ();
 sg13g2_fill_2 FILLER_26_552 ();
 sg13g2_fill_1 FILLER_26_554 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_4 FILLER_26_586 ();
 sg13g2_decap_8 FILLER_26_614 ();
 sg13g2_decap_8 FILLER_26_621 ();
 sg13g2_decap_8 FILLER_26_628 ();
 sg13g2_decap_8 FILLER_26_635 ();
 sg13g2_decap_8 FILLER_26_642 ();
 sg13g2_decap_8 FILLER_26_649 ();
 sg13g2_decap_8 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_decap_8 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_698 ();
 sg13g2_decap_8 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_712 ();
 sg13g2_decap_8 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_747 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_fill_2 FILLER_26_859 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_38 ();
 sg13g2_fill_2 FILLER_27_45 ();
 sg13g2_fill_1 FILLER_27_47 ();
 sg13g2_fill_2 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_79 ();
 sg13g2_decap_8 FILLER_27_96 ();
 sg13g2_decap_4 FILLER_27_103 ();
 sg13g2_decap_8 FILLER_27_134 ();
 sg13g2_decap_4 FILLER_27_141 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_223 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_decap_8 FILLER_27_244 ();
 sg13g2_decap_4 FILLER_27_251 ();
 sg13g2_decap_8 FILLER_27_268 ();
 sg13g2_fill_2 FILLER_27_275 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_decap_4 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_fill_2 FILLER_27_323 ();
 sg13g2_decap_4 FILLER_27_330 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_fill_2 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_1 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_27_417 ();
 sg13g2_fill_1 FILLER_27_424 ();
 sg13g2_fill_1 FILLER_27_444 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_fill_2 FILLER_27_475 ();
 sg13g2_decap_8 FILLER_27_507 ();
 sg13g2_decap_8 FILLER_27_514 ();
 sg13g2_fill_2 FILLER_27_521 ();
 sg13g2_fill_2 FILLER_27_531 ();
 sg13g2_decap_4 FILLER_27_541 ();
 sg13g2_fill_1 FILLER_27_545 ();
 sg13g2_fill_2 FILLER_27_563 ();
 sg13g2_fill_1 FILLER_27_565 ();
 sg13g2_decap_8 FILLER_27_578 ();
 sg13g2_fill_1 FILLER_27_585 ();
 sg13g2_fill_1 FILLER_27_598 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_20 ();
 sg13g2_fill_1 FILLER_28_33 ();
 sg13g2_decap_8 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_53 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_fill_1 FILLER_28_69 ();
 sg13g2_fill_2 FILLER_28_78 ();
 sg13g2_fill_1 FILLER_28_80 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_decap_8 FILLER_28_129 ();
 sg13g2_decap_4 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_fill_2 FILLER_28_190 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_decap_4 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_decap_4 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_decap_4 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_fill_2 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_fill_2 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_fill_2 FILLER_28_390 ();
 sg13g2_fill_2 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_411 ();
 sg13g2_fill_2 FILLER_28_418 ();
 sg13g2_decap_4 FILLER_28_428 ();
 sg13g2_fill_1 FILLER_28_432 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_fill_2 FILLER_28_448 ();
 sg13g2_fill_2 FILLER_28_464 ();
 sg13g2_fill_1 FILLER_28_466 ();
 sg13g2_decap_8 FILLER_28_472 ();
 sg13g2_decap_4 FILLER_28_479 ();
 sg13g2_fill_1 FILLER_28_483 ();
 sg13g2_fill_2 FILLER_28_488 ();
 sg13g2_fill_1 FILLER_28_517 ();
 sg13g2_decap_4 FILLER_28_537 ();
 sg13g2_fill_2 FILLER_28_552 ();
 sg13g2_fill_1 FILLER_28_554 ();
 sg13g2_decap_4 FILLER_28_568 ();
 sg13g2_fill_2 FILLER_28_590 ();
 sg13g2_fill_2 FILLER_28_605 ();
 sg13g2_fill_1 FILLER_28_607 ();
 sg13g2_decap_8 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_decap_8 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_20 ();
 sg13g2_decap_8 FILLER_29_51 ();
 sg13g2_fill_2 FILLER_29_58 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_decap_4 FILLER_29_101 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_187 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_263 ();
 sg13g2_decap_4 FILLER_29_270 ();
 sg13g2_fill_2 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_decap_4 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_4 FILLER_29_364 ();
 sg13g2_fill_1 FILLER_29_372 ();
 sg13g2_fill_2 FILLER_29_386 ();
 sg13g2_fill_1 FILLER_29_388 ();
 sg13g2_fill_2 FILLER_29_416 ();
 sg13g2_fill_1 FILLER_29_418 ();
 sg13g2_fill_2 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_452 ();
 sg13g2_fill_2 FILLER_29_459 ();
 sg13g2_decap_8 FILLER_29_506 ();
 sg13g2_decap_8 FILLER_29_513 ();
 sg13g2_decap_8 FILLER_29_540 ();
 sg13g2_fill_2 FILLER_29_547 ();
 sg13g2_fill_1 FILLER_29_549 ();
 sg13g2_fill_1 FILLER_29_563 ();
 sg13g2_fill_2 FILLER_29_585 ();
 sg13g2_fill_2 FILLER_29_599 ();
 sg13g2_fill_1 FILLER_29_601 ();
 sg13g2_decap_8 FILLER_29_618 ();
 sg13g2_decap_8 FILLER_29_625 ();
 sg13g2_decap_8 FILLER_29_632 ();
 sg13g2_decap_8 FILLER_29_639 ();
 sg13g2_decap_8 FILLER_29_646 ();
 sg13g2_decap_8 FILLER_29_653 ();
 sg13g2_decap_8 FILLER_29_660 ();
 sg13g2_decap_8 FILLER_29_667 ();
 sg13g2_decap_8 FILLER_29_674 ();
 sg13g2_decap_8 FILLER_29_681 ();
 sg13g2_decap_8 FILLER_29_688 ();
 sg13g2_decap_8 FILLER_29_695 ();
 sg13g2_decap_8 FILLER_29_702 ();
 sg13g2_decap_8 FILLER_29_709 ();
 sg13g2_decap_8 FILLER_29_716 ();
 sg13g2_decap_8 FILLER_29_723 ();
 sg13g2_decap_8 FILLER_29_730 ();
 sg13g2_decap_8 FILLER_29_737 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_decap_8 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_758 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_8 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_8 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_828 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_842 ();
 sg13g2_decap_8 FILLER_29_849 ();
 sg13g2_decap_4 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_41 ();
 sg13g2_fill_2 FILLER_30_48 ();
 sg13g2_decap_4 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_82 ();
 sg13g2_decap_4 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_106 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_fill_2 FILLER_30_120 ();
 sg13g2_decap_4 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_decap_4 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_216 ();
 sg13g2_fill_2 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_2 FILLER_30_319 ();
 sg13g2_fill_1 FILLER_30_321 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_376 ();
 sg13g2_decap_4 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_fill_2 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_458 ();
 sg13g2_decap_4 FILLER_30_465 ();
 sg13g2_fill_2 FILLER_30_469 ();
 sg13g2_decap_4 FILLER_30_476 ();
 sg13g2_fill_2 FILLER_30_480 ();
 sg13g2_fill_2 FILLER_30_493 ();
 sg13g2_fill_2 FILLER_30_507 ();
 sg13g2_decap_4 FILLER_30_521 ();
 sg13g2_fill_2 FILLER_30_525 ();
 sg13g2_fill_2 FILLER_30_539 ();
 sg13g2_fill_2 FILLER_30_546 ();
 sg13g2_fill_1 FILLER_30_548 ();
 sg13g2_decap_4 FILLER_30_554 ();
 sg13g2_decap_8 FILLER_30_571 ();
 sg13g2_decap_4 FILLER_30_590 ();
 sg13g2_fill_1 FILLER_30_594 ();
 sg13g2_decap_8 FILLER_30_600 ();
 sg13g2_decap_8 FILLER_30_607 ();
 sg13g2_decap_8 FILLER_30_614 ();
 sg13g2_decap_8 FILLER_30_621 ();
 sg13g2_decap_8 FILLER_30_628 ();
 sg13g2_decap_8 FILLER_30_635 ();
 sg13g2_decap_8 FILLER_30_642 ();
 sg13g2_decap_8 FILLER_30_649 ();
 sg13g2_decap_8 FILLER_30_656 ();
 sg13g2_decap_8 FILLER_30_663 ();
 sg13g2_decap_8 FILLER_30_670 ();
 sg13g2_decap_8 FILLER_30_677 ();
 sg13g2_decap_8 FILLER_30_684 ();
 sg13g2_decap_8 FILLER_30_691 ();
 sg13g2_decap_8 FILLER_30_698 ();
 sg13g2_decap_8 FILLER_30_705 ();
 sg13g2_decap_8 FILLER_30_712 ();
 sg13g2_decap_8 FILLER_30_719 ();
 sg13g2_decap_8 FILLER_30_726 ();
 sg13g2_decap_8 FILLER_30_733 ();
 sg13g2_decap_8 FILLER_30_740 ();
 sg13g2_decap_8 FILLER_30_747 ();
 sg13g2_decap_8 FILLER_30_754 ();
 sg13g2_decap_8 FILLER_30_761 ();
 sg13g2_decap_8 FILLER_30_768 ();
 sg13g2_decap_8 FILLER_30_775 ();
 sg13g2_decap_8 FILLER_30_782 ();
 sg13g2_decap_8 FILLER_30_789 ();
 sg13g2_decap_8 FILLER_30_796 ();
 sg13g2_decap_8 FILLER_30_803 ();
 sg13g2_decap_8 FILLER_30_810 ();
 sg13g2_decap_8 FILLER_30_817 ();
 sg13g2_decap_8 FILLER_30_824 ();
 sg13g2_decap_8 FILLER_30_831 ();
 sg13g2_decap_8 FILLER_30_838 ();
 sg13g2_decap_8 FILLER_30_845 ();
 sg13g2_decap_8 FILLER_30_852 ();
 sg13g2_fill_2 FILLER_30_859 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_44 ();
 sg13g2_fill_1 FILLER_31_46 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_decap_8 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_108 ();
 sg13g2_decap_4 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_137 ();
 sg13g2_decap_4 FILLER_31_144 ();
 sg13g2_fill_1 FILLER_31_148 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_4 FILLER_31_224 ();
 sg13g2_fill_2 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_250 ();
 sg13g2_decap_4 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_271 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_decap_4 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_decap_8 FILLER_31_328 ();
 sg13g2_fill_1 FILLER_31_335 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_fill_2 FILLER_31_363 ();
 sg13g2_fill_2 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_31_384 ();
 sg13g2_fill_2 FILLER_31_401 ();
 sg13g2_decap_4 FILLER_31_411 ();
 sg13g2_fill_1 FILLER_31_415 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_31_508 ();
 sg13g2_decap_4 FILLER_31_559 ();
 sg13g2_fill_2 FILLER_31_563 ();
 sg13g2_fill_2 FILLER_31_577 ();
 sg13g2_fill_1 FILLER_31_579 ();
 sg13g2_fill_2 FILLER_31_593 ();
 sg13g2_decap_8 FILLER_31_603 ();
 sg13g2_decap_8 FILLER_31_610 ();
 sg13g2_decap_8 FILLER_31_617 ();
 sg13g2_decap_4 FILLER_31_624 ();
 sg13g2_fill_2 FILLER_31_628 ();
 sg13g2_decap_8 FILLER_31_634 ();
 sg13g2_decap_8 FILLER_31_641 ();
 sg13g2_decap_8 FILLER_31_648 ();
 sg13g2_decap_8 FILLER_31_655 ();
 sg13g2_decap_8 FILLER_31_662 ();
 sg13g2_decap_8 FILLER_31_669 ();
 sg13g2_decap_4 FILLER_31_676 ();
 sg13g2_fill_2 FILLER_31_680 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_decap_4 FILLER_32_23 ();
 sg13g2_decap_4 FILLER_32_43 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_decap_4 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_fill_1 FILLER_32_90 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_decap_4 FILLER_32_175 ();
 sg13g2_fill_2 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_185 ();
 sg13g2_decap_4 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_decap_4 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_241 ();
 sg13g2_decap_4 FILLER_32_247 ();
 sg13g2_decap_4 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_decap_4 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_fill_2 FILLER_32_361 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_377 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_1 FILLER_32_426 ();
 sg13g2_fill_1 FILLER_32_431 ();
 sg13g2_decap_8 FILLER_32_436 ();
 sg13g2_fill_2 FILLER_32_443 ();
 sg13g2_fill_1 FILLER_32_445 ();
 sg13g2_decap_8 FILLER_32_452 ();
 sg13g2_decap_8 FILLER_32_459 ();
 sg13g2_decap_4 FILLER_32_466 ();
 sg13g2_fill_1 FILLER_32_470 ();
 sg13g2_decap_4 FILLER_32_475 ();
 sg13g2_fill_1 FILLER_32_487 ();
 sg13g2_decap_8 FILLER_32_509 ();
 sg13g2_fill_1 FILLER_32_516 ();
 sg13g2_decap_8 FILLER_32_537 ();
 sg13g2_fill_2 FILLER_32_544 ();
 sg13g2_decap_8 FILLER_32_556 ();
 sg13g2_decap_4 FILLER_32_563 ();
 sg13g2_fill_1 FILLER_32_567 ();
 sg13g2_decap_8 FILLER_32_585 ();
 sg13g2_fill_1 FILLER_32_592 ();
 sg13g2_decap_8 FILLER_32_610 ();
 sg13g2_decap_8 FILLER_32_642 ();
 sg13g2_decap_8 FILLER_32_649 ();
 sg13g2_decap_4 FILLER_32_656 ();
 sg13g2_decap_4 FILLER_32_665 ();
 sg13g2_fill_2 FILLER_32_669 ();
 sg13g2_decap_8 FILLER_32_696 ();
 sg13g2_decap_4 FILLER_32_703 ();
 sg13g2_fill_1 FILLER_32_707 ();
 sg13g2_fill_2 FILLER_32_713 ();
 sg13g2_decap_8 FILLER_32_723 ();
 sg13g2_decap_4 FILLER_32_730 ();
 sg13g2_fill_2 FILLER_32_734 ();
 sg13g2_decap_8 FILLER_32_741 ();
 sg13g2_fill_2 FILLER_32_748 ();
 sg13g2_fill_1 FILLER_32_750 ();
 sg13g2_decap_8 FILLER_32_776 ();
 sg13g2_decap_8 FILLER_32_783 ();
 sg13g2_decap_8 FILLER_32_790 ();
 sg13g2_decap_8 FILLER_32_797 ();
 sg13g2_decap_8 FILLER_32_804 ();
 sg13g2_decap_8 FILLER_32_811 ();
 sg13g2_decap_8 FILLER_32_818 ();
 sg13g2_decap_8 FILLER_32_825 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_839 ();
 sg13g2_decap_8 FILLER_32_846 ();
 sg13g2_decap_8 FILLER_32_853 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_31 ();
 sg13g2_fill_1 FILLER_33_38 ();
 sg13g2_decap_8 FILLER_33_44 ();
 sg13g2_fill_2 FILLER_33_51 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_86 ();
 sg13g2_decap_4 FILLER_33_107 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_260 ();
 sg13g2_decap_8 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_decap_4 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_decap_4 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_410 ();
 sg13g2_fill_1 FILLER_33_422 ();
 sg13g2_decap_8 FILLER_33_450 ();
 sg13g2_fill_2 FILLER_33_457 ();
 sg13g2_fill_1 FILLER_33_468 ();
 sg13g2_fill_1 FILLER_33_484 ();
 sg13g2_fill_2 FILLER_33_498 ();
 sg13g2_fill_1 FILLER_33_515 ();
 sg13g2_decap_4 FILLER_33_538 ();
 sg13g2_fill_1 FILLER_33_542 ();
 sg13g2_decap_8 FILLER_33_561 ();
 sg13g2_fill_2 FILLER_33_568 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_fill_2 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_fill_1 FILLER_33_623 ();
 sg13g2_decap_4 FILLER_33_649 ();
 sg13g2_fill_1 FILLER_33_653 ();
 sg13g2_fill_2 FILLER_33_700 ();
 sg13g2_decap_4 FILLER_33_726 ();
 sg13g2_fill_1 FILLER_33_730 ();
 sg13g2_decap_8 FILLER_33_747 ();
 sg13g2_fill_1 FILLER_33_754 ();
 sg13g2_decap_8 FILLER_33_764 ();
 sg13g2_decap_8 FILLER_33_771 ();
 sg13g2_decap_4 FILLER_33_778 ();
 sg13g2_fill_2 FILLER_33_782 ();
 sg13g2_decap_8 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_16 ();
 sg13g2_decap_4 FILLER_34_30 ();
 sg13g2_decap_8 FILLER_34_55 ();
 sg13g2_decap_4 FILLER_34_72 ();
 sg13g2_fill_2 FILLER_34_76 ();
 sg13g2_decap_8 FILLER_34_97 ();
 sg13g2_decap_8 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_177 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_decap_4 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_decap_4 FILLER_34_205 ();
 sg13g2_decap_4 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_fill_2 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_fill_1 FILLER_34_264 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_fill_1 FILLER_34_314 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_decap_4 FILLER_34_356 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_405 ();
 sg13g2_fill_2 FILLER_34_412 ();
 sg13g2_fill_2 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_482 ();
 sg13g2_fill_1 FILLER_34_489 ();
 sg13g2_decap_8 FILLER_34_495 ();
 sg13g2_fill_1 FILLER_34_502 ();
 sg13g2_decap_4 FILLER_34_513 ();
 sg13g2_fill_1 FILLER_34_517 ();
 sg13g2_decap_8 FILLER_34_535 ();
 sg13g2_fill_2 FILLER_34_542 ();
 sg13g2_fill_1 FILLER_34_544 ();
 sg13g2_decap_4 FILLER_34_570 ();
 sg13g2_decap_8 FILLER_34_584 ();
 sg13g2_fill_2 FILLER_34_591 ();
 sg13g2_fill_1 FILLER_34_593 ();
 sg13g2_decap_4 FILLER_34_614 ();
 sg13g2_decap_8 FILLER_34_643 ();
 sg13g2_decap_4 FILLER_34_650 ();
 sg13g2_fill_1 FILLER_34_654 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_4 FILLER_34_679 ();
 sg13g2_fill_1 FILLER_34_683 ();
 sg13g2_decap_8 FILLER_34_689 ();
 sg13g2_decap_8 FILLER_34_696 ();
 sg13g2_fill_2 FILLER_34_703 ();
 sg13g2_fill_1 FILLER_34_705 ();
 sg13g2_fill_1 FILLER_34_716 ();
 sg13g2_decap_8 FILLER_34_729 ();
 sg13g2_fill_1 FILLER_34_736 ();
 sg13g2_decap_4 FILLER_34_742 ();
 sg13g2_fill_2 FILLER_34_746 ();
 sg13g2_fill_1 FILLER_34_768 ();
 sg13g2_fill_1 FILLER_34_790 ();
 sg13g2_fill_1 FILLER_34_814 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_fill_2 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_62 ();
 sg13g2_decap_8 FILLER_35_69 ();
 sg13g2_decap_8 FILLER_35_76 ();
 sg13g2_decap_4 FILLER_35_83 ();
 sg13g2_decap_4 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_104 ();
 sg13g2_decap_8 FILLER_35_115 ();
 sg13g2_decap_8 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_180 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_decap_8 FILLER_35_209 ();
 sg13g2_decap_8 FILLER_35_216 ();
 sg13g2_fill_1 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_315 ();
 sg13g2_fill_1 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_2 FILLER_35_357 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_decap_4 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_4 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_410 ();
 sg13g2_decap_4 FILLER_35_416 ();
 sg13g2_fill_1 FILLER_35_420 ();
 sg13g2_decap_4 FILLER_35_431 ();
 sg13g2_fill_2 FILLER_35_435 ();
 sg13g2_decap_8 FILLER_35_442 ();
 sg13g2_decap_8 FILLER_35_449 ();
 sg13g2_fill_2 FILLER_35_456 ();
 sg13g2_fill_1 FILLER_35_458 ();
 sg13g2_decap_8 FILLER_35_468 ();
 sg13g2_decap_8 FILLER_35_475 ();
 sg13g2_fill_1 FILLER_35_482 ();
 sg13g2_fill_1 FILLER_35_499 ();
 sg13g2_decap_8 FILLER_35_508 ();
 sg13g2_decap_8 FILLER_35_515 ();
 sg13g2_decap_4 FILLER_35_522 ();
 sg13g2_decap_8 FILLER_35_531 ();
 sg13g2_fill_1 FILLER_35_538 ();
 sg13g2_fill_1 FILLER_35_556 ();
 sg13g2_decap_4 FILLER_35_561 ();
 sg13g2_fill_2 FILLER_35_565 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_4 FILLER_35_620 ();
 sg13g2_decap_4 FILLER_35_640 ();
 sg13g2_fill_2 FILLER_35_644 ();
 sg13g2_fill_1 FILLER_35_675 ();
 sg13g2_decap_8 FILLER_35_697 ();
 sg13g2_decap_4 FILLER_35_726 ();
 sg13g2_fill_2 FILLER_35_730 ();
 sg13g2_decap_8 FILLER_35_765 ();
 sg13g2_decap_4 FILLER_35_772 ();
 sg13g2_fill_1 FILLER_35_795 ();
 sg13g2_fill_2 FILLER_35_801 ();
 sg13g2_fill_1 FILLER_35_803 ();
 sg13g2_fill_1 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_834 ();
 sg13g2_decap_8 FILLER_35_841 ();
 sg13g2_decap_8 FILLER_35_848 ();
 sg13g2_decap_8 FILLER_35_855 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_16 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_25 ();
 sg13g2_decap_8 FILLER_36_39 ();
 sg13g2_fill_2 FILLER_36_46 ();
 sg13g2_fill_2 FILLER_36_64 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_180 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_decap_4 FILLER_36_201 ();
 sg13g2_fill_2 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_decap_4 FILLER_36_226 ();
 sg13g2_decap_4 FILLER_36_234 ();
 sg13g2_decap_4 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_decap_4 FILLER_36_326 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_decap_4 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_1 FILLER_36_407 ();
 sg13g2_fill_2 FILLER_36_441 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_fill_2 FILLER_36_474 ();
 sg13g2_fill_1 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_502 ();
 sg13g2_decap_4 FILLER_36_509 ();
 sg13g2_fill_1 FILLER_36_517 ();
 sg13g2_fill_2 FILLER_36_526 ();
 sg13g2_fill_2 FILLER_36_536 ();
 sg13g2_fill_1 FILLER_36_538 ();
 sg13g2_decap_8 FILLER_36_563 ();
 sg13g2_decap_4 FILLER_36_591 ();
 sg13g2_fill_2 FILLER_36_612 ();
 sg13g2_decap_4 FILLER_36_624 ();
 sg13g2_decap_4 FILLER_36_653 ();
 sg13g2_decap_4 FILLER_36_681 ();
 sg13g2_fill_1 FILLER_36_701 ();
 sg13g2_fill_2 FILLER_36_720 ();
 sg13g2_fill_2 FILLER_36_726 ();
 sg13g2_decap_4 FILLER_36_750 ();
 sg13g2_decap_8 FILLER_36_759 ();
 sg13g2_fill_2 FILLER_36_766 ();
 sg13g2_fill_1 FILLER_36_768 ();
 sg13g2_fill_2 FILLER_36_777 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_fill_2 FILLER_36_803 ();
 sg13g2_fill_1 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_811 ();
 sg13g2_decap_4 FILLER_36_818 ();
 sg13g2_fill_1 FILLER_36_822 ();
 sg13g2_decap_8 FILLER_36_841 ();
 sg13g2_decap_8 FILLER_36_848 ();
 sg13g2_decap_8 FILLER_36_855 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_53 ();
 sg13g2_decap_4 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_94 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_decap_4 FILLER_37_139 ();
 sg13g2_fill_2 FILLER_37_143 ();
 sg13g2_decap_4 FILLER_37_155 ();
 sg13g2_fill_1 FILLER_37_159 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_187 ();
 sg13g2_decap_4 FILLER_37_192 ();
 sg13g2_fill_2 FILLER_37_196 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_decap_4 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_257 ();
 sg13g2_decap_4 FILLER_37_271 ();
 sg13g2_fill_2 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_288 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_320 ();
 sg13g2_decap_4 FILLER_37_333 ();
 sg13g2_decap_4 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_4 FILLER_37_379 ();
 sg13g2_decap_4 FILLER_37_399 ();
 sg13g2_fill_1 FILLER_37_403 ();
 sg13g2_decap_8 FILLER_37_409 ();
 sg13g2_fill_2 FILLER_37_416 ();
 sg13g2_fill_1 FILLER_37_418 ();
 sg13g2_decap_8 FILLER_37_450 ();
 sg13g2_decap_8 FILLER_37_457 ();
 sg13g2_fill_2 FILLER_37_464 ();
 sg13g2_fill_1 FILLER_37_466 ();
 sg13g2_fill_1 FILLER_37_481 ();
 sg13g2_decap_4 FILLER_37_502 ();
 sg13g2_fill_1 FILLER_37_506 ();
 sg13g2_fill_2 FILLER_37_538 ();
 sg13g2_decap_4 FILLER_37_550 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_fill_1 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_579 ();
 sg13g2_decap_4 FILLER_37_586 ();
 sg13g2_fill_2 FILLER_37_590 ();
 sg13g2_decap_8 FILLER_37_608 ();
 sg13g2_fill_1 FILLER_37_615 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_fill_2 FILLER_37_651 ();
 sg13g2_decap_4 FILLER_37_682 ();
 sg13g2_fill_2 FILLER_37_696 ();
 sg13g2_decap_4 FILLER_37_707 ();
 sg13g2_fill_2 FILLER_37_711 ();
 sg13g2_fill_1 FILLER_37_730 ();
 sg13g2_fill_1 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_744 ();
 sg13g2_decap_4 FILLER_37_751 ();
 sg13g2_fill_1 FILLER_37_755 ();
 sg13g2_decap_4 FILLER_37_764 ();
 sg13g2_fill_1 FILLER_37_768 ();
 sg13g2_decap_4 FILLER_37_787 ();
 sg13g2_decap_8 FILLER_37_806 ();
 sg13g2_fill_1 FILLER_37_813 ();
 sg13g2_fill_2 FILLER_37_842 ();
 sg13g2_decap_8 FILLER_37_852 ();
 sg13g2_fill_2 FILLER_37_859 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_25 ();
 sg13g2_decap_4 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_71 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_decap_8 FILLER_38_93 ();
 sg13g2_fill_2 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_122 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_146 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_4 FILLER_38_186 ();
 sg13g2_decap_4 FILLER_38_202 ();
 sg13g2_fill_2 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_2 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_361 ();
 sg13g2_decap_4 FILLER_38_385 ();
 sg13g2_fill_1 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_403 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_440 ();
 sg13g2_fill_1 FILLER_38_447 ();
 sg13g2_decap_8 FILLER_38_461 ();
 sg13g2_decap_8 FILLER_38_468 ();
 sg13g2_fill_2 FILLER_38_475 ();
 sg13g2_fill_1 FILLER_38_477 ();
 sg13g2_fill_2 FILLER_38_498 ();
 sg13g2_decap_8 FILLER_38_537 ();
 sg13g2_fill_2 FILLER_38_544 ();
 sg13g2_fill_1 FILLER_38_546 ();
 sg13g2_decap_8 FILLER_38_557 ();
 sg13g2_fill_1 FILLER_38_564 ();
 sg13g2_decap_4 FILLER_38_577 ();
 sg13g2_fill_1 FILLER_38_581 ();
 sg13g2_decap_4 FILLER_38_611 ();
 sg13g2_fill_1 FILLER_38_615 ();
 sg13g2_fill_1 FILLER_38_620 ();
 sg13g2_decap_8 FILLER_38_635 ();
 sg13g2_decap_4 FILLER_38_642 ();
 sg13g2_fill_2 FILLER_38_646 ();
 sg13g2_fill_1 FILLER_38_653 ();
 sg13g2_fill_2 FILLER_38_658 ();
 sg13g2_fill_1 FILLER_38_660 ();
 sg13g2_decap_8 FILLER_38_673 ();
 sg13g2_fill_1 FILLER_38_680 ();
 sg13g2_fill_2 FILLER_38_687 ();
 sg13g2_fill_2 FILLER_38_693 ();
 sg13g2_fill_1 FILLER_38_695 ();
 sg13g2_fill_1 FILLER_38_712 ();
 sg13g2_decap_4 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_721 ();
 sg13g2_fill_1 FILLER_38_734 ();
 sg13g2_fill_2 FILLER_38_776 ();
 sg13g2_fill_2 FILLER_38_783 ();
 sg13g2_fill_1 FILLER_38_785 ();
 sg13g2_decap_4 FILLER_38_809 ();
 sg13g2_fill_1 FILLER_38_826 ();
 sg13g2_fill_2 FILLER_38_839 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_42 ();
 sg13g2_fill_1 FILLER_39_44 ();
 sg13g2_decap_8 FILLER_39_67 ();
 sg13g2_fill_1 FILLER_39_74 ();
 sg13g2_decap_8 FILLER_39_95 ();
 sg13g2_fill_2 FILLER_39_102 ();
 sg13g2_decap_8 FILLER_39_117 ();
 sg13g2_decap_8 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_131 ();
 sg13g2_decap_8 FILLER_39_143 ();
 sg13g2_fill_2 FILLER_39_183 ();
 sg13g2_fill_1 FILLER_39_185 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_fill_2 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_236 ();
 sg13g2_decap_4 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_247 ();
 sg13g2_decap_8 FILLER_39_265 ();
 sg13g2_fill_2 FILLER_39_272 ();
 sg13g2_decap_4 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_4 FILLER_39_355 ();
 sg13g2_fill_2 FILLER_39_359 ();
 sg13g2_decap_4 FILLER_39_369 ();
 sg13g2_fill_2 FILLER_39_373 ();
 sg13g2_decap_4 FILLER_39_383 ();
 sg13g2_fill_1 FILLER_39_387 ();
 sg13g2_fill_1 FILLER_39_393 ();
 sg13g2_fill_2 FILLER_39_408 ();
 sg13g2_decap_4 FILLER_39_422 ();
 sg13g2_fill_2 FILLER_39_448 ();
 sg13g2_fill_1 FILLER_39_450 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_decap_4 FILLER_39_477 ();
 sg13g2_fill_2 FILLER_39_481 ();
 sg13g2_decap_4 FILLER_39_516 ();
 sg13g2_fill_2 FILLER_39_520 ();
 sg13g2_decap_4 FILLER_39_541 ();
 sg13g2_fill_1 FILLER_39_553 ();
 sg13g2_decap_4 FILLER_39_584 ();
 sg13g2_fill_2 FILLER_39_609 ();
 sg13g2_fill_1 FILLER_39_611 ();
 sg13g2_fill_2 FILLER_39_632 ();
 sg13g2_fill_2 FILLER_39_660 ();
 sg13g2_fill_2 FILLER_39_667 ();
 sg13g2_decap_8 FILLER_39_673 ();
 sg13g2_fill_2 FILLER_39_680 ();
 sg13g2_fill_1 FILLER_39_682 ();
 sg13g2_fill_2 FILLER_39_695 ();
 sg13g2_fill_1 FILLER_39_697 ();
 sg13g2_decap_8 FILLER_39_706 ();
 sg13g2_decap_8 FILLER_39_713 ();
 sg13g2_decap_8 FILLER_39_720 ();
 sg13g2_fill_1 FILLER_39_727 ();
 sg13g2_fill_1 FILLER_39_732 ();
 sg13g2_fill_2 FILLER_39_737 ();
 sg13g2_fill_1 FILLER_39_743 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_fill_2 FILLER_39_756 ();
 sg13g2_fill_1 FILLER_39_758 ();
 sg13g2_fill_1 FILLER_39_763 ();
 sg13g2_fill_2 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_804 ();
 sg13g2_decap_4 FILLER_39_811 ();
 sg13g2_decap_8 FILLER_39_822 ();
 sg13g2_fill_2 FILLER_39_829 ();
 sg13g2_decap_4 FILLER_39_842 ();
 sg13g2_fill_2 FILLER_39_846 ();
 sg13g2_decap_8 FILLER_39_852 ();
 sg13g2_fill_2 FILLER_39_859 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_14 ();
 sg13g2_fill_2 FILLER_40_18 ();
 sg13g2_decap_4 FILLER_40_40 ();
 sg13g2_fill_1 FILLER_40_44 ();
 sg13g2_decap_8 FILLER_40_64 ();
 sg13g2_fill_1 FILLER_40_71 ();
 sg13g2_fill_1 FILLER_40_86 ();
 sg13g2_decap_4 FILLER_40_95 ();
 sg13g2_fill_2 FILLER_40_127 ();
 sg13g2_fill_1 FILLER_40_146 ();
 sg13g2_fill_2 FILLER_40_156 ();
 sg13g2_decap_8 FILLER_40_163 ();
 sg13g2_fill_2 FILLER_40_183 ();
 sg13g2_fill_2 FILLER_40_198 ();
 sg13g2_fill_1 FILLER_40_200 ();
 sg13g2_fill_2 FILLER_40_222 ();
 sg13g2_fill_2 FILLER_40_254 ();
 sg13g2_fill_1 FILLER_40_256 ();
 sg13g2_decap_8 FILLER_40_265 ();
 sg13g2_fill_2 FILLER_40_272 ();
 sg13g2_decap_8 FILLER_40_300 ();
 sg13g2_fill_2 FILLER_40_307 ();
 sg13g2_fill_1 FILLER_40_309 ();
 sg13g2_decap_8 FILLER_40_331 ();
 sg13g2_fill_2 FILLER_40_338 ();
 sg13g2_decap_8 FILLER_40_345 ();
 sg13g2_decap_8 FILLER_40_352 ();
 sg13g2_fill_2 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_decap_8 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_40_415 ();
 sg13g2_decap_8 FILLER_40_428 ();
 sg13g2_decap_8 FILLER_40_440 ();
 sg13g2_decap_8 FILLER_40_447 ();
 sg13g2_decap_4 FILLER_40_454 ();
 sg13g2_decap_4 FILLER_40_478 ();
 sg13g2_decap_8 FILLER_40_512 ();
 sg13g2_fill_2 FILLER_40_519 ();
 sg13g2_decap_8 FILLER_40_541 ();
 sg13g2_fill_1 FILLER_40_548 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_fill_2 FILLER_40_581 ();
 sg13g2_fill_1 FILLER_40_583 ();
 sg13g2_decap_8 FILLER_40_589 ();
 sg13g2_decap_8 FILLER_40_596 ();
 sg13g2_fill_1 FILLER_40_603 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_fill_1 FILLER_40_623 ();
 sg13g2_decap_4 FILLER_40_634 ();
 sg13g2_fill_2 FILLER_40_638 ();
 sg13g2_decap_4 FILLER_40_648 ();
 sg13g2_fill_1 FILLER_40_652 ();
 sg13g2_fill_2 FILLER_40_673 ();
 sg13g2_decap_8 FILLER_40_680 ();
 sg13g2_decap_4 FILLER_40_687 ();
 sg13g2_fill_2 FILLER_40_691 ();
 sg13g2_fill_1 FILLER_40_698 ();
 sg13g2_fill_2 FILLER_40_716 ();
 sg13g2_decap_8 FILLER_40_759 ();
 sg13g2_fill_2 FILLER_40_766 ();
 sg13g2_fill_1 FILLER_40_768 ();
 sg13g2_decap_8 FILLER_40_785 ();
 sg13g2_fill_2 FILLER_40_792 ();
 sg13g2_fill_1 FILLER_40_794 ();
 sg13g2_fill_1 FILLER_40_818 ();
 sg13g2_fill_1 FILLER_40_827 ();
 sg13g2_fill_2 FILLER_40_846 ();
 sg13g2_decap_8 FILLER_40_855 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_16 ();
 sg13g2_fill_2 FILLER_41_30 ();
 sg13g2_decap_4 FILLER_41_37 ();
 sg13g2_fill_2 FILLER_41_41 ();
 sg13g2_decap_8 FILLER_41_55 ();
 sg13g2_fill_2 FILLER_41_62 ();
 sg13g2_fill_1 FILLER_41_64 ();
 sg13g2_decap_4 FILLER_41_91 ();
 sg13g2_fill_1 FILLER_41_95 ();
 sg13g2_fill_2 FILLER_41_108 ();
 sg13g2_fill_1 FILLER_41_110 ();
 sg13g2_decap_8 FILLER_41_124 ();
 sg13g2_decap_4 FILLER_41_131 ();
 sg13g2_fill_2 FILLER_41_135 ();
 sg13g2_fill_2 FILLER_41_149 ();
 sg13g2_decap_8 FILLER_41_167 ();
 sg13g2_decap_4 FILLER_41_174 ();
 sg13g2_fill_2 FILLER_41_178 ();
 sg13g2_decap_8 FILLER_41_198 ();
 sg13g2_fill_2 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_225 ();
 sg13g2_fill_1 FILLER_41_232 ();
 sg13g2_decap_4 FILLER_41_254 ();
 sg13g2_fill_2 FILLER_41_258 ();
 sg13g2_fill_2 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_288 ();
 sg13g2_decap_8 FILLER_41_302 ();
 sg13g2_fill_1 FILLER_41_324 ();
 sg13g2_decap_8 FILLER_41_333 ();
 sg13g2_fill_1 FILLER_41_340 ();
 sg13g2_fill_1 FILLER_41_344 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_fill_1 FILLER_41_364 ();
 sg13g2_decap_4 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_385 ();
 sg13g2_decap_4 FILLER_41_391 ();
 sg13g2_fill_1 FILLER_41_395 ();
 sg13g2_fill_2 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_444 ();
 sg13g2_fill_2 FILLER_41_451 ();
 sg13g2_fill_1 FILLER_41_453 ();
 sg13g2_fill_2 FILLER_41_480 ();
 sg13g2_fill_1 FILLER_41_482 ();
 sg13g2_fill_2 FILLER_41_497 ();
 sg13g2_fill_1 FILLER_41_499 ();
 sg13g2_fill_1 FILLER_41_513 ();
 sg13g2_decap_8 FILLER_41_552 ();
 sg13g2_fill_2 FILLER_41_568 ();
 sg13g2_fill_1 FILLER_41_570 ();
 sg13g2_fill_2 FILLER_41_592 ();
 sg13g2_fill_1 FILLER_41_594 ();
 sg13g2_fill_1 FILLER_41_621 ();
 sg13g2_decap_8 FILLER_41_628 ();
 sg13g2_decap_8 FILLER_41_640 ();
 sg13g2_decap_8 FILLER_41_647 ();
 sg13g2_decap_8 FILLER_41_668 ();
 sg13g2_decap_4 FILLER_41_675 ();
 sg13g2_fill_1 FILLER_41_697 ();
 sg13g2_decap_8 FILLER_41_711 ();
 sg13g2_fill_1 FILLER_41_718 ();
 sg13g2_decap_8 FILLER_41_723 ();
 sg13g2_fill_2 FILLER_41_730 ();
 sg13g2_fill_1 FILLER_41_732 ();
 sg13g2_fill_2 FILLER_41_752 ();
 sg13g2_fill_2 FILLER_41_809 ();
 sg13g2_decap_4 FILLER_41_816 ();
 sg13g2_fill_1 FILLER_41_820 ();
 sg13g2_decap_4 FILLER_41_829 ();
 sg13g2_fill_1 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_837 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_4 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_25 ();
 sg13g2_fill_1 FILLER_42_39 ();
 sg13g2_decap_8 FILLER_42_52 ();
 sg13g2_decap_4 FILLER_42_59 ();
 sg13g2_decap_8 FILLER_42_81 ();
 sg13g2_decap_4 FILLER_42_92 ();
 sg13g2_fill_1 FILLER_42_96 ();
 sg13g2_decap_8 FILLER_42_110 ();
 sg13g2_fill_2 FILLER_42_117 ();
 sg13g2_fill_1 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_136 ();
 sg13g2_fill_2 FILLER_42_143 ();
 sg13g2_decap_4 FILLER_42_158 ();
 sg13g2_fill_2 FILLER_42_162 ();
 sg13g2_fill_2 FILLER_42_169 ();
 sg13g2_fill_1 FILLER_42_171 ();
 sg13g2_fill_2 FILLER_42_193 ();
 sg13g2_fill_1 FILLER_42_195 ();
 sg13g2_decap_8 FILLER_42_201 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_fill_2 FILLER_42_238 ();
 sg13g2_fill_1 FILLER_42_240 ();
 sg13g2_decap_8 FILLER_42_263 ();
 sg13g2_fill_2 FILLER_42_270 ();
 sg13g2_fill_1 FILLER_42_272 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_4 FILLER_42_301 ();
 sg13g2_fill_2 FILLER_42_305 ();
 sg13g2_fill_1 FILLER_42_334 ();
 sg13g2_fill_2 FILLER_42_360 ();
 sg13g2_decap_4 FILLER_42_389 ();
 sg13g2_fill_2 FILLER_42_393 ();
 sg13g2_fill_2 FILLER_42_400 ();
 sg13g2_fill_1 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_fill_2 FILLER_42_455 ();
 sg13g2_fill_1 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_479 ();
 sg13g2_decap_8 FILLER_42_492 ();
 sg13g2_fill_1 FILLER_42_499 ();
 sg13g2_decap_8 FILLER_42_525 ();
 sg13g2_fill_2 FILLER_42_532 ();
 sg13g2_fill_2 FILLER_42_546 ();
 sg13g2_decap_4 FILLER_42_571 ();
 sg13g2_fill_2 FILLER_42_575 ();
 sg13g2_decap_8 FILLER_42_591 ();
 sg13g2_decap_8 FILLER_42_615 ();
 sg13g2_decap_4 FILLER_42_622 ();
 sg13g2_fill_2 FILLER_42_651 ();
 sg13g2_decap_4 FILLER_42_674 ();
 sg13g2_fill_1 FILLER_42_678 ();
 sg13g2_fill_2 FILLER_42_683 ();
 sg13g2_fill_1 FILLER_42_689 ();
 sg13g2_fill_1 FILLER_42_706 ();
 sg13g2_fill_2 FILLER_42_729 ();
 sg13g2_fill_1 FILLER_42_731 ();
 sg13g2_fill_2 FILLER_42_751 ();
 sg13g2_fill_1 FILLER_42_753 ();
 sg13g2_decap_8 FILLER_42_774 ();
 sg13g2_decap_4 FILLER_42_781 ();
 sg13g2_fill_1 FILLER_42_785 ();
 sg13g2_decap_8 FILLER_42_801 ();
 sg13g2_fill_1 FILLER_42_808 ();
 sg13g2_fill_2 FILLER_42_813 ();
 sg13g2_fill_1 FILLER_42_827 ();
 sg13g2_decap_8 FILLER_42_844 ();
 sg13g2_decap_8 FILLER_42_851 ();
 sg13g2_decap_4 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_4 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_25 ();
 sg13g2_decap_4 FILLER_43_47 ();
 sg13g2_fill_2 FILLER_43_69 ();
 sg13g2_fill_1 FILLER_43_71 ();
 sg13g2_decap_4 FILLER_43_77 ();
 sg13g2_fill_1 FILLER_43_81 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_117 ();
 sg13g2_fill_2 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_141 ();
 sg13g2_decap_8 FILLER_43_151 ();
 sg13g2_fill_2 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_176 ();
 sg13g2_decap_8 FILLER_43_206 ();
 sg13g2_decap_4 FILLER_43_213 ();
 sg13g2_fill_2 FILLER_43_217 ();
 sg13g2_fill_1 FILLER_43_228 ();
 sg13g2_decap_8 FILLER_43_241 ();
 sg13g2_decap_4 FILLER_43_248 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_fill_2 FILLER_43_317 ();
 sg13g2_fill_1 FILLER_43_319 ();
 sg13g2_decap_4 FILLER_43_328 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_decap_8 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_43_415 ();
 sg13g2_fill_1 FILLER_43_422 ();
 sg13g2_fill_1 FILLER_43_441 ();
 sg13g2_fill_2 FILLER_43_457 ();
 sg13g2_fill_1 FILLER_43_473 ();
 sg13g2_decap_8 FILLER_43_502 ();
 sg13g2_decap_4 FILLER_43_518 ();
 sg13g2_fill_1 FILLER_43_522 ();
 sg13g2_decap_8 FILLER_43_527 ();
 sg13g2_fill_2 FILLER_43_534 ();
 sg13g2_fill_1 FILLER_43_536 ();
 sg13g2_decap_8 FILLER_43_547 ();
 sg13g2_fill_1 FILLER_43_554 ();
 sg13g2_fill_2 FILLER_43_603 ();
 sg13g2_fill_1 FILLER_43_646 ();
 sg13g2_decap_8 FILLER_43_659 ();
 sg13g2_decap_4 FILLER_43_666 ();
 sg13g2_fill_2 FILLER_43_670 ();
 sg13g2_fill_2 FILLER_43_684 ();
 sg13g2_decap_8 FILLER_43_702 ();
 sg13g2_fill_2 FILLER_43_709 ();
 sg13g2_fill_1 FILLER_43_711 ();
 sg13g2_fill_2 FILLER_43_738 ();
 sg13g2_fill_1 FILLER_43_740 ();
 sg13g2_decap_8 FILLER_43_746 ();
 sg13g2_fill_1 FILLER_43_753 ();
 sg13g2_fill_2 FILLER_43_759 ();
 sg13g2_fill_2 FILLER_43_766 ();
 sg13g2_fill_1 FILLER_43_768 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_792 ();
 sg13g2_fill_1 FILLER_43_799 ();
 sg13g2_fill_2 FILLER_43_826 ();
 sg13g2_fill_1 FILLER_43_832 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_fill_1 FILLER_43_845 ();
 sg13g2_fill_2 FILLER_43_859 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_4 FILLER_44_21 ();
 sg13g2_fill_1 FILLER_44_25 ();
 sg13g2_fill_1 FILLER_44_53 ();
 sg13g2_decap_8 FILLER_44_61 ();
 sg13g2_fill_2 FILLER_44_68 ();
 sg13g2_fill_2 FILLER_44_83 ();
 sg13g2_decap_8 FILLER_44_97 ();
 sg13g2_decap_8 FILLER_44_117 ();
 sg13g2_decap_4 FILLER_44_124 ();
 sg13g2_fill_2 FILLER_44_150 ();
 sg13g2_fill_1 FILLER_44_152 ();
 sg13g2_fill_1 FILLER_44_165 ();
 sg13g2_decap_4 FILLER_44_171 ();
 sg13g2_fill_1 FILLER_44_175 ();
 sg13g2_decap_4 FILLER_44_196 ();
 sg13g2_fill_2 FILLER_44_200 ();
 sg13g2_fill_1 FILLER_44_215 ();
 sg13g2_decap_4 FILLER_44_249 ();
 sg13g2_fill_2 FILLER_44_253 ();
 sg13g2_decap_8 FILLER_44_272 ();
 sg13g2_decap_8 FILLER_44_292 ();
 sg13g2_decap_8 FILLER_44_299 ();
 sg13g2_fill_1 FILLER_44_306 ();
 sg13g2_decap_4 FILLER_44_323 ();
 sg13g2_decap_4 FILLER_44_331 ();
 sg13g2_fill_2 FILLER_44_335 ();
 sg13g2_fill_1 FILLER_44_342 ();
 sg13g2_decap_4 FILLER_44_351 ();
 sg13g2_fill_2 FILLER_44_355 ();
 sg13g2_fill_2 FILLER_44_379 ();
 sg13g2_decap_4 FILLER_44_388 ();
 sg13g2_fill_2 FILLER_44_392 ();
 sg13g2_decap_4 FILLER_44_409 ();
 sg13g2_fill_2 FILLER_44_413 ();
 sg13g2_decap_4 FILLER_44_441 ();
 sg13g2_fill_2 FILLER_44_497 ();
 sg13g2_fill_2 FILLER_44_509 ();
 sg13g2_fill_1 FILLER_44_511 ();
 sg13g2_fill_2 FILLER_44_543 ();
 sg13g2_fill_2 FILLER_44_585 ();
 sg13g2_decap_4 FILLER_44_591 ();
 sg13g2_fill_1 FILLER_44_595 ();
 sg13g2_decap_4 FILLER_44_610 ();
 sg13g2_fill_2 FILLER_44_614 ();
 sg13g2_decap_8 FILLER_44_620 ();
 sg13g2_decap_4 FILLER_44_627 ();
 sg13g2_fill_1 FILLER_44_635 ();
 sg13g2_fill_2 FILLER_44_639 ();
 sg13g2_fill_1 FILLER_44_641 ();
 sg13g2_fill_2 FILLER_44_647 ();
 sg13g2_decap_8 FILLER_44_658 ();
 sg13g2_fill_2 FILLER_44_665 ();
 sg13g2_fill_1 FILLER_44_667 ();
 sg13g2_decap_8 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_711 ();
 sg13g2_fill_2 FILLER_44_718 ();
 sg13g2_fill_1 FILLER_44_720 ();
 sg13g2_fill_2 FILLER_44_743 ();
 sg13g2_fill_1 FILLER_44_745 ();
 sg13g2_fill_2 FILLER_44_778 ();
 sg13g2_fill_1 FILLER_44_780 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_fill_1 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_fill_2 FILLER_44_830 ();
 sg13g2_fill_1 FILLER_44_832 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_fill_2 FILLER_44_859 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_43 ();
 sg13g2_decap_4 FILLER_45_50 ();
 sg13g2_fill_2 FILLER_45_54 ();
 sg13g2_decap_8 FILLER_45_81 ();
 sg13g2_decap_4 FILLER_45_88 ();
 sg13g2_fill_2 FILLER_45_92 ();
 sg13g2_fill_1 FILLER_45_106 ();
 sg13g2_decap_8 FILLER_45_124 ();
 sg13g2_fill_1 FILLER_45_131 ();
 sg13g2_decap_8 FILLER_45_136 ();
 sg13g2_decap_4 FILLER_45_143 ();
 sg13g2_fill_2 FILLER_45_147 ();
 sg13g2_fill_1 FILLER_45_157 ();
 sg13g2_decap_8 FILLER_45_170 ();
 sg13g2_fill_1 FILLER_45_177 ();
 sg13g2_fill_2 FILLER_45_192 ();
 sg13g2_fill_1 FILLER_45_194 ();
 sg13g2_fill_2 FILLER_45_205 ();
 sg13g2_fill_1 FILLER_45_207 ();
 sg13g2_decap_8 FILLER_45_216 ();
 sg13g2_decap_4 FILLER_45_241 ();
 sg13g2_decap_4 FILLER_45_258 ();
 sg13g2_fill_2 FILLER_45_270 ();
 sg13g2_decap_4 FILLER_45_301 ();
 sg13g2_fill_1 FILLER_45_305 ();
 sg13g2_fill_2 FILLER_45_345 ();
 sg13g2_fill_1 FILLER_45_347 ();
 sg13g2_fill_1 FILLER_45_361 ();
 sg13g2_decap_4 FILLER_45_370 ();
 sg13g2_decap_4 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_405 ();
 sg13g2_decap_4 FILLER_45_410 ();
 sg13g2_fill_2 FILLER_45_414 ();
 sg13g2_fill_2 FILLER_45_420 ();
 sg13g2_fill_2 FILLER_45_435 ();
 sg13g2_fill_2 FILLER_45_441 ();
 sg13g2_fill_1 FILLER_45_443 ();
 sg13g2_fill_1 FILLER_45_449 ();
 sg13g2_decap_4 FILLER_45_477 ();
 sg13g2_fill_1 FILLER_45_481 ();
 sg13g2_fill_2 FILLER_45_492 ();
 sg13g2_fill_2 FILLER_45_512 ();
 sg13g2_fill_1 FILLER_45_522 ();
 sg13g2_fill_1 FILLER_45_537 ();
 sg13g2_fill_2 FILLER_45_571 ();
 sg13g2_fill_1 FILLER_45_573 ();
 sg13g2_fill_2 FILLER_45_600 ();
 sg13g2_fill_1 FILLER_45_664 ();
 sg13g2_decap_4 FILLER_45_681 ();
 sg13g2_fill_1 FILLER_45_685 ();
 sg13g2_decap_8 FILLER_45_691 ();
 sg13g2_fill_1 FILLER_45_702 ();
 sg13g2_fill_2 FILLER_45_716 ();
 sg13g2_decap_8 FILLER_45_724 ();
 sg13g2_decap_4 FILLER_45_748 ();
 sg13g2_fill_1 FILLER_45_752 ();
 sg13g2_decap_4 FILLER_45_768 ();
 sg13g2_fill_1 FILLER_45_772 ();
 sg13g2_fill_2 FILLER_45_777 ();
 sg13g2_fill_1 FILLER_45_779 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_fill_2 FILLER_45_845 ();
 sg13g2_fill_1 FILLER_45_847 ();
 sg13g2_decap_4 FILLER_45_856 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_fill_2 FILLER_46_35 ();
 sg13g2_fill_2 FILLER_46_66 ();
 sg13g2_decap_8 FILLER_46_86 ();
 sg13g2_fill_2 FILLER_46_108 ();
 sg13g2_fill_1 FILLER_46_110 ();
 sg13g2_decap_8 FILLER_46_141 ();
 sg13g2_fill_2 FILLER_46_148 ();
 sg13g2_decap_4 FILLER_46_179 ();
 sg13g2_fill_2 FILLER_46_192 ();
 sg13g2_fill_1 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_200 ();
 sg13g2_fill_2 FILLER_46_225 ();
 sg13g2_decap_8 FILLER_46_246 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_decap_4 FILLER_46_275 ();
 sg13g2_fill_2 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_293 ();
 sg13g2_fill_1 FILLER_46_295 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_4 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_321 ();
 sg13g2_fill_2 FILLER_46_328 ();
 sg13g2_fill_1 FILLER_46_330 ();
 sg13g2_decap_8 FILLER_46_351 ();
 sg13g2_fill_2 FILLER_46_358 ();
 sg13g2_fill_1 FILLER_46_360 ();
 sg13g2_decap_8 FILLER_46_374 ();
 sg13g2_fill_2 FILLER_46_381 ();
 sg13g2_fill_1 FILLER_46_388 ();
 sg13g2_fill_2 FILLER_46_446 ();
 sg13g2_fill_2 FILLER_46_474 ();
 sg13g2_fill_1 FILLER_46_476 ();
 sg13g2_decap_4 FILLER_46_589 ();
 sg13g2_fill_2 FILLER_46_593 ();
 sg13g2_decap_4 FILLER_46_598 ();
 sg13g2_fill_2 FILLER_46_602 ();
 sg13g2_fill_2 FILLER_46_616 ();
 sg13g2_decap_4 FILLER_46_622 ();
 sg13g2_decap_8 FILLER_46_643 ();
 sg13g2_decap_8 FILLER_46_650 ();
 sg13g2_fill_1 FILLER_46_657 ();
 sg13g2_decap_8 FILLER_46_662 ();
 sg13g2_fill_1 FILLER_46_669 ();
 sg13g2_decap_4 FILLER_46_682 ();
 sg13g2_fill_1 FILLER_46_686 ();
 sg13g2_decap_4 FILLER_46_695 ();
 sg13g2_decap_4 FILLER_46_720 ();
 sg13g2_decap_8 FILLER_46_750 ();
 sg13g2_decap_8 FILLER_46_757 ();
 sg13g2_decap_8 FILLER_46_764 ();
 sg13g2_fill_2 FILLER_46_771 ();
 sg13g2_fill_1 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_790 ();
 sg13g2_fill_2 FILLER_46_797 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_4 FILLER_46_829 ();
 sg13g2_fill_1 FILLER_46_833 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_4 FILLER_47_35 ();
 sg13g2_fill_2 FILLER_47_64 ();
 sg13g2_fill_2 FILLER_47_71 ();
 sg13g2_decap_8 FILLER_47_81 ();
 sg13g2_decap_4 FILLER_47_91 ();
 sg13g2_fill_1 FILLER_47_95 ();
 sg13g2_decap_8 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_141 ();
 sg13g2_decap_4 FILLER_47_176 ();
 sg13g2_fill_2 FILLER_47_195 ();
 sg13g2_fill_1 FILLER_47_202 ();
 sg13g2_fill_1 FILLER_47_222 ();
 sg13g2_decap_8 FILLER_47_242 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_decap_8 FILLER_47_254 ();
 sg13g2_fill_1 FILLER_47_261 ();
 sg13g2_decap_4 FILLER_47_267 ();
 sg13g2_decap_8 FILLER_47_274 ();
 sg13g2_decap_4 FILLER_47_281 ();
 sg13g2_fill_2 FILLER_47_285 ();
 sg13g2_decap_4 FILLER_47_304 ();
 sg13g2_fill_2 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_441 ();
 sg13g2_fill_2 FILLER_47_451 ();
 sg13g2_fill_1 FILLER_47_453 ();
 sg13g2_fill_2 FILLER_47_470 ();
 sg13g2_fill_1 FILLER_47_472 ();
 sg13g2_decap_8 FILLER_47_482 ();
 sg13g2_fill_2 FILLER_47_516 ();
 sg13g2_fill_1 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_531 ();
 sg13g2_fill_1 FILLER_47_548 ();
 sg13g2_decap_8 FILLER_47_562 ();
 sg13g2_fill_1 FILLER_47_569 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_fill_2 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_620 ();
 sg13g2_fill_2 FILLER_47_627 ();
 sg13g2_fill_1 FILLER_47_629 ();
 sg13g2_fill_2 FILLER_47_692 ();
 sg13g2_fill_1 FILLER_47_694 ();
 sg13g2_decap_4 FILLER_47_720 ();
 sg13g2_decap_4 FILLER_47_728 ();
 sg13g2_fill_2 FILLER_47_732 ();
 sg13g2_decap_8 FILLER_47_750 ();
 sg13g2_fill_2 FILLER_47_757 ();
 sg13g2_fill_1 FILLER_47_759 ();
 sg13g2_decap_4 FILLER_47_778 ();
 sg13g2_fill_1 FILLER_47_782 ();
 sg13g2_fill_1 FILLER_47_799 ();
 sg13g2_decap_8 FILLER_47_813 ();
 sg13g2_decap_8 FILLER_47_820 ();
 sg13g2_fill_2 FILLER_47_831 ();
 sg13g2_fill_1 FILLER_47_833 ();
 sg13g2_fill_2 FILLER_47_859 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_4 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_58 ();
 sg13g2_fill_2 FILLER_48_65 ();
 sg13g2_decap_4 FILLER_48_75 ();
 sg13g2_fill_1 FILLER_48_84 ();
 sg13g2_fill_1 FILLER_48_102 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_fill_1 FILLER_48_123 ();
 sg13g2_decap_8 FILLER_48_129 ();
 sg13g2_decap_8 FILLER_48_136 ();
 sg13g2_decap_8 FILLER_48_143 ();
 sg13g2_fill_2 FILLER_48_150 ();
 sg13g2_fill_1 FILLER_48_165 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_decap_4 FILLER_48_183 ();
 sg13g2_fill_1 FILLER_48_194 ();
 sg13g2_fill_2 FILLER_48_223 ();
 sg13g2_fill_2 FILLER_48_230 ();
 sg13g2_fill_1 FILLER_48_232 ();
 sg13g2_fill_2 FILLER_48_239 ();
 sg13g2_fill_1 FILLER_48_286 ();
 sg13g2_fill_2 FILLER_48_303 ();
 sg13g2_fill_2 FILLER_48_315 ();
 sg13g2_fill_1 FILLER_48_317 ();
 sg13g2_decap_8 FILLER_48_331 ();
 sg13g2_fill_2 FILLER_48_338 ();
 sg13g2_fill_1 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_346 ();
 sg13g2_fill_2 FILLER_48_351 ();
 sg13g2_fill_1 FILLER_48_356 ();
 sg13g2_fill_2 FILLER_48_362 ();
 sg13g2_fill_1 FILLER_48_364 ();
 sg13g2_decap_4 FILLER_48_369 ();
 sg13g2_fill_2 FILLER_48_378 ();
 sg13g2_fill_1 FILLER_48_380 ();
 sg13g2_fill_2 FILLER_48_396 ();
 sg13g2_fill_2 FILLER_48_495 ();
 sg13g2_decap_8 FILLER_48_531 ();
 sg13g2_decap_8 FILLER_48_538 ();
 sg13g2_fill_2 FILLER_48_545 ();
 sg13g2_decap_8 FILLER_48_565 ();
 sg13g2_fill_1 FILLER_48_572 ();
 sg13g2_decap_4 FILLER_48_599 ();
 sg13g2_fill_2 FILLER_48_620 ();
 sg13g2_fill_1 FILLER_48_622 ();
 sg13g2_fill_2 FILLER_48_635 ();
 sg13g2_decap_4 FILLER_48_641 ();
 sg13g2_fill_2 FILLER_48_645 ();
 sg13g2_fill_1 FILLER_48_651 ();
 sg13g2_fill_1 FILLER_48_658 ();
 sg13g2_fill_2 FILLER_48_664 ();
 sg13g2_fill_1 FILLER_48_666 ();
 sg13g2_decap_8 FILLER_48_690 ();
 sg13g2_decap_4 FILLER_48_697 ();
 sg13g2_decap_8 FILLER_48_713 ();
 sg13g2_decap_4 FILLER_48_720 ();
 sg13g2_fill_1 FILLER_48_724 ();
 sg13g2_fill_2 FILLER_48_735 ();
 sg13g2_fill_1 FILLER_48_737 ();
 sg13g2_decap_4 FILLER_48_743 ();
 sg13g2_fill_1 FILLER_48_747 ();
 sg13g2_fill_1 FILLER_48_784 ();
 sg13g2_fill_2 FILLER_48_791 ();
 sg13g2_fill_2 FILLER_48_806 ();
 sg13g2_fill_1 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_4 FILLER_48_856 ();
 sg13g2_fill_2 FILLER_48_860 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_44 ();
 sg13g2_fill_1 FILLER_49_58 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_107 ();
 sg13g2_decap_4 FILLER_49_114 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_fill_2 FILLER_49_141 ();
 sg13g2_fill_1 FILLER_49_143 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_fill_2 FILLER_49_200 ();
 sg13g2_fill_1 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_226 ();
 sg13g2_decap_4 FILLER_49_233 ();
 sg13g2_decap_8 FILLER_49_241 ();
 sg13g2_fill_2 FILLER_49_248 ();
 sg13g2_fill_1 FILLER_49_250 ();
 sg13g2_fill_2 FILLER_49_255 ();
 sg13g2_fill_1 FILLER_49_265 ();
 sg13g2_decap_8 FILLER_49_283 ();
 sg13g2_decap_8 FILLER_49_290 ();
 sg13g2_decap_8 FILLER_49_314 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_354 ();
 sg13g2_decap_4 FILLER_49_365 ();
 sg13g2_fill_2 FILLER_49_369 ();
 sg13g2_fill_2 FILLER_49_396 ();
 sg13g2_fill_2 FILLER_49_416 ();
 sg13g2_fill_1 FILLER_49_418 ();
 sg13g2_decap_4 FILLER_49_423 ();
 sg13g2_fill_2 FILLER_49_427 ();
 sg13g2_decap_4 FILLER_49_437 ();
 sg13g2_fill_2 FILLER_49_453 ();
 sg13g2_fill_1 FILLER_49_455 ();
 sg13g2_fill_2 FILLER_49_493 ();
 sg13g2_fill_1 FILLER_49_495 ();
 sg13g2_fill_2 FILLER_49_501 ();
 sg13g2_fill_1 FILLER_49_503 ();
 sg13g2_decap_4 FILLER_49_517 ();
 sg13g2_fill_1 FILLER_49_521 ();
 sg13g2_fill_1 FILLER_49_540 ();
 sg13g2_fill_1 FILLER_49_576 ();
 sg13g2_fill_2 FILLER_49_607 ();
 sg13g2_fill_1 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_619 ();
 sg13g2_decap_4 FILLER_49_626 ();
 sg13g2_fill_1 FILLER_49_630 ();
 sg13g2_decap_4 FILLER_49_635 ();
 sg13g2_fill_1 FILLER_49_664 ();
 sg13g2_decap_4 FILLER_49_674 ();
 sg13g2_decap_8 FILLER_49_697 ();
 sg13g2_fill_2 FILLER_49_704 ();
 sg13g2_fill_2 FILLER_49_725 ();
 sg13g2_fill_1 FILLER_49_727 ();
 sg13g2_decap_4 FILLER_49_753 ();
 sg13g2_decap_8 FILLER_49_765 ();
 sg13g2_decap_8 FILLER_49_772 ();
 sg13g2_fill_2 FILLER_49_798 ();
 sg13g2_fill_1 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_817 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_841 ();
 sg13g2_decap_8 FILLER_49_848 ();
 sg13g2_decap_8 FILLER_49_855 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_49 ();
 sg13g2_fill_2 FILLER_50_65 ();
 sg13g2_fill_1 FILLER_50_67 ();
 sg13g2_decap_4 FILLER_50_78 ();
 sg13g2_fill_2 FILLER_50_82 ();
 sg13g2_decap_4 FILLER_50_105 ();
 sg13g2_fill_2 FILLER_50_121 ();
 sg13g2_fill_1 FILLER_50_123 ();
 sg13g2_decap_8 FILLER_50_129 ();
 sg13g2_fill_1 FILLER_50_152 ();
 sg13g2_decap_4 FILLER_50_162 ();
 sg13g2_fill_1 FILLER_50_179 ();
 sg13g2_decap_8 FILLER_50_190 ();
 sg13g2_fill_2 FILLER_50_197 ();
 sg13g2_fill_2 FILLER_50_212 ();
 sg13g2_decap_8 FILLER_50_227 ();
 sg13g2_fill_2 FILLER_50_269 ();
 sg13g2_decap_8 FILLER_50_287 ();
 sg13g2_fill_2 FILLER_50_294 ();
 sg13g2_decap_4 FILLER_50_322 ();
 sg13g2_fill_2 FILLER_50_326 ();
 sg13g2_decap_4 FILLER_50_372 ();
 sg13g2_fill_2 FILLER_50_376 ();
 sg13g2_decap_8 FILLER_50_407 ();
 sg13g2_decap_4 FILLER_50_414 ();
 sg13g2_fill_2 FILLER_50_427 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_decap_8 FILLER_50_469 ();
 sg13g2_fill_2 FILLER_50_476 ();
 sg13g2_decap_4 FILLER_50_487 ();
 sg13g2_fill_2 FILLER_50_511 ();
 sg13g2_fill_1 FILLER_50_513 ();
 sg13g2_fill_2 FILLER_50_526 ();
 sg13g2_fill_2 FILLER_50_597 ();
 sg13g2_fill_2 FILLER_50_604 ();
 sg13g2_decap_4 FILLER_50_614 ();
 sg13g2_fill_1 FILLER_50_618 ();
 sg13g2_decap_4 FILLER_50_636 ();
 sg13g2_fill_1 FILLER_50_640 ();
 sg13g2_fill_1 FILLER_50_649 ();
 sg13g2_fill_1 FILLER_50_660 ();
 sg13g2_decap_4 FILLER_50_675 ();
 sg13g2_fill_1 FILLER_50_679 ();
 sg13g2_fill_2 FILLER_50_695 ();
 sg13g2_fill_1 FILLER_50_697 ();
 sg13g2_decap_8 FILLER_50_726 ();
 sg13g2_decap_8 FILLER_50_741 ();
 sg13g2_decap_4 FILLER_50_748 ();
 sg13g2_fill_2 FILLER_50_772 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_decap_8 FILLER_50_846 ();
 sg13g2_decap_8 FILLER_50_853 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_4 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_87 ();
 sg13g2_fill_1 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_103 ();
 sg13g2_decap_4 FILLER_51_138 ();
 sg13g2_decap_4 FILLER_51_173 ();
 sg13g2_decap_4 FILLER_51_194 ();
 sg13g2_fill_2 FILLER_51_198 ();
 sg13g2_decap_8 FILLER_51_217 ();
 sg13g2_fill_2 FILLER_51_224 ();
 sg13g2_decap_4 FILLER_51_241 ();
 sg13g2_fill_2 FILLER_51_249 ();
 sg13g2_fill_1 FILLER_51_251 ();
 sg13g2_decap_4 FILLER_51_257 ();
 sg13g2_fill_1 FILLER_51_271 ();
 sg13g2_decap_8 FILLER_51_279 ();
 sg13g2_decap_4 FILLER_51_286 ();
 sg13g2_fill_2 FILLER_51_290 ();
 sg13g2_decap_4 FILLER_51_300 ();
 sg13g2_fill_2 FILLER_51_304 ();
 sg13g2_decap_8 FILLER_51_314 ();
 sg13g2_decap_4 FILLER_51_334 ();
 sg13g2_fill_1 FILLER_51_346 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_decap_8 FILLER_51_364 ();
 sg13g2_decap_8 FILLER_51_371 ();
 sg13g2_decap_4 FILLER_51_378 ();
 sg13g2_fill_2 FILLER_51_382 ();
 sg13g2_fill_1 FILLER_51_389 ();
 sg13g2_fill_2 FILLER_51_418 ();
 sg13g2_fill_1 FILLER_51_432 ();
 sg13g2_fill_2 FILLER_51_438 ();
 sg13g2_fill_1 FILLER_51_440 ();
 sg13g2_decap_8 FILLER_51_454 ();
 sg13g2_fill_2 FILLER_51_461 ();
 sg13g2_decap_4 FILLER_51_484 ();
 sg13g2_fill_2 FILLER_51_513 ();
 sg13g2_decap_4 FILLER_51_539 ();
 sg13g2_decap_8 FILLER_51_552 ();
 sg13g2_decap_8 FILLER_51_559 ();
 sg13g2_decap_8 FILLER_51_566 ();
 sg13g2_fill_1 FILLER_51_616 ();
 sg13g2_decap_4 FILLER_51_638 ();
 sg13g2_fill_2 FILLER_51_642 ();
 sg13g2_decap_8 FILLER_51_662 ();
 sg13g2_decap_8 FILLER_51_669 ();
 sg13g2_fill_2 FILLER_51_676 ();
 sg13g2_fill_1 FILLER_51_678 ();
 sg13g2_fill_2 FILLER_51_703 ();
 sg13g2_fill_1 FILLER_51_705 ();
 sg13g2_decap_8 FILLER_51_717 ();
 sg13g2_decap_4 FILLER_51_724 ();
 sg13g2_fill_2 FILLER_51_748 ();
 sg13g2_decap_8 FILLER_51_767 ();
 sg13g2_decap_4 FILLER_51_774 ();
 sg13g2_decap_8 FILLER_51_795 ();
 sg13g2_fill_2 FILLER_51_802 ();
 sg13g2_fill_1 FILLER_51_804 ();
 sg13g2_decap_4 FILLER_51_810 ();
 sg13g2_fill_2 FILLER_51_838 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_fill_2 FILLER_52_49 ();
 sg13g2_decap_4 FILLER_52_54 ();
 sg13g2_fill_2 FILLER_52_58 ();
 sg13g2_fill_2 FILLER_52_68 ();
 sg13g2_decap_4 FILLER_52_88 ();
 sg13g2_fill_1 FILLER_52_104 ();
 sg13g2_fill_2 FILLER_52_110 ();
 sg13g2_fill_2 FILLER_52_117 ();
 sg13g2_fill_1 FILLER_52_119 ();
 sg13g2_fill_1 FILLER_52_124 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_fill_2 FILLER_52_154 ();
 sg13g2_fill_1 FILLER_52_156 ();
 sg13g2_decap_8 FILLER_52_171 ();
 sg13g2_fill_1 FILLER_52_178 ();
 sg13g2_decap_8 FILLER_52_194 ();
 sg13g2_fill_2 FILLER_52_201 ();
 sg13g2_decap_8 FILLER_52_207 ();
 sg13g2_fill_2 FILLER_52_218 ();
 sg13g2_decap_4 FILLER_52_238 ();
 sg13g2_decap_4 FILLER_52_283 ();
 sg13g2_decap_8 FILLER_52_305 ();
 sg13g2_fill_2 FILLER_52_312 ();
 sg13g2_fill_1 FILLER_52_314 ();
 sg13g2_fill_1 FILLER_52_319 ();
 sg13g2_fill_1 FILLER_52_355 ();
 sg13g2_decap_8 FILLER_52_393 ();
 sg13g2_decap_8 FILLER_52_400 ();
 sg13g2_fill_1 FILLER_52_407 ();
 sg13g2_decap_4 FILLER_52_416 ();
 sg13g2_fill_2 FILLER_52_433 ();
 sg13g2_decap_8 FILLER_52_448 ();
 sg13g2_fill_1 FILLER_52_455 ();
 sg13g2_decap_8 FILLER_52_461 ();
 sg13g2_decap_4 FILLER_52_468 ();
 sg13g2_fill_1 FILLER_52_482 ();
 sg13g2_fill_1 FILLER_52_505 ();
 sg13g2_fill_2 FILLER_52_514 ();
 sg13g2_fill_1 FILLER_52_516 ();
 sg13g2_decap_4 FILLER_52_522 ();
 sg13g2_fill_2 FILLER_52_551 ();
 sg13g2_fill_1 FILLER_52_579 ();
 sg13g2_decap_8 FILLER_52_589 ();
 sg13g2_decap_4 FILLER_52_596 ();
 sg13g2_decap_8 FILLER_52_608 ();
 sg13g2_decap_8 FILLER_52_615 ();
 sg13g2_fill_2 FILLER_52_622 ();
 sg13g2_fill_1 FILLER_52_624 ();
 sg13g2_decap_8 FILLER_52_633 ();
 sg13g2_fill_1 FILLER_52_640 ();
 sg13g2_fill_2 FILLER_52_648 ();
 sg13g2_fill_1 FILLER_52_650 ();
 sg13g2_decap_8 FILLER_52_664 ();
 sg13g2_fill_2 FILLER_52_671 ();
 sg13g2_decap_8 FILLER_52_690 ();
 sg13g2_decap_4 FILLER_52_697 ();
 sg13g2_decap_4 FILLER_52_721 ();
 sg13g2_fill_1 FILLER_52_725 ();
 sg13g2_decap_8 FILLER_52_750 ();
 sg13g2_decap_4 FILLER_52_757 ();
 sg13g2_fill_1 FILLER_52_761 ();
 sg13g2_decap_8 FILLER_52_770 ();
 sg13g2_fill_2 FILLER_52_777 ();
 sg13g2_fill_1 FILLER_52_779 ();
 sg13g2_decap_8 FILLER_52_798 ();
 sg13g2_fill_2 FILLER_52_805 ();
 sg13g2_fill_1 FILLER_52_807 ();
 sg13g2_fill_2 FILLER_52_813 ();
 sg13g2_fill_1 FILLER_52_815 ();
 sg13g2_decap_8 FILLER_52_823 ();
 sg13g2_decap_4 FILLER_52_830 ();
 sg13g2_decap_4 FILLER_52_839 ();
 sg13g2_decap_8 FILLER_52_851 ();
 sg13g2_decap_4 FILLER_52_858 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_59 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_4 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_95 ();
 sg13g2_fill_2 FILLER_53_109 ();
 sg13g2_fill_1 FILLER_53_111 ();
 sg13g2_fill_2 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_124 ();
 sg13g2_fill_2 FILLER_53_130 ();
 sg13g2_fill_1 FILLER_53_132 ();
 sg13g2_decap_8 FILLER_53_159 ();
 sg13g2_fill_2 FILLER_53_265 ();
 sg13g2_fill_2 FILLER_53_280 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_fill_2 FILLER_53_291 ();
 sg13g2_fill_1 FILLER_53_293 ();
 sg13g2_decap_8 FILLER_53_330 ();
 sg13g2_decap_8 FILLER_53_337 ();
 sg13g2_fill_1 FILLER_53_344 ();
 sg13g2_fill_1 FILLER_53_355 ();
 sg13g2_decap_8 FILLER_53_372 ();
 sg13g2_fill_1 FILLER_53_379 ();
 sg13g2_decap_4 FILLER_53_394 ();
 sg13g2_fill_1 FILLER_53_398 ();
 sg13g2_decap_4 FILLER_53_424 ();
 sg13g2_fill_2 FILLER_53_428 ();
 sg13g2_fill_2 FILLER_53_447 ();
 sg13g2_fill_2 FILLER_53_501 ();
 sg13g2_fill_1 FILLER_53_503 ();
 sg13g2_fill_1 FILLER_53_509 ();
 sg13g2_decap_8 FILLER_53_519 ();
 sg13g2_fill_2 FILLER_53_526 ();
 sg13g2_fill_1 FILLER_53_539 ();
 sg13g2_decap_4 FILLER_53_554 ();
 sg13g2_fill_1 FILLER_53_558 ();
 sg13g2_fill_1 FILLER_53_573 ();
 sg13g2_decap_4 FILLER_53_579 ();
 sg13g2_fill_2 FILLER_53_583 ();
 sg13g2_fill_1 FILLER_53_600 ();
 sg13g2_fill_1 FILLER_53_619 ();
 sg13g2_fill_1 FILLER_53_633 ();
 sg13g2_decap_4 FILLER_53_646 ();
 sg13g2_fill_2 FILLER_53_650 ();
 sg13g2_fill_1 FILLER_53_665 ();
 sg13g2_fill_2 FILLER_53_698 ();
 sg13g2_fill_1 FILLER_53_700 ();
 sg13g2_decap_8 FILLER_53_726 ();
 sg13g2_fill_2 FILLER_53_733 ();
 sg13g2_fill_1 FILLER_53_735 ();
 sg13g2_decap_4 FILLER_53_745 ();
 sg13g2_fill_2 FILLER_53_749 ();
 sg13g2_decap_4 FILLER_53_777 ();
 sg13g2_fill_2 FILLER_53_795 ();
 sg13g2_fill_1 FILLER_53_797 ();
 sg13g2_decap_8 FILLER_53_850 ();
 sg13g2_decap_4 FILLER_53_857 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_4 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_79 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_fill_2 FILLER_54_119 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_decap_4 FILLER_54_138 ();
 sg13g2_fill_1 FILLER_54_142 ();
 sg13g2_decap_8 FILLER_54_156 ();
 sg13g2_decap_8 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_190 ();
 sg13g2_decap_8 FILLER_54_201 ();
 sg13g2_decap_4 FILLER_54_208 ();
 sg13g2_fill_1 FILLER_54_242 ();
 sg13g2_fill_1 FILLER_54_272 ();
 sg13g2_decap_4 FILLER_54_277 ();
 sg13g2_decap_4 FILLER_54_286 ();
 sg13g2_fill_1 FILLER_54_290 ();
 sg13g2_decap_8 FILLER_54_300 ();
 sg13g2_decap_8 FILLER_54_307 ();
 sg13g2_decap_4 FILLER_54_328 ();
 sg13g2_fill_2 FILLER_54_332 ();
 sg13g2_decap_8 FILLER_54_338 ();
 sg13g2_fill_2 FILLER_54_397 ();
 sg13g2_decap_4 FILLER_54_429 ();
 sg13g2_fill_1 FILLER_54_433 ();
 sg13g2_decap_8 FILLER_54_449 ();
 sg13g2_decap_4 FILLER_54_456 ();
 sg13g2_fill_2 FILLER_54_464 ();
 sg13g2_fill_2 FILLER_54_469 ();
 sg13g2_decap_8 FILLER_54_474 ();
 sg13g2_fill_1 FILLER_54_485 ();
 sg13g2_fill_2 FILLER_54_525 ();
 sg13g2_fill_1 FILLER_54_550 ();
 sg13g2_decap_8 FILLER_54_559 ();
 sg13g2_decap_4 FILLER_54_566 ();
 sg13g2_fill_2 FILLER_54_570 ();
 sg13g2_fill_2 FILLER_54_602 ();
 sg13g2_fill_2 FILLER_54_617 ();
 sg13g2_fill_2 FILLER_54_632 ();
 sg13g2_fill_2 FILLER_54_653 ();
 sg13g2_decap_8 FILLER_54_667 ();
 sg13g2_fill_2 FILLER_54_674 ();
 sg13g2_fill_1 FILLER_54_676 ();
 sg13g2_decap_8 FILLER_54_693 ();
 sg13g2_fill_2 FILLER_54_700 ();
 sg13g2_fill_1 FILLER_54_702 ();
 sg13g2_decap_8 FILLER_54_719 ();
 sg13g2_fill_1 FILLER_54_726 ();
 sg13g2_fill_2 FILLER_54_747 ();
 sg13g2_fill_1 FILLER_54_757 ();
 sg13g2_decap_8 FILLER_54_798 ();
 sg13g2_fill_2 FILLER_54_814 ();
 sg13g2_fill_1 FILLER_54_816 ();
 sg13g2_decap_8 FILLER_54_822 ();
 sg13g2_decap_4 FILLER_54_829 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_decap_4 FILLER_54_856 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_fill_2 FILLER_55_49 ();
 sg13g2_fill_1 FILLER_55_82 ();
 sg13g2_decap_4 FILLER_55_109 ();
 sg13g2_fill_1 FILLER_55_113 ();
 sg13g2_fill_2 FILLER_55_129 ();
 sg13g2_fill_1 FILLER_55_131 ();
 sg13g2_fill_2 FILLER_55_184 ();
 sg13g2_decap_4 FILLER_55_220 ();
 sg13g2_fill_1 FILLER_55_242 ();
 sg13g2_decap_8 FILLER_55_349 ();
 sg13g2_fill_1 FILLER_55_356 ();
 sg13g2_fill_1 FILLER_55_366 ();
 sg13g2_fill_2 FILLER_55_377 ();
 sg13g2_fill_1 FILLER_55_379 ();
 sg13g2_decap_4 FILLER_55_424 ();
 sg13g2_fill_1 FILLER_55_428 ();
 sg13g2_fill_2 FILLER_55_469 ();
 sg13g2_fill_2 FILLER_55_508 ();
 sg13g2_fill_1 FILLER_55_514 ();
 sg13g2_decap_8 FILLER_55_524 ();
 sg13g2_decap_8 FILLER_55_531 ();
 sg13g2_decap_8 FILLER_55_538 ();
 sg13g2_fill_2 FILLER_55_545 ();
 sg13g2_fill_2 FILLER_55_569 ();
 sg13g2_fill_1 FILLER_55_571 ();
 sg13g2_fill_2 FILLER_55_581 ();
 sg13g2_decap_8 FILLER_55_602 ();
 sg13g2_decap_8 FILLER_55_630 ();
 sg13g2_fill_2 FILLER_55_637 ();
 sg13g2_decap_4 FILLER_55_644 ();
 sg13g2_fill_1 FILLER_55_648 ();
 sg13g2_fill_2 FILLER_55_670 ();
 sg13g2_decap_4 FILLER_55_701 ();
 sg13g2_fill_1 FILLER_55_705 ();
 sg13g2_decap_8 FILLER_55_723 ();
 sg13g2_fill_2 FILLER_55_730 ();
 sg13g2_decap_8 FILLER_55_748 ();
 sg13g2_fill_2 FILLER_55_755 ();
 sg13g2_fill_1 FILLER_55_757 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_4 FILLER_55_777 ();
 sg13g2_fill_2 FILLER_55_781 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_fill_1 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_820 ();
 sg13g2_decap_8 FILLER_55_827 ();
 sg13g2_decap_8 FILLER_55_846 ();
 sg13g2_decap_8 FILLER_55_853 ();
 sg13g2_fill_2 FILLER_55_860 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_4 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_60 ();
 sg13g2_fill_2 FILLER_56_119 ();
 sg13g2_decap_4 FILLER_56_129 ();
 sg13g2_fill_1 FILLER_56_133 ();
 sg13g2_fill_1 FILLER_56_139 ();
 sg13g2_decap_8 FILLER_56_164 ();
 sg13g2_fill_1 FILLER_56_171 ();
 sg13g2_decap_4 FILLER_56_191 ();
 sg13g2_fill_2 FILLER_56_202 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_fill_1 FILLER_56_214 ();
 sg13g2_decap_4 FILLER_56_236 ();
 sg13g2_fill_1 FILLER_56_240 ();
 sg13g2_fill_1 FILLER_56_263 ();
 sg13g2_decap_4 FILLER_56_268 ();
 sg13g2_fill_1 FILLER_56_272 ();
 sg13g2_fill_2 FILLER_56_280 ();
 sg13g2_fill_1 FILLER_56_286 ();
 sg13g2_fill_1 FILLER_56_301 ();
 sg13g2_decap_4 FILLER_56_357 ();
 sg13g2_fill_2 FILLER_56_361 ();
 sg13g2_fill_2 FILLER_56_372 ();
 sg13g2_fill_1 FILLER_56_374 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_fill_1 FILLER_56_397 ();
 sg13g2_fill_1 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_420 ();
 sg13g2_decap_8 FILLER_56_426 ();
 sg13g2_fill_2 FILLER_56_433 ();
 sg13g2_decap_8 FILLER_56_454 ();
 sg13g2_fill_2 FILLER_56_461 ();
 sg13g2_decap_8 FILLER_56_501 ();
 sg13g2_fill_1 FILLER_56_508 ();
 sg13g2_fill_2 FILLER_56_543 ();
 sg13g2_decap_8 FILLER_56_550 ();
 sg13g2_fill_2 FILLER_56_575 ();
 sg13g2_fill_1 FILLER_56_577 ();
 sg13g2_fill_1 FILLER_56_585 ();
 sg13g2_decap_8 FILLER_56_607 ();
 sg13g2_decap_8 FILLER_56_614 ();
 sg13g2_decap_8 FILLER_56_621 ();
 sg13g2_fill_1 FILLER_56_628 ();
 sg13g2_fill_1 FILLER_56_650 ();
 sg13g2_decap_8 FILLER_56_667 ();
 sg13g2_decap_4 FILLER_56_674 ();
 sg13g2_fill_1 FILLER_56_678 ();
 sg13g2_decap_8 FILLER_56_695 ();
 sg13g2_decap_4 FILLER_56_729 ();
 sg13g2_fill_1 FILLER_56_733 ();
 sg13g2_decap_8 FILLER_56_750 ();
 sg13g2_decap_4 FILLER_56_765 ();
 sg13g2_decap_8 FILLER_56_794 ();
 sg13g2_fill_2 FILLER_56_801 ();
 sg13g2_fill_2 FILLER_56_821 ();
 sg13g2_fill_1 FILLER_56_823 ();
 sg13g2_decap_8 FILLER_56_845 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_fill_2 FILLER_57_68 ();
 sg13g2_decap_4 FILLER_57_77 ();
 sg13g2_fill_2 FILLER_57_88 ();
 sg13g2_fill_1 FILLER_57_90 ();
 sg13g2_fill_2 FILLER_57_101 ();
 sg13g2_fill_1 FILLER_57_103 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_decap_4 FILLER_57_162 ();
 sg13g2_fill_1 FILLER_57_166 ();
 sg13g2_decap_4 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_198 ();
 sg13g2_fill_2 FILLER_57_222 ();
 sg13g2_fill_1 FILLER_57_238 ();
 sg13g2_decap_8 FILLER_57_246 ();
 sg13g2_decap_8 FILLER_57_253 ();
 sg13g2_fill_2 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_decap_8 FILLER_57_267 ();
 sg13g2_fill_1 FILLER_57_274 ();
 sg13g2_fill_1 FILLER_57_288 ();
 sg13g2_fill_1 FILLER_57_302 ();
 sg13g2_fill_1 FILLER_57_328 ();
 sg13g2_fill_2 FILLER_57_380 ();
 sg13g2_decap_4 FILLER_57_462 ();
 sg13g2_fill_2 FILLER_57_466 ();
 sg13g2_fill_2 FILLER_57_472 ();
 sg13g2_fill_2 FILLER_57_489 ();
 sg13g2_fill_1 FILLER_57_491 ();
 sg13g2_decap_4 FILLER_57_516 ();
 sg13g2_decap_4 FILLER_57_524 ();
 sg13g2_fill_1 FILLER_57_528 ();
 sg13g2_fill_1 FILLER_57_558 ();
 sg13g2_decap_8 FILLER_57_586 ();
 sg13g2_fill_2 FILLER_57_593 ();
 sg13g2_fill_1 FILLER_57_595 ();
 sg13g2_fill_2 FILLER_57_621 ();
 sg13g2_fill_1 FILLER_57_637 ();
 sg13g2_decap_8 FILLER_57_643 ();
 sg13g2_decap_8 FILLER_57_650 ();
 sg13g2_decap_4 FILLER_57_657 ();
 sg13g2_decap_4 FILLER_57_677 ();
 sg13g2_decap_8 FILLER_57_702 ();
 sg13g2_fill_1 FILLER_57_709 ();
 sg13g2_decap_4 FILLER_57_723 ();
 sg13g2_decap_4 FILLER_57_745 ();
 sg13g2_fill_1 FILLER_57_749 ();
 sg13g2_decap_4 FILLER_57_789 ();
 sg13g2_fill_2 FILLER_57_801 ();
 sg13g2_fill_1 FILLER_57_803 ();
 sg13g2_decap_4 FILLER_57_829 ();
 sg13g2_decap_8 FILLER_57_838 ();
 sg13g2_decap_8 FILLER_57_845 ();
 sg13g2_decap_8 FILLER_57_852 ();
 sg13g2_fill_2 FILLER_57_859 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_4 FILLER_58_35 ();
 sg13g2_fill_2 FILLER_58_39 ();
 sg13g2_fill_1 FILLER_58_76 ();
 sg13g2_fill_1 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_90 ();
 sg13g2_fill_1 FILLER_58_92 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_4 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_109 ();
 sg13g2_decap_8 FILLER_58_130 ();
 sg13g2_decap_4 FILLER_58_137 ();
 sg13g2_fill_2 FILLER_58_141 ();
 sg13g2_decap_4 FILLER_58_165 ();
 sg13g2_fill_1 FILLER_58_224 ();
 sg13g2_fill_2 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_decap_4 FILLER_58_273 ();
 sg13g2_fill_1 FILLER_58_277 ();
 sg13g2_fill_2 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_307 ();
 sg13g2_decap_8 FILLER_58_326 ();
 sg13g2_fill_1 FILLER_58_333 ();
 sg13g2_decap_8 FILLER_58_341 ();
 sg13g2_decap_8 FILLER_58_348 ();
 sg13g2_decap_8 FILLER_58_355 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_377 ();
 sg13g2_decap_4 FILLER_58_400 ();
 sg13g2_fill_2 FILLER_58_417 ();
 sg13g2_fill_2 FILLER_58_439 ();
 sg13g2_decap_8 FILLER_58_456 ();
 sg13g2_decap_4 FILLER_58_463 ();
 sg13g2_fill_1 FILLER_58_490 ();
 sg13g2_fill_1 FILLER_58_510 ();
 sg13g2_fill_2 FILLER_58_546 ();
 sg13g2_fill_2 FILLER_58_574 ();
 sg13g2_fill_1 FILLER_58_576 ();
 sg13g2_decap_4 FILLER_58_585 ();
 sg13g2_decap_4 FILLER_58_593 ();
 sg13g2_fill_1 FILLER_58_620 ();
 sg13g2_fill_2 FILLER_58_624 ();
 sg13g2_decap_8 FILLER_58_647 ();
 sg13g2_decap_4 FILLER_58_654 ();
 sg13g2_decap_8 FILLER_58_669 ();
 sg13g2_decap_4 FILLER_58_676 ();
 sg13g2_fill_2 FILLER_58_693 ();
 sg13g2_fill_1 FILLER_58_708 ();
 sg13g2_decap_8 FILLER_58_727 ();
 sg13g2_fill_2 FILLER_58_734 ();
 sg13g2_fill_1 FILLER_58_736 ();
 sg13g2_decap_4 FILLER_58_753 ();
 sg13g2_decap_8 FILLER_58_765 ();
 sg13g2_fill_2 FILLER_58_793 ();
 sg13g2_decap_8 FILLER_58_821 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_fill_2 FILLER_59_42 ();
 sg13g2_fill_1 FILLER_59_44 ();
 sg13g2_fill_2 FILLER_59_71 ();
 sg13g2_fill_1 FILLER_59_107 ();
 sg13g2_fill_1 FILLER_59_113 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_fill_2 FILLER_59_156 ();
 sg13g2_decap_8 FILLER_59_170 ();
 sg13g2_fill_2 FILLER_59_187 ();
 sg13g2_fill_1 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_200 ();
 sg13g2_fill_2 FILLER_59_207 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_decap_4 FILLER_59_225 ();
 sg13g2_fill_2 FILLER_59_229 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_decap_8 FILLER_59_260 ();
 sg13g2_fill_2 FILLER_59_271 ();
 sg13g2_fill_1 FILLER_59_273 ();
 sg13g2_fill_2 FILLER_59_280 ();
 sg13g2_fill_1 FILLER_59_282 ();
 sg13g2_fill_2 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_304 ();
 sg13g2_fill_2 FILLER_59_310 ();
 sg13g2_fill_1 FILLER_59_312 ();
 sg13g2_decap_8 FILLER_59_359 ();
 sg13g2_fill_2 FILLER_59_366 ();
 sg13g2_fill_1 FILLER_59_394 ();
 sg13g2_decap_8 FILLER_59_410 ();
 sg13g2_fill_2 FILLER_59_417 ();
 sg13g2_decap_8 FILLER_59_438 ();
 sg13g2_fill_2 FILLER_59_471 ();
 sg13g2_fill_2 FILLER_59_514 ();
 sg13g2_fill_1 FILLER_59_516 ();
 sg13g2_decap_8 FILLER_59_530 ();
 sg13g2_decap_8 FILLER_59_537 ();
 sg13g2_decap_4 FILLER_59_544 ();
 sg13g2_fill_2 FILLER_59_567 ();
 sg13g2_decap_8 FILLER_59_604 ();
 sg13g2_fill_2 FILLER_59_619 ();
 sg13g2_fill_2 FILLER_59_625 ();
 sg13g2_fill_1 FILLER_59_627 ();
 sg13g2_fill_2 FILLER_59_641 ();
 sg13g2_fill_1 FILLER_59_651 ();
 sg13g2_fill_2 FILLER_59_657 ();
 sg13g2_fill_1 FILLER_59_659 ();
 sg13g2_fill_2 FILLER_59_673 ();
 sg13g2_fill_2 FILLER_59_683 ();
 sg13g2_fill_1 FILLER_59_685 ();
 sg13g2_fill_2 FILLER_59_712 ();
 sg13g2_fill_1 FILLER_59_714 ();
 sg13g2_fill_2 FILLER_59_741 ();
 sg13g2_fill_1 FILLER_59_743 ();
 sg13g2_fill_2 FILLER_59_749 ();
 sg13g2_decap_8 FILLER_59_779 ();
 sg13g2_fill_1 FILLER_59_786 ();
 sg13g2_decap_8 FILLER_59_792 ();
 sg13g2_decap_8 FILLER_59_799 ();
 sg13g2_decap_8 FILLER_59_806 ();
 sg13g2_decap_8 FILLER_59_813 ();
 sg13g2_decap_8 FILLER_59_820 ();
 sg13g2_decap_8 FILLER_59_827 ();
 sg13g2_decap_8 FILLER_59_834 ();
 sg13g2_decap_8 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_855 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_4 FILLER_60_35 ();
 sg13g2_decap_4 FILLER_60_118 ();
 sg13g2_decap_8 FILLER_60_132 ();
 sg13g2_decap_4 FILLER_60_139 ();
 sg13g2_fill_2 FILLER_60_147 ();
 sg13g2_fill_1 FILLER_60_161 ();
 sg13g2_decap_4 FILLER_60_167 ();
 sg13g2_fill_2 FILLER_60_171 ();
 sg13g2_fill_2 FILLER_60_194 ();
 sg13g2_fill_1 FILLER_60_196 ();
 sg13g2_fill_2 FILLER_60_202 ();
 sg13g2_fill_2 FILLER_60_253 ();
 sg13g2_fill_1 FILLER_60_255 ();
 sg13g2_fill_2 FILLER_60_317 ();
 sg13g2_fill_1 FILLER_60_324 ();
 sg13g2_fill_2 FILLER_60_354 ();
 sg13g2_fill_2 FILLER_60_366 ();
 sg13g2_fill_2 FILLER_60_394 ();
 sg13g2_fill_1 FILLER_60_396 ();
 sg13g2_fill_2 FILLER_60_405 ();
 sg13g2_fill_1 FILLER_60_407 ();
 sg13g2_fill_1 FILLER_60_436 ();
 sg13g2_fill_2 FILLER_60_476 ();
 sg13g2_fill_1 FILLER_60_486 ();
 sg13g2_decap_4 FILLER_60_507 ();
 sg13g2_fill_2 FILLER_60_511 ();
 sg13g2_decap_4 FILLER_60_517 ();
 sg13g2_decap_4 FILLER_60_544 ();
 sg13g2_fill_1 FILLER_60_548 ();
 sg13g2_decap_4 FILLER_60_583 ();
 sg13g2_fill_1 FILLER_60_596 ();
 sg13g2_decap_4 FILLER_60_623 ();
 sg13g2_fill_1 FILLER_60_627 ();
 sg13g2_decap_8 FILLER_60_679 ();
 sg13g2_decap_8 FILLER_60_686 ();
 sg13g2_decap_4 FILLER_60_693 ();
 sg13g2_fill_1 FILLER_60_697 ();
 sg13g2_decap_8 FILLER_60_714 ();
 sg13g2_fill_1 FILLER_60_721 ();
 sg13g2_decap_4 FILLER_60_742 ();
 sg13g2_decap_8 FILLER_60_751 ();
 sg13g2_fill_1 FILLER_60_758 ();
 sg13g2_decap_8 FILLER_60_767 ();
 sg13g2_decap_8 FILLER_60_774 ();
 sg13g2_decap_8 FILLER_60_781 ();
 sg13g2_decap_8 FILLER_60_788 ();
 sg13g2_decap_8 FILLER_60_795 ();
 sg13g2_decap_8 FILLER_60_802 ();
 sg13g2_decap_8 FILLER_60_809 ();
 sg13g2_decap_8 FILLER_60_816 ();
 sg13g2_decap_8 FILLER_60_823 ();
 sg13g2_decap_8 FILLER_60_830 ();
 sg13g2_decap_8 FILLER_60_837 ();
 sg13g2_decap_8 FILLER_60_844 ();
 sg13g2_decap_8 FILLER_60_851 ();
 sg13g2_decap_4 FILLER_60_858 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_4 FILLER_61_35 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_fill_1 FILLER_61_67 ();
 sg13g2_fill_2 FILLER_61_73 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_fill_2 FILLER_61_105 ();
 sg13g2_fill_1 FILLER_61_177 ();
 sg13g2_decap_8 FILLER_61_201 ();
 sg13g2_decap_8 FILLER_61_213 ();
 sg13g2_fill_2 FILLER_61_227 ();
 sg13g2_fill_1 FILLER_61_229 ();
 sg13g2_decap_4 FILLER_61_239 ();
 sg13g2_fill_1 FILLER_61_253 ();
 sg13g2_decap_4 FILLER_61_269 ();
 sg13g2_fill_2 FILLER_61_273 ();
 sg13g2_fill_1 FILLER_61_308 ();
 sg13g2_decap_4 FILLER_61_324 ();
 sg13g2_decap_4 FILLER_61_340 ();
 sg13g2_fill_1 FILLER_61_344 ();
 sg13g2_decap_4 FILLER_61_413 ();
 sg13g2_decap_4 FILLER_61_422 ();
 sg13g2_decap_8 FILLER_61_435 ();
 sg13g2_decap_4 FILLER_61_442 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_fill_1 FILLER_61_466 ();
 sg13g2_fill_2 FILLER_61_479 ();
 sg13g2_fill_1 FILLER_61_490 ();
 sg13g2_decap_4 FILLER_61_561 ();
 sg13g2_fill_1 FILLER_61_565 ();
 sg13g2_fill_2 FILLER_61_581 ();
 sg13g2_fill_1 FILLER_61_593 ();
 sg13g2_fill_1 FILLER_61_608 ();
 sg13g2_decap_4 FILLER_61_622 ();
 sg13g2_fill_2 FILLER_61_626 ();
 sg13g2_fill_1 FILLER_61_633 ();
 sg13g2_decap_8 FILLER_61_639 ();
 sg13g2_fill_2 FILLER_61_646 ();
 sg13g2_fill_2 FILLER_61_656 ();
 sg13g2_decap_8 FILLER_61_684 ();
 sg13g2_decap_8 FILLER_61_691 ();
 sg13g2_fill_2 FILLER_61_698 ();
 sg13g2_fill_1 FILLER_61_700 ();
 sg13g2_decap_8 FILLER_61_714 ();
 sg13g2_decap_8 FILLER_61_721 ();
 sg13g2_decap_8 FILLER_61_728 ();
 sg13g2_decap_8 FILLER_61_735 ();
 sg13g2_decap_8 FILLER_61_742 ();
 sg13g2_decap_8 FILLER_61_749 ();
 sg13g2_decap_8 FILLER_61_756 ();
 sg13g2_decap_8 FILLER_61_763 ();
 sg13g2_decap_8 FILLER_61_770 ();
 sg13g2_decap_8 FILLER_61_777 ();
 sg13g2_decap_8 FILLER_61_784 ();
 sg13g2_decap_8 FILLER_61_791 ();
 sg13g2_decap_8 FILLER_61_798 ();
 sg13g2_decap_8 FILLER_61_805 ();
 sg13g2_decap_8 FILLER_61_812 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_decap_8 FILLER_61_826 ();
 sg13g2_decap_8 FILLER_61_833 ();
 sg13g2_decap_8 FILLER_61_840 ();
 sg13g2_decap_8 FILLER_61_847 ();
 sg13g2_decap_8 FILLER_61_854 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_fill_2 FILLER_62_49 ();
 sg13g2_fill_1 FILLER_62_51 ();
 sg13g2_fill_2 FILLER_62_56 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_fill_2 FILLER_62_93 ();
 sg13g2_fill_2 FILLER_62_113 ();
 sg13g2_fill_1 FILLER_62_168 ();
 sg13g2_fill_2 FILLER_62_174 ();
 sg13g2_decap_8 FILLER_62_184 ();
 sg13g2_decap_8 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_198 ();
 sg13g2_fill_2 FILLER_62_213 ();
 sg13g2_fill_2 FILLER_62_232 ();
 sg13g2_fill_1 FILLER_62_234 ();
 sg13g2_fill_2 FILLER_62_256 ();
 sg13g2_fill_1 FILLER_62_275 ();
 sg13g2_fill_1 FILLER_62_320 ();
 sg13g2_fill_1 FILLER_62_343 ();
 sg13g2_fill_1 FILLER_62_369 ();
 sg13g2_fill_1 FILLER_62_379 ();
 sg13g2_decap_8 FILLER_62_387 ();
 sg13g2_decap_4 FILLER_62_394 ();
 sg13g2_decap_4 FILLER_62_454 ();
 sg13g2_fill_1 FILLER_62_458 ();
 sg13g2_fill_2 FILLER_62_504 ();
 sg13g2_decap_8 FILLER_62_509 ();
 sg13g2_decap_8 FILLER_62_516 ();
 sg13g2_decap_4 FILLER_62_523 ();
 sg13g2_decap_4 FILLER_62_561 ();
 sg13g2_fill_1 FILLER_62_565 ();
 sg13g2_fill_1 FILLER_62_607 ();
 sg13g2_decap_8 FILLER_62_612 ();
 sg13g2_fill_1 FILLER_62_619 ();
 sg13g2_fill_1 FILLER_62_649 ();
 sg13g2_decap_8 FILLER_62_659 ();
 sg13g2_fill_2 FILLER_62_666 ();
 sg13g2_fill_1 FILLER_62_668 ();
 sg13g2_decap_8 FILLER_62_686 ();
 sg13g2_decap_8 FILLER_62_693 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_707 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_decap_8 FILLER_62_721 ();
 sg13g2_decap_8 FILLER_62_728 ();
 sg13g2_decap_8 FILLER_62_735 ();
 sg13g2_decap_8 FILLER_62_742 ();
 sg13g2_decap_8 FILLER_62_749 ();
 sg13g2_decap_8 FILLER_62_756 ();
 sg13g2_decap_8 FILLER_62_763 ();
 sg13g2_decap_8 FILLER_62_770 ();
 sg13g2_decap_8 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_791 ();
 sg13g2_decap_8 FILLER_62_798 ();
 sg13g2_decap_8 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_62_812 ();
 sg13g2_decap_8 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_826 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_decap_8 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_fill_1 FILLER_63_49 ();
 sg13g2_fill_2 FILLER_63_76 ();
 sg13g2_fill_1 FILLER_63_78 ();
 sg13g2_fill_2 FILLER_63_93 ();
 sg13g2_fill_2 FILLER_63_111 ();
 sg13g2_fill_2 FILLER_63_121 ();
 sg13g2_fill_1 FILLER_63_128 ();
 sg13g2_fill_2 FILLER_63_139 ();
 sg13g2_fill_1 FILLER_63_141 ();
 sg13g2_fill_2 FILLER_63_146 ();
 sg13g2_fill_1 FILLER_63_148 ();
 sg13g2_fill_2 FILLER_63_178 ();
 sg13g2_fill_1 FILLER_63_180 ();
 sg13g2_decap_4 FILLER_63_189 ();
 sg13g2_fill_1 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_227 ();
 sg13g2_fill_2 FILLER_63_243 ();
 sg13g2_fill_2 FILLER_63_271 ();
 sg13g2_decap_4 FILLER_63_299 ();
 sg13g2_decap_8 FILLER_63_306 ();
 sg13g2_decap_4 FILLER_63_330 ();
 sg13g2_decap_4 FILLER_63_339 ();
 sg13g2_fill_1 FILLER_63_343 ();
 sg13g2_fill_2 FILLER_63_348 ();
 sg13g2_decap_4 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_398 ();
 sg13g2_fill_1 FILLER_63_405 ();
 sg13g2_decap_8 FILLER_63_414 ();
 sg13g2_decap_8 FILLER_63_421 ();
 sg13g2_decap_8 FILLER_63_428 ();
 sg13g2_decap_8 FILLER_63_435 ();
 sg13g2_fill_2 FILLER_63_442 ();
 sg13g2_fill_2 FILLER_63_457 ();
 sg13g2_fill_1 FILLER_63_459 ();
 sg13g2_decap_8 FILLER_63_482 ();
 sg13g2_fill_1 FILLER_63_494 ();
 sg13g2_fill_2 FILLER_63_510 ();
 sg13g2_fill_1 FILLER_63_512 ();
 sg13g2_decap_4 FILLER_63_527 ();
 sg13g2_fill_2 FILLER_63_549 ();
 sg13g2_fill_1 FILLER_63_551 ();
 sg13g2_fill_2 FILLER_63_579 ();
 sg13g2_fill_1 FILLER_63_585 ();
 sg13g2_fill_1 FILLER_63_603 ();
 sg13g2_decap_4 FILLER_63_617 ();
 sg13g2_fill_2 FILLER_63_621 ();
 sg13g2_fill_2 FILLER_63_661 ();
 sg13g2_decap_8 FILLER_63_689 ();
 sg13g2_decap_8 FILLER_63_696 ();
 sg13g2_decap_8 FILLER_63_703 ();
 sg13g2_decap_8 FILLER_63_710 ();
 sg13g2_decap_8 FILLER_63_717 ();
 sg13g2_decap_8 FILLER_63_724 ();
 sg13g2_decap_8 FILLER_63_731 ();
 sg13g2_decap_8 FILLER_63_738 ();
 sg13g2_decap_8 FILLER_63_745 ();
 sg13g2_decap_8 FILLER_63_752 ();
 sg13g2_decap_8 FILLER_63_759 ();
 sg13g2_decap_8 FILLER_63_766 ();
 sg13g2_decap_8 FILLER_63_773 ();
 sg13g2_decap_8 FILLER_63_780 ();
 sg13g2_decap_8 FILLER_63_787 ();
 sg13g2_decap_8 FILLER_63_794 ();
 sg13g2_decap_8 FILLER_63_801 ();
 sg13g2_decap_8 FILLER_63_808 ();
 sg13g2_decap_8 FILLER_63_815 ();
 sg13g2_decap_8 FILLER_63_822 ();
 sg13g2_decap_8 FILLER_63_829 ();
 sg13g2_decap_8 FILLER_63_836 ();
 sg13g2_decap_8 FILLER_63_843 ();
 sg13g2_decap_8 FILLER_63_850 ();
 sg13g2_decap_4 FILLER_63_857 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_fill_1 FILLER_64_109 ();
 sg13g2_decap_4 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_165 ();
 sg13g2_fill_2 FILLER_64_190 ();
 sg13g2_fill_1 FILLER_64_192 ();
 sg13g2_fill_2 FILLER_64_202 ();
 sg13g2_fill_1 FILLER_64_204 ();
 sg13g2_fill_1 FILLER_64_222 ();
 sg13g2_fill_2 FILLER_64_228 ();
 sg13g2_fill_1 FILLER_64_230 ();
 sg13g2_fill_2 FILLER_64_247 ();
 sg13g2_fill_1 FILLER_64_249 ();
 sg13g2_decap_4 FILLER_64_263 ();
 sg13g2_fill_2 FILLER_64_267 ();
 sg13g2_decap_8 FILLER_64_299 ();
 sg13g2_fill_2 FILLER_64_323 ();
 sg13g2_fill_1 FILLER_64_325 ();
 sg13g2_fill_1 FILLER_64_364 ();
 sg13g2_decap_4 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_403 ();
 sg13g2_fill_1 FILLER_64_422 ();
 sg13g2_decap_8 FILLER_64_445 ();
 sg13g2_fill_1 FILLER_64_452 ();
 sg13g2_decap_8 FILLER_64_499 ();
 sg13g2_fill_2 FILLER_64_528 ();
 sg13g2_fill_2 FILLER_64_535 ();
 sg13g2_decap_8 FILLER_64_540 ();
 sg13g2_decap_8 FILLER_64_547 ();
 sg13g2_decap_4 FILLER_64_572 ();
 sg13g2_fill_1 FILLER_64_576 ();
 sg13g2_decap_8 FILLER_64_587 ();
 sg13g2_decap_4 FILLER_64_594 ();
 sg13g2_fill_1 FILLER_64_598 ();
 sg13g2_fill_1 FILLER_64_604 ();
 sg13g2_fill_2 FILLER_64_614 ();
 sg13g2_fill_2 FILLER_64_653 ();
 sg13g2_fill_2 FILLER_64_671 ();
 sg13g2_decap_8 FILLER_64_682 ();
 sg13g2_decap_8 FILLER_64_689 ();
 sg13g2_decap_8 FILLER_64_696 ();
 sg13g2_decap_8 FILLER_64_703 ();
 sg13g2_decap_8 FILLER_64_710 ();
 sg13g2_decap_8 FILLER_64_717 ();
 sg13g2_decap_8 FILLER_64_724 ();
 sg13g2_decap_8 FILLER_64_731 ();
 sg13g2_decap_8 FILLER_64_738 ();
 sg13g2_decap_8 FILLER_64_745 ();
 sg13g2_decap_8 FILLER_64_752 ();
 sg13g2_decap_8 FILLER_64_759 ();
 sg13g2_decap_8 FILLER_64_766 ();
 sg13g2_decap_8 FILLER_64_773 ();
 sg13g2_decap_8 FILLER_64_780 ();
 sg13g2_decap_8 FILLER_64_787 ();
 sg13g2_decap_8 FILLER_64_794 ();
 sg13g2_decap_8 FILLER_64_801 ();
 sg13g2_decap_8 FILLER_64_808 ();
 sg13g2_decap_8 FILLER_64_815 ();
 sg13g2_decap_8 FILLER_64_822 ();
 sg13g2_decap_8 FILLER_64_829 ();
 sg13g2_decap_8 FILLER_64_836 ();
 sg13g2_decap_8 FILLER_64_843 ();
 sg13g2_decap_8 FILLER_64_850 ();
 sg13g2_decap_4 FILLER_64_857 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_4 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_60 ();
 sg13g2_fill_1 FILLER_65_88 ();
 sg13g2_decap_4 FILLER_65_102 ();
 sg13g2_fill_1 FILLER_65_128 ();
 sg13g2_decap_8 FILLER_65_146 ();
 sg13g2_decap_8 FILLER_65_153 ();
 sg13g2_decap_8 FILLER_65_277 ();
 sg13g2_decap_8 FILLER_65_284 ();
 sg13g2_decap_8 FILLER_65_291 ();
 sg13g2_fill_1 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_fill_2 FILLER_65_350 ();
 sg13g2_decap_4 FILLER_65_386 ();
 sg13g2_fill_2 FILLER_65_390 ();
 sg13g2_decap_4 FILLER_65_397 ();
 sg13g2_decap_4 FILLER_65_405 ();
 sg13g2_decap_4 FILLER_65_431 ();
 sg13g2_fill_2 FILLER_65_435 ();
 sg13g2_decap_4 FILLER_65_450 ();
 sg13g2_fill_1 FILLER_65_454 ();
 sg13g2_fill_1 FILLER_65_460 ();
 sg13g2_fill_2 FILLER_65_471 ();
 sg13g2_fill_1 FILLER_65_473 ();
 sg13g2_decap_8 FILLER_65_499 ();
 sg13g2_fill_2 FILLER_65_511 ();
 sg13g2_fill_1 FILLER_65_513 ();
 sg13g2_decap_4 FILLER_65_547 ();
 sg13g2_decap_4 FILLER_65_564 ();
 sg13g2_fill_1 FILLER_65_579 ();
 sg13g2_fill_2 FILLER_65_601 ();
 sg13g2_fill_2 FILLER_65_623 ();
 sg13g2_fill_1 FILLER_65_645 ();
 sg13g2_fill_2 FILLER_65_650 ();
 sg13g2_fill_1 FILLER_65_652 ();
 sg13g2_decap_8 FILLER_65_676 ();
 sg13g2_decap_8 FILLER_65_683 ();
 sg13g2_decap_8 FILLER_65_690 ();
 sg13g2_decap_8 FILLER_65_697 ();
 sg13g2_decap_8 FILLER_65_704 ();
 sg13g2_decap_8 FILLER_65_711 ();
 sg13g2_decap_8 FILLER_65_718 ();
 sg13g2_decap_8 FILLER_65_725 ();
 sg13g2_decap_8 FILLER_65_732 ();
 sg13g2_decap_8 FILLER_65_739 ();
 sg13g2_decap_8 FILLER_65_746 ();
 sg13g2_decap_8 FILLER_65_753 ();
 sg13g2_decap_8 FILLER_65_760 ();
 sg13g2_decap_8 FILLER_65_767 ();
 sg13g2_decap_8 FILLER_65_774 ();
 sg13g2_decap_8 FILLER_65_781 ();
 sg13g2_decap_8 FILLER_65_788 ();
 sg13g2_decap_8 FILLER_65_795 ();
 sg13g2_decap_8 FILLER_65_802 ();
 sg13g2_decap_8 FILLER_65_809 ();
 sg13g2_decap_8 FILLER_65_816 ();
 sg13g2_decap_8 FILLER_65_823 ();
 sg13g2_decap_8 FILLER_65_830 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_8 FILLER_65_844 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_fill_2 FILLER_66_53 ();
 sg13g2_fill_2 FILLER_66_104 ();
 sg13g2_decap_4 FILLER_66_110 ();
 sg13g2_fill_2 FILLER_66_118 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_decap_8 FILLER_66_124 ();
 sg13g2_fill_2 FILLER_66_131 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_decap_4 FILLER_66_146 ();
 sg13g2_fill_1 FILLER_66_150 ();
 sg13g2_fill_2 FILLER_66_176 ();
 sg13g2_fill_1 FILLER_66_178 ();
 sg13g2_decap_4 FILLER_66_192 ();
 sg13g2_decap_4 FILLER_66_281 ();
 sg13g2_fill_2 FILLER_66_285 ();
 sg13g2_decap_8 FILLER_66_304 ();
 sg13g2_fill_2 FILLER_66_324 ();
 sg13g2_fill_2 FILLER_66_360 ();
 sg13g2_fill_1 FILLER_66_362 ();
 sg13g2_fill_2 FILLER_66_373 ();
 sg13g2_decap_4 FILLER_66_380 ();
 sg13g2_fill_1 FILLER_66_384 ();
 sg13g2_decap_8 FILLER_66_418 ();
 sg13g2_fill_2 FILLER_66_425 ();
 sg13g2_fill_2 FILLER_66_513 ();
 sg13g2_fill_1 FILLER_66_515 ();
 sg13g2_decap_8 FILLER_66_520 ();
 sg13g2_fill_1 FILLER_66_537 ();
 sg13g2_decap_8 FILLER_66_548 ();
 sg13g2_fill_1 FILLER_66_600 ();
 sg13g2_fill_2 FILLER_66_610 ();
 sg13g2_decap_4 FILLER_66_646 ();
 sg13g2_fill_2 FILLER_66_650 ();
 sg13g2_decap_8 FILLER_66_674 ();
 sg13g2_decap_8 FILLER_66_681 ();
 sg13g2_decap_8 FILLER_66_688 ();
 sg13g2_decap_8 FILLER_66_695 ();
 sg13g2_decap_8 FILLER_66_702 ();
 sg13g2_decap_8 FILLER_66_709 ();
 sg13g2_decap_8 FILLER_66_716 ();
 sg13g2_decap_8 FILLER_66_723 ();
 sg13g2_decap_8 FILLER_66_730 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_744 ();
 sg13g2_decap_8 FILLER_66_751 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_fill_2 FILLER_67_35 ();
 sg13g2_fill_1 FILLER_67_37 ();
 sg13g2_fill_1 FILLER_67_64 ();
 sg13g2_fill_2 FILLER_67_79 ();
 sg13g2_fill_2 FILLER_67_109 ();
 sg13g2_fill_1 FILLER_67_163 ();
 sg13g2_decap_4 FILLER_67_188 ();
 sg13g2_fill_2 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_260 ();
 sg13g2_fill_1 FILLER_67_327 ();
 sg13g2_fill_2 FILLER_67_368 ();
 sg13g2_decap_4 FILLER_67_416 ();
 sg13g2_fill_2 FILLER_67_420 ();
 sg13g2_decap_8 FILLER_67_426 ();
 sg13g2_decap_4 FILLER_67_433 ();
 sg13g2_decap_4 FILLER_67_442 ();
 sg13g2_fill_2 FILLER_67_450 ();
 sg13g2_decap_4 FILLER_67_457 ();
 sg13g2_fill_2 FILLER_67_461 ();
 sg13g2_decap_4 FILLER_67_473 ();
 sg13g2_decap_4 FILLER_67_486 ();
 sg13g2_decap_8 FILLER_67_507 ();
 sg13g2_decap_8 FILLER_67_514 ();
 sg13g2_decap_8 FILLER_67_521 ();
 sg13g2_fill_2 FILLER_67_528 ();
 sg13g2_fill_2 FILLER_67_553 ();
 sg13g2_decap_8 FILLER_67_565 ();
 sg13g2_decap_4 FILLER_67_572 ();
 sg13g2_decap_4 FILLER_67_589 ();
 sg13g2_decap_8 FILLER_67_606 ();
 sg13g2_decap_4 FILLER_67_613 ();
 sg13g2_fill_2 FILLER_67_638 ();
 sg13g2_fill_1 FILLER_67_640 ();
 sg13g2_fill_1 FILLER_67_652 ();
 sg13g2_fill_2 FILLER_67_658 ();
 sg13g2_fill_1 FILLER_67_660 ();
 sg13g2_decap_8 FILLER_67_675 ();
 sg13g2_decap_8 FILLER_67_682 ();
 sg13g2_decap_8 FILLER_67_689 ();
 sg13g2_decap_8 FILLER_67_696 ();
 sg13g2_decap_8 FILLER_67_703 ();
 sg13g2_decap_8 FILLER_67_710 ();
 sg13g2_decap_8 FILLER_67_717 ();
 sg13g2_decap_8 FILLER_67_724 ();
 sg13g2_decap_8 FILLER_67_731 ();
 sg13g2_decap_8 FILLER_67_738 ();
 sg13g2_decap_8 FILLER_67_745 ();
 sg13g2_decap_8 FILLER_67_752 ();
 sg13g2_decap_8 FILLER_67_759 ();
 sg13g2_decap_8 FILLER_67_766 ();
 sg13g2_decap_8 FILLER_67_773 ();
 sg13g2_decap_8 FILLER_67_780 ();
 sg13g2_decap_8 FILLER_67_787 ();
 sg13g2_decap_8 FILLER_67_794 ();
 sg13g2_decap_8 FILLER_67_801 ();
 sg13g2_decap_8 FILLER_67_808 ();
 sg13g2_decap_8 FILLER_67_815 ();
 sg13g2_decap_8 FILLER_67_822 ();
 sg13g2_decap_8 FILLER_67_829 ();
 sg13g2_decap_8 FILLER_67_836 ();
 sg13g2_decap_8 FILLER_67_843 ();
 sg13g2_decap_8 FILLER_67_850 ();
 sg13g2_decap_4 FILLER_67_857 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_fill_1 FILLER_68_28 ();
 sg13g2_fill_2 FILLER_68_46 ();
 sg13g2_fill_1 FILLER_68_48 ();
 sg13g2_fill_2 FILLER_68_102 ();
 sg13g2_fill_2 FILLER_68_145 ();
 sg13g2_decap_8 FILLER_68_152 ();
 sg13g2_decap_4 FILLER_68_159 ();
 sg13g2_decap_4 FILLER_68_175 ();
 sg13g2_fill_2 FILLER_68_179 ();
 sg13g2_fill_2 FILLER_68_212 ();
 sg13g2_fill_1 FILLER_68_214 ();
 sg13g2_fill_2 FILLER_68_250 ();
 sg13g2_decap_4 FILLER_68_278 ();
 sg13g2_fill_1 FILLER_68_282 ();
 sg13g2_decap_8 FILLER_68_305 ();
 sg13g2_decap_4 FILLER_68_312 ();
 sg13g2_fill_1 FILLER_68_316 ();
 sg13g2_fill_1 FILLER_68_332 ();
 sg13g2_fill_1 FILLER_68_349 ();
 sg13g2_fill_2 FILLER_68_380 ();
 sg13g2_decap_8 FILLER_68_387 ();
 sg13g2_decap_4 FILLER_68_406 ();
 sg13g2_fill_2 FILLER_68_410 ();
 sg13g2_fill_2 FILLER_68_473 ();
 sg13g2_fill_1 FILLER_68_475 ();
 sg13g2_fill_2 FILLER_68_496 ();
 sg13g2_fill_1 FILLER_68_498 ();
 sg13g2_fill_1 FILLER_68_511 ();
 sg13g2_decap_8 FILLER_68_535 ();
 sg13g2_decap_4 FILLER_68_557 ();
 sg13g2_fill_1 FILLER_68_578 ();
 sg13g2_fill_2 FILLER_68_592 ();
 sg13g2_fill_1 FILLER_68_594 ();
 sg13g2_fill_2 FILLER_68_616 ();
 sg13g2_fill_2 FILLER_68_635 ();
 sg13g2_fill_2 FILLER_68_657 ();
 sg13g2_decap_8 FILLER_68_669 ();
 sg13g2_decap_8 FILLER_68_676 ();
 sg13g2_decap_8 FILLER_68_683 ();
 sg13g2_decap_8 FILLER_68_690 ();
 sg13g2_decap_8 FILLER_68_697 ();
 sg13g2_decap_8 FILLER_68_704 ();
 sg13g2_decap_8 FILLER_68_711 ();
 sg13g2_decap_8 FILLER_68_718 ();
 sg13g2_decap_8 FILLER_68_725 ();
 sg13g2_decap_8 FILLER_68_732 ();
 sg13g2_decap_8 FILLER_68_739 ();
 sg13g2_decap_8 FILLER_68_746 ();
 sg13g2_decap_8 FILLER_68_753 ();
 sg13g2_decap_8 FILLER_68_760 ();
 sg13g2_decap_8 FILLER_68_767 ();
 sg13g2_decap_8 FILLER_68_774 ();
 sg13g2_decap_8 FILLER_68_781 ();
 sg13g2_decap_8 FILLER_68_788 ();
 sg13g2_decap_8 FILLER_68_795 ();
 sg13g2_decap_8 FILLER_68_802 ();
 sg13g2_decap_8 FILLER_68_809 ();
 sg13g2_decap_8 FILLER_68_816 ();
 sg13g2_decap_8 FILLER_68_823 ();
 sg13g2_decap_8 FILLER_68_830 ();
 sg13g2_decap_8 FILLER_68_837 ();
 sg13g2_decap_8 FILLER_68_844 ();
 sg13g2_decap_8 FILLER_68_851 ();
 sg13g2_decap_4 FILLER_68_858 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_4 FILLER_69_21 ();
 sg13g2_fill_2 FILLER_69_25 ();
 sg13g2_fill_2 FILLER_69_57 ();
 sg13g2_fill_1 FILLER_69_76 ();
 sg13g2_fill_1 FILLER_69_97 ();
 sg13g2_decap_8 FILLER_69_131 ();
 sg13g2_fill_2 FILLER_69_138 ();
 sg13g2_decap_8 FILLER_69_157 ();
 sg13g2_fill_2 FILLER_69_164 ();
 sg13g2_decap_4 FILLER_69_175 ();
 sg13g2_fill_1 FILLER_69_179 ();
 sg13g2_decap_4 FILLER_69_188 ();
 sg13g2_fill_1 FILLER_69_192 ();
 sg13g2_fill_2 FILLER_69_212 ();
 sg13g2_fill_1 FILLER_69_214 ();
 sg13g2_fill_2 FILLER_69_223 ();
 sg13g2_fill_1 FILLER_69_225 ();
 sg13g2_fill_2 FILLER_69_230 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_2 FILLER_69_262 ();
 sg13g2_fill_1 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_283 ();
 sg13g2_decap_8 FILLER_69_290 ();
 sg13g2_decap_8 FILLER_69_297 ();
 sg13g2_decap_4 FILLER_69_321 ();
 sg13g2_fill_2 FILLER_69_325 ();
 sg13g2_fill_2 FILLER_69_337 ();
 sg13g2_fill_1 FILLER_69_356 ();
 sg13g2_fill_2 FILLER_69_375 ();
 sg13g2_fill_1 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_decap_4 FILLER_69_408 ();
 sg13g2_fill_1 FILLER_69_422 ();
 sg13g2_fill_2 FILLER_69_427 ();
 sg13g2_decap_4 FILLER_69_439 ();
 sg13g2_fill_1 FILLER_69_452 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_decap_4 FILLER_69_467 ();
 sg13g2_fill_2 FILLER_69_479 ();
 sg13g2_decap_8 FILLER_69_518 ();
 sg13g2_fill_1 FILLER_69_525 ();
 sg13g2_decap_4 FILLER_69_531 ();
 sg13g2_decap_4 FILLER_69_543 ();
 sg13g2_fill_2 FILLER_69_547 ();
 sg13g2_fill_1 FILLER_69_555 ();
 sg13g2_decap_8 FILLER_69_571 ();
 sg13g2_decap_8 FILLER_69_578 ();
 sg13g2_decap_8 FILLER_69_585 ();
 sg13g2_fill_2 FILLER_69_597 ();
 sg13g2_fill_2 FILLER_69_604 ();
 sg13g2_decap_8 FILLER_69_614 ();
 sg13g2_fill_1 FILLER_69_621 ();
 sg13g2_fill_2 FILLER_69_627 ();
 sg13g2_fill_1 FILLER_69_635 ();
 sg13g2_fill_1 FILLER_69_641 ();
 sg13g2_decap_4 FILLER_69_650 ();
 sg13g2_fill_1 FILLER_69_654 ();
 sg13g2_fill_2 FILLER_69_660 ();
 sg13g2_fill_1 FILLER_69_662 ();
 sg13g2_decap_8 FILLER_69_676 ();
 sg13g2_decap_8 FILLER_69_683 ();
 sg13g2_decap_8 FILLER_69_690 ();
 sg13g2_decap_8 FILLER_69_697 ();
 sg13g2_decap_8 FILLER_69_704 ();
 sg13g2_decap_8 FILLER_69_711 ();
 sg13g2_decap_8 FILLER_69_718 ();
 sg13g2_decap_8 FILLER_69_725 ();
 sg13g2_decap_8 FILLER_69_732 ();
 sg13g2_decap_8 FILLER_69_739 ();
 sg13g2_decap_8 FILLER_69_746 ();
 sg13g2_decap_8 FILLER_69_753 ();
 sg13g2_decap_8 FILLER_69_760 ();
 sg13g2_decap_8 FILLER_69_767 ();
 sg13g2_decap_8 FILLER_69_774 ();
 sg13g2_decap_8 FILLER_69_781 ();
 sg13g2_decap_8 FILLER_69_788 ();
 sg13g2_decap_8 FILLER_69_795 ();
 sg13g2_decap_8 FILLER_69_802 ();
 sg13g2_decap_8 FILLER_69_809 ();
 sg13g2_decap_8 FILLER_69_816 ();
 sg13g2_decap_8 FILLER_69_823 ();
 sg13g2_decap_8 FILLER_69_830 ();
 sg13g2_decap_8 FILLER_69_837 ();
 sg13g2_decap_8 FILLER_69_844 ();
 sg13g2_decap_8 FILLER_69_851 ();
 sg13g2_decap_4 FILLER_69_858 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_11 ();
 sg13g2_fill_2 FILLER_70_38 ();
 sg13g2_fill_1 FILLER_70_40 ();
 sg13g2_fill_2 FILLER_70_55 ();
 sg13g2_fill_2 FILLER_70_97 ();
 sg13g2_fill_1 FILLER_70_127 ();
 sg13g2_decap_8 FILLER_70_157 ();
 sg13g2_decap_4 FILLER_70_164 ();
 sg13g2_fill_1 FILLER_70_168 ();
 sg13g2_fill_1 FILLER_70_217 ();
 sg13g2_decap_4 FILLER_70_244 ();
 sg13g2_fill_1 FILLER_70_248 ();
 sg13g2_decap_8 FILLER_70_290 ();
 sg13g2_decap_4 FILLER_70_314 ();
 sg13g2_fill_2 FILLER_70_318 ();
 sg13g2_decap_8 FILLER_70_346 ();
 sg13g2_fill_1 FILLER_70_353 ();
 sg13g2_decap_8 FILLER_70_363 ();
 sg13g2_fill_2 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_386 ();
 sg13g2_fill_2 FILLER_70_393 ();
 sg13g2_decap_8 FILLER_70_412 ();
 sg13g2_fill_2 FILLER_70_419 ();
 sg13g2_fill_2 FILLER_70_472 ();
 sg13g2_decap_4 FILLER_70_500 ();
 sg13g2_fill_2 FILLER_70_527 ();
 sg13g2_fill_1 FILLER_70_569 ();
 sg13g2_fill_2 FILLER_70_587 ();
 sg13g2_fill_2 FILLER_70_621 ();
 sg13g2_decap_8 FILLER_70_681 ();
 sg13g2_decap_8 FILLER_70_688 ();
 sg13g2_decap_8 FILLER_70_695 ();
 sg13g2_decap_8 FILLER_70_702 ();
 sg13g2_decap_8 FILLER_70_709 ();
 sg13g2_decap_8 FILLER_70_716 ();
 sg13g2_decap_8 FILLER_70_723 ();
 sg13g2_decap_8 FILLER_70_730 ();
 sg13g2_decap_8 FILLER_70_737 ();
 sg13g2_decap_8 FILLER_70_744 ();
 sg13g2_decap_8 FILLER_70_751 ();
 sg13g2_decap_8 FILLER_70_758 ();
 sg13g2_decap_8 FILLER_70_765 ();
 sg13g2_decap_8 FILLER_70_772 ();
 sg13g2_decap_8 FILLER_70_779 ();
 sg13g2_decap_8 FILLER_70_786 ();
 sg13g2_decap_8 FILLER_70_793 ();
 sg13g2_decap_8 FILLER_70_800 ();
 sg13g2_decap_8 FILLER_70_807 ();
 sg13g2_decap_8 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_821 ();
 sg13g2_decap_8 FILLER_70_828 ();
 sg13g2_decap_8 FILLER_70_835 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_4 FILLER_70_856 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_39 ();
 sg13g2_fill_2 FILLER_71_70 ();
 sg13g2_fill_2 FILLER_71_92 ();
 sg13g2_fill_2 FILLER_71_177 ();
 sg13g2_fill_1 FILLER_71_179 ();
 sg13g2_decap_4 FILLER_71_184 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_205 ();
 sg13g2_fill_1 FILLER_71_214 ();
 sg13g2_fill_1 FILLER_71_233 ();
 sg13g2_fill_2 FILLER_71_243 ();
 sg13g2_fill_1 FILLER_71_245 ();
 sg13g2_fill_2 FILLER_71_270 ();
 sg13g2_fill_2 FILLER_71_281 ();
 sg13g2_fill_1 FILLER_71_283 ();
 sg13g2_decap_8 FILLER_71_309 ();
 sg13g2_decap_4 FILLER_71_316 ();
 sg13g2_fill_2 FILLER_71_320 ();
 sg13g2_fill_1 FILLER_71_327 ();
 sg13g2_fill_1 FILLER_71_336 ();
 sg13g2_decap_4 FILLER_71_346 ();
 sg13g2_fill_2 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_71_389 ();
 sg13g2_fill_1 FILLER_71_396 ();
 sg13g2_decap_4 FILLER_71_422 ();
 sg13g2_fill_2 FILLER_71_426 ();
 sg13g2_fill_2 FILLER_71_437 ();
 sg13g2_fill_1 FILLER_71_439 ();
 sg13g2_fill_1 FILLER_71_444 ();
 sg13g2_decap_4 FILLER_71_450 ();
 sg13g2_decap_4 FILLER_71_458 ();
 sg13g2_fill_1 FILLER_71_472 ();
 sg13g2_decap_4 FILLER_71_499 ();
 sg13g2_fill_2 FILLER_71_514 ();
 sg13g2_fill_1 FILLER_71_530 ();
 sg13g2_decap_4 FILLER_71_535 ();
 sg13g2_decap_8 FILLER_71_548 ();
 sg13g2_decap_4 FILLER_71_555 ();
 sg13g2_fill_1 FILLER_71_559 ();
 sg13g2_fill_2 FILLER_71_592 ();
 sg13g2_fill_2 FILLER_71_600 ();
 sg13g2_decap_4 FILLER_71_631 ();
 sg13g2_fill_2 FILLER_71_635 ();
 sg13g2_fill_2 FILLER_71_655 ();
 sg13g2_fill_1 FILLER_71_657 ();
 sg13g2_decap_8 FILLER_71_676 ();
 sg13g2_decap_8 FILLER_71_683 ();
 sg13g2_decap_8 FILLER_71_690 ();
 sg13g2_decap_8 FILLER_71_697 ();
 sg13g2_decap_8 FILLER_71_704 ();
 sg13g2_decap_8 FILLER_71_711 ();
 sg13g2_decap_8 FILLER_71_718 ();
 sg13g2_decap_8 FILLER_71_725 ();
 sg13g2_decap_8 FILLER_71_732 ();
 sg13g2_decap_8 FILLER_71_739 ();
 sg13g2_decap_8 FILLER_71_746 ();
 sg13g2_decap_8 FILLER_71_753 ();
 sg13g2_decap_8 FILLER_71_760 ();
 sg13g2_decap_8 FILLER_71_767 ();
 sg13g2_decap_8 FILLER_71_774 ();
 sg13g2_decap_8 FILLER_71_781 ();
 sg13g2_decap_8 FILLER_71_788 ();
 sg13g2_decap_8 FILLER_71_795 ();
 sg13g2_decap_8 FILLER_71_802 ();
 sg13g2_decap_8 FILLER_71_809 ();
 sg13g2_decap_8 FILLER_71_816 ();
 sg13g2_decap_8 FILLER_71_823 ();
 sg13g2_decap_8 FILLER_71_830 ();
 sg13g2_decap_8 FILLER_71_837 ();
 sg13g2_decap_8 FILLER_71_844 ();
 sg13g2_decap_8 FILLER_71_851 ();
 sg13g2_decap_4 FILLER_71_858 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_35 ();
 sg13g2_fill_1 FILLER_72_104 ();
 sg13g2_fill_2 FILLER_72_146 ();
 sg13g2_decap_8 FILLER_72_165 ();
 sg13g2_decap_8 FILLER_72_172 ();
 sg13g2_decap_4 FILLER_72_210 ();
 sg13g2_decap_4 FILLER_72_233 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_1 FILLER_72_330 ();
 sg13g2_decap_8 FILLER_72_341 ();
 sg13g2_decap_4 FILLER_72_348 ();
 sg13g2_fill_2 FILLER_72_352 ();
 sg13g2_fill_2 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_366 ();
 sg13g2_fill_2 FILLER_72_384 ();
 sg13g2_fill_1 FILLER_72_386 ();
 sg13g2_decap_4 FILLER_72_414 ();
 sg13g2_fill_1 FILLER_72_418 ();
 sg13g2_fill_1 FILLER_72_510 ();
 sg13g2_fill_2 FILLER_72_520 ();
 sg13g2_fill_1 FILLER_72_522 ();
 sg13g2_fill_1 FILLER_72_538 ();
 sg13g2_fill_1 FILLER_72_553 ();
 sg13g2_fill_2 FILLER_72_579 ();
 sg13g2_fill_1 FILLER_72_581 ();
 sg13g2_fill_1 FILLER_72_609 ();
 sg13g2_fill_1 FILLER_72_636 ();
 sg13g2_decap_4 FILLER_72_653 ();
 sg13g2_decap_8 FILLER_72_683 ();
 sg13g2_decap_8 FILLER_72_690 ();
 sg13g2_decap_8 FILLER_72_697 ();
 sg13g2_decap_8 FILLER_72_704 ();
 sg13g2_decap_8 FILLER_72_711 ();
 sg13g2_decap_8 FILLER_72_718 ();
 sg13g2_decap_8 FILLER_72_725 ();
 sg13g2_decap_8 FILLER_72_732 ();
 sg13g2_decap_8 FILLER_72_739 ();
 sg13g2_decap_8 FILLER_72_746 ();
 sg13g2_decap_8 FILLER_72_753 ();
 sg13g2_decap_8 FILLER_72_760 ();
 sg13g2_decap_8 FILLER_72_767 ();
 sg13g2_decap_8 FILLER_72_774 ();
 sg13g2_decap_8 FILLER_72_781 ();
 sg13g2_decap_8 FILLER_72_788 ();
 sg13g2_decap_8 FILLER_72_795 ();
 sg13g2_decap_8 FILLER_72_802 ();
 sg13g2_decap_8 FILLER_72_809 ();
 sg13g2_decap_8 FILLER_72_816 ();
 sg13g2_decap_8 FILLER_72_823 ();
 sg13g2_decap_8 FILLER_72_830 ();
 sg13g2_decap_8 FILLER_72_837 ();
 sg13g2_decap_8 FILLER_72_844 ();
 sg13g2_decap_8 FILLER_72_851 ();
 sg13g2_decap_4 FILLER_72_858 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_4 FILLER_73_14 ();
 sg13g2_fill_1 FILLER_73_44 ();
 sg13g2_fill_1 FILLER_73_53 ();
 sg13g2_fill_2 FILLER_73_115 ();
 sg13g2_decap_4 FILLER_73_166 ();
 sg13g2_fill_2 FILLER_73_269 ();
 sg13g2_fill_1 FILLER_73_271 ();
 sg13g2_decap_8 FILLER_73_281 ();
 sg13g2_decap_8 FILLER_73_293 ();
 sg13g2_fill_1 FILLER_73_300 ();
 sg13g2_decap_4 FILLER_73_349 ();
 sg13g2_fill_1 FILLER_73_353 ();
 sg13g2_fill_1 FILLER_73_370 ();
 sg13g2_decap_8 FILLER_73_390 ();
 sg13g2_fill_2 FILLER_73_397 ();
 sg13g2_decap_8 FILLER_73_414 ();
 sg13g2_decap_8 FILLER_73_421 ();
 sg13g2_fill_1 FILLER_73_428 ();
 sg13g2_decap_8 FILLER_73_433 ();
 sg13g2_decap_4 FILLER_73_440 ();
 sg13g2_fill_1 FILLER_73_485 ();
 sg13g2_fill_1 FILLER_73_490 ();
 sg13g2_fill_2 FILLER_73_495 ();
 sg13g2_fill_2 FILLER_73_519 ();
 sg13g2_fill_1 FILLER_73_521 ();
 sg13g2_fill_2 FILLER_73_582 ();
 sg13g2_fill_1 FILLER_73_584 ();
 sg13g2_fill_2 FILLER_73_603 ();
 sg13g2_decap_4 FILLER_73_631 ();
 sg13g2_fill_2 FILLER_73_653 ();
 sg13g2_decap_8 FILLER_73_669 ();
 sg13g2_decap_8 FILLER_73_676 ();
 sg13g2_decap_8 FILLER_73_683 ();
 sg13g2_decap_8 FILLER_73_690 ();
 sg13g2_decap_8 FILLER_73_697 ();
 sg13g2_decap_8 FILLER_73_704 ();
 sg13g2_decap_8 FILLER_73_711 ();
 sg13g2_decap_8 FILLER_73_718 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_decap_8 FILLER_73_732 ();
 sg13g2_decap_8 FILLER_73_739 ();
 sg13g2_decap_8 FILLER_73_746 ();
 sg13g2_decap_8 FILLER_73_753 ();
 sg13g2_decap_8 FILLER_73_760 ();
 sg13g2_decap_8 FILLER_73_767 ();
 sg13g2_decap_8 FILLER_73_774 ();
 sg13g2_decap_8 FILLER_73_781 ();
 sg13g2_decap_8 FILLER_73_788 ();
 sg13g2_decap_8 FILLER_73_795 ();
 sg13g2_decap_8 FILLER_73_802 ();
 sg13g2_decap_8 FILLER_73_809 ();
 sg13g2_decap_8 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_830 ();
 sg13g2_decap_8 FILLER_73_837 ();
 sg13g2_decap_8 FILLER_73_844 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_decap_4 FILLER_73_858 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_fill_2 FILLER_74_50 ();
 sg13g2_fill_2 FILLER_74_69 ();
 sg13g2_fill_2 FILLER_74_104 ();
 sg13g2_fill_2 FILLER_74_166 ();
 sg13g2_fill_2 FILLER_74_213 ();
 sg13g2_fill_1 FILLER_74_215 ();
 sg13g2_decap_4 FILLER_74_239 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_fill_1 FILLER_74_299 ();
 sg13g2_fill_2 FILLER_74_326 ();
 sg13g2_fill_1 FILLER_74_328 ();
 sg13g2_fill_2 FILLER_74_333 ();
 sg13g2_fill_2 FILLER_74_368 ();
 sg13g2_fill_1 FILLER_74_370 ();
 sg13g2_fill_2 FILLER_74_444 ();
 sg13g2_fill_1 FILLER_74_496 ();
 sg13g2_fill_2 FILLER_74_531 ();
 sg13g2_fill_2 FILLER_74_577 ();
 sg13g2_fill_2 FILLER_74_583 ();
 sg13g2_fill_1 FILLER_74_585 ();
 sg13g2_fill_2 FILLER_74_594 ();
 sg13g2_fill_2 FILLER_74_631 ();
 sg13g2_fill_1 FILLER_74_633 ();
 sg13g2_decap_8 FILLER_74_669 ();
 sg13g2_decap_8 FILLER_74_676 ();
 sg13g2_decap_8 FILLER_74_683 ();
 sg13g2_decap_8 FILLER_74_690 ();
 sg13g2_decap_8 FILLER_74_697 ();
 sg13g2_decap_8 FILLER_74_704 ();
 sg13g2_decap_8 FILLER_74_711 ();
 sg13g2_decap_8 FILLER_74_718 ();
 sg13g2_decap_8 FILLER_74_725 ();
 sg13g2_decap_8 FILLER_74_732 ();
 sg13g2_decap_8 FILLER_74_739 ();
 sg13g2_decap_8 FILLER_74_746 ();
 sg13g2_decap_8 FILLER_74_753 ();
 sg13g2_decap_8 FILLER_74_760 ();
 sg13g2_decap_8 FILLER_74_767 ();
 sg13g2_decap_8 FILLER_74_774 ();
 sg13g2_decap_8 FILLER_74_781 ();
 sg13g2_decap_8 FILLER_74_788 ();
 sg13g2_decap_8 FILLER_74_795 ();
 sg13g2_decap_8 FILLER_74_802 ();
 sg13g2_decap_8 FILLER_74_809 ();
 sg13g2_decap_8 FILLER_74_816 ();
 sg13g2_decap_8 FILLER_74_823 ();
 sg13g2_decap_8 FILLER_74_830 ();
 sg13g2_decap_8 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_844 ();
 sg13g2_decap_8 FILLER_74_851 ();
 sg13g2_decap_4 FILLER_74_858 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_fill_2 FILLER_75_28 ();
 sg13g2_fill_1 FILLER_75_30 ();
 sg13g2_fill_1 FILLER_75_75 ();
 sg13g2_decap_4 FILLER_75_229 ();
 sg13g2_fill_1 FILLER_75_233 ();
 sg13g2_fill_2 FILLER_75_261 ();
 sg13g2_fill_1 FILLER_75_263 ();
 sg13g2_decap_4 FILLER_75_274 ();
 sg13g2_fill_1 FILLER_75_278 ();
 sg13g2_decap_4 FILLER_75_283 ();
 sg13g2_decap_8 FILLER_75_318 ();
 sg13g2_decap_8 FILLER_75_325 ();
 sg13g2_decap_4 FILLER_75_332 ();
 sg13g2_fill_1 FILLER_75_336 ();
 sg13g2_fill_2 FILLER_75_361 ();
 sg13g2_fill_1 FILLER_75_363 ();
 sg13g2_fill_2 FILLER_75_377 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_fill_1 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_402 ();
 sg13g2_fill_2 FILLER_75_409 ();
 sg13g2_fill_1 FILLER_75_411 ();
 sg13g2_decap_8 FILLER_75_438 ();
 sg13g2_fill_2 FILLER_75_445 ();
 sg13g2_fill_1 FILLER_75_480 ();
 sg13g2_fill_2 FILLER_75_489 ();
 sg13g2_fill_1 FILLER_75_491 ();
 sg13g2_fill_2 FILLER_75_501 ();
 sg13g2_fill_1 FILLER_75_503 ();
 sg13g2_fill_2 FILLER_75_560 ();
 sg13g2_decap_8 FILLER_75_618 ();
 sg13g2_decap_8 FILLER_75_625 ();
 sg13g2_decap_8 FILLER_75_632 ();
 sg13g2_decap_8 FILLER_75_644 ();
 sg13g2_fill_2 FILLER_75_651 ();
 sg13g2_decap_8 FILLER_75_657 ();
 sg13g2_decap_8 FILLER_75_664 ();
 sg13g2_decap_8 FILLER_75_671 ();
 sg13g2_decap_8 FILLER_75_678 ();
 sg13g2_decap_8 FILLER_75_685 ();
 sg13g2_decap_8 FILLER_75_692 ();
 sg13g2_decap_8 FILLER_75_699 ();
 sg13g2_decap_8 FILLER_75_706 ();
 sg13g2_decap_8 FILLER_75_713 ();
 sg13g2_decap_8 FILLER_75_720 ();
 sg13g2_decap_8 FILLER_75_727 ();
 sg13g2_decap_8 FILLER_75_734 ();
 sg13g2_decap_8 FILLER_75_741 ();
 sg13g2_decap_8 FILLER_75_748 ();
 sg13g2_decap_8 FILLER_75_755 ();
 sg13g2_decap_8 FILLER_75_762 ();
 sg13g2_decap_8 FILLER_75_769 ();
 sg13g2_decap_8 FILLER_75_776 ();
 sg13g2_decap_8 FILLER_75_783 ();
 sg13g2_decap_8 FILLER_75_790 ();
 sg13g2_decap_8 FILLER_75_797 ();
 sg13g2_decap_8 FILLER_75_804 ();
 sg13g2_decap_8 FILLER_75_811 ();
 sg13g2_decap_8 FILLER_75_818 ();
 sg13g2_decap_8 FILLER_75_825 ();
 sg13g2_decap_8 FILLER_75_832 ();
 sg13g2_decap_8 FILLER_75_839 ();
 sg13g2_decap_8 FILLER_75_846 ();
 sg13g2_decap_8 FILLER_75_853 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_fill_1 FILLER_76_85 ();
 sg13g2_fill_2 FILLER_76_111 ();
 sg13g2_fill_2 FILLER_76_170 ();
 sg13g2_fill_2 FILLER_76_222 ();
 sg13g2_decap_8 FILLER_76_278 ();
 sg13g2_fill_1 FILLER_76_285 ();
 sg13g2_decap_8 FILLER_76_290 ();
 sg13g2_fill_2 FILLER_76_297 ();
 sg13g2_fill_2 FILLER_76_304 ();
 sg13g2_fill_1 FILLER_76_306 ();
 sg13g2_decap_8 FILLER_76_316 ();
 sg13g2_decap_4 FILLER_76_323 ();
 sg13g2_fill_1 FILLER_76_353 ();
 sg13g2_fill_2 FILLER_76_380 ();
 sg13g2_fill_1 FILLER_76_382 ();
 sg13g2_decap_8 FILLER_76_409 ();
 sg13g2_fill_2 FILLER_76_416 ();
 sg13g2_fill_1 FILLER_76_418 ();
 sg13g2_fill_1 FILLER_76_432 ();
 sg13g2_fill_2 FILLER_76_459 ();
 sg13g2_fill_2 FILLER_76_483 ();
 sg13g2_fill_1 FILLER_76_485 ();
 sg13g2_fill_2 FILLER_76_512 ();
 sg13g2_fill_1 FILLER_76_514 ();
 sg13g2_decap_8 FILLER_76_519 ();
 sg13g2_decap_4 FILLER_76_526 ();
 sg13g2_fill_1 FILLER_76_530 ();
 sg13g2_decap_8 FILLER_76_539 ();
 sg13g2_decap_8 FILLER_76_546 ();
 sg13g2_decap_8 FILLER_76_553 ();
 sg13g2_decap_8 FILLER_76_560 ();
 sg13g2_decap_8 FILLER_76_567 ();
 sg13g2_decap_8 FILLER_76_574 ();
 sg13g2_decap_8 FILLER_76_581 ();
 sg13g2_decap_8 FILLER_76_588 ();
 sg13g2_decap_8 FILLER_76_595 ();
 sg13g2_decap_8 FILLER_76_602 ();
 sg13g2_decap_8 FILLER_76_609 ();
 sg13g2_decap_8 FILLER_76_616 ();
 sg13g2_decap_8 FILLER_76_623 ();
 sg13g2_decap_8 FILLER_76_630 ();
 sg13g2_decap_8 FILLER_76_637 ();
 sg13g2_decap_8 FILLER_76_644 ();
 sg13g2_decap_8 FILLER_76_651 ();
 sg13g2_decap_8 FILLER_76_658 ();
 sg13g2_decap_8 FILLER_76_665 ();
 sg13g2_decap_8 FILLER_76_672 ();
 sg13g2_decap_8 FILLER_76_679 ();
 sg13g2_decap_8 FILLER_76_686 ();
 sg13g2_decap_8 FILLER_76_693 ();
 sg13g2_decap_8 FILLER_76_700 ();
 sg13g2_decap_8 FILLER_76_707 ();
 sg13g2_decap_8 FILLER_76_714 ();
 sg13g2_decap_8 FILLER_76_721 ();
 sg13g2_decap_8 FILLER_76_728 ();
 sg13g2_decap_8 FILLER_76_735 ();
 sg13g2_decap_8 FILLER_76_742 ();
 sg13g2_decap_8 FILLER_76_749 ();
 sg13g2_decap_8 FILLER_76_756 ();
 sg13g2_decap_8 FILLER_76_763 ();
 sg13g2_decap_8 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_784 ();
 sg13g2_decap_8 FILLER_76_791 ();
 sg13g2_decap_8 FILLER_76_798 ();
 sg13g2_decap_8 FILLER_76_805 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_decap_8 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_833 ();
 sg13g2_decap_8 FILLER_76_840 ();
 sg13g2_decap_8 FILLER_76_847 ();
 sg13g2_decap_8 FILLER_76_854 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_fill_2 FILLER_77_28 ();
 sg13g2_fill_1 FILLER_77_30 ();
 sg13g2_fill_2 FILLER_77_61 ();
 sg13g2_fill_1 FILLER_77_110 ();
 sg13g2_fill_1 FILLER_77_120 ();
 sg13g2_fill_2 FILLER_77_147 ();
 sg13g2_fill_2 FILLER_77_179 ();
 sg13g2_fill_1 FILLER_77_245 ();
 sg13g2_fill_2 FILLER_77_272 ();
 sg13g2_fill_1 FILLER_77_274 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_fill_2 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_342 ();
 sg13g2_decap_8 FILLER_77_349 ();
 sg13g2_decap_8 FILLER_77_356 ();
 sg13g2_fill_2 FILLER_77_363 ();
 sg13g2_decap_8 FILLER_77_369 ();
 sg13g2_decap_8 FILLER_77_376 ();
 sg13g2_decap_8 FILLER_77_383 ();
 sg13g2_decap_4 FILLER_77_390 ();
 sg13g2_decap_8 FILLER_77_398 ();
 sg13g2_decap_8 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_77_412 ();
 sg13g2_decap_8 FILLER_77_419 ();
 sg13g2_decap_8 FILLER_77_426 ();
 sg13g2_decap_8 FILLER_77_433 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_fill_1 FILLER_77_442 ();
 sg13g2_decap_8 FILLER_77_447 ();
 sg13g2_fill_1 FILLER_77_454 ();
 sg13g2_decap_8 FILLER_77_481 ();
 sg13g2_decap_4 FILLER_77_488 ();
 sg13g2_fill_2 FILLER_77_492 ();
 sg13g2_decap_8 FILLER_77_503 ();
 sg13g2_decap_8 FILLER_77_510 ();
 sg13g2_decap_8 FILLER_77_517 ();
 sg13g2_decap_8 FILLER_77_524 ();
 sg13g2_decap_8 FILLER_77_531 ();
 sg13g2_decap_8 FILLER_77_538 ();
 sg13g2_decap_8 FILLER_77_545 ();
 sg13g2_decap_8 FILLER_77_552 ();
 sg13g2_decap_8 FILLER_77_559 ();
 sg13g2_decap_8 FILLER_77_566 ();
 sg13g2_decap_8 FILLER_77_573 ();
 sg13g2_decap_8 FILLER_77_580 ();
 sg13g2_decap_8 FILLER_77_587 ();
 sg13g2_decap_8 FILLER_77_594 ();
 sg13g2_decap_8 FILLER_77_601 ();
 sg13g2_decap_8 FILLER_77_608 ();
 sg13g2_decap_8 FILLER_77_615 ();
 sg13g2_decap_8 FILLER_77_622 ();
 sg13g2_decap_8 FILLER_77_629 ();
 sg13g2_decap_8 FILLER_77_636 ();
 sg13g2_decap_8 FILLER_77_643 ();
 sg13g2_decap_8 FILLER_77_650 ();
 sg13g2_decap_8 FILLER_77_657 ();
 sg13g2_decap_8 FILLER_77_664 ();
 sg13g2_decap_8 FILLER_77_671 ();
 sg13g2_decap_8 FILLER_77_678 ();
 sg13g2_decap_8 FILLER_77_685 ();
 sg13g2_decap_8 FILLER_77_692 ();
 sg13g2_decap_8 FILLER_77_699 ();
 sg13g2_decap_8 FILLER_77_706 ();
 sg13g2_decap_8 FILLER_77_713 ();
 sg13g2_decap_8 FILLER_77_720 ();
 sg13g2_decap_8 FILLER_77_727 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_decap_8 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_755 ();
 sg13g2_decap_8 FILLER_77_762 ();
 sg13g2_decap_8 FILLER_77_769 ();
 sg13g2_decap_8 FILLER_77_776 ();
 sg13g2_decap_8 FILLER_77_783 ();
 sg13g2_decap_8 FILLER_77_790 ();
 sg13g2_decap_8 FILLER_77_797 ();
 sg13g2_decap_8 FILLER_77_804 ();
 sg13g2_decap_8 FILLER_77_811 ();
 sg13g2_decap_8 FILLER_77_818 ();
 sg13g2_decap_8 FILLER_77_825 ();
 sg13g2_decap_8 FILLER_77_832 ();
 sg13g2_decap_8 FILLER_77_839 ();
 sg13g2_decap_8 FILLER_77_846 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_4 FILLER_78_35 ();
 sg13g2_fill_1 FILLER_78_149 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_182 ();
 sg13g2_decap_4 FILLER_78_187 ();
 sg13g2_fill_1 FILLER_78_191 ();
 sg13g2_fill_1 FILLER_78_196 ();
 sg13g2_fill_1 FILLER_78_233 ();
 sg13g2_decap_8 FILLER_78_265 ();
 sg13g2_decap_8 FILLER_78_272 ();
 sg13g2_decap_8 FILLER_78_279 ();
 sg13g2_decap_8 FILLER_78_286 ();
 sg13g2_decap_8 FILLER_78_293 ();
 sg13g2_decap_8 FILLER_78_300 ();
 sg13g2_decap_8 FILLER_78_307 ();
 sg13g2_decap_8 FILLER_78_314 ();
 sg13g2_decap_8 FILLER_78_321 ();
 sg13g2_decap_8 FILLER_78_328 ();
 sg13g2_decap_8 FILLER_78_335 ();
 sg13g2_decap_8 FILLER_78_342 ();
 sg13g2_decap_8 FILLER_78_349 ();
 sg13g2_decap_8 FILLER_78_356 ();
 sg13g2_decap_8 FILLER_78_363 ();
 sg13g2_decap_8 FILLER_78_370 ();
 sg13g2_decap_8 FILLER_78_377 ();
 sg13g2_decap_8 FILLER_78_384 ();
 sg13g2_decap_8 FILLER_78_391 ();
 sg13g2_decap_8 FILLER_78_398 ();
 sg13g2_decap_8 FILLER_78_405 ();
 sg13g2_decap_8 FILLER_78_412 ();
 sg13g2_decap_8 FILLER_78_419 ();
 sg13g2_decap_8 FILLER_78_426 ();
 sg13g2_decap_8 FILLER_78_433 ();
 sg13g2_decap_8 FILLER_78_440 ();
 sg13g2_decap_8 FILLER_78_447 ();
 sg13g2_decap_8 FILLER_78_454 ();
 sg13g2_decap_4 FILLER_78_461 ();
 sg13g2_fill_1 FILLER_78_465 ();
 sg13g2_decap_8 FILLER_78_470 ();
 sg13g2_decap_8 FILLER_78_477 ();
 sg13g2_decap_8 FILLER_78_484 ();
 sg13g2_decap_8 FILLER_78_491 ();
 sg13g2_decap_8 FILLER_78_498 ();
 sg13g2_decap_8 FILLER_78_505 ();
 sg13g2_decap_8 FILLER_78_512 ();
 sg13g2_decap_8 FILLER_78_519 ();
 sg13g2_decap_8 FILLER_78_526 ();
 sg13g2_decap_8 FILLER_78_533 ();
 sg13g2_decap_8 FILLER_78_540 ();
 sg13g2_decap_8 FILLER_78_547 ();
 sg13g2_decap_8 FILLER_78_554 ();
 sg13g2_decap_8 FILLER_78_561 ();
 sg13g2_decap_8 FILLER_78_568 ();
 sg13g2_decap_8 FILLER_78_575 ();
 sg13g2_decap_8 FILLER_78_582 ();
 sg13g2_decap_8 FILLER_78_589 ();
 sg13g2_decap_8 FILLER_78_596 ();
 sg13g2_decap_8 FILLER_78_603 ();
 sg13g2_decap_8 FILLER_78_610 ();
 sg13g2_decap_8 FILLER_78_617 ();
 sg13g2_decap_8 FILLER_78_624 ();
 sg13g2_decap_8 FILLER_78_631 ();
 sg13g2_decap_8 FILLER_78_638 ();
 sg13g2_decap_8 FILLER_78_645 ();
 sg13g2_decap_8 FILLER_78_652 ();
 sg13g2_decap_8 FILLER_78_659 ();
 sg13g2_decap_8 FILLER_78_666 ();
 sg13g2_decap_8 FILLER_78_673 ();
 sg13g2_decap_8 FILLER_78_680 ();
 sg13g2_decap_8 FILLER_78_687 ();
 sg13g2_decap_8 FILLER_78_694 ();
 sg13g2_decap_8 FILLER_78_701 ();
 sg13g2_decap_8 FILLER_78_708 ();
 sg13g2_decap_8 FILLER_78_715 ();
 sg13g2_decap_8 FILLER_78_722 ();
 sg13g2_decap_8 FILLER_78_729 ();
 sg13g2_decap_8 FILLER_78_736 ();
 sg13g2_decap_8 FILLER_78_743 ();
 sg13g2_decap_8 FILLER_78_750 ();
 sg13g2_decap_8 FILLER_78_757 ();
 sg13g2_decap_8 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_771 ();
 sg13g2_decap_8 FILLER_78_778 ();
 sg13g2_decap_8 FILLER_78_785 ();
 sg13g2_decap_8 FILLER_78_792 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_806 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_8 FILLER_78_820 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_4 FILLER_79_42 ();
 sg13g2_fill_1 FILLER_79_46 ();
 sg13g2_fill_2 FILLER_79_55 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_fill_2 FILLER_79_84 ();
 sg13g2_fill_2 FILLER_79_109 ();
 sg13g2_fill_1 FILLER_79_111 ();
 sg13g2_fill_2 FILLER_79_129 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_fill_2 FILLER_79_196 ();
 sg13g2_fill_1 FILLER_79_198 ();
 sg13g2_decap_4 FILLER_79_202 ();
 sg13g2_fill_1 FILLER_79_206 ();
 sg13g2_decap_8 FILLER_79_211 ();
 sg13g2_decap_8 FILLER_79_222 ();
 sg13g2_decap_8 FILLER_79_229 ();
 sg13g2_decap_8 FILLER_79_236 ();
 sg13g2_fill_2 FILLER_79_243 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_decap_8 FILLER_79_511 ();
 sg13g2_decap_8 FILLER_79_518 ();
 sg13g2_decap_8 FILLER_79_525 ();
 sg13g2_decap_8 FILLER_79_532 ();
 sg13g2_decap_8 FILLER_79_539 ();
 sg13g2_decap_8 FILLER_79_546 ();
 sg13g2_decap_8 FILLER_79_553 ();
 sg13g2_decap_8 FILLER_79_560 ();
 sg13g2_decap_8 FILLER_79_567 ();
 sg13g2_decap_8 FILLER_79_574 ();
 sg13g2_decap_8 FILLER_79_581 ();
 sg13g2_decap_8 FILLER_79_588 ();
 sg13g2_decap_8 FILLER_79_595 ();
 sg13g2_decap_8 FILLER_79_602 ();
 sg13g2_decap_8 FILLER_79_609 ();
 sg13g2_decap_8 FILLER_79_616 ();
 sg13g2_decap_8 FILLER_79_623 ();
 sg13g2_decap_8 FILLER_79_630 ();
 sg13g2_decap_8 FILLER_79_637 ();
 sg13g2_decap_8 FILLER_79_644 ();
 sg13g2_decap_8 FILLER_79_651 ();
 sg13g2_decap_8 FILLER_79_658 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_8 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_679 ();
 sg13g2_decap_8 FILLER_79_686 ();
 sg13g2_decap_8 FILLER_79_693 ();
 sg13g2_decap_8 FILLER_79_700 ();
 sg13g2_decap_8 FILLER_79_707 ();
 sg13g2_decap_8 FILLER_79_714 ();
 sg13g2_decap_8 FILLER_79_721 ();
 sg13g2_decap_8 FILLER_79_728 ();
 sg13g2_decap_8 FILLER_79_735 ();
 sg13g2_decap_8 FILLER_79_742 ();
 sg13g2_decap_8 FILLER_79_749 ();
 sg13g2_decap_8 FILLER_79_756 ();
 sg13g2_decap_8 FILLER_79_763 ();
 sg13g2_decap_8 FILLER_79_770 ();
 sg13g2_decap_8 FILLER_79_777 ();
 sg13g2_decap_8 FILLER_79_784 ();
 sg13g2_decap_8 FILLER_79_791 ();
 sg13g2_decap_8 FILLER_79_798 ();
 sg13g2_decap_8 FILLER_79_805 ();
 sg13g2_decap_8 FILLER_79_812 ();
 sg13g2_decap_8 FILLER_79_819 ();
 sg13g2_decap_8 FILLER_79_826 ();
 sg13g2_decap_8 FILLER_79_833 ();
 sg13g2_decap_8 FILLER_79_840 ();
 sg13g2_decap_8 FILLER_79_847 ();
 sg13g2_decap_8 FILLER_79_854 ();
 sg13g2_fill_1 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_fill_2 FILLER_80_92 ();
 sg13g2_fill_2 FILLER_80_118 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_4 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_fill_2 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_decap_4 FILLER_80_276 ();
 sg13g2_decap_4 FILLER_80_284 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_295 ();
 sg13g2_fill_2 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_303 ();
 sg13g2_fill_2 FILLER_80_309 ();
 sg13g2_fill_1 FILLER_80_311 ();
 sg13g2_decap_4 FILLER_80_316 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_decap_8 FILLER_80_429 ();
 sg13g2_decap_8 FILLER_80_436 ();
 sg13g2_decap_8 FILLER_80_443 ();
 sg13g2_decap_8 FILLER_80_450 ();
 sg13g2_decap_8 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_464 ();
 sg13g2_decap_8 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_478 ();
 sg13g2_decap_8 FILLER_80_485 ();
 sg13g2_decap_8 FILLER_80_492 ();
 sg13g2_decap_8 FILLER_80_499 ();
 sg13g2_decap_8 FILLER_80_506 ();
 sg13g2_decap_8 FILLER_80_513 ();
 sg13g2_decap_8 FILLER_80_520 ();
 sg13g2_decap_8 FILLER_80_527 ();
 sg13g2_decap_8 FILLER_80_534 ();
 sg13g2_decap_8 FILLER_80_541 ();
 sg13g2_decap_8 FILLER_80_548 ();
 sg13g2_decap_8 FILLER_80_555 ();
 sg13g2_decap_8 FILLER_80_562 ();
 sg13g2_decap_8 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_576 ();
 sg13g2_decap_8 FILLER_80_583 ();
 sg13g2_decap_8 FILLER_80_590 ();
 sg13g2_decap_8 FILLER_80_597 ();
 sg13g2_decap_8 FILLER_80_604 ();
 sg13g2_decap_8 FILLER_80_611 ();
 sg13g2_decap_8 FILLER_80_618 ();
 sg13g2_decap_8 FILLER_80_625 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_8 FILLER_80_639 ();
 sg13g2_decap_8 FILLER_80_646 ();
 sg13g2_decap_8 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_660 ();
 sg13g2_decap_8 FILLER_80_667 ();
 sg13g2_decap_8 FILLER_80_674 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_695 ();
 sg13g2_decap_8 FILLER_80_702 ();
 sg13g2_decap_8 FILLER_80_709 ();
 sg13g2_decap_8 FILLER_80_716 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_4 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule

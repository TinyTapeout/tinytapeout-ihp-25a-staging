module tt_um_wokwi_group_12 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire \proj_10.net10 ;
 wire \proj_10.net100 ;
 wire \proj_10.net101 ;
 wire \proj_10.net102 ;
 wire \proj_10.net103 ;
 wire \proj_10.net104 ;
 wire \proj_10.net105 ;
 wire \proj_10.net106 ;
 wire \proj_10.net107 ;
 wire \proj_10.net108 ;
 wire \proj_10.net109 ;
 wire \proj_10.net11 ;
 wire \proj_10.net110 ;
 wire \proj_10.net111 ;
 wire \proj_10.net112 ;
 wire \proj_10.net113 ;
 wire \proj_10.net114 ;
 wire \proj_10.net115 ;
 wire \proj_10.net116 ;
 wire \proj_10.net117 ;
 wire \proj_10.net118 ;
 wire \proj_10.net119 ;
 wire \proj_10.net12 ;
 wire \proj_10.net120 ;
 wire \proj_10.net121 ;
 wire \proj_10.net122 ;
 wire \proj_10.net123 ;
 wire \proj_10.net124 ;
 wire \proj_10.net125 ;
 wire \proj_10.net126 ;
 wire \proj_10.net127 ;
 wire \proj_10.net128 ;
 wire \proj_10.net129 ;
 wire \proj_10.net13 ;
 wire \proj_10.net130 ;
 wire \proj_10.net131 ;
 wire \proj_10.net132 ;
 wire \proj_10.net133 ;
 wire \proj_10.net134 ;
 wire \proj_10.net135 ;
 wire \proj_10.net136 ;
 wire \proj_10.net137 ;
 wire \proj_10.net138 ;
 wire \proj_10.net139 ;
 wire \proj_10.net14 ;
 wire \proj_10.net140 ;
 wire \proj_10.net141 ;
 wire \proj_10.net142 ;
 wire \proj_10.net143 ;
 wire \proj_10.net144 ;
 wire \proj_10.net145 ;
 wire \proj_10.net146 ;
 wire \proj_10.net147 ;
 wire \proj_10.net148 ;
 wire \proj_10.net149 ;
 wire \proj_10.net15 ;
 wire \proj_10.net150 ;
 wire \proj_10.net151 ;
 wire \proj_10.net152 ;
 wire \proj_10.net153 ;
 wire \proj_10.net154 ;
 wire \proj_10.net155 ;
 wire \proj_10.net156 ;
 wire \proj_10.net157 ;
 wire \proj_10.net158 ;
 wire \proj_10.net159 ;
 wire \proj_10.net16 ;
 wire \proj_10.net160 ;
 wire \proj_10.net161 ;
 wire \proj_10.net162 ;
 wire \proj_10.net163 ;
 wire \proj_10.net164 ;
 wire \proj_10.net165 ;
 wire \proj_10.net166 ;
 wire \proj_10.net167 ;
 wire \proj_10.net168 ;
 wire \proj_10.net169 ;
 wire \proj_10.net17 ;
 wire \proj_10.net170 ;
 wire \proj_10.net171 ;
 wire \proj_10.net172 ;
 wire \proj_10.net173 ;
 wire \proj_10.net174 ;
 wire \proj_10.net175 ;
 wire \proj_10.net176 ;
 wire \proj_10.net177 ;
 wire \proj_10.net178 ;
 wire \proj_10.net179 ;
 wire \proj_10.net180 ;
 wire \proj_10.net181 ;
 wire \proj_10.net182 ;
 wire \proj_10.net183 ;
 wire \proj_10.net184 ;
 wire \proj_10.net185 ;
 wire \proj_10.net186 ;
 wire \proj_10.net187 ;
 wire \proj_10.net188 ;
 wire \proj_10.net189 ;
 wire \proj_10.net190 ;
 wire \proj_10.net191 ;
 wire \proj_10.net192 ;
 wire \proj_10.net193 ;
 wire \proj_10.net194 ;
 wire \proj_10.net195 ;
 wire \proj_10.net196 ;
 wire \proj_10.net197 ;
 wire \proj_10.net198 ;
 wire \proj_10.net199 ;
 wire \proj_10.net200 ;
 wire \proj_10.net201 ;
 wire \proj_10.net202 ;
 wire \proj_10.net203 ;
 wire \proj_10.net204 ;
 wire \proj_10.net205 ;
 wire \proj_10.net206 ;
 wire \proj_10.net207 ;
 wire \proj_10.net208 ;
 wire \proj_10.net209 ;
 wire \proj_10.net210 ;
 wire \proj_10.net211 ;
 wire \proj_10.net212 ;
 wire \proj_10.net214 ;
 wire \proj_10.net215 ;
 wire \proj_10.net216 ;
 wire \proj_10.net217 ;
 wire \proj_10.net218 ;
 wire \proj_10.net219 ;
 wire \proj_10.net220 ;
 wire \proj_10.net23 ;
 wire \proj_10.net24 ;
 wire \proj_10.net25 ;
 wire \proj_10.net26 ;
 wire \proj_10.net27 ;
 wire \proj_10.net28 ;
 wire \proj_10.net29 ;
 wire \proj_10.net30 ;
 wire \proj_10.net31 ;
 wire \proj_10.net32 ;
 wire \proj_10.net33 ;
 wire \proj_10.net34 ;
 wire \proj_10.net35 ;
 wire \proj_10.net36 ;
 wire \proj_10.net37 ;
 wire \proj_10.net38 ;
 wire \proj_10.net39 ;
 wire \proj_10.net40 ;
 wire \proj_10.net41 ;
 wire \proj_10.net42 ;
 wire \proj_10.net43 ;
 wire \proj_10.net44 ;
 wire \proj_10.net45 ;
 wire \proj_10.net46 ;
 wire \proj_10.net47 ;
 wire \proj_10.net48 ;
 wire \proj_10.net49 ;
 wire \proj_10.net50 ;
 wire \proj_10.net51 ;
 wire \proj_10.net52 ;
 wire \proj_10.net53 ;
 wire \proj_10.net54 ;
 wire \proj_10.net55 ;
 wire \proj_10.net56 ;
 wire \proj_10.net57 ;
 wire \proj_10.net58 ;
 wire \proj_10.net59 ;
 wire \proj_10.net60 ;
 wire \proj_10.net61 ;
 wire \proj_10.net62 ;
 wire \proj_10.net63 ;
 wire \proj_10.net64 ;
 wire \proj_10.net65 ;
 wire \proj_10.net66 ;
 wire \proj_10.net67 ;
 wire \proj_10.net68 ;
 wire \proj_10.net69 ;
 wire \proj_10.net70 ;
 wire \proj_10.net71 ;
 wire \proj_10.net72 ;
 wire \proj_10.net73 ;
 wire \proj_10.net74 ;
 wire \proj_10.net76 ;
 wire \proj_10.net78 ;
 wire \proj_10.net79 ;
 wire \proj_10.net80 ;
 wire \proj_10.net81 ;
 wire \proj_10.net82 ;
 wire \proj_10.net83 ;
 wire \proj_10.net84 ;
 wire \proj_10.net85 ;
 wire \proj_10.net86 ;
 wire \proj_10.net87 ;
 wire \proj_10.net88 ;
 wire \proj_10.net89 ;
 wire \proj_10.net90 ;
 wire \proj_10.net91 ;
 wire \proj_10.net92 ;
 wire \proj_10.net93 ;
 wire \proj_10.net94 ;
 wire \proj_10.net95 ;
 wire \proj_10.net96 ;
 wire \proj_10.net97 ;
 wire \proj_10.net98 ;
 wire \proj_10.net99 ;
 wire \proj_11.net3 ;
 wire \proj_11.net4 ;
 wire \proj_11.net5 ;
 wire \proj_12.net10 ;
 wire \proj_12.net16 ;
 wire \proj_12.net17 ;
 wire \proj_12.net18 ;
 wire \proj_12.net19 ;
 wire \proj_12.net20 ;
 wire \proj_12.net21 ;
 wire \proj_12.net22 ;
 wire \proj_12.net23 ;
 wire \proj_12.net24 ;
 wire \proj_12.net25 ;
 wire \proj_12.net26 ;
 wire \proj_12.net27 ;
 wire \proj_12.net9 ;
 wire \proj_13.net11 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net14 ;
 wire \proj_13.net15 ;
 wire \proj_13.net16 ;
 wire \proj_13.net17 ;
 wire \proj_13.net18 ;
 wire \proj_13.net20 ;
 wire \proj_13.net9 ;
 wire \proj__0.net15 ;
 wire \proj__0.net16 ;
 wire \proj__0.net17 ;
 wire \proj__0.net18 ;
 wire \proj__0.net19 ;
 wire \proj__0.net20 ;
 wire \proj__0.net21 ;
 wire \proj__0.net22 ;
 wire \proj__0.net23 ;
 wire \proj__0.net24 ;
 wire \proj__0.net25 ;
 wire \proj__0.net26 ;
 wire \proj__0.net27 ;
 wire \proj__0.net28 ;
 wire \proj__0.net29 ;
 wire \proj__0.net30 ;
 wire \proj__0.net9 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net9 ;
 wire \proj__2.net10 ;
 wire \proj__2.net11 ;
 wire \proj__2.net12 ;
 wire \proj__2.net13 ;
 wire \proj__2.net19 ;
 wire \proj__2.net20 ;
 wire \proj__2.net21 ;
 wire \proj__2.net22 ;
 wire \proj__2.net23 ;
 wire \proj__2.net24 ;
 wire \proj__2.net25 ;
 wire \proj__2.net26 ;
 wire \proj__2.net27 ;
 wire \proj__2.net28 ;
 wire \proj__2.net29 ;
 wire \proj__2.net30 ;
 wire \proj__2.net9 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net14 ;
 wire \proj__3.net15 ;
 wire \proj__3.net21 ;
 wire \proj__3.net22 ;
 wire \proj__3.net23 ;
 wire \proj__3.net24 ;
 wire \proj__3.net25 ;
 wire \proj__3.net26 ;
 wire \proj__4.net10 ;
 wire \proj__4.net9 ;
 wire \proj__5.net6 ;
 wire \proj__5.net7 ;
 wire \proj__5.net8 ;
 wire \proj__6.net10 ;
 wire \proj__6.net16 ;
 wire \proj__6.net17 ;
 wire \proj__6.net18 ;
 wire \proj__6.net19 ;
 wire \proj__6.net20 ;
 wire \proj__6.net21 ;
 wire \proj__6.net22 ;
 wire \proj__6.net23 ;
 wire \proj__6.net7 ;
 wire \proj__6.net8 ;
 wire \proj__6.net9 ;
 wire \proj__7.net10 ;
 wire \proj__7.net11 ;
 wire \proj__7.net12 ;
 wire \proj__7.net9 ;
 wire \proj__8.net7 ;
 wire \proj__9.net10 ;
 wire \proj__9.net100 ;
 wire \proj__9.net101 ;
 wire \proj__9.net102 ;
 wire \proj__9.net103 ;
 wire \proj__9.net104 ;
 wire \proj__9.net105 ;
 wire \proj__9.net106 ;
 wire \proj__9.net107 ;
 wire \proj__9.net108 ;
 wire \proj__9.net109 ;
 wire \proj__9.net11 ;
 wire \proj__9.net110 ;
 wire \proj__9.net111 ;
 wire \proj__9.net112 ;
 wire \proj__9.net113 ;
 wire \proj__9.net114 ;
 wire \proj__9.net12 ;
 wire \proj__9.net13 ;
 wire \proj__9.net14 ;
 wire \proj__9.net15 ;
 wire \proj__9.net16 ;
 wire \proj__9.net22 ;
 wire \proj__9.net23 ;
 wire \proj__9.net24 ;
 wire \proj__9.net25 ;
 wire \proj__9.net26 ;
 wire \proj__9.net27 ;
 wire \proj__9.net28 ;
 wire \proj__9.net29 ;
 wire \proj__9.net30 ;
 wire \proj__9.net31 ;
 wire \proj__9.net32 ;
 wire \proj__9.net33 ;
 wire \proj__9.net34 ;
 wire \proj__9.net35 ;
 wire \proj__9.net36 ;
 wire \proj__9.net37 ;
 wire \proj__9.net38 ;
 wire \proj__9.net39 ;
 wire \proj__9.net40 ;
 wire \proj__9.net41 ;
 wire \proj__9.net42 ;
 wire \proj__9.net43 ;
 wire \proj__9.net44 ;
 wire \proj__9.net45 ;
 wire \proj__9.net46 ;
 wire \proj__9.net47 ;
 wire \proj__9.net48 ;
 wire \proj__9.net49 ;
 wire \proj__9.net50 ;
 wire \proj__9.net51 ;
 wire \proj__9.net52 ;
 wire \proj__9.net53 ;
 wire \proj__9.net54 ;
 wire \proj__9.net55 ;
 wire \proj__9.net56 ;
 wire \proj__9.net57 ;
 wire \proj__9.net58 ;
 wire \proj__9.net59 ;
 wire \proj__9.net60 ;
 wire \proj__9.net61 ;
 wire \proj__9.net62 ;
 wire \proj__9.net64 ;
 wire \proj__9.net65 ;
 wire \proj__9.net66 ;
 wire \proj__9.net67 ;
 wire \proj__9.net68 ;
 wire \proj__9.net69 ;
 wire \proj__9.net70 ;
 wire \proj__9.net71 ;
 wire \proj__9.net72 ;
 wire \proj__9.net73 ;
 wire \proj__9.net74 ;
 wire \proj__9.net75 ;
 wire \proj__9.net76 ;
 wire \proj__9.net77 ;
 wire \proj__9.net78 ;
 wire \proj__9.net79 ;
 wire \proj__9.net80 ;
 wire \proj__9.net81 ;
 wire \proj__9.net82 ;
 wire \proj__9.net83 ;
 wire \proj__9.net84 ;
 wire \proj__9.net85 ;
 wire \proj__9.net86 ;
 wire \proj__9.net87 ;
 wire \proj__9.net88 ;
 wire \proj__9.net89 ;
 wire \proj__9.net9 ;
 wire \proj__9.net90 ;
 wire \proj__9.net91 ;
 wire \proj__9.net92 ;
 wire \proj__9.net93 ;
 wire \proj__9.net94 ;
 wire \proj__9.net95 ;
 wire \proj__9.net96 ;
 wire \proj__9.net97 ;
 wire \proj__9.net98 ;
 wire \proj__9.net99 ;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire \proj_10.flop1/notq ;
 wire net59;
 wire \proj_10.flop10/notq ;
 wire net60;
 wire \proj_10.flop11/notq ;
 wire net61;
 wire \proj_10.flop12/notq ;
 wire net62;
 wire \proj_10.flop13/notq ;
 wire net63;
 wire \proj_10.flop14/notq ;
 wire net64;
 wire \proj_10.flop15/notq ;
 wire net65;
 wire \proj_10.flop16/notq ;
 wire net66;
 wire \proj_10.flop17/notq ;
 wire net67;
 wire \proj_10.flop18/notq ;
 wire net68;
 wire \proj_10.flop19/notq ;
 wire net69;
 wire \proj_10.flop2/notq ;
 wire net70;
 wire \proj_10.flop20/notq ;
 wire net71;
 wire \proj_10.flop21/notq ;
 wire net72;
 wire \proj_10.flop22/notq ;
 wire net73;
 wire \proj_10.flop23/notq ;
 wire net74;
 wire \proj_10.flop24/notq ;
 wire net75;
 wire \proj_10.flop3/notq ;
 wire net76;
 wire \proj_10.flop4/notq ;
 wire net77;
 wire \proj_10.flop5/notq ;
 wire net78;
 wire \proj_10.flop6/notq ;
 wire net79;
 wire \proj_10.flop7/notq ;
 wire net80;
 wire \proj_10.flop8/notq ;
 wire \proj_10.flop9/notq ;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;

 sg13g2_a221oi_1 _098_ (.B2(\proj__3.net11 ),
    .C1(_046_),
    .B1(_048_),
    .A1(\proj__1.net9 ),
    .Y(_049_),
    .A2(_047_));
 sg13g2_and2_2 _099_ (.A(_033_),
    .B(_039_),
    .X(_050_));
 sg13g2_and2_1 _100_ (.A(_033_),
    .B(_041_),
    .X(_051_));
 sg13g2_nand2_1 _101_ (.Y(_052_),
    .A(_033_),
    .B(_041_));
 sg13g2_and4_1 _102_ (.A(net3),
    .B(net4),
    .C(\proj_12.net9 ),
    .D(_041_),
    .X(_053_));
 sg13g2_a221oi_1 _103_ (.B2(\proj__8.net7 ),
    .C1(_053_),
    .B1(_051_),
    .A1(\proj__9.net9 ),
    .Y(_054_),
    .A2(_050_));
 sg13g2_and3_2 _104_ (.X(_055_),
    .A(net2),
    .B(_032_),
    .C(_033_));
 sg13g2_and3_2 _105_ (.X(_056_),
    .A(net2),
    .B(_032_),
    .C(_045_));
 sg13g2_a22oi_1 _106_ (.Y(_057_),
    .B1(_056_),
    .B2(\proj__2.net9 ),
    .A2(_055_),
    .A1(\proj_10.net10 ));
 sg13g2_and3_1 _107_ (.X(_058_),
    .A(_049_),
    .B(_054_),
    .C(_057_));
 sg13g2_nand3_1 _108_ (.B(_044_),
    .C(_058_),
    .A(_037_),
    .Y(uo_out[0]));
 sg13g2_a22oi_1 _109_ (.Y(_059_),
    .B1(_056_),
    .B2(\proj__2.net10 ),
    .A2(_055_),
    .A1(\proj_10.net11 ));
 sg13g2_a22oi_1 _110_ (.Y(_060_),
    .B1(_043_),
    .B2(net131),
    .A2(_036_),
    .A1(\proj__6.net8 ));
 sg13g2_and4_1 _111_ (.A(net3),
    .B(net4),
    .C(\proj_12.net10 ),
    .D(_041_),
    .X(_061_));
 sg13g2_a221oi_1 _112_ (.B2(\proj__9.net10 ),
    .C1(_061_),
    .B1(_050_),
    .A1(\proj__7.net10 ),
    .Y(_000_),
    .A2(_038_));
 sg13g2_nand4_1 _113_ (.B(_059_),
    .C(_060_),
    .A(_049_),
    .Y(uo_out[1]),
    .D(_000_));
 sg13g2_a22oi_1 _114_ (.Y(_001_),
    .B1(_056_),
    .B2(\proj__2.net11 ),
    .A2(_055_),
    .A1(\proj_10.net12 ));
 sg13g2_or2_1 _115_ (.X(_002_),
    .B(_047_),
    .A(_040_));
 sg13g2_a22oi_1 _116_ (.Y(_003_),
    .B1(_002_),
    .B2(net127),
    .A2(_038_),
    .A1(\proj__7.net11 ));
 sg13g2_a21o_1 _117_ (.A2(_048_),
    .A1(\proj__3.net12 ),
    .B1(_046_),
    .X(_004_));
 sg13g2_a221oi_1 _118_ (.B2(\proj__9.net11 ),
    .C1(_004_),
    .B1(_050_),
    .A1(\proj__6.net9 ),
    .Y(_005_),
    .A2(_036_));
 sg13g2_nand3_1 _119_ (.B(_003_),
    .C(_005_),
    .A(_001_),
    .Y(uo_out[2]));
 sg13g2_nand2_1 _120_ (.Y(_006_),
    .A(\proj__7.net12 ),
    .B(_038_));
 sg13g2_nand2_1 _121_ (.Y(_007_),
    .A(\proj__9.net12 ),
    .B(_050_));
 sg13g2_nand3_1 _122_ (.B(_035_),
    .C(_041_),
    .A(\proj__4.net9 ),
    .Y(_008_));
 sg13g2_and2_1 _123_ (.A(_035_),
    .B(_039_),
    .X(_009_));
 sg13g2_nand2_1 _124_ (.Y(_010_),
    .A(\proj__5.net6 ),
    .B(_009_));
 sg13g2_nand2_1 _125_ (.Y(_011_),
    .A(\proj__6.net10 ),
    .B(_036_));
 sg13g2_and2_1 _126_ (.A(net126),
    .B(_002_),
    .X(_012_));
 sg13g2_a22oi_1 _127_ (.Y(_013_),
    .B1(_056_),
    .B2(\proj__2.net12 ),
    .A2(_055_),
    .A1(\proj_10.net13 ));
 sg13g2_nand3_1 _128_ (.B(_010_),
    .C(_013_),
    .A(_006_),
    .Y(_014_));
 sg13g2_nand3_1 _129_ (.B(_008_),
    .C(_011_),
    .A(_007_),
    .Y(_015_));
 sg13g2_or4_1 _130_ (.A(_004_),
    .B(_012_),
    .C(_014_),
    .D(_015_),
    .X(uo_out[3]));
 sg13g2_nand3b_1 _131_ (.B(_042_),
    .C(_052_),
    .Y(_016_),
    .A_N(_038_));
 sg13g2_o21ai_1 _132_ (.B1(net123),
    .Y(_017_),
    .A1(_002_),
    .A2(_016_));
 sg13g2_a21oi_1 _133_ (.A1(\proj__3.net13 ),
    .A2(_048_),
    .Y(_018_),
    .B1(_046_));
 sg13g2_a22oi_1 _134_ (.Y(_019_),
    .B1(_056_),
    .B2(\proj__2.net13 ),
    .A2(_034_),
    .A1(net130));
 sg13g2_a22oi_1 _135_ (.Y(_020_),
    .B1(_055_),
    .B2(\proj_10.net14 ),
    .A2(_050_),
    .A1(\proj__9.net13 ));
 sg13g2_nand4_1 _136_ (.B(_018_),
    .C(_019_),
    .A(_017_),
    .Y(uo_out[4]),
    .D(_020_));
 sg13g2_o21ai_1 _137_ (.B1(net119),
    .Y(_021_),
    .A1(_040_),
    .A2(_016_));
 sg13g2_a22oi_1 _138_ (.Y(_022_),
    .B1(_055_),
    .B2(\proj_10.net15 ),
    .A2(_047_),
    .A1(\proj__1.net10 ));
 sg13g2_a22oi_1 _139_ (.Y(_023_),
    .B1(_009_),
    .B2(\proj__5.net7 ),
    .A2(_050_),
    .A1(\proj__9.net14 ));
 sg13g2_nand4_1 _140_ (.B(_021_),
    .C(_022_),
    .A(_018_),
    .Y(uo_out[5]),
    .D(_023_));
 sg13g2_o21ai_1 _141_ (.B1(net115),
    .Y(_024_),
    .A1(_040_),
    .A2(_016_));
 sg13g2_a21oi_1 _142_ (.A1(\proj__1.net11 ),
    .A2(_047_),
    .Y(_025_),
    .B1(_046_));
 sg13g2_nand2_1 _143_ (.Y(_026_),
    .A(\proj_10.net16 ),
    .B(_055_));
 sg13g2_a22oi_1 _144_ (.Y(_027_),
    .B1(_050_),
    .B2(\proj__9.net15 ),
    .A2(_048_),
    .A1(\proj__3.net14 ));
 sg13g2_nand4_1 _145_ (.B(_025_),
    .C(_026_),
    .A(_024_),
    .Y(uo_out[6]),
    .D(_027_));
 sg13g2_a22oi_1 _146_ (.Y(_028_),
    .B1(_040_),
    .B2(\proj_13.net9 ),
    .A2(_034_),
    .A1(\proj_11.net4 ));
 sg13g2_a22oi_1 _147_ (.Y(_029_),
    .B1(_055_),
    .B2(\proj_10.net17 ),
    .A2(_050_),
    .A1(\proj__9.net16 ));
 sg13g2_a22oi_1 _148_ (.Y(_030_),
    .B1(_009_),
    .B2(\proj__5.net8 ),
    .A2(_048_),
    .A1(\proj__3.net15 ));
 sg13g2_nand4_1 _149_ (.B(_028_),
    .C(_029_),
    .A(_025_),
    .Y(_031_),
    .D(_030_));
 sg13g2_a21o_2 _150_ (.A2(_016_),
    .A1(net108),
    .B1(_031_),
    .X(uo_out[7]));
 sg13g2_inv_1 _151_ (.Y(_032_),
    .A(net1));
 sg13g2_nor2b_2 _152_ (.A(net3),
    .B_N(net4),
    .Y(_033_));
 sg13g2_and3_1 _153_ (.X(_034_),
    .A(net2),
    .B(net1),
    .C(_033_));
 sg13g2_nor2b_2 _154_ (.A(net4),
    .B_N(net3),
    .Y(_035_));
 sg13g2_and3_2 _155_ (.X(_036_),
    .A(net2),
    .B(_032_),
    .C(_035_));
 sg13g2_a22oi_1 _156_ (.Y(_037_),
    .B1(_036_),
    .B2(\proj__6.net7 ),
    .A2(_034_),
    .A1(\proj_11.net3 ));
 sg13g2_and3_2 _157_ (.X(_038_),
    .A(net2),
    .B(net1),
    .C(_035_));
 sg13g2_nor2b_1 _158_ (.A(net2),
    .B_N(net1),
    .Y(_039_));
 sg13g2_and3_2 _159_ (.X(_040_),
    .A(net3),
    .B(net4),
    .C(_039_));
 sg13g2_nor2_2 _160_ (.A(net2),
    .B(net1),
    .Y(_041_));
 sg13g2_nand2_1 _161_ (.Y(_042_),
    .A(_035_),
    .B(_041_));
 sg13g2_nand2b_1 _162_ (.Y(_043_),
    .B(_042_),
    .A_N(_040_));
 sg13g2_a22oi_1 _163_ (.Y(_044_),
    .B1(_043_),
    .B2(net136),
    .A2(_038_),
    .A1(\proj__7.net9 ));
 sg13g2_nor2_1 _164_ (.A(net3),
    .B(net4),
    .Y(_045_));
 sg13g2_and3_1 _165_ (.X(_046_),
    .A(\proj__0.net9 ),
    .B(_041_),
    .C(_045_));
 sg13g2_and2_1 _166_ (.A(_039_),
    .B(_045_),
    .X(_047_));
 sg13g2_and3_2 _167_ (.X(_048_),
    .A(net2),
    .B(net1),
    .C(_045_));
 sg13g2_tielo \proj_10.flop10/_1__6  (.L_LO(net6));
 sg13g2_tielo \proj_10.flop11/_1__7  (.L_LO(net7));
 sg13g2_tielo \proj_10.flop12/_1__8  (.L_LO(net8));
 sg13g2_tielo \proj_10.flop13/_1__9  (.L_LO(net9));
 sg13g2_tielo \proj_10.flop14/_1__10  (.L_LO(net10));
 sg13g2_tielo \proj_10.flop15/_1__11  (.L_LO(net11));
 sg13g2_tielo \proj_10.flop16/_1__12  (.L_LO(net12));
 sg13g2_tielo \proj_10.flop17/_1__13  (.L_LO(net13));
 sg13g2_tielo \proj_10.flop18/_1__14  (.L_LO(net14));
 sg13g2_tielo \proj_10.flop19/_1__15  (.L_LO(net15));
 sg13g2_tielo \proj_10.flop2/_1__16  (.L_LO(net16));
 sg13g2_tielo \proj_10.flop20/_1__17  (.L_LO(net17));
 sg13g2_tielo \proj_10.flop21/_1__18  (.L_LO(net18));
 sg13g2_tielo \proj_10.flop22/_1__19  (.L_LO(net19));
 sg13g2_tielo \proj_10.flop23/_1__20  (.L_LO(net20));
 sg13g2_tielo \proj_10.flop24/_1__21  (.L_LO(net21));
 sg13g2_tielo \proj_10.flop3/_1__22  (.L_LO(net22));
 sg13g2_tielo \proj_10.flop4/_1__23  (.L_LO(net23));
 sg13g2_tielo \proj_10.flop5/_1__24  (.L_LO(net24));
 sg13g2_tielo \proj_10.flop6/_1__25  (.L_LO(net25));
 sg13g2_tielo \proj_10.flop7/_1__26  (.L_LO(net26));
 sg13g2_tielo \proj_10.flop8/_1__27  (.L_LO(net27));
 sg13g2_tielo \proj_10.flop9/_1__28  (.L_LO(net28));
 sg13g2_tielo \proj_10.or49/_0__29  (.L_LO(net29));
 sg13g2_tielo \proj_10.or50/_0__30  (.L_LO(net30));
 sg13g2_tielo \proj_10.or51/_0__31  (.L_LO(net31));
 sg13g2_tielo \proj_10.or52/_0__32  (.L_LO(net32));
 sg13g2_tielo \proj_10.or53/_0__33  (.L_LO(net33));
 sg13g2_tielo \proj_10.or54/_0__34  (.L_LO(net34));
 sg13g2_tielo \proj_10.or55/_0__35  (.L_LO(net35));
 sg13g2_tielo \proj_10.or56/_0__36  (.L_LO(net36));
 sg13g2_tielo \proj__3.not1/_0__37  (.L_LO(net37));
 sg13g2_tielo \proj__3.xor1/_0__38  (.L_LO(net38));
 sg13g2_tielo \proj__9.and19/_0__39  (.L_LO(net39));
 sg13g2_tielo \proj__9.xor4/_0__40  (.L_LO(net40));
 sg13g2_tielo tt_um_wokwi_group_12_41 (.L_LO(net41));
 sg13g2_tielo tt_um_wokwi_group_12_42 (.L_LO(net42));
 sg13g2_tielo tt_um_wokwi_group_12_43 (.L_LO(net43));
 sg13g2_tielo tt_um_wokwi_group_12_44 (.L_LO(net44));
 sg13g2_tielo tt_um_wokwi_group_12_45 (.L_LO(net45));
 sg13g2_tielo tt_um_wokwi_group_12_46 (.L_LO(net46));
 sg13g2_tielo tt_um_wokwi_group_12_47 (.L_LO(net47));
 sg13g2_tielo tt_um_wokwi_group_12_48 (.L_LO(net48));
 sg13g2_tielo tt_um_wokwi_group_12_49 (.L_LO(net49));
 sg13g2_tielo tt_um_wokwi_group_12_50 (.L_LO(net50));
 sg13g2_tielo tt_um_wokwi_group_12_51 (.L_LO(net51));
 sg13g2_tielo tt_um_wokwi_group_12_52 (.L_LO(net52));
 sg13g2_tielo tt_um_wokwi_group_12_53 (.L_LO(net53));
 sg13g2_tielo tt_um_wokwi_group_12_54 (.L_LO(net54));
 sg13g2_tielo tt_um_wokwi_group_12_55 (.L_LO(net55));
 sg13g2_tielo tt_um_wokwi_group_12_56 (.L_LO(net56));
 sg13g2_tiehi \proj_10.flop1/_1__57  (.L_HI(net57));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(net105),
    .B(\proj_10.net10 ),
    .X(\proj_10.net111 ));
 sg13g2_and2_1 \proj_10.and10/_0_  (.A(\proj_10.net46 ),
    .B(\proj_10.net43 ),
    .X(\proj_10.net49 ));
 sg13g2_and2_1 \proj_10.and11/_0_  (.A(\proj_10.net52 ),
    .B(\proj_10.net51 ),
    .X(\proj_10.net54 ));
 sg13g2_and2_1 \proj_10.and12/_0_  (.A(\proj_10.net53 ),
    .B(\proj_10.net50 ),
    .X(\proj_10.net56 ));
 sg13g2_and2_1 \proj_10.and13/_0_  (.A(\proj_10.net59 ),
    .B(\proj_10.net58 ),
    .X(\proj_10.net61 ));
 sg13g2_and2_1 \proj_10.and14/_0_  (.A(\proj_10.net60 ),
    .B(\proj_10.net57 ),
    .X(\proj_10.net63 ));
 sg13g2_and2_1 \proj_10.and15/_0_  (.A(\proj_10.net66 ),
    .B(\proj_10.net65 ),
    .X(\proj_10.net68 ));
 sg13g2_and2_1 \proj_10.and16/_0_  (.A(\proj_10.net67 ),
    .B(\proj_10.net64 ),
    .X(\proj_10.net70 ));
 sg13g2_and2_1 \proj_10.and19/_0_  (.A(net105),
    .B(\proj_10.net12 ),
    .X(\proj_10.net113 ));
 sg13g2_and2_1 \proj_10.and2/_0_  (.A(net105),
    .B(\proj_10.net11 ),
    .X(\proj_10.net112 ));
 sg13g2_and2_1 \proj_10.and20/_0_  (.A(net105),
    .B(\proj_10.net13 ),
    .X(\proj_10.net114 ));
 sg13g2_and2_1 \proj_10.and21/_0_  (.A(\proj_10.net110 ),
    .B(\proj_10.net14 ),
    .X(\proj_10.net115 ));
 sg13g2_and2_1 \proj_10.and22/_0_  (.A(net105),
    .B(\proj_10.net15 ),
    .X(\proj_10.net116 ));
 sg13g2_and2_1 \proj_10.and23/_0_  (.A(net105),
    .B(\proj_10.net16 ),
    .X(\proj_10.net117 ));
 sg13g2_and2_1 \proj_10.and24/_0_  (.A(net105),
    .B(\proj_10.net17 ),
    .X(\proj_10.net118 ));
 sg13g2_and2_1 \proj_10.and25/_0_  (.A(\proj_10.net119 ),
    .B(\proj_10.net23 ),
    .X(\proj_10.net120 ));
 sg13g2_and2_1 \proj_10.and26/_0_  (.A(\proj_10.net119 ),
    .B(\proj_10.net30 ),
    .X(\proj_10.net121 ));
 sg13g2_and2_1 \proj_10.and27/_0_  (.A(\proj_10.net119 ),
    .B(\proj_10.net37 ),
    .X(\proj_10.net122 ));
 sg13g2_and2_1 \proj_10.and28/_0_  (.A(\proj_10.net119 ),
    .B(\proj_10.net44 ),
    .X(\proj_10.net123 ));
 sg13g2_and2_1 \proj_10.and29/_0_  (.A(\proj_10.net119 ),
    .B(\proj_10.net51 ),
    .X(\proj_10.net124 ));
 sg13g2_and2_1 \proj_10.and3/_0_  (.A(\proj_10.net24 ),
    .B(\proj_10.net23 ),
    .X(\proj_10.net26 ));
 sg13g2_and2_1 \proj_10.and30/_0_  (.A(\proj_10.net119 ),
    .B(\proj_10.net58 ),
    .X(\proj_10.net125 ));
 sg13g2_and2_1 \proj_10.and31/_0_  (.A(\proj_10.net119 ),
    .B(\proj_10.net65 ),
    .X(\proj_10.net126 ));
 sg13g2_and2_1 \proj_10.and32/_0_  (.A(\proj_10.net119 ),
    .B(\proj_10.net72 ),
    .X(\proj_10.net127 ));
 sg13g2_and2_1 \proj_10.and33/_0_  (.A(net131),
    .B(\proj_10.net102 ),
    .X(\proj_10.net136 ));
 sg13g2_and2_1 \proj_10.and34/_0_  (.A(net131),
    .B(\proj_10.net103 ),
    .X(\proj_10.net137 ));
 sg13g2_and2_1 \proj_10.and35/_0_  (.A(net131),
    .B(\proj_10.net104 ),
    .X(\proj_10.net138 ));
 sg13g2_and2_1 \proj_10.and36/_0_  (.A(net131),
    .B(\proj_10.net105 ),
    .X(\proj_10.net139 ));
 sg13g2_and2_1 \proj_10.and37/_0_  (.A(net133),
    .B(\proj_10.net106 ),
    .X(\proj_10.net140 ));
 sg13g2_and2_1 \proj_10.and38/_0_  (.A(net133),
    .B(\proj_10.net107 ),
    .X(\proj_10.net141 ));
 sg13g2_and2_1 \proj_10.and39/_0_  (.A(net133),
    .B(\proj_10.net108 ),
    .X(\proj_10.net142 ));
 sg13g2_and2_1 \proj_10.and4/_0_  (.A(\proj_10.net25 ),
    .B(net107),
    .X(\proj_10.net28 ));
 sg13g2_and2_1 \proj_10.and40/_0_  (.A(net133),
    .B(\proj_10.net109 ),
    .X(\proj_10.net143 ));
 sg13g2_and2_1 \proj_10.and41/_0_  (.A(net106),
    .B(\proj_10.net10 ),
    .X(\proj_10.net145 ));
 sg13g2_and2_1 \proj_10.and42/_0_  (.A(net106),
    .B(\proj_10.net11 ),
    .X(\proj_10.net146 ));
 sg13g2_and2_1 \proj_10.and43/_0_  (.A(net106),
    .B(\proj_10.net12 ),
    .X(\proj_10.net147 ));
 sg13g2_and2_1 \proj_10.and44/_0_  (.A(\proj_10.net144 ),
    .B(\proj_10.net13 ),
    .X(\proj_10.net148 ));
 sg13g2_and2_1 \proj_10.and45/_0_  (.A(net106),
    .B(\proj_10.net14 ),
    .X(\proj_10.net149 ));
 sg13g2_and2_1 \proj_10.and46/_0_  (.A(net106),
    .B(\proj_10.net15 ),
    .X(\proj_10.net150 ));
 sg13g2_and2_1 \proj_10.and47/_0_  (.A(net106),
    .B(\proj_10.net16 ),
    .X(\proj_10.net151 ));
 sg13g2_and2_1 \proj_10.and48/_0_  (.A(net106),
    .B(\proj_10.net17 ),
    .X(\proj_10.net152 ));
 sg13g2_and2_1 \proj_10.and49/_0_  (.A(\proj_10.net153 ),
    .B(\proj_10.net87 ),
    .X(\proj_10.net154 ));
 sg13g2_and2_1 \proj_10.and5/_0_  (.A(\proj_10.net31 ),
    .B(\proj_10.net30 ),
    .X(\proj_10.net33 ));
 sg13g2_and2_1 \proj_10.and50/_0_  (.A(\proj_10.net153 ),
    .B(\proj_10.net89 ),
    .X(\proj_10.net155 ));
 sg13g2_and2_1 \proj_10.and51/_0_  (.A(\proj_10.net153 ),
    .B(\proj_10.net91 ),
    .X(\proj_10.net156 ));
 sg13g2_and2_1 \proj_10.and52/_0_  (.A(\proj_10.net153 ),
    .B(\proj_10.net93 ),
    .X(\proj_10.net157 ));
 sg13g2_and2_1 \proj_10.and53/_0_  (.A(\proj_10.net153 ),
    .B(\proj_10.net95 ),
    .X(\proj_10.net158 ));
 sg13g2_and2_1 \proj_10.and54/_0_  (.A(\proj_10.net153 ),
    .B(\proj_10.net97 ),
    .X(\proj_10.net159 ));
 sg13g2_and2_1 \proj_10.and55/_0_  (.A(\proj_10.net153 ),
    .B(\proj_10.net99 ),
    .X(\proj_10.net160 ));
 sg13g2_and2_1 \proj_10.and56/_0_  (.A(\proj_10.net153 ),
    .B(\proj_10.net101 ),
    .X(\proj_10.net161 ));
 sg13g2_and2_1 \proj_10.and57/_0_  (.A(net112),
    .B(\proj_10.net145 ),
    .X(\proj_10.net170 ));
 sg13g2_and2_1 \proj_10.and58/_0_  (.A(\proj_10.net87 ),
    .B(\proj_10.net172 ),
    .X(\proj_10.net171 ));
 sg13g2_and2_1 \proj_10.and59/_0_  (.A(net112),
    .B(\proj_10.net146 ),
    .X(\proj_10.net173 ));
 sg13g2_and2_1 \proj_10.and6/_0_  (.A(\proj_10.net32 ),
    .B(\proj_10.net29 ),
    .X(\proj_10.net35 ));
 sg13g2_and2_1 \proj_10.and60/_0_  (.A(\proj_10.net89 ),
    .B(\proj_10.net172 ),
    .X(\proj_10.net174 ));
 sg13g2_and2_1 \proj_10.and61/_0_  (.A(net112),
    .B(\proj_10.net147 ),
    .X(\proj_10.net175 ));
 sg13g2_and2_1 \proj_10.and62/_0_  (.A(\proj_10.net91 ),
    .B(\proj_10.net172 ),
    .X(\proj_10.net176 ));
 sg13g2_and2_1 \proj_10.and63/_0_  (.A(net112),
    .B(\proj_10.net148 ),
    .X(\proj_10.net177 ));
 sg13g2_and2_1 \proj_10.and64/_0_  (.A(\proj_10.net93 ),
    .B(\proj_10.net172 ),
    .X(\proj_10.net178 ));
 sg13g2_and2_1 \proj_10.and65/_0_  (.A(net114),
    .B(\proj_10.net149 ),
    .X(\proj_10.net179 ));
 sg13g2_and2_1 \proj_10.and66/_0_  (.A(\proj_10.net95 ),
    .B(\proj_10.net172 ),
    .X(\proj_10.net180 ));
 sg13g2_and2_1 \proj_10.and67/_0_  (.A(net114),
    .B(\proj_10.net150 ),
    .X(\proj_10.net181 ));
 sg13g2_and2_1 \proj_10.and68/_0_  (.A(\proj_10.net97 ),
    .B(\proj_10.net172 ),
    .X(\proj_10.net182 ));
 sg13g2_and2_1 \proj_10.and69/_0_  (.A(net114),
    .B(\proj_10.net151 ),
    .X(\proj_10.net183 ));
 sg13g2_and2_1 \proj_10.and7/_0_  (.A(\proj_10.net38 ),
    .B(\proj_10.net37 ),
    .X(\proj_10.net40 ));
 sg13g2_and2_1 \proj_10.and70/_0_  (.A(\proj_10.net99 ),
    .B(\proj_10.net172 ),
    .X(\proj_10.net184 ));
 sg13g2_and2_1 \proj_10.and71/_0_  (.A(net114),
    .B(\proj_10.net152 ),
    .X(\proj_10.net185 ));
 sg13g2_and2_1 \proj_10.and72/_0_  (.A(\proj_10.net101 ),
    .B(\proj_10.net172 ),
    .X(\proj_10.net186 ));
 sg13g2_and2_1 \proj_10.and73/_0_  (.A(net116),
    .B(\proj_10.net111 ),
    .X(\proj_10.net187 ));
 sg13g2_and2_1 \proj_10.and74/_0_  (.A(\proj_10.net23 ),
    .B(\proj_10.net188 ),
    .X(\proj_10.net189 ));
 sg13g2_and2_1 \proj_10.and75/_0_  (.A(net116),
    .B(\proj_10.net112 ),
    .X(\proj_10.net190 ));
 sg13g2_and2_1 \proj_10.and76/_0_  (.A(\proj_10.net30 ),
    .B(\proj_10.net188 ),
    .X(\proj_10.net191 ));
 sg13g2_and2_1 \proj_10.and77/_0_  (.A(net116),
    .B(\proj_10.net113 ),
    .X(\proj_10.net192 ));
 sg13g2_and2_1 \proj_10.and78/_0_  (.A(\proj_10.net37 ),
    .B(\proj_10.net188 ),
    .X(\proj_10.net193 ));
 sg13g2_and2_1 \proj_10.and79/_0_  (.A(net116),
    .B(\proj_10.net114 ),
    .X(\proj_10.net194 ));
 sg13g2_and2_1 \proj_10.and8/_0_  (.A(\proj_10.net39 ),
    .B(\proj_10.net36 ),
    .X(\proj_10.net42 ));
 sg13g2_and2_1 \proj_10.and80/_0_  (.A(\proj_10.net44 ),
    .B(\proj_10.net188 ),
    .X(\proj_10.net195 ));
 sg13g2_and2_1 \proj_10.and81/_0_  (.A(net118),
    .B(\proj_10.net115 ),
    .X(\proj_10.net196 ));
 sg13g2_and2_1 \proj_10.and82/_0_  (.A(\proj_10.net51 ),
    .B(\proj_10.net188 ),
    .X(\proj_10.net197 ));
 sg13g2_and2_1 \proj_10.and83/_0_  (.A(net118),
    .B(\proj_10.net116 ),
    .X(\proj_10.net198 ));
 sg13g2_and2_1 \proj_10.and84/_0_  (.A(\proj_10.net58 ),
    .B(\proj_10.net188 ),
    .X(\proj_10.net199 ));
 sg13g2_and2_1 \proj_10.and85/_0_  (.A(net118),
    .B(\proj_10.net117 ),
    .X(\proj_10.net200 ));
 sg13g2_and2_1 \proj_10.and86/_0_  (.A(\proj_10.net65 ),
    .B(\proj_10.net188 ),
    .X(\proj_10.net201 ));
 sg13g2_and2_1 \proj_10.and87/_0_  (.A(net118),
    .B(\proj_10.net118 ),
    .X(\proj_10.net202 ));
 sg13g2_and2_1 \proj_10.and88/_0_  (.A(\proj_10.net72 ),
    .B(\proj_10.net188 ),
    .X(\proj_10.net203 ));
 sg13g2_and2_1 \proj_10.and89/_0_  (.A(\proj_10.net27 ),
    .B(net120),
    .X(\proj_10.net212 ));
 sg13g2_and2_1 \proj_10.and9/_0_  (.A(\proj_10.net45 ),
    .B(\proj_10.net44 ),
    .X(\proj_10.net47 ));
 sg13g2_and2_1 \proj_10.and90/_0_  (.A(\proj_10.net34 ),
    .B(net120),
    .X(\proj_10.net214 ));
 sg13g2_and2_1 \proj_10.and91/_0_  (.A(\proj_10.net41 ),
    .B(net120),
    .X(\proj_10.net215 ));
 sg13g2_and2_1 \proj_10.and92/_0_  (.A(\proj_10.net48 ),
    .B(net120),
    .X(\proj_10.net216 ));
 sg13g2_and2_1 \proj_10.and93/_0_  (.A(\proj_10.net55 ),
    .B(net122),
    .X(\proj_10.net217 ));
 sg13g2_and2_1 \proj_10.and94/_0_  (.A(\proj_10.net62 ),
    .B(net122),
    .X(\proj_10.net218 ));
 sg13g2_and2_1 \proj_10.and95/_0_  (.A(\proj_10.net69 ),
    .B(net122),
    .X(\proj_10.net219 ));
 sg13g2_and2_1 \proj_10.and96/_0_  (.A(\proj_10.net76 ),
    .B(net122),
    .X(\proj_10.net220 ));
 sg13g2_dfrbp_1 \proj_10.flop1/_1_  (.CLK(net5),
    .RESET_B(net57),
    .D(\proj_10.net78 ),
    .Q_N(\proj_10.flop1/notq ),
    .Q(\proj_10.net23 ));
 sg13g2_tiehi \proj_10.flop10/_1__58  (.L_HI(net58));
 sg13g2_dfrbp_1 \proj_10.flop10/_1_  (.CLK(net6),
    .RESET_B(net58),
    .D(\proj_10.net88 ),
    .Q_N(\proj_10.flop10/notq ),
    .Q(\proj_10.net89 ));
 sg13g2_tiehi \proj_10.flop11/_1__59  (.L_HI(net59));
 sg13g2_dfrbp_1 \proj_10.flop11/_1_  (.CLK(net7),
    .RESET_B(net59),
    .D(\proj_10.net90 ),
    .Q_N(\proj_10.flop11/notq ),
    .Q(\proj_10.net91 ));
 sg13g2_tiehi \proj_10.flop12/_1__60  (.L_HI(net60));
 sg13g2_dfrbp_1 \proj_10.flop12/_1_  (.CLK(net8),
    .RESET_B(net60),
    .D(\proj_10.net92 ),
    .Q_N(\proj_10.flop12/notq ),
    .Q(\proj_10.net93 ));
 sg13g2_tiehi \proj_10.flop13/_1__61  (.L_HI(net61));
 sg13g2_dfrbp_1 \proj_10.flop13/_1_  (.CLK(net9),
    .RESET_B(net61),
    .D(\proj_10.net94 ),
    .Q_N(\proj_10.flop13/notq ),
    .Q(\proj_10.net95 ));
 sg13g2_tiehi \proj_10.flop14/_1__62  (.L_HI(net62));
 sg13g2_dfrbp_1 \proj_10.flop14/_1_  (.CLK(net10),
    .RESET_B(net62),
    .D(\proj_10.net96 ),
    .Q_N(\proj_10.flop14/notq ),
    .Q(\proj_10.net97 ));
 sg13g2_tiehi \proj_10.flop15/_1__63  (.L_HI(net63));
 sg13g2_dfrbp_1 \proj_10.flop15/_1_  (.CLK(net11),
    .RESET_B(net63),
    .D(\proj_10.net98 ),
    .Q_N(\proj_10.flop15/notq ),
    .Q(\proj_10.net99 ));
 sg13g2_tiehi \proj_10.flop16/_1__64  (.L_HI(net64));
 sg13g2_dfrbp_1 \proj_10.flop16/_1_  (.CLK(net12),
    .RESET_B(net64),
    .D(\proj_10.net100 ),
    .Q_N(\proj_10.flop16/notq ),
    .Q(\proj_10.net101 ));
 sg13g2_tiehi \proj_10.flop17/_1__65  (.L_HI(net65));
 sg13g2_dfrbp_1 \proj_10.flop17/_1_  (.CLK(net13),
    .RESET_B(net65),
    .D(net134),
    .Q_N(\proj_10.flop17/notq ),
    .Q(\proj_10.net102 ));
 sg13g2_tiehi \proj_10.flop18/_1__66  (.L_HI(net66));
 sg13g2_dfrbp_1 \proj_10.flop18/_1_  (.CLK(net14),
    .RESET_B(net66),
    .D(\proj_10.net102 ),
    .Q_N(\proj_10.flop18/notq ),
    .Q(\proj_10.net103 ));
 sg13g2_tiehi \proj_10.flop19/_1__67  (.L_HI(net67));
 sg13g2_dfrbp_1 \proj_10.flop19/_1_  (.CLK(net15),
    .RESET_B(net67),
    .D(\proj_10.net103 ),
    .Q_N(\proj_10.flop19/notq ),
    .Q(\proj_10.net104 ));
 sg13g2_tiehi \proj_10.flop2/_1__68  (.L_HI(net68));
 sg13g2_dfrbp_1 \proj_10.flop2/_1_  (.CLK(net16),
    .RESET_B(net68),
    .D(\proj_10.net79 ),
    .Q_N(\proj_10.flop2/notq ),
    .Q(\proj_10.net30 ));
 sg13g2_tiehi \proj_10.flop20/_1__69  (.L_HI(net69));
 sg13g2_dfrbp_1 \proj_10.flop20/_1_  (.CLK(net17),
    .RESET_B(net69),
    .D(\proj_10.net104 ),
    .Q_N(\proj_10.flop20/notq ),
    .Q(\proj_10.net105 ));
 sg13g2_tiehi \proj_10.flop21/_1__70  (.L_HI(net70));
 sg13g2_dfrbp_1 \proj_10.flop21/_1_  (.CLK(net18),
    .RESET_B(net70),
    .D(\proj_10.net105 ),
    .Q_N(\proj_10.flop21/notq ),
    .Q(\proj_10.net106 ));
 sg13g2_tiehi \proj_10.flop22/_1__71  (.L_HI(net71));
 sg13g2_dfrbp_1 \proj_10.flop22/_1_  (.CLK(net19),
    .RESET_B(net71),
    .D(\proj_10.net106 ),
    .Q_N(\proj_10.flop22/notq ),
    .Q(\proj_10.net107 ));
 sg13g2_tiehi \proj_10.flop23/_1__72  (.L_HI(net72));
 sg13g2_dfrbp_1 \proj_10.flop23/_1_  (.CLK(net20),
    .RESET_B(net72),
    .D(\proj_10.net107 ),
    .Q_N(\proj_10.flop23/notq ),
    .Q(\proj_10.net108 ));
 sg13g2_tiehi \proj_10.flop24/_1__73  (.L_HI(net73));
 sg13g2_dfrbp_1 \proj_10.flop24/_1_  (.CLK(net21),
    .RESET_B(net73),
    .D(\proj_10.net108 ),
    .Q_N(\proj_10.flop24/notq ),
    .Q(\proj_10.net109 ));
 sg13g2_tiehi \proj_10.flop3/_1__74  (.L_HI(net74));
 sg13g2_dfrbp_1 \proj_10.flop3/_1_  (.CLK(net22),
    .RESET_B(net74),
    .D(\proj_10.net80 ),
    .Q_N(\proj_10.flop3/notq ),
    .Q(\proj_10.net37 ));
 sg13g2_tiehi \proj_10.flop4/_1__75  (.L_HI(net75));
 sg13g2_dfrbp_1 \proj_10.flop4/_1_  (.CLK(net23),
    .RESET_B(net75),
    .D(\proj_10.net81 ),
    .Q_N(\proj_10.flop4/notq ),
    .Q(\proj_10.net44 ));
 sg13g2_tiehi \proj_10.flop5/_1__76  (.L_HI(net76));
 sg13g2_dfrbp_1 \proj_10.flop5/_1_  (.CLK(net24),
    .RESET_B(net76),
    .D(\proj_10.net82 ),
    .Q_N(\proj_10.flop5/notq ),
    .Q(\proj_10.net51 ));
 sg13g2_tiehi \proj_10.flop6/_1__77  (.L_HI(net77));
 sg13g2_dfrbp_1 \proj_10.flop6/_1_  (.CLK(net25),
    .RESET_B(net77),
    .D(\proj_10.net83 ),
    .Q_N(\proj_10.flop6/notq ),
    .Q(\proj_10.net58 ));
 sg13g2_tiehi \proj_10.flop7/_1__78  (.L_HI(net78));
 sg13g2_dfrbp_1 \proj_10.flop7/_1_  (.CLK(net26),
    .RESET_B(net78),
    .D(\proj_10.net84 ),
    .Q_N(\proj_10.flop7/notq ),
    .Q(\proj_10.net65 ));
 sg13g2_tiehi \proj_10.flop8/_1__79  (.L_HI(net79));
 sg13g2_dfrbp_1 \proj_10.flop8/_1_  (.CLK(net27),
    .RESET_B(net79),
    .D(\proj_10.net85 ),
    .Q_N(\proj_10.flop8/notq ),
    .Q(\proj_10.net72 ));
 sg13g2_tiehi \proj_10.flop9/_1__80  (.L_HI(net80));
 sg13g2_dfrbp_1 \proj_10.flop9/_1_  (.CLK(net28),
    .RESET_B(net80),
    .D(\proj_10.net86 ),
    .Q_N(\proj_10.flop9/notq ),
    .Q(\proj_10.net87 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_inv_2 \proj_10.not1/_0_  (.Y(\proj_10.net119 ),
    .A(net105));
 sg13g2_inv_2 \proj_10.not2/_0_  (.Y(\proj_10.net153 ),
    .A(net106));
 sg13g2_inv_1 \proj_10.not3/_0_  (.Y(\proj_10.net144 ),
    .A(net124));
 sg13g2_inv_1 \proj_10.not4/_0_  (.Y(\proj_10.net110 ),
    .A(net127));
 sg13g2_inv_2 \proj_10.not5/_0_  (.Y(\proj_10.net172 ),
    .A(net114));
 sg13g2_inv_2 \proj_10.not6/_0_  (.Y(\proj_10.net188 ),
    .A(net116));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net10 ),
    .B(\proj_10.net128 ),
    .A(\proj_10.net120 ));
 sg13g2_or2_1 \proj_10.or10/_0_  (.X(\proj_10.net11 ),
    .B(\proj_10.net129 ),
    .A(\proj_10.net121 ));
 sg13g2_or2_1 \proj_10.or11/_0_  (.X(\proj_10.net12 ),
    .B(\proj_10.net130 ),
    .A(\proj_10.net122 ));
 sg13g2_or2_1 \proj_10.or12/_0_  (.X(\proj_10.net13 ),
    .B(\proj_10.net131 ),
    .A(\proj_10.net123 ));
 sg13g2_or2_1 \proj_10.or13/_0_  (.X(\proj_10.net14 ),
    .B(\proj_10.net132 ),
    .A(\proj_10.net124 ));
 sg13g2_or2_1 \proj_10.or14/_0_  (.X(\proj_10.net15 ),
    .B(\proj_10.net133 ),
    .A(\proj_10.net125 ));
 sg13g2_or2_1 \proj_10.or15/_0_  (.X(\proj_10.net16 ),
    .B(\proj_10.net134 ),
    .A(\proj_10.net126 ));
 sg13g2_or2_1 \proj_10.or16/_0_  (.X(\proj_10.net17 ),
    .B(\proj_10.net135 ),
    .A(\proj_10.net127 ));
 sg13g2_or2_1 \proj_10.or17/_0_  (.X(\proj_10.net128 ),
    .B(\proj_10.net162 ),
    .A(\proj_10.net136 ));
 sg13g2_or2_1 \proj_10.or18/_0_  (.X(\proj_10.net129 ),
    .B(\proj_10.net163 ),
    .A(\proj_10.net137 ));
 sg13g2_or2_1 \proj_10.or19/_0_  (.X(\proj_10.net130 ),
    .B(\proj_10.net164 ),
    .A(\proj_10.net138 ));
 sg13g2_or2_1 \proj_10.or2/_0_  (.X(\proj_10.net29 ),
    .B(\proj_10.net26 ),
    .A(\proj_10.net28 ));
 sg13g2_or2_1 \proj_10.or20/_0_  (.X(\proj_10.net131 ),
    .B(\proj_10.net165 ),
    .A(\proj_10.net139 ));
 sg13g2_or2_1 \proj_10.or21/_0_  (.X(\proj_10.net132 ),
    .B(\proj_10.net166 ),
    .A(\proj_10.net140 ));
 sg13g2_or2_1 \proj_10.or22/_0_  (.X(\proj_10.net133 ),
    .B(\proj_10.net167 ),
    .A(\proj_10.net141 ));
 sg13g2_or2_1 \proj_10.or23/_0_  (.X(\proj_10.net134 ),
    .B(\proj_10.net168 ),
    .A(\proj_10.net142 ));
 sg13g2_or2_1 \proj_10.or24/_0_  (.X(\proj_10.net135 ),
    .B(\proj_10.net169 ),
    .A(\proj_10.net143 ));
 sg13g2_or2_1 \proj_10.or25/_0_  (.X(\proj_10.net86 ),
    .B(\proj_10.net171 ),
    .A(\proj_10.net170 ));
 sg13g2_or2_1 \proj_10.or26/_0_  (.X(\proj_10.net88 ),
    .B(\proj_10.net174 ),
    .A(\proj_10.net173 ));
 sg13g2_or2_1 \proj_10.or27/_0_  (.X(\proj_10.net90 ),
    .B(\proj_10.net176 ),
    .A(\proj_10.net175 ));
 sg13g2_or2_1 \proj_10.or28/_0_  (.X(\proj_10.net92 ),
    .B(\proj_10.net178 ),
    .A(\proj_10.net177 ));
 sg13g2_or2_1 \proj_10.or29/_0_  (.X(\proj_10.net94 ),
    .B(\proj_10.net180 ),
    .A(\proj_10.net179 ));
 sg13g2_or2_1 \proj_10.or3/_0_  (.X(\proj_10.net36 ),
    .B(\proj_10.net33 ),
    .A(\proj_10.net35 ));
 sg13g2_or2_1 \proj_10.or30/_0_  (.X(\proj_10.net96 ),
    .B(\proj_10.net182 ),
    .A(\proj_10.net181 ));
 sg13g2_or2_1 \proj_10.or31/_0_  (.X(\proj_10.net98 ),
    .B(\proj_10.net184 ),
    .A(\proj_10.net183 ));
 sg13g2_or2_1 \proj_10.or32/_0_  (.X(\proj_10.net100 ),
    .B(\proj_10.net186 ),
    .A(\proj_10.net185 ));
 sg13g2_or2_1 \proj_10.or33/_0_  (.X(\proj_10.net78 ),
    .B(\proj_10.net189 ),
    .A(\proj_10.net187 ));
 sg13g2_or2_1 \proj_10.or34/_0_  (.X(\proj_10.net79 ),
    .B(\proj_10.net191 ),
    .A(\proj_10.net190 ));
 sg13g2_or2_1 \proj_10.or35/_0_  (.X(\proj_10.net80 ),
    .B(\proj_10.net193 ),
    .A(\proj_10.net192 ));
 sg13g2_or2_1 \proj_10.or36/_0_  (.X(\proj_10.net81 ),
    .B(\proj_10.net195 ),
    .A(\proj_10.net194 ));
 sg13g2_or2_1 \proj_10.or37/_0_  (.X(\proj_10.net82 ),
    .B(\proj_10.net197 ),
    .A(\proj_10.net196 ));
 sg13g2_or2_1 \proj_10.or38/_0_  (.X(\proj_10.net83 ),
    .B(\proj_10.net199 ),
    .A(\proj_10.net198 ));
 sg13g2_or2_1 \proj_10.or39/_0_  (.X(\proj_10.net84 ),
    .B(\proj_10.net201 ),
    .A(\proj_10.net200 ));
 sg13g2_or2_1 \proj_10.or4/_0_  (.X(\proj_10.net43 ),
    .B(\proj_10.net40 ),
    .A(\proj_10.net42 ));
 sg13g2_or2_1 \proj_10.or40/_0_  (.X(\proj_10.net85 ),
    .B(\proj_10.net203 ),
    .A(\proj_10.net202 ));
 sg13g2_or2_1 \proj_10.or41/_0_  (.X(\proj_10.net162 ),
    .B(\proj_10.net154 ),
    .A(\proj_10.net204 ));
 sg13g2_or2_1 \proj_10.or42/_0_  (.X(\proj_10.net163 ),
    .B(\proj_10.net155 ),
    .A(\proj_10.net205 ));
 sg13g2_or2_1 \proj_10.or43/_0_  (.X(\proj_10.net164 ),
    .B(\proj_10.net156 ),
    .A(\proj_10.net206 ));
 sg13g2_or2_1 \proj_10.or44/_0_  (.X(\proj_10.net165 ),
    .B(\proj_10.net157 ),
    .A(\proj_10.net207 ));
 sg13g2_or2_1 \proj_10.or45/_0_  (.X(\proj_10.net166 ),
    .B(\proj_10.net158 ),
    .A(\proj_10.net208 ));
 sg13g2_or2_1 \proj_10.or46/_0_  (.X(\proj_10.net167 ),
    .B(\proj_10.net159 ),
    .A(\proj_10.net209 ));
 sg13g2_or2_1 \proj_10.or47/_0_  (.X(\proj_10.net168 ),
    .B(\proj_10.net160 ),
    .A(\proj_10.net210 ));
 sg13g2_or2_1 \proj_10.or48/_0_  (.X(\proj_10.net169 ),
    .B(\proj_10.net161 ),
    .A(\proj_10.net211 ));
 sg13g2_or2_1 \proj_10.or49/_0_  (.X(\proj_10.net204 ),
    .B(\proj_10.net212 ),
    .A(net29));
 sg13g2_or2_1 \proj_10.or5/_0_  (.X(\proj_10.net50 ),
    .B(\proj_10.net47 ),
    .A(\proj_10.net49 ));
 sg13g2_or2_1 \proj_10.or50/_0_  (.X(\proj_10.net205 ),
    .B(\proj_10.net214 ),
    .A(net30));
 sg13g2_or2_1 \proj_10.or51/_0_  (.X(\proj_10.net206 ),
    .B(\proj_10.net215 ),
    .A(net31));
 sg13g2_or2_1 \proj_10.or52/_0_  (.X(\proj_10.net207 ),
    .B(\proj_10.net216 ),
    .A(net32));
 sg13g2_or2_1 \proj_10.or53/_0_  (.X(\proj_10.net208 ),
    .B(\proj_10.net217 ),
    .A(net33));
 sg13g2_or2_1 \proj_10.or54/_0_  (.X(\proj_10.net209 ),
    .B(\proj_10.net218 ),
    .A(net34));
 sg13g2_or2_1 \proj_10.or55/_0_  (.X(\proj_10.net210 ),
    .B(\proj_10.net219 ),
    .A(net35));
 sg13g2_or2_1 \proj_10.or56/_0_  (.X(\proj_10.net211 ),
    .B(\proj_10.net220 ),
    .A(net36));
 sg13g2_or2_1 \proj_10.or6/_0_  (.X(\proj_10.net57 ),
    .B(\proj_10.net54 ),
    .A(\proj_10.net56 ));
 sg13g2_or2_1 \proj_10.or7/_0_  (.X(\proj_10.net64 ),
    .B(\proj_10.net61 ),
    .A(\proj_10.net63 ));
 sg13g2_or2_1 \proj_10.or8/_0_  (.X(\proj_10.net71 ),
    .B(\proj_10.net68 ),
    .A(\proj_10.net70 ));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(net107),
    .A(\proj_10.net87 ),
    .X(\proj_10.net24 ));
 sg13g2_xor2_1 \proj_10.xor10/_0_  (.B(\proj_10.net43 ),
    .A(\proj_10.net46 ),
    .X(\proj_10.net48 ));
 sg13g2_xor2_1 \proj_10.xor11/_0_  (.B(\proj_10.net51 ),
    .A(\proj_10.net52 ),
    .X(\proj_10.net53 ));
 sg13g2_xor2_1 \proj_10.xor12/_0_  (.B(\proj_10.net50 ),
    .A(\proj_10.net53 ),
    .X(\proj_10.net55 ));
 sg13g2_xor2_1 \proj_10.xor13/_0_  (.B(\proj_10.net58 ),
    .A(\proj_10.net59 ),
    .X(\proj_10.net60 ));
 sg13g2_xor2_1 \proj_10.xor14/_0_  (.B(\proj_10.net57 ),
    .A(\proj_10.net60 ),
    .X(\proj_10.net62 ));
 sg13g2_xor2_1 \proj_10.xor15/_0_  (.B(\proj_10.net65 ),
    .A(\proj_10.net66 ),
    .X(\proj_10.net67 ));
 sg13g2_xor2_1 \proj_10.xor16/_0_  (.B(\proj_10.net64 ),
    .A(\proj_10.net67 ),
    .X(\proj_10.net69 ));
 sg13g2_xor2_1 \proj_10.xor17/_0_  (.B(\proj_10.net72 ),
    .A(\proj_10.net73 ),
    .X(\proj_10.net74 ));
 sg13g2_xor2_1 \proj_10.xor18/_0_  (.B(\proj_10.net71 ),
    .A(\proj_10.net74 ),
    .X(\proj_10.net76 ));
 sg13g2_xor2_1 \proj_10.xor19/_0_  (.B(net107),
    .A(\proj_10.net91 ),
    .X(\proj_10.net38 ));
 sg13g2_xor2_1 \proj_10.xor2/_0_  (.B(net107),
    .A(\proj_10.net89 ),
    .X(\proj_10.net31 ));
 sg13g2_xor2_1 \proj_10.xor20/_0_  (.B(net107),
    .A(\proj_10.net93 ),
    .X(\proj_10.net45 ));
 sg13g2_xor2_1 \proj_10.xor21/_0_  (.B(net109),
    .A(\proj_10.net95 ),
    .X(\proj_10.net52 ));
 sg13g2_xor2_1 \proj_10.xor22/_0_  (.B(net109),
    .A(\proj_10.net97 ),
    .X(\proj_10.net59 ));
 sg13g2_xor2_1 \proj_10.xor23/_0_  (.B(net109),
    .A(\proj_10.net99 ),
    .X(\proj_10.net66 ));
 sg13g2_xor2_1 \proj_10.xor24/_0_  (.B(net109),
    .A(\proj_10.net101 ),
    .X(\proj_10.net73 ));
 sg13g2_xor2_1 \proj_10.xor3/_0_  (.B(\proj_10.net23 ),
    .A(\proj_10.net24 ),
    .X(\proj_10.net25 ));
 sg13g2_xor2_1 \proj_10.xor4/_0_  (.B(net107),
    .A(\proj_10.net25 ),
    .X(\proj_10.net27 ));
 sg13g2_xor2_1 \proj_10.xor5/_0_  (.B(\proj_10.net30 ),
    .A(\proj_10.net31 ),
    .X(\proj_10.net32 ));
 sg13g2_xor2_1 \proj_10.xor6/_0_  (.B(\proj_10.net29 ),
    .A(\proj_10.net32 ),
    .X(\proj_10.net34 ));
 sg13g2_xor2_1 \proj_10.xor7/_0_  (.B(\proj_10.net37 ),
    .A(\proj_10.net38 ),
    .X(\proj_10.net39 ));
 sg13g2_xor2_1 \proj_10.xor8/_0_  (.B(\proj_10.net36 ),
    .A(\proj_10.net39 ),
    .X(\proj_10.net41 ));
 sg13g2_xor2_1 \proj_10.xor9/_0_  (.B(\proj_10.net44 ),
    .A(\proj_10.net45 ),
    .X(\proj_10.net46 ));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(\proj_11.net5 ),
    .B(net135),
    .X(\proj_11.net4 ));
 sg13g2_inv_1 \proj_11.not5/_0_  (.Y(\proj_11.net3 ),
    .A(net134));
 sg13g2_inv_1 \proj_11.not6/_0_  (.Y(\proj_11.net5 ),
    .A(net131));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net117),
    .B(net121),
    .X(\proj_12.net22 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(net132),
    .B(net135),
    .X(\proj_12.net23 ));
 sg13g2_and2_1 \proj_12.and3/_0_  (.A(net125),
    .B(net129),
    .X(\proj_12.net24 ));
 sg13g2_and2_1 \proj_12.and4/_0_  (.A(net110),
    .B(net113),
    .X(\proj_12.net25 ));
 sg13g2_and2_1 \proj_12.and5/_0_  (.A(\proj_12.net24 ),
    .B(\proj_12.net23 ),
    .X(\proj_12.net26 ));
 sg13g2_and2_1 \proj_12.and6/_0_  (.A(\proj_12.net25 ),
    .B(\proj_12.net22 ),
    .X(\proj_12.net27 ));
 sg13g2_and2_1 \proj_12.and7/_0_  (.A(\proj_12.net27 ),
    .B(\proj_12.net26 ),
    .X(\proj_12.net10 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net128),
    .A(net125),
    .X(\proj_12.net16 ));
 sg13g2_xor2_1 \proj_12.xor2/_0_  (.B(net121),
    .A(net117),
    .X(\proj_12.net17 ));
 sg13g2_xor2_1 \proj_12.xor3/_0_  (.B(net113),
    .A(net110),
    .X(\proj_12.net18 ));
 sg13g2_xor2_1 \proj_12.xor4/_0_  (.B(net136),
    .A(net133),
    .X(\proj_12.net19 ));
 sg13g2_xor2_1 \proj_12.xor5/_0_  (.B(\proj_12.net19 ),
    .A(\proj_12.net16 ),
    .X(\proj_12.net20 ));
 sg13g2_xor2_1 \proj_12.xor6/_0_  (.B(\proj_12.net17 ),
    .A(\proj_12.net18 ),
    .X(\proj_12.net21 ));
 sg13g2_xor2_1 \proj_12.xor7/_0_  (.B(\proj_12.net20 ),
    .A(\proj_12.net21 ),
    .X(\proj_12.net9 ));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(net133),
    .B(\proj_13.net11 ),
    .X(\proj_13.net12 ));
 sg13g2_and2_1 \proj_13.and3/_0_  (.A(net129),
    .B(\proj_13.net12 ),
    .X(\proj_13.net13 ));
 sg13g2_and2_1 \proj_13.and4/_0_  (.A(\proj_13.net14 ),
    .B(\proj_13.net13 ),
    .X(\proj_13.net15 ));
 sg13g2_and2_1 \proj_13.and5/_0_  (.A(net122),
    .B(\proj_13.net15 ),
    .X(\proj_13.net16 ));
 sg13g2_and2_1 \proj_13.and6/_0_  (.A(net117),
    .B(\proj_13.net16 ),
    .X(\proj_13.net17 ));
 sg13g2_and2_1 \proj_13.and7/_0_  (.A(net113),
    .B(\proj_13.net17 ),
    .X(\proj_13.net18 ));
 sg13g2_and2_1 \proj_13.and8/_0_  (.A(\proj_13.net18 ),
    .B(\proj_13.net20 ),
    .X(\proj_13.net9 ));
 sg13g2_inv_1 \proj_13.not1/_0_  (.Y(\proj_13.net11 ),
    .A(net136));
 sg13g2_inv_1 \proj_13.not2/_0_  (.Y(\proj_13.net20 ),
    .A(net110));
 sg13g2_inv_1 \proj_13.not3/_0_  (.Y(\proj_13.net14 ),
    .A(net126));
 sg13g2_and2_1 \proj__0.and1/_0_  (.A(net132),
    .B(net135),
    .X(\proj__0.net15 ));
 sg13g2_and2_1 \proj__0.and10/_0_  (.A(\proj__0.net26 ),
    .B(\proj__0.net25 ),
    .X(\proj__0.net28 ));
 sg13g2_and2_1 \proj__0.and11/_0_  (.A(\proj__0.net27 ),
    .B(\proj__0.net26 ),
    .X(\proj__0.net29 ));
 sg13g2_and2_1 \proj__0.and12/_0_  (.A(\proj__0.net29 ),
    .B(\proj__0.net28 ),
    .X(\proj__0.net30 ));
 sg13g2_and2_1 \proj__0.and13/_0_  (.A(\proj__0.net30 ),
    .B(\proj__0.net20 ),
    .X(\proj__0.net9 ));
 sg13g2_and2_1 \proj__0.and2/_0_  (.A(net128),
    .B(net132),
    .X(\proj__0.net16 ));
 sg13g2_and2_1 \proj__0.and3/_0_  (.A(net125),
    .B(net128),
    .X(\proj__0.net17 ));
 sg13g2_and2_1 \proj__0.and4/_0_  (.A(\proj__0.net16 ),
    .B(\proj__0.net15 ),
    .X(\proj__0.net18 ));
 sg13g2_and2_1 \proj__0.and5/_0_  (.A(\proj__0.net17 ),
    .B(\proj__0.net16 ),
    .X(\proj__0.net19 ));
 sg13g2_and2_1 \proj__0.and6/_0_  (.A(\proj__0.net19 ),
    .B(\proj__0.net18 ),
    .X(\proj__0.net20 ));
 sg13g2_and2_1 \proj__0.and7/_0_  (.A(\proj__0.net22 ),
    .B(\proj__0.net21 ),
    .X(\proj__0.net25 ));
 sg13g2_and2_1 \proj__0.and8/_0_  (.A(\proj__0.net23 ),
    .B(\proj__0.net22 ),
    .X(\proj__0.net26 ));
 sg13g2_and2_1 \proj__0.and9/_0_  (.A(\proj__0.net24 ),
    .B(\proj__0.net23 ),
    .X(\proj__0.net27 ));
 sg13g2_inv_1 \proj__0.not1/_0_  (.Y(\proj__0.net21 ),
    .A(net121));
 sg13g2_inv_1 \proj__0.not2/_0_  (.Y(\proj__0.net22 ),
    .A(net118));
 sg13g2_inv_1 \proj__0.not3/_0_  (.Y(\proj__0.net23 ),
    .A(net114));
 sg13g2_inv_1 \proj__0.not4/_0_  (.Y(\proj__0.net24 ),
    .A(net110));
 sg13g2_and2_1 \proj__1.and1/_0_  (.A(net130),
    .B(net134),
    .X(\proj__1.net9 ));
 sg13g2_inv_1 \proj__1.not1/_0_  (.Y(\proj__1.net11 ),
    .A(net108));
 sg13g2_xor2_1 \proj__1.xor1/_0_  (.B(net119),
    .A(net115),
    .X(\proj__1.net10 ));
 sg13g2_and2_1 \proj__2.and1/_0_  (.A(net120),
    .B(net134),
    .X(\proj__2.net19 ));
 sg13g2_and2_1 \proj__2.and2/_0_  (.A(net116),
    .B(net130),
    .X(\proj__2.net21 ));
 sg13g2_and2_1 \proj__2.and3/_0_  (.A(\proj__2.net19 ),
    .B(\proj__2.net20 ),
    .X(\proj__2.net22 ));
 sg13g2_and2_1 \proj__2.and4/_0_  (.A(net112),
    .B(net127),
    .X(\proj__2.net24 ));
 sg13g2_and2_1 \proj__2.and5/_0_  (.A(\proj__2.net23 ),
    .B(\proj__2.net25 ),
    .X(\proj__2.net26 ));
 sg13g2_and2_1 \proj__2.and6/_0_  (.A(\proj__2.net28 ),
    .B(\proj__2.net27 ),
    .X(\proj__2.net29 ));
 sg13g2_and2_1 \proj__2.and7/_0_  (.A(net108),
    .B(net124),
    .X(\proj__2.net30 ));
 sg13g2_or2_1 \proj__2.or1/_0_  (.X(\proj__2.net23 ),
    .B(\proj__2.net21 ),
    .A(\proj__2.net22 ));
 sg13g2_or2_1 \proj__2.or2/_0_  (.X(\proj__2.net27 ),
    .B(\proj__2.net26 ),
    .A(\proj__2.net24 ));
 sg13g2_or2_1 \proj__2.or3/_0_  (.X(\proj__2.net13 ),
    .B(\proj__2.net30 ),
    .A(\proj__2.net29 ));
 sg13g2_xor2_1 \proj__2.xor1/_0_  (.B(net134),
    .A(net120),
    .X(\proj__2.net9 ));
 sg13g2_xor2_1 \proj__2.xor2/_0_  (.B(\proj__2.net20 ),
    .A(\proj__2.net19 ),
    .X(\proj__2.net10 ));
 sg13g2_xor2_1 \proj__2.xor3/_0_  (.B(net130),
    .A(net116),
    .X(\proj__2.net20 ));
 sg13g2_xor2_1 \proj__2.xor4/_0_  (.B(net127),
    .A(net112),
    .X(\proj__2.net25 ));
 sg13g2_xor2_1 \proj__2.xor5/_0_  (.B(\proj__2.net27 ),
    .A(\proj__2.net28 ),
    .X(\proj__2.net12 ));
 sg13g2_xor2_1 \proj__2.xor6/_0_  (.B(net124),
    .A(net108),
    .X(\proj__2.net28 ));
 sg13g2_xor2_1 \proj__2.xor7/_0_  (.B(\proj__2.net25 ),
    .A(\proj__2.net23 ),
    .X(\proj__2.net11 ));
 sg13g2_and2_1 \proj__3.and1/_0_  (.A(\proj__3.net22 ),
    .B(\proj__3.net21 ),
    .X(\proj__3.net12 ));
 sg13g2_and2_1 \proj__3.and2/_0_  (.A(\proj__3.net22 ),
    .B(\proj__3.net21 ),
    .X(\proj__3.net25 ));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net26 ),
    .B(\proj__3.net25 ),
    .X(\proj__3.net13 ));
 sg13g2_nand2_1 \proj__3.nand1/_0_  (.Y(\proj__3.net11 ),
    .A(\proj__3.net22 ),
    .B(\proj__3.net24 ));
 sg13g2_nand2_1 \proj__3.nand2/_0_  (.Y(\proj__3.net26 ),
    .A(\proj__3.net15 ),
    .B(\proj__3.net24 ));
 sg13g2_nand2_1 \proj__3.nand3/_0_  (.Y(\proj__3.net14 ),
    .A(\proj__3.net26 ),
    .B(\proj__3.net25 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net23 ),
    .A(net37));
 sg13g2_or2_1 \proj__3.or1/_0_  (.X(\proj__3.net15 ),
    .B(net112),
    .A(net107));
 sg13g2_or2_1 \proj__3.or3/_0_  (.X(\proj__3.net21 ),
    .B(net129),
    .A(net126));
 sg13g2_or2_1 \proj__3.or4/_0_  (.X(\proj__3.net22 ),
    .B(net134),
    .A(net130));
 sg13g2_xor2_1 \proj__3.xor1/_0_  (.B(\proj__3.net23 ),
    .A(net38),
    .X(\proj__3.net24 ));
 sg13g2_nand2_1 \proj__4.nand1/_0_  (.Y(\proj__4.net9 ),
    .A(net124),
    .B(\proj__4.net10 ));
 sg13g2_inv_1 \proj__4.not3/_0_  (.Y(\proj__4.net10 ),
    .A(net127));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net107),
    .B(net112),
    .X(\proj__5.net8 ));
 sg13g2_inv_1 \proj__5.not1/_0_  (.Y(\proj__5.net7 ),
    .A(net123));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net6 ),
    .B(net130),
    .A(net124));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(\proj__6.net17 ),
    .B(\proj__6.net16 ),
    .X(\proj__6.net18 ));
 sg13g2_and2_1 \proj__6.and3/_0_  (.A(\proj__6.net20 ),
    .B(\proj__6.net21 ),
    .X(\proj__6.net22 ));
 sg13g2_and2_1 \proj__6.and4/_0_  (.A(net131),
    .B(net136),
    .X(\proj__6.net17 ));
 sg13g2_and2_1 \proj__6.and5/_0_  (.A(net124),
    .B(net127),
    .X(\proj__6.net19 ));
 sg13g2_and2_1 \proj__6.and6/_0_  (.A(net116),
    .B(net120),
    .X(\proj__6.net23 ));
 sg13g2_or2_1 \proj__6.or2/_0_  (.X(\proj__6.net20 ),
    .B(\proj__6.net18 ),
    .A(\proj__6.net19 ));
 sg13g2_or2_1 \proj__6.or3/_0_  (.X(\proj__6.net10 ),
    .B(\proj__6.net22 ),
    .A(\proj__6.net23 ));
 sg13g2_xor2_1 \proj__6.xor2/_0_  (.B(net134),
    .A(net130),
    .X(\proj__6.net7 ));
 sg13g2_xor2_1 \proj__6.xor3/_0_  (.B(\proj__6.net17 ),
    .A(\proj__6.net16 ),
    .X(\proj__6.net8 ));
 sg13g2_xor2_1 \proj__6.xor4/_0_  (.B(net127),
    .A(net124),
    .X(\proj__6.net16 ));
 sg13g2_xor2_1 \proj__6.xor5/_0_  (.B(\proj__6.net20 ),
    .A(\proj__6.net21 ),
    .X(\proj__6.net9 ));
 sg13g2_xor2_1 \proj__6.xor6/_0_  (.B(net120),
    .A(net119),
    .X(\proj__6.net21 ));
 sg13g2_inv_1 \proj__7.not1/_0_  (.Y(\proj__7.net9 ),
    .A(net134));
 sg13g2_inv_1 \proj__7.not2/_0_  (.Y(\proj__7.net10 ),
    .A(net132));
 sg13g2_inv_1 \proj__7.not3/_0_  (.Y(\proj__7.net11 ),
    .A(net127));
 sg13g2_inv_1 \proj__7.not4/_0_  (.Y(\proj__7.net12 ),
    .A(net124));
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(net130),
    .B(net135),
    .X(\proj__8.net7 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(net132),
    .B(\proj__9.net22 ),
    .X(\proj__9.net23 ));
 sg13g2_and2_1 \proj__9.and10/_0_  (.A(\proj__9.net26 ),
    .B(\proj__9.net52 ),
    .X(\proj__9.net32 ));
 sg13g2_and2_1 \proj__9.and11/_0_  (.A(\proj__9.net56 ),
    .B(\proj__9.net51 ),
    .X(\proj__9.net37 ));
 sg13g2_and2_1 \proj__9.and12/_0_  (.A(\proj__9.net23 ),
    .B(\proj__9.net27 ),
    .X(\proj__9.net36 ));
 sg13g2_and2_1 \proj__9.and13/_0_  (.A(\proj__9.net57 ),
    .B(\proj__9.net54 ),
    .X(\proj__9.net40 ));
 sg13g2_and2_1 \proj__9.and14/_0_  (.A(\proj__9.net58 ),
    .B(\proj__9.net52 ),
    .X(\proj__9.net39 ));
 sg13g2_and2_1 \proj__9.and15/_0_  (.A(\proj__9.net59 ),
    .B(\proj__9.net51 ),
    .X(\proj__9.net44 ));
 sg13g2_and2_1 \proj__9.and16/_0_  (.A(\proj__9.net23 ),
    .B(\proj__9.net28 ),
    .X(\proj__9.net43 ));
 sg13g2_and2_1 \proj__9.and17/_0_  (.A(\proj__9.net60 ),
    .B(\proj__9.net54 ),
    .X(\proj__9.net47 ));
 sg13g2_and2_1 \proj__9.and18/_0_  (.A(\proj__9.net61 ),
    .B(\proj__9.net52 ),
    .X(\proj__9.net46 ));
 sg13g2_and2_1 \proj__9.and19/_0_  (.A(net39),
    .B(\proj__9.net62 ),
    .X(\proj__9.net64 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(\proj__9.net50 ),
    .B(net135),
    .X(\proj__9.net51 ));
 sg13g2_and2_1 \proj__9.and20/_0_  (.A(net109),
    .B(net121),
    .X(\proj__9.net65 ));
 sg13g2_and2_1 \proj__9.and21/_0_  (.A(\proj__9.net66 ),
    .B(\proj__9.net67 ),
    .X(\proj__9.net68 ));
 sg13g2_and2_1 \proj__9.and22/_0_  (.A(net113),
    .B(net125),
    .X(\proj__9.net69 ));
 sg13g2_and2_1 \proj__9.and23/_0_  (.A(\proj__9.net70 ),
    .B(\proj__9.net71 ),
    .X(\proj__9.net72 ));
 sg13g2_and2_1 \proj__9.and24/_0_  (.A(net117),
    .B(net128),
    .X(\proj__9.net73 ));
 sg13g2_and2_1 \proj__9.and25/_0_  (.A(\proj__9.net74 ),
    .B(\proj__9.net54 ),
    .X(\proj__9.net16 ));
 sg13g2_and2_1 \proj__9.and26/_0_  (.A(\proj__9.net75 ),
    .B(\proj__9.net35 ),
    .X(\proj__9.net76 ));
 sg13g2_and2_1 \proj__9.and27/_0_  (.A(\proj__9.net79 ),
    .B(\proj__9.net42 ),
    .X(\proj__9.net80 ));
 sg13g2_and2_1 \proj__9.and28/_0_  (.A(\proj__9.net78 ),
    .B(\proj__9.net77 ),
    .X(\proj__9.net79 ));
 sg13g2_and2_1 \proj__9.and29/_0_  (.A(\proj__9.net81 ),
    .B(net104),
    .X(\proj__9.net82 ));
 sg13g2_and2_1 \proj__9.and3/_0_  (.A(net132),
    .B(net135),
    .X(\proj__9.net52 ));
 sg13g2_and2_1 \proj__9.and30/_0_  (.A(\proj__9.net84 ),
    .B(\proj__9.net83 ),
    .X(\proj__9.net81 ));
 sg13g2_and2_1 \proj__9.and31/_0_  (.A(\proj__9.net90 ),
    .B(\proj__9.net89 ),
    .X(\proj__9.net91 ));
 sg13g2_and2_1 \proj__9.and32/_0_  (.A(net102),
    .B(\proj__9.net91 ),
    .X(\proj__9.net87 ));
 sg13g2_and2_1 \proj__9.and33/_0_  (.A(net103),
    .B(net102),
    .X(\proj__9.net92 ));
 sg13g2_and2_1 \proj__9.and34/_0_  (.A(net104),
    .B(\proj__9.net92 ),
    .X(\proj__9.net88 ));
 sg13g2_and2_1 \proj__9.and35/_0_  (.A(\proj__9.net94 ),
    .B(\proj__9.net93 ),
    .X(\proj__9.net95 ));
 sg13g2_and2_1 \proj__9.and36/_0_  (.A(net103),
    .B(\proj__9.net100 ),
    .X(\proj__9.net97 ));
 sg13g2_and2_1 \proj__9.and37/_0_  (.A(net103),
    .B(net102),
    .X(\proj__9.net102 ));
 sg13g2_and2_1 \proj__9.and38/_0_  (.A(\proj__9.net103 ),
    .B(\proj__9.net102 ),
    .X(\proj__9.net99 ));
 sg13g2_and2_1 \proj__9.and39/_0_  (.A(net104),
    .B(net102),
    .X(\proj__9.net107 ));
 sg13g2_and2_1 \proj__9.and4/_0_  (.A(net117),
    .B(net128),
    .X(\proj__9.net53 ));
 sg13g2_and2_1 \proj__9.and40/_0_  (.A(\proj__9.net108 ),
    .B(\proj__9.net107 ),
    .X(\proj__9.net105 ));
 sg13g2_and2_1 \proj__9.and41/_0_  (.A(net104),
    .B(\proj__9.net112 ),
    .X(\proj__9.net109 ));
 sg13g2_and2_1 \proj__9.and5/_0_  (.A(net113),
    .B(net125),
    .X(\proj__9.net56 ));
 sg13g2_and2_1 \proj__9.and6/_0_  (.A(net109),
    .B(net121),
    .X(\proj__9.net59 ));
 sg13g2_and2_1 \proj__9.and7/_0_  (.A(\proj__9.net53 ),
    .B(\proj__9.net51 ),
    .X(\proj__9.net30 ));
 sg13g2_and2_1 \proj__9.and8/_0_  (.A(\proj__9.net25 ),
    .B(\proj__9.net23 ),
    .X(\proj__9.net29 ));
 sg13g2_and2_1 \proj__9.and9/_0_  (.A(\proj__9.net55 ),
    .B(\proj__9.net54 ),
    .X(\proj__9.net33 ));
 sg13g2_or2_1 \proj__9.nand1/_0_  (.X(\proj__9.net24 ),
    .B(net132),
    .A(net135));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net22 ),
    .A(net135));
 sg13g2_inv_1 \proj__9.not10/_0_  (.Y(\proj__9.net10 ),
    .A(\proj__9.net76 ));
 sg13g2_inv_1 \proj__9.not11/_0_  (.Y(\proj__9.net11 ),
    .A(\proj__9.net80 ));
 sg13g2_inv_1 \proj__9.not12/_0_  (.Y(\proj__9.net12 ),
    .A(\proj__9.net86 ));
 sg13g2_inv_1 \proj__9.not13/_0_  (.Y(\proj__9.net94 ),
    .A(net104));
 sg13g2_inv_1 \proj__9.not14/_0_  (.Y(\proj__9.net93 ),
    .A(\proj__9.net96 ));
 sg13g2_inv_1 \proj__9.not15/_0_  (.Y(\proj__9.net100 ),
    .A(\proj__9.net101 ));
 sg13g2_inv_1 \proj__9.not16/_0_  (.Y(\proj__9.net103 ),
    .A(net104));
 sg13g2_inv_1 \proj__9.not17/_0_  (.Y(\proj__9.net108 ),
    .A(net103));
 sg13g2_inv_1 \proj__9.not18/_0_  (.Y(\proj__9.net9 ),
    .A(\proj__9.net110 ));
 sg13g2_inv_1 \proj__9.not19/_0_  (.Y(\proj__9.net112 ),
    .A(\proj__9.net111 ));
 sg13g2_inv_1 \proj__9.not2/_0_  (.Y(\proj__9.net50 ),
    .A(net132));
 sg13g2_inv_1 \proj__9.not20/_0_  (.Y(\proj__9.net15 ),
    .A(\proj__9.net114 ));
 sg13g2_inv_1 \proj__9.not3/_0_  (.Y(\proj__9.net54 ),
    .A(\proj__9.net24 ));
 sg13g2_inv_1 \proj__9.not4/_0_  (.Y(\proj__9.net77 ),
    .A(\proj__9.net35 ));
 sg13g2_inv_1 \proj__9.not5/_0_  (.Y(\proj__9.net78 ),
    .A(\proj__9.net49 ));
 sg13g2_inv_1 \proj__9.not6/_0_  (.Y(\proj__9.net89 ),
    .A(net103));
 sg13g2_inv_1 \proj__9.not7/_0_  (.Y(\proj__9.net90 ),
    .A(net104));
 sg13g2_inv_1 \proj__9.not8/_0_  (.Y(\proj__9.net83 ),
    .A(net102));
 sg13g2_inv_1 \proj__9.not9/_0_  (.Y(\proj__9.net84 ),
    .A(net103));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net25 ),
    .B(net128),
    .A(net117));
 sg13g2_or2_1 \proj__9.or10/_0_  (.X(\proj__9.net45 ),
    .B(\proj__9.net43 ),
    .A(\proj__9.net44 ));
 sg13g2_or2_1 \proj__9.or11/_0_  (.X(\proj__9.net48 ),
    .B(\proj__9.net46 ),
    .A(\proj__9.net47 ));
 sg13g2_or2_2 \proj__9.or12/_0_  (.X(\proj__9.net49 ),
    .B(\proj__9.net45 ),
    .A(\proj__9.net48 ));
 sg13g2_or2_1 \proj__9.or13/_0_  (.X(\proj__9.net66 ),
    .B(\proj__9.net64 ),
    .A(\proj__9.net65 ));
 sg13g2_or2_1 \proj__9.or14/_0_  (.X(\proj__9.net70 ),
    .B(\proj__9.net68 ),
    .A(\proj__9.net69 ));
 sg13g2_or2_1 \proj__9.or15/_0_  (.X(\proj__9.net74 ),
    .B(\proj__9.net72 ),
    .A(\proj__9.net73 ));
 sg13g2_or2_1 \proj__9.or16/_0_  (.X(\proj__9.net86 ),
    .B(\proj__9.net82 ),
    .A(\proj__9.net85 ));
 sg13g2_or2_1 \proj__9.or17/_0_  (.X(\proj__9.net85 ),
    .B(\proj__9.net87 ),
    .A(\proj__9.net88 ));
 sg13g2_or2_1 \proj__9.or18/_0_  (.X(\proj__9.net96 ),
    .B(net102),
    .A(net103));
 sg13g2_or2_1 \proj__9.or19/_0_  (.X(\proj__9.net98 ),
    .B(\proj__9.net95 ),
    .A(\proj__9.net97 ));
 sg13g2_or2_1 \proj__9.or2/_0_  (.X(\proj__9.net27 ),
    .B(net125),
    .A(net113));
 sg13g2_or2_1 \proj__9.or20/_0_  (.X(\proj__9.net13 ),
    .B(\proj__9.net98 ),
    .A(\proj__9.net99 ));
 sg13g2_or2_1 \proj__9.or21/_0_  (.X(\proj__9.net101 ),
    .B(net104),
    .A(net102));
 sg13g2_or2_1 \proj__9.or22/_0_  (.X(\proj__9.net104 ),
    .B(\proj__9.net95 ),
    .A(\proj__9.net87 ));
 sg13g2_or2_1 \proj__9.or23/_0_  (.X(\proj__9.net106 ),
    .B(\proj__9.net99 ),
    .A(\proj__9.net105 ));
 sg13g2_or2_1 \proj__9.or24/_0_  (.X(\proj__9.net14 ),
    .B(\proj__9.net104 ),
    .A(\proj__9.net106 ));
 sg13g2_or2_1 \proj__9.or25/_0_  (.X(\proj__9.net110 ),
    .B(\proj__9.net109 ),
    .A(\proj__9.net87 ));
 sg13g2_or2_1 \proj__9.or26/_0_  (.X(\proj__9.net111 ),
    .B(net102),
    .A(net103));
 sg13g2_or2_1 \proj__9.or27/_0_  (.X(\proj__9.net113 ),
    .B(\proj__9.net109 ),
    .A(\proj__9.net95 ));
 sg13g2_or2_1 \proj__9.or28/_0_  (.X(\proj__9.net114 ),
    .B(\proj__9.net113 ),
    .A(\proj__9.net88 ));
 sg13g2_or2_1 \proj__9.or3/_0_  (.X(\proj__9.net28 ),
    .B(net121),
    .A(net110));
 sg13g2_or2_1 \proj__9.or4/_0_  (.X(\proj__9.net31 ),
    .B(\proj__9.net29 ),
    .A(\proj__9.net30 ));
 sg13g2_or2_1 \proj__9.or5/_0_  (.X(\proj__9.net34 ),
    .B(\proj__9.net32 ),
    .A(\proj__9.net33 ));
 sg13g2_or2_2 \proj__9.or6/_0_  (.X(\proj__9.net35 ),
    .B(\proj__9.net31 ),
    .A(\proj__9.net34 ));
 sg13g2_or2_1 \proj__9.or7/_0_  (.X(\proj__9.net38 ),
    .B(\proj__9.net36 ),
    .A(\proj__9.net37 ));
 sg13g2_or2_1 \proj__9.or8/_0_  (.X(\proj__9.net41 ),
    .B(\proj__9.net39 ),
    .A(\proj__9.net40 ));
 sg13g2_or2_2 \proj__9.or9/_0_  (.X(\proj__9.net42 ),
    .B(\proj__9.net38 ),
    .A(\proj__9.net41 ));
 sg13g2_xor2_1 \proj__9.xor1/_0_  (.B(net128),
    .A(net117),
    .X(\proj__9.net26 ));
 sg13g2_xor2_1 \proj__9.xor10/_0_  (.B(\proj__9.net42 ),
    .A(\proj__9.net49 ),
    .X(\proj__9.net75 ));
 sg13g2_xor2_1 \proj__9.xor2/_0_  (.B(net125),
    .A(net113),
    .X(\proj__9.net58 ));
 sg13g2_xor2_1 \proj__9.xor3/_0_  (.B(net121),
    .A(net109),
    .X(\proj__9.net61 ));
 sg13g2_xor2_1 \proj__9.xor4/_0_  (.B(\proj__9.net62 ),
    .A(net40),
    .X(\proj__9.net60 ));
 sg13g2_xor2_1 \proj__9.xor5/_0_  (.B(net121),
    .A(net109),
    .X(\proj__9.net62 ));
 sg13g2_xor2_1 \proj__9.xor6/_0_  (.B(\proj__9.net67 ),
    .A(\proj__9.net66 ),
    .X(\proj__9.net57 ));
 sg13g2_xor2_1 \proj__9.xor7/_0_  (.B(net125),
    .A(net113),
    .X(\proj__9.net67 ));
 sg13g2_xor2_1 \proj__9.xor8/_0_  (.B(net128),
    .A(net117),
    .X(\proj__9.net71 ));
 sg13g2_xor2_1 \proj__9.xor9/_0_  (.B(\proj__9.net71 ),
    .A(\proj__9.net70 ),
    .X(\proj__9.net55 ));
 sg13g2_buf_2 fanout102 (.A(\proj__9.net35 ),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(\proj__9.net42 ),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(\proj__9.net49 ),
    .X(net104));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(\proj_10.net110 ));
 sg13g2_buf_2 fanout106 (.A(\proj_10.net144 ),
    .X(net106));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net111));
 sg13g2_buf_1 fanout108 (.A(net111),
    .X(net108));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(net111));
 sg13g2_buf_2 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(ui_in[7]),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net115),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(net115),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(ui_in[6]),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(net119),
    .X(net116));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(net118));
 sg13g2_buf_2 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(ui_in[5]),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(net123));
 sg13g2_buf_2 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(ui_in[4]),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(net126),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(ui_in[3]),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net129),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(net129),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(ui_in[2]),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(ui_in[1]));
 sg13g2_buf_2 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(ui_in[1]),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net136),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(ui_in[0]),
    .X(net136));
 sg13g2_buf_2 input1 (.A(uio_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(uio_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(uio_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(uio_in[3]),
    .X(net4));
 sg13g2_tielo \proj_10.flop1/_1__5  (.L_LO(net5));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_fill_2 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_fill_2 FILLER_19_316 ();
 sg13g2_fill_1 FILLER_19_318 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_350 ();
 sg13g2_fill_2 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_185 ();
 sg13g2_decap_8 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_fill_2 FILLER_20_204 ();
 sg13g2_fill_2 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_decap_4 FILLER_20_282 ();
 sg13g2_decap_4 FILLER_20_299 ();
 sg13g2_decap_4 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_decap_4 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_4 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_fill_2 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_4 FILLER_21_327 ();
 sg13g2_fill_1 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_fill_2 FILLER_21_360 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_fill_2 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_4 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_decap_4 FILLER_22_151 ();
 sg13g2_fill_2 FILLER_22_155 ();
 sg13g2_decap_8 FILLER_22_162 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_204 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_250 ();
 sg13g2_fill_2 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_decap_4 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_118 ();
 sg13g2_decap_8 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_decap_4 FILLER_23_164 ();
 sg13g2_fill_2 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_4 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_241 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_fill_2 FILLER_23_318 ();
 sg13g2_fill_1 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_4 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_4 FILLER_23_376 ();
 sg13g2_fill_2 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_129 ();
 sg13g2_decap_4 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_decap_4 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_fill_2 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_328 ();
 sg13g2_decap_4 FILLER_24_335 ();
 sg13g2_fill_1 FILLER_24_339 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_2 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_118 ();
 sg13g2_fill_1 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_decap_4 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_210 ();
 sg13g2_decap_4 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_4 FILLER_25_291 ();
 sg13g2_fill_2 FILLER_25_300 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_decap_4 FILLER_25_308 ();
 sg13g2_fill_2 FILLER_25_316 ();
 sg13g2_decap_4 FILLER_25_322 ();
 sg13g2_fill_2 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_fill_2 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_decap_4 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_4 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_decap_4 FILLER_26_202 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_237 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_fill_2 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_decap_4 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_334 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_380 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_4 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_decap_8 FILLER_27_118 ();
 sg13g2_decap_4 FILLER_27_143 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_167 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_decap_4 FILLER_27_213 ();
 sg13g2_decap_4 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_decap_4 FILLER_27_255 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_275 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_293 ();
 sg13g2_decap_4 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_304 ();
 sg13g2_decap_4 FILLER_27_315 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_2 FILLER_27_325 ();
 sg13g2_decap_4 FILLER_27_331 ();
 sg13g2_fill_2 FILLER_27_335 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_decap_4 FILLER_27_349 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_4 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_384 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_decap_8 FILLER_28_164 ();
 sg13g2_fill_2 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_fill_2 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_246 ();
 sg13g2_decap_4 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_decap_4 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_297 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_107 ();
 sg13g2_decap_8 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_decap_4 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_decap_8 FILLER_29_208 ();
 sg13g2_decap_4 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_decap_4 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_2 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_4 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_311 ();
 sg13g2_decap_4 FILLER_29_322 ();
 sg13g2_decap_4 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_decap_4 FILLER_29_337 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_346 ();
 sg13g2_decap_8 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_365 ();
 sg13g2_fill_2 FILLER_29_381 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_117 ();
 sg13g2_decap_8 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_fill_2 FILLER_30_135 ();
 sg13g2_decap_4 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_174 ();
 sg13g2_decap_4 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_decap_4 FILLER_30_190 ();
 sg13g2_fill_2 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_fill_2 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_decap_8 FILLER_30_239 ();
 sg13g2_fill_2 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_248 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_decap_4 FILLER_30_272 ();
 sg13g2_fill_2 FILLER_30_276 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_336 ();
 sg13g2_fill_1 FILLER_30_353 ();
 sg13g2_decap_4 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_4 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_172 ();
 sg13g2_decap_4 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_decap_4 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_fill_2 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_decap_4 FILLER_31_331 ();
 sg13g2_fill_2 FILLER_31_338 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_fill_1 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_decap_4 FILLER_32_170 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_4 FILLER_32_186 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_2 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_238 ();
 sg13g2_fill_2 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_271 ();
 sg13g2_decap_4 FILLER_32_302 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_decap_4 FILLER_32_339 ();
 sg13g2_fill_2 FILLER_32_343 ();
 sg13g2_decap_4 FILLER_32_348 ();
 sg13g2_fill_2 FILLER_32_352 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_4 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_144 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_194 ();
 sg13g2_decap_8 FILLER_33_219 ();
 sg13g2_decap_4 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_230 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_decap_4 FILLER_33_258 ();
 sg13g2_decap_4 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_decap_4 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_313 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_decap_4 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_decap_4 FILLER_33_365 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_165 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_decap_4 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_294 ();
 sg13g2_decap_4 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_fill_1 FILLER_34_352 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_2 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_239 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_decap_4 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_fill_2 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_35_383 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_159 ();
 sg13g2_decap_8 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_176 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_decap_4 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_211 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_decap_8 FILLER_36_225 ();
 sg13g2_decap_8 FILLER_36_232 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_293 ();
 sg13g2_decap_4 FILLER_36_300 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_decap_4 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_fill_2 FILLER_36_365 ();
 sg13g2_decap_4 FILLER_36_372 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_fill_1 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_261 ();
 sg13g2_decap_8 FILLER_37_268 ();
 sg13g2_decap_8 FILLER_37_275 ();
 sg13g2_decap_8 FILLER_37_282 ();
 sg13g2_decap_8 FILLER_37_289 ();
 sg13g2_decap_8 FILLER_37_296 ();
 sg13g2_fill_2 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_4 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_decap_8 FILLER_38_321 ();
 sg13g2_decap_8 FILLER_38_328 ();
 sg13g2_decap_8 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_342 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_decap_8 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net41;
 assign uio_oe[1] = net42;
 assign uio_oe[2] = net43;
 assign uio_oe[3] = net44;
 assign uio_oe[4] = net45;
 assign uio_oe[5] = net46;
 assign uio_oe[6] = net47;
 assign uio_oe[7] = net48;
 assign uio_out[0] = net49;
 assign uio_out[1] = net50;
 assign uio_out[2] = net51;
 assign uio_out[3] = net52;
 assign uio_out[4] = net53;
 assign uio_out[5] = net54;
 assign uio_out[6] = net55;
 assign uio_out[7] = net56;
endmodule

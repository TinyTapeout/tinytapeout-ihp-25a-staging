module tt_um_branch_pred (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire clk_regs;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire \abs_sum[0] ;
 wire \cnt[0] ;
 wire \cnt[1] ;
 wire \cnt[2] ;
 wire \cnt[3] ;
 wire \history_buffer[0] ;
 wire \history_buffer[1] ;
 wire \history_buffer[2] ;
 wire \history_buffer[3] ;
 wire \history_buffer[4] ;
 wire \history_buffer[5] ;
 wire \history_buffer[6] ;
 wire \history_buffer[7] ;
 wire history_buffer_empty_state;
 wire \history_buffer_index[0] ;
 wire \history_buffer_index[1] ;
 wire \history_buffer_index[2] ;
 wire history_buffer_output;
 wire history_buffer_request_prev;
 wire \latch_mem.RAM[0][0] ;
 wire \latch_mem.RAM[0][1] ;
 wire \latch_mem.RAM[0][2] ;
 wire \latch_mem.RAM[0][3] ;
 wire \latch_mem.RAM[0][4] ;
 wire \latch_mem.RAM[0][5] ;
 wire \latch_mem.RAM[0][6] ;
 wire \latch_mem.RAM[0][7] ;
 wire \latch_mem.RAM[10][0] ;
 wire \latch_mem.RAM[10][1] ;
 wire \latch_mem.RAM[10][2] ;
 wire \latch_mem.RAM[10][3] ;
 wire \latch_mem.RAM[10][4] ;
 wire \latch_mem.RAM[10][5] ;
 wire \latch_mem.RAM[10][6] ;
 wire \latch_mem.RAM[10][7] ;
 wire \latch_mem.RAM[11][0] ;
 wire \latch_mem.RAM[11][1] ;
 wire \latch_mem.RAM[11][2] ;
 wire \latch_mem.RAM[11][3] ;
 wire \latch_mem.RAM[11][4] ;
 wire \latch_mem.RAM[11][5] ;
 wire \latch_mem.RAM[11][6] ;
 wire \latch_mem.RAM[11][7] ;
 wire \latch_mem.RAM[12][0] ;
 wire \latch_mem.RAM[12][1] ;
 wire \latch_mem.RAM[12][2] ;
 wire \latch_mem.RAM[12][3] ;
 wire \latch_mem.RAM[12][4] ;
 wire \latch_mem.RAM[12][5] ;
 wire \latch_mem.RAM[12][6] ;
 wire \latch_mem.RAM[12][7] ;
 wire \latch_mem.RAM[13][0] ;
 wire \latch_mem.RAM[13][1] ;
 wire \latch_mem.RAM[13][2] ;
 wire \latch_mem.RAM[13][3] ;
 wire \latch_mem.RAM[13][4] ;
 wire \latch_mem.RAM[13][5] ;
 wire \latch_mem.RAM[13][6] ;
 wire \latch_mem.RAM[13][7] ;
 wire \latch_mem.RAM[14][0] ;
 wire \latch_mem.RAM[14][1] ;
 wire \latch_mem.RAM[14][2] ;
 wire \latch_mem.RAM[14][3] ;
 wire \latch_mem.RAM[14][4] ;
 wire \latch_mem.RAM[14][5] ;
 wire \latch_mem.RAM[14][6] ;
 wire \latch_mem.RAM[14][7] ;
 wire \latch_mem.RAM[15][0] ;
 wire \latch_mem.RAM[15][1] ;
 wire \latch_mem.RAM[15][2] ;
 wire \latch_mem.RAM[15][3] ;
 wire \latch_mem.RAM[15][4] ;
 wire \latch_mem.RAM[15][5] ;
 wire \latch_mem.RAM[15][6] ;
 wire \latch_mem.RAM[15][7] ;
 wire \latch_mem.RAM[16][0] ;
 wire \latch_mem.RAM[16][1] ;
 wire \latch_mem.RAM[16][2] ;
 wire \latch_mem.RAM[16][3] ;
 wire \latch_mem.RAM[16][4] ;
 wire \latch_mem.RAM[16][5] ;
 wire \latch_mem.RAM[16][6] ;
 wire \latch_mem.RAM[16][7] ;
 wire \latch_mem.RAM[17][0] ;
 wire \latch_mem.RAM[17][1] ;
 wire \latch_mem.RAM[17][2] ;
 wire \latch_mem.RAM[17][3] ;
 wire \latch_mem.RAM[17][4] ;
 wire \latch_mem.RAM[17][5] ;
 wire \latch_mem.RAM[17][6] ;
 wire \latch_mem.RAM[17][7] ;
 wire \latch_mem.RAM[18][0] ;
 wire \latch_mem.RAM[18][1] ;
 wire \latch_mem.RAM[18][2] ;
 wire \latch_mem.RAM[18][3] ;
 wire \latch_mem.RAM[18][4] ;
 wire \latch_mem.RAM[18][5] ;
 wire \latch_mem.RAM[18][6] ;
 wire \latch_mem.RAM[18][7] ;
 wire \latch_mem.RAM[19][0] ;
 wire \latch_mem.RAM[19][1] ;
 wire \latch_mem.RAM[19][2] ;
 wire \latch_mem.RAM[19][3] ;
 wire \latch_mem.RAM[19][4] ;
 wire \latch_mem.RAM[19][5] ;
 wire \latch_mem.RAM[19][6] ;
 wire \latch_mem.RAM[19][7] ;
 wire \latch_mem.RAM[1][0] ;
 wire \latch_mem.RAM[1][1] ;
 wire \latch_mem.RAM[1][2] ;
 wire \latch_mem.RAM[1][3] ;
 wire \latch_mem.RAM[1][4] ;
 wire \latch_mem.RAM[1][5] ;
 wire \latch_mem.RAM[1][6] ;
 wire \latch_mem.RAM[1][7] ;
 wire \latch_mem.RAM[20][0] ;
 wire \latch_mem.RAM[20][1] ;
 wire \latch_mem.RAM[20][2] ;
 wire \latch_mem.RAM[20][3] ;
 wire \latch_mem.RAM[20][4] ;
 wire \latch_mem.RAM[20][5] ;
 wire \latch_mem.RAM[20][6] ;
 wire \latch_mem.RAM[20][7] ;
 wire \latch_mem.RAM[21][0] ;
 wire \latch_mem.RAM[21][1] ;
 wire \latch_mem.RAM[21][2] ;
 wire \latch_mem.RAM[21][3] ;
 wire \latch_mem.RAM[21][4] ;
 wire \latch_mem.RAM[21][5] ;
 wire \latch_mem.RAM[21][6] ;
 wire \latch_mem.RAM[21][7] ;
 wire \latch_mem.RAM[22][0] ;
 wire \latch_mem.RAM[22][1] ;
 wire \latch_mem.RAM[22][2] ;
 wire \latch_mem.RAM[22][3] ;
 wire \latch_mem.RAM[22][4] ;
 wire \latch_mem.RAM[22][5] ;
 wire \latch_mem.RAM[22][6] ;
 wire \latch_mem.RAM[22][7] ;
 wire \latch_mem.RAM[23][0] ;
 wire \latch_mem.RAM[23][1] ;
 wire \latch_mem.RAM[23][2] ;
 wire \latch_mem.RAM[23][3] ;
 wire \latch_mem.RAM[23][4] ;
 wire \latch_mem.RAM[23][5] ;
 wire \latch_mem.RAM[23][6] ;
 wire \latch_mem.RAM[23][7] ;
 wire \latch_mem.RAM[24][0] ;
 wire \latch_mem.RAM[24][1] ;
 wire \latch_mem.RAM[24][2] ;
 wire \latch_mem.RAM[24][3] ;
 wire \latch_mem.RAM[24][4] ;
 wire \latch_mem.RAM[24][5] ;
 wire \latch_mem.RAM[24][6] ;
 wire \latch_mem.RAM[24][7] ;
 wire \latch_mem.RAM[25][0] ;
 wire \latch_mem.RAM[25][1] ;
 wire \latch_mem.RAM[25][2] ;
 wire \latch_mem.RAM[25][3] ;
 wire \latch_mem.RAM[25][4] ;
 wire \latch_mem.RAM[25][5] ;
 wire \latch_mem.RAM[25][6] ;
 wire \latch_mem.RAM[25][7] ;
 wire \latch_mem.RAM[26][0] ;
 wire \latch_mem.RAM[26][1] ;
 wire \latch_mem.RAM[26][2] ;
 wire \latch_mem.RAM[26][3] ;
 wire \latch_mem.RAM[26][4] ;
 wire \latch_mem.RAM[26][5] ;
 wire \latch_mem.RAM[26][6] ;
 wire \latch_mem.RAM[26][7] ;
 wire \latch_mem.RAM[27][0] ;
 wire \latch_mem.RAM[27][1] ;
 wire \latch_mem.RAM[27][2] ;
 wire \latch_mem.RAM[27][3] ;
 wire \latch_mem.RAM[27][4] ;
 wire \latch_mem.RAM[27][5] ;
 wire \latch_mem.RAM[27][6] ;
 wire \latch_mem.RAM[27][7] ;
 wire \latch_mem.RAM[28][0] ;
 wire \latch_mem.RAM[28][1] ;
 wire \latch_mem.RAM[28][2] ;
 wire \latch_mem.RAM[28][3] ;
 wire \latch_mem.RAM[28][4] ;
 wire \latch_mem.RAM[28][5] ;
 wire \latch_mem.RAM[28][6] ;
 wire \latch_mem.RAM[28][7] ;
 wire \latch_mem.RAM[29][0] ;
 wire \latch_mem.RAM[29][1] ;
 wire \latch_mem.RAM[29][2] ;
 wire \latch_mem.RAM[29][3] ;
 wire \latch_mem.RAM[29][4] ;
 wire \latch_mem.RAM[29][5] ;
 wire \latch_mem.RAM[29][6] ;
 wire \latch_mem.RAM[29][7] ;
 wire \latch_mem.RAM[2][0] ;
 wire \latch_mem.RAM[2][1] ;
 wire \latch_mem.RAM[2][2] ;
 wire \latch_mem.RAM[2][3] ;
 wire \latch_mem.RAM[2][4] ;
 wire \latch_mem.RAM[2][5] ;
 wire \latch_mem.RAM[2][6] ;
 wire \latch_mem.RAM[2][7] ;
 wire \latch_mem.RAM[30][0] ;
 wire \latch_mem.RAM[30][1] ;
 wire \latch_mem.RAM[30][2] ;
 wire \latch_mem.RAM[30][3] ;
 wire \latch_mem.RAM[30][4] ;
 wire \latch_mem.RAM[30][5] ;
 wire \latch_mem.RAM[30][6] ;
 wire \latch_mem.RAM[30][7] ;
 wire \latch_mem.RAM[31][0] ;
 wire \latch_mem.RAM[31][1] ;
 wire \latch_mem.RAM[31][2] ;
 wire \latch_mem.RAM[31][3] ;
 wire \latch_mem.RAM[31][4] ;
 wire \latch_mem.RAM[31][5] ;
 wire \latch_mem.RAM[31][6] ;
 wire \latch_mem.RAM[31][7] ;
 wire \latch_mem.RAM[32][0] ;
 wire \latch_mem.RAM[32][1] ;
 wire \latch_mem.RAM[32][2] ;
 wire \latch_mem.RAM[32][3] ;
 wire \latch_mem.RAM[32][4] ;
 wire \latch_mem.RAM[32][5] ;
 wire \latch_mem.RAM[32][6] ;
 wire \latch_mem.RAM[32][7] ;
 wire \latch_mem.RAM[33][0] ;
 wire \latch_mem.RAM[33][1] ;
 wire \latch_mem.RAM[33][2] ;
 wire \latch_mem.RAM[33][3] ;
 wire \latch_mem.RAM[33][4] ;
 wire \latch_mem.RAM[33][5] ;
 wire \latch_mem.RAM[33][6] ;
 wire \latch_mem.RAM[33][7] ;
 wire \latch_mem.RAM[34][0] ;
 wire \latch_mem.RAM[34][1] ;
 wire \latch_mem.RAM[34][2] ;
 wire \latch_mem.RAM[34][3] ;
 wire \latch_mem.RAM[34][4] ;
 wire \latch_mem.RAM[34][5] ;
 wire \latch_mem.RAM[34][6] ;
 wire \latch_mem.RAM[34][7] ;
 wire \latch_mem.RAM[35][0] ;
 wire \latch_mem.RAM[35][1] ;
 wire \latch_mem.RAM[35][2] ;
 wire \latch_mem.RAM[35][3] ;
 wire \latch_mem.RAM[35][4] ;
 wire \latch_mem.RAM[35][5] ;
 wire \latch_mem.RAM[35][6] ;
 wire \latch_mem.RAM[35][7] ;
 wire \latch_mem.RAM[36][0] ;
 wire \latch_mem.RAM[36][1] ;
 wire \latch_mem.RAM[36][2] ;
 wire \latch_mem.RAM[36][3] ;
 wire \latch_mem.RAM[36][4] ;
 wire \latch_mem.RAM[36][5] ;
 wire \latch_mem.RAM[36][6] ;
 wire \latch_mem.RAM[36][7] ;
 wire \latch_mem.RAM[37][0] ;
 wire \latch_mem.RAM[37][1] ;
 wire \latch_mem.RAM[37][2] ;
 wire \latch_mem.RAM[37][3] ;
 wire \latch_mem.RAM[37][4] ;
 wire \latch_mem.RAM[37][5] ;
 wire \latch_mem.RAM[37][6] ;
 wire \latch_mem.RAM[37][7] ;
 wire \latch_mem.RAM[38][0] ;
 wire \latch_mem.RAM[38][1] ;
 wire \latch_mem.RAM[38][2] ;
 wire \latch_mem.RAM[38][3] ;
 wire \latch_mem.RAM[38][4] ;
 wire \latch_mem.RAM[38][5] ;
 wire \latch_mem.RAM[38][6] ;
 wire \latch_mem.RAM[38][7] ;
 wire \latch_mem.RAM[39][0] ;
 wire \latch_mem.RAM[39][1] ;
 wire \latch_mem.RAM[39][2] ;
 wire \latch_mem.RAM[39][3] ;
 wire \latch_mem.RAM[39][4] ;
 wire \latch_mem.RAM[39][5] ;
 wire \latch_mem.RAM[39][6] ;
 wire \latch_mem.RAM[39][7] ;
 wire \latch_mem.RAM[3][0] ;
 wire \latch_mem.RAM[3][1] ;
 wire \latch_mem.RAM[3][2] ;
 wire \latch_mem.RAM[3][3] ;
 wire \latch_mem.RAM[3][4] ;
 wire \latch_mem.RAM[3][5] ;
 wire \latch_mem.RAM[3][6] ;
 wire \latch_mem.RAM[3][7] ;
 wire \latch_mem.RAM[40][0] ;
 wire \latch_mem.RAM[40][1] ;
 wire \latch_mem.RAM[40][2] ;
 wire \latch_mem.RAM[40][3] ;
 wire \latch_mem.RAM[40][4] ;
 wire \latch_mem.RAM[40][5] ;
 wire \latch_mem.RAM[40][6] ;
 wire \latch_mem.RAM[40][7] ;
 wire \latch_mem.RAM[41][0] ;
 wire \latch_mem.RAM[41][1] ;
 wire \latch_mem.RAM[41][2] ;
 wire \latch_mem.RAM[41][3] ;
 wire \latch_mem.RAM[41][4] ;
 wire \latch_mem.RAM[41][5] ;
 wire \latch_mem.RAM[41][6] ;
 wire \latch_mem.RAM[41][7] ;
 wire \latch_mem.RAM[42][0] ;
 wire \latch_mem.RAM[42][1] ;
 wire \latch_mem.RAM[42][2] ;
 wire \latch_mem.RAM[42][3] ;
 wire \latch_mem.RAM[42][4] ;
 wire \latch_mem.RAM[42][5] ;
 wire \latch_mem.RAM[42][6] ;
 wire \latch_mem.RAM[42][7] ;
 wire \latch_mem.RAM[43][0] ;
 wire \latch_mem.RAM[43][1] ;
 wire \latch_mem.RAM[43][2] ;
 wire \latch_mem.RAM[43][3] ;
 wire \latch_mem.RAM[43][4] ;
 wire \latch_mem.RAM[43][5] ;
 wire \latch_mem.RAM[43][6] ;
 wire \latch_mem.RAM[43][7] ;
 wire \latch_mem.RAM[44][0] ;
 wire \latch_mem.RAM[44][1] ;
 wire \latch_mem.RAM[44][2] ;
 wire \latch_mem.RAM[44][3] ;
 wire \latch_mem.RAM[44][4] ;
 wire \latch_mem.RAM[44][5] ;
 wire \latch_mem.RAM[44][6] ;
 wire \latch_mem.RAM[44][7] ;
 wire \latch_mem.RAM[45][0] ;
 wire \latch_mem.RAM[45][1] ;
 wire \latch_mem.RAM[45][2] ;
 wire \latch_mem.RAM[45][3] ;
 wire \latch_mem.RAM[45][4] ;
 wire \latch_mem.RAM[45][5] ;
 wire \latch_mem.RAM[45][6] ;
 wire \latch_mem.RAM[45][7] ;
 wire \latch_mem.RAM[46][0] ;
 wire \latch_mem.RAM[46][1] ;
 wire \latch_mem.RAM[46][2] ;
 wire \latch_mem.RAM[46][3] ;
 wire \latch_mem.RAM[46][4] ;
 wire \latch_mem.RAM[46][5] ;
 wire \latch_mem.RAM[46][6] ;
 wire \latch_mem.RAM[46][7] ;
 wire \latch_mem.RAM[47][0] ;
 wire \latch_mem.RAM[47][1] ;
 wire \latch_mem.RAM[47][2] ;
 wire \latch_mem.RAM[47][3] ;
 wire \latch_mem.RAM[47][4] ;
 wire \latch_mem.RAM[47][5] ;
 wire \latch_mem.RAM[47][6] ;
 wire \latch_mem.RAM[47][7] ;
 wire \latch_mem.RAM[48][0] ;
 wire \latch_mem.RAM[48][1] ;
 wire \latch_mem.RAM[48][2] ;
 wire \latch_mem.RAM[48][3] ;
 wire \latch_mem.RAM[48][4] ;
 wire \latch_mem.RAM[48][5] ;
 wire \latch_mem.RAM[48][6] ;
 wire \latch_mem.RAM[48][7] ;
 wire \latch_mem.RAM[49][0] ;
 wire \latch_mem.RAM[49][1] ;
 wire \latch_mem.RAM[49][2] ;
 wire \latch_mem.RAM[49][3] ;
 wire \latch_mem.RAM[49][4] ;
 wire \latch_mem.RAM[49][5] ;
 wire \latch_mem.RAM[49][6] ;
 wire \latch_mem.RAM[49][7] ;
 wire \latch_mem.RAM[4][0] ;
 wire \latch_mem.RAM[4][1] ;
 wire \latch_mem.RAM[4][2] ;
 wire \latch_mem.RAM[4][3] ;
 wire \latch_mem.RAM[4][4] ;
 wire \latch_mem.RAM[4][5] ;
 wire \latch_mem.RAM[4][6] ;
 wire \latch_mem.RAM[4][7] ;
 wire \latch_mem.RAM[50][0] ;
 wire \latch_mem.RAM[50][1] ;
 wire \latch_mem.RAM[50][2] ;
 wire \latch_mem.RAM[50][3] ;
 wire \latch_mem.RAM[50][4] ;
 wire \latch_mem.RAM[50][5] ;
 wire \latch_mem.RAM[50][6] ;
 wire \latch_mem.RAM[50][7] ;
 wire \latch_mem.RAM[51][0] ;
 wire \latch_mem.RAM[51][1] ;
 wire \latch_mem.RAM[51][2] ;
 wire \latch_mem.RAM[51][3] ;
 wire \latch_mem.RAM[51][4] ;
 wire \latch_mem.RAM[51][5] ;
 wire \latch_mem.RAM[51][6] ;
 wire \latch_mem.RAM[51][7] ;
 wire \latch_mem.RAM[52][0] ;
 wire \latch_mem.RAM[52][1] ;
 wire \latch_mem.RAM[52][2] ;
 wire \latch_mem.RAM[52][3] ;
 wire \latch_mem.RAM[52][4] ;
 wire \latch_mem.RAM[52][5] ;
 wire \latch_mem.RAM[52][6] ;
 wire \latch_mem.RAM[52][7] ;
 wire \latch_mem.RAM[53][0] ;
 wire \latch_mem.RAM[53][1] ;
 wire \latch_mem.RAM[53][2] ;
 wire \latch_mem.RAM[53][3] ;
 wire \latch_mem.RAM[53][4] ;
 wire \latch_mem.RAM[53][5] ;
 wire \latch_mem.RAM[53][6] ;
 wire \latch_mem.RAM[53][7] ;
 wire \latch_mem.RAM[54][0] ;
 wire \latch_mem.RAM[54][1] ;
 wire \latch_mem.RAM[54][2] ;
 wire \latch_mem.RAM[54][3] ;
 wire \latch_mem.RAM[54][4] ;
 wire \latch_mem.RAM[54][5] ;
 wire \latch_mem.RAM[54][6] ;
 wire \latch_mem.RAM[54][7] ;
 wire \latch_mem.RAM[55][0] ;
 wire \latch_mem.RAM[55][1] ;
 wire \latch_mem.RAM[55][2] ;
 wire \latch_mem.RAM[55][3] ;
 wire \latch_mem.RAM[55][4] ;
 wire \latch_mem.RAM[55][5] ;
 wire \latch_mem.RAM[55][6] ;
 wire \latch_mem.RAM[55][7] ;
 wire \latch_mem.RAM[56][0] ;
 wire \latch_mem.RAM[56][1] ;
 wire \latch_mem.RAM[56][2] ;
 wire \latch_mem.RAM[56][3] ;
 wire \latch_mem.RAM[56][4] ;
 wire \latch_mem.RAM[56][5] ;
 wire \latch_mem.RAM[56][6] ;
 wire \latch_mem.RAM[56][7] ;
 wire \latch_mem.RAM[57][0] ;
 wire \latch_mem.RAM[57][1] ;
 wire \latch_mem.RAM[57][2] ;
 wire \latch_mem.RAM[57][3] ;
 wire \latch_mem.RAM[57][4] ;
 wire \latch_mem.RAM[57][5] ;
 wire \latch_mem.RAM[57][6] ;
 wire \latch_mem.RAM[57][7] ;
 wire \latch_mem.RAM[58][0] ;
 wire \latch_mem.RAM[58][1] ;
 wire \latch_mem.RAM[58][2] ;
 wire \latch_mem.RAM[58][3] ;
 wire \latch_mem.RAM[58][4] ;
 wire \latch_mem.RAM[58][5] ;
 wire \latch_mem.RAM[58][6] ;
 wire \latch_mem.RAM[58][7] ;
 wire \latch_mem.RAM[59][0] ;
 wire \latch_mem.RAM[59][1] ;
 wire \latch_mem.RAM[59][2] ;
 wire \latch_mem.RAM[59][3] ;
 wire \latch_mem.RAM[59][4] ;
 wire \latch_mem.RAM[59][5] ;
 wire \latch_mem.RAM[59][6] ;
 wire \latch_mem.RAM[59][7] ;
 wire \latch_mem.RAM[5][0] ;
 wire \latch_mem.RAM[5][1] ;
 wire \latch_mem.RAM[5][2] ;
 wire \latch_mem.RAM[5][3] ;
 wire \latch_mem.RAM[5][4] ;
 wire \latch_mem.RAM[5][5] ;
 wire \latch_mem.RAM[5][6] ;
 wire \latch_mem.RAM[5][7] ;
 wire \latch_mem.RAM[60][0] ;
 wire \latch_mem.RAM[60][1] ;
 wire \latch_mem.RAM[60][2] ;
 wire \latch_mem.RAM[60][3] ;
 wire \latch_mem.RAM[60][4] ;
 wire \latch_mem.RAM[60][5] ;
 wire \latch_mem.RAM[60][6] ;
 wire \latch_mem.RAM[60][7] ;
 wire \latch_mem.RAM[61][0] ;
 wire \latch_mem.RAM[61][1] ;
 wire \latch_mem.RAM[61][2] ;
 wire \latch_mem.RAM[61][3] ;
 wire \latch_mem.RAM[61][4] ;
 wire \latch_mem.RAM[61][5] ;
 wire \latch_mem.RAM[61][6] ;
 wire \latch_mem.RAM[61][7] ;
 wire \latch_mem.RAM[62][0] ;
 wire \latch_mem.RAM[62][1] ;
 wire \latch_mem.RAM[62][2] ;
 wire \latch_mem.RAM[62][3] ;
 wire \latch_mem.RAM[62][4] ;
 wire \latch_mem.RAM[62][5] ;
 wire \latch_mem.RAM[62][6] ;
 wire \latch_mem.RAM[62][7] ;
 wire \latch_mem.RAM[63][0] ;
 wire \latch_mem.RAM[63][1] ;
 wire \latch_mem.RAM[63][2] ;
 wire \latch_mem.RAM[63][3] ;
 wire \latch_mem.RAM[63][4] ;
 wire \latch_mem.RAM[63][5] ;
 wire \latch_mem.RAM[63][6] ;
 wire \latch_mem.RAM[63][7] ;
 wire \latch_mem.RAM[6][0] ;
 wire \latch_mem.RAM[6][1] ;
 wire \latch_mem.RAM[6][2] ;
 wire \latch_mem.RAM[6][3] ;
 wire \latch_mem.RAM[6][4] ;
 wire \latch_mem.RAM[6][5] ;
 wire \latch_mem.RAM[6][6] ;
 wire \latch_mem.RAM[6][7] ;
 wire \latch_mem.RAM[7][0] ;
 wire \latch_mem.RAM[7][1] ;
 wire \latch_mem.RAM[7][2] ;
 wire \latch_mem.RAM[7][3] ;
 wire \latch_mem.RAM[7][4] ;
 wire \latch_mem.RAM[7][5] ;
 wire \latch_mem.RAM[7][6] ;
 wire \latch_mem.RAM[7][7] ;
 wire \latch_mem.RAM[8][0] ;
 wire \latch_mem.RAM[8][1] ;
 wire \latch_mem.RAM[8][2] ;
 wire \latch_mem.RAM[8][3] ;
 wire \latch_mem.RAM[8][4] ;
 wire \latch_mem.RAM[8][5] ;
 wire \latch_mem.RAM[8][6] ;
 wire \latch_mem.RAM[8][7] ;
 wire \latch_mem.RAM[9][0] ;
 wire \latch_mem.RAM[9][1] ;
 wire \latch_mem.RAM[9][2] ;
 wire \latch_mem.RAM[9][3] ;
 wire \latch_mem.RAM[9][4] ;
 wire \latch_mem.RAM[9][5] ;
 wire \latch_mem.RAM[9][6] ;
 wire \latch_mem.RAM[9][7] ;
 wire \latch_mem.addr_in[0] ;
 wire \latch_mem.addr_in[1] ;
 wire \latch_mem.addr_in[2] ;
 wire \latch_mem.addr_in[3] ;
 wire \latch_mem.addr_in[4] ;
 wire \latch_mem.addr_in[5] ;
 wire \latch_mem.addr_read[0] ;
 wire \latch_mem.addr_read[1] ;
 wire \latch_mem.addr_read[2] ;
 wire \latch_mem.addr_read[3] ;
 wire \latch_mem.addr_write[0] ;
 wire \latch_mem.addr_write[1] ;
 wire \latch_mem.addr_write[2] ;
 wire \latch_mem.addr_write[3] ;
 wire \latch_mem.addr_write[4] ;
 wire \latch_mem.addr_write[5] ;
 wire \latch_mem.combined_out[0] ;
 wire \latch_mem.combined_out[1] ;
 wire \latch_mem.combined_out[2] ;
 wire \latch_mem.combined_out[3] ;
 wire \latch_mem.combined_out[4] ;
 wire \latch_mem.combined_out[5] ;
 wire \latch_mem.combined_out[6] ;
 wire \latch_mem.combined_out[7] ;
 wire \latch_mem.data_to_write[0] ;
 wire \latch_mem.data_to_write[1] ;
 wire \latch_mem.data_to_write[2] ;
 wire \latch_mem.data_to_write[3] ;
 wire \latch_mem.data_to_write[4] ;
 wire \latch_mem.data_to_write[5] ;
 wire \latch_mem.data_to_write[6] ;
 wire \latch_mem.data_to_write[7] ;
 wire \latch_mem.genblk1[0].sel_byte ;
 wire \latch_mem.genblk1[0].wr_en_this_byte ;
 wire \latch_mem.genblk1[10].sel_byte ;
 wire \latch_mem.genblk1[10].wr_en_this_byte ;
 wire \latch_mem.genblk1[11].sel_byte ;
 wire \latch_mem.genblk1[11].wr_en_this_byte ;
 wire \latch_mem.genblk1[12].sel_byte ;
 wire \latch_mem.genblk1[12].wr_en_this_byte ;
 wire \latch_mem.genblk1[13].sel_byte ;
 wire \latch_mem.genblk1[13].wr_en_this_byte ;
 wire \latch_mem.genblk1[14].sel_byte ;
 wire \latch_mem.genblk1[14].wr_en_this_byte ;
 wire \latch_mem.genblk1[15].sel_byte ;
 wire \latch_mem.genblk1[15].wr_en_this_byte ;
 wire \latch_mem.genblk1[16].sel_byte ;
 wire \latch_mem.genblk1[16].wr_en_this_byte ;
 wire \latch_mem.genblk1[17].sel_byte ;
 wire \latch_mem.genblk1[17].wr_en_this_byte ;
 wire \latch_mem.genblk1[18].sel_byte ;
 wire \latch_mem.genblk1[18].wr_en_this_byte ;
 wire \latch_mem.genblk1[19].sel_byte ;
 wire \latch_mem.genblk1[19].wr_en_this_byte ;
 wire \latch_mem.genblk1[1].sel_byte ;
 wire \latch_mem.genblk1[1].wr_en_this_byte ;
 wire \latch_mem.genblk1[20].sel_byte ;
 wire \latch_mem.genblk1[20].wr_en_this_byte ;
 wire \latch_mem.genblk1[21].sel_byte ;
 wire \latch_mem.genblk1[21].wr_en_this_byte ;
 wire \latch_mem.genblk1[22].sel_byte ;
 wire \latch_mem.genblk1[22].wr_en_this_byte ;
 wire \latch_mem.genblk1[23].sel_byte ;
 wire \latch_mem.genblk1[23].wr_en_this_byte ;
 wire \latch_mem.genblk1[24].sel_byte ;
 wire \latch_mem.genblk1[24].wr_en_this_byte ;
 wire \latch_mem.genblk1[25].sel_byte ;
 wire \latch_mem.genblk1[25].wr_en_this_byte ;
 wire \latch_mem.genblk1[26].sel_byte ;
 wire \latch_mem.genblk1[26].wr_en_this_byte ;
 wire \latch_mem.genblk1[27].sel_byte ;
 wire \latch_mem.genblk1[27].wr_en_this_byte ;
 wire \latch_mem.genblk1[28].sel_byte ;
 wire \latch_mem.genblk1[28].wr_en_this_byte ;
 wire \latch_mem.genblk1[29].sel_byte ;
 wire \latch_mem.genblk1[29].wr_en_this_byte ;
 wire \latch_mem.genblk1[2].sel_byte ;
 wire \latch_mem.genblk1[2].wr_en_this_byte ;
 wire \latch_mem.genblk1[30].sel_byte ;
 wire \latch_mem.genblk1[30].wr_en_this_byte ;
 wire \latch_mem.genblk1[31].sel_byte ;
 wire \latch_mem.genblk1[31].wr_en_this_byte ;
 wire \latch_mem.genblk1[32].sel_byte ;
 wire \latch_mem.genblk1[32].wr_en_this_byte ;
 wire \latch_mem.genblk1[33].sel_byte ;
 wire \latch_mem.genblk1[33].wr_en_this_byte ;
 wire \latch_mem.genblk1[34].sel_byte ;
 wire \latch_mem.genblk1[34].wr_en_this_byte ;
 wire \latch_mem.genblk1[35].sel_byte ;
 wire \latch_mem.genblk1[35].wr_en_this_byte ;
 wire \latch_mem.genblk1[36].sel_byte ;
 wire \latch_mem.genblk1[36].wr_en_this_byte ;
 wire \latch_mem.genblk1[37].sel_byte ;
 wire \latch_mem.genblk1[37].wr_en_this_byte ;
 wire \latch_mem.genblk1[38].sel_byte ;
 wire \latch_mem.genblk1[38].wr_en_this_byte ;
 wire \latch_mem.genblk1[39].sel_byte ;
 wire \latch_mem.genblk1[39].wr_en_this_byte ;
 wire \latch_mem.genblk1[3].sel_byte ;
 wire \latch_mem.genblk1[3].wr_en_this_byte ;
 wire \latch_mem.genblk1[40].sel_byte ;
 wire \latch_mem.genblk1[40].wr_en_this_byte ;
 wire \latch_mem.genblk1[41].sel_byte ;
 wire \latch_mem.genblk1[41].wr_en_this_byte ;
 wire \latch_mem.genblk1[42].sel_byte ;
 wire \latch_mem.genblk1[42].wr_en_this_byte ;
 wire \latch_mem.genblk1[43].sel_byte ;
 wire \latch_mem.genblk1[43].wr_en_this_byte ;
 wire \latch_mem.genblk1[44].sel_byte ;
 wire \latch_mem.genblk1[44].wr_en_this_byte ;
 wire \latch_mem.genblk1[45].sel_byte ;
 wire \latch_mem.genblk1[45].wr_en_this_byte ;
 wire \latch_mem.genblk1[46].sel_byte ;
 wire \latch_mem.genblk1[46].wr_en_this_byte ;
 wire \latch_mem.genblk1[47].sel_byte ;
 wire \latch_mem.genblk1[47].wr_en_this_byte ;
 wire \latch_mem.genblk1[48].sel_byte ;
 wire \latch_mem.genblk1[48].wr_en_this_byte ;
 wire \latch_mem.genblk1[49].sel_byte ;
 wire \latch_mem.genblk1[49].wr_en_this_byte ;
 wire \latch_mem.genblk1[4].sel_byte ;
 wire \latch_mem.genblk1[4].wr_en_this_byte ;
 wire \latch_mem.genblk1[50].sel_byte ;
 wire \latch_mem.genblk1[50].wr_en_this_byte ;
 wire \latch_mem.genblk1[51].sel_byte ;
 wire \latch_mem.genblk1[51].wr_en_this_byte ;
 wire \latch_mem.genblk1[52].sel_byte ;
 wire \latch_mem.genblk1[52].wr_en_this_byte ;
 wire \latch_mem.genblk1[53].sel_byte ;
 wire \latch_mem.genblk1[53].wr_en_this_byte ;
 wire \latch_mem.genblk1[54].sel_byte ;
 wire \latch_mem.genblk1[54].wr_en_this_byte ;
 wire \latch_mem.genblk1[55].sel_byte ;
 wire \latch_mem.genblk1[55].wr_en_this_byte ;
 wire \latch_mem.genblk1[56].sel_byte ;
 wire \latch_mem.genblk1[56].wr_en_this_byte ;
 wire \latch_mem.genblk1[57].sel_byte ;
 wire \latch_mem.genblk1[57].wr_en_this_byte ;
 wire \latch_mem.genblk1[58].sel_byte ;
 wire \latch_mem.genblk1[58].wr_en_this_byte ;
 wire \latch_mem.genblk1[59].sel_byte ;
 wire \latch_mem.genblk1[59].wr_en_this_byte ;
 wire \latch_mem.genblk1[5].sel_byte ;
 wire \latch_mem.genblk1[5].wr_en_this_byte ;
 wire \latch_mem.genblk1[60].sel_byte ;
 wire \latch_mem.genblk1[60].wr_en_this_byte ;
 wire \latch_mem.genblk1[61].sel_byte ;
 wire \latch_mem.genblk1[61].wr_en_this_byte ;
 wire \latch_mem.genblk1[62].sel_byte ;
 wire \latch_mem.genblk1[62].wr_en_this_byte ;
 wire \latch_mem.genblk1[63].sel_byte ;
 wire \latch_mem.genblk1[63].wr_en_this_byte ;
 wire \latch_mem.genblk1[6].sel_byte ;
 wire \latch_mem.genblk1[6].wr_en_this_byte ;
 wire \latch_mem.genblk1[7].sel_byte ;
 wire \latch_mem.genblk1[7].wr_en_this_byte ;
 wire \latch_mem.genblk1[8].sel_byte ;
 wire \latch_mem.genblk1[8].wr_en_this_byte ;
 wire \latch_mem.genblk1[9].sel_byte ;
 wire \latch_mem.genblk1[9].wr_en_this_byte ;
 wire \latch_mem.genblk2[0].partition_sel_n ;
 wire \latch_mem.genblk2[0].selected_out[0] ;
 wire \latch_mem.genblk2[0].selected_out[1] ;
 wire \latch_mem.genblk2[0].selected_out[2] ;
 wire \latch_mem.genblk2[0].selected_out[3] ;
 wire \latch_mem.genblk2[0].selected_out[4] ;
 wire \latch_mem.genblk2[0].selected_out[5] ;
 wire \latch_mem.genblk2[0].selected_out[6] ;
 wire \latch_mem.genblk2[0].selected_out[7] ;
 wire \latch_mem.genblk2[1].partition_sel_n ;
 wire \latch_mem.genblk2[1].selected_out[0] ;
 wire \latch_mem.genblk2[1].selected_out[1] ;
 wire \latch_mem.genblk2[1].selected_out[2] ;
 wire \latch_mem.genblk2[1].selected_out[3] ;
 wire \latch_mem.genblk2[1].selected_out[4] ;
 wire \latch_mem.genblk2[1].selected_out[5] ;
 wire \latch_mem.genblk2[1].selected_out[6] ;
 wire \latch_mem.genblk2[1].selected_out[7] ;
 wire \latch_mem.genblk2[2].partition_sel_n ;
 wire \latch_mem.genblk2[2].selected_out[0] ;
 wire \latch_mem.genblk2[2].selected_out[1] ;
 wire \latch_mem.genblk2[2].selected_out[2] ;
 wire \latch_mem.genblk2[2].selected_out[3] ;
 wire \latch_mem.genblk2[2].selected_out[4] ;
 wire \latch_mem.genblk2[2].selected_out[5] ;
 wire \latch_mem.genblk2[2].selected_out[6] ;
 wire \latch_mem.genblk2[2].selected_out[7] ;
 wire \latch_mem.genblk2[3].partition_sel_n ;
 wire \latch_mem.genblk2[3].selected_out[0] ;
 wire \latch_mem.genblk2[3].selected_out[1] ;
 wire \latch_mem.genblk2[3].selected_out[2] ;
 wire \latch_mem.genblk2[3].selected_out[3] ;
 wire \latch_mem.genblk2[3].selected_out[4] ;
 wire \latch_mem.genblk2[3].selected_out[5] ;
 wire \latch_mem.genblk2[3].selected_out[6] ;
 wire \latch_mem.genblk2[3].selected_out[7] ;
 wire \latch_mem.uio_in[0] ;
 wire \latch_mem.uio_in[1] ;
 wire \latch_mem.uio_in[2] ;
 wire \latch_mem.uio_in[3] ;
 wire \latch_mem.uio_in[4] ;
 wire \latch_mem.uio_in[5] ;
 wire \latch_mem.uio_in[6] ;
 wire \latch_mem.uio_in[7] ;
 wire \latch_mem.uo_out[0] ;
 wire \latch_mem.uo_out[1] ;
 wire \latch_mem.uo_out[2] ;
 wire \latch_mem.uo_out[3] ;
 wire \latch_mem.uo_out[4] ;
 wire \latch_mem.uo_out[5] ;
 wire \latch_mem.uo_out[6] ;
 wire \latch_mem.uo_out[7] ;
 wire \latch_mem.wr_en ;
 wire \latch_mem.wr_en_in ;
 wire \latch_mem.wr_en_next ;
 wire \latch_mem.wr_en_ok ;
 wire \latch_mem.wr_en_valid ;
 wire mem_reset_done;
 wire new_data_avail_posedge;
 wire new_data_avail_prev;
 wire pred_ready;
 wire prediction;
 wire state_rst_memory;
 wire \substate[0] ;
 wire \substate[1] ;
 wire \substate[2] ;
 wire \substate[3] ;
 wire \sum[1] ;
 wire \sum[2] ;
 wire \sum[3] ;
 wire \sum[4] ;
 wire \sum[5] ;
 wire \sum[6] ;
 wire \sum[7] ;
 wire \sum[8] ;
 wire \sum[9] ;
 wire training_done;
 wire net8;
 wire net9;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire delaynet_0_clk;
 wire delaynet_1_clk;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;

 sg13g2_nand2_1 _0917_ (.Y(_0702_),
    .A(\latch_mem.addr_write[4] ),
    .B(\latch_mem.addr_write[5] ));
 sg13g2_nor2_1 _0918_ (.A(_0701_),
    .B(net794),
    .Y(\latch_mem.genblk1[63].sel_byte ));
 sg13g2_nor2_1 _0919_ (.A(\latch_mem.addr_write[0] ),
    .B(_0661_),
    .Y(_0703_));
 sg13g2_nand3_1 _0920_ (.B(net803),
    .C(_0703_),
    .A(net805),
    .Y(_0704_));
 sg13g2_nor2_1 _0921_ (.A(_0702_),
    .B(_0704_),
    .Y(\latch_mem.genblk1[62].sel_byte ));
 sg13g2_nor2_1 _0922_ (.A(_0660_),
    .B(\latch_mem.addr_write[1] ),
    .Y(_0705_));
 sg13g2_nand3_1 _0923_ (.B(net803),
    .C(_0705_),
    .A(net805),
    .Y(_0706_));
 sg13g2_nor2_1 _0924_ (.A(net795),
    .B(_0706_),
    .Y(\latch_mem.genblk1[61].sel_byte ));
 sg13g2_nor2_1 _0925_ (.A(\latch_mem.addr_write[0] ),
    .B(\latch_mem.addr_write[1] ),
    .Y(_0707_));
 sg13g2_nand3_1 _0926_ (.B(net803),
    .C(_0707_),
    .A(net805),
    .Y(_0708_));
 sg13g2_nor2_1 _0927_ (.A(net794),
    .B(_0708_),
    .Y(\latch_mem.genblk1[60].sel_byte ));
 sg13g2_nand4_1 _0928_ (.B(\latch_mem.addr_write[1] ),
    .C(_0662_),
    .A(\latch_mem.addr_write[0] ),
    .Y(_0709_),
    .D(net804));
 sg13g2_nor2_1 _0929_ (.A(net795),
    .B(_0709_),
    .Y(\latch_mem.genblk1[59].sel_byte ));
 sg13g2_nand3_1 _0930_ (.B(net804),
    .C(_0703_),
    .A(_0662_),
    .Y(_0710_));
 sg13g2_nor2_1 _0931_ (.A(net795),
    .B(_0710_),
    .Y(\latch_mem.genblk1[58].sel_byte ));
 sg13g2_nand3_1 _0932_ (.B(net803),
    .C(_0705_),
    .A(_0662_),
    .Y(_0711_));
 sg13g2_nor2_1 _0933_ (.A(net794),
    .B(_0711_),
    .Y(\latch_mem.genblk1[57].sel_byte ));
 sg13g2_nor3_2 _0934_ (.A(\latch_mem.addr_write[0] ),
    .B(\latch_mem.addr_write[1] ),
    .C(\latch_mem.addr_write[2] ),
    .Y(_0712_));
 sg13g2_nand2_2 _0935_ (.Y(_0713_),
    .A(net804),
    .B(_0712_));
 sg13g2_nor2_1 _0936_ (.A(net794),
    .B(_0713_),
    .Y(\latch_mem.genblk1[56].sel_byte ));
 sg13g2_nor2_2 _0937_ (.A(_0662_),
    .B(net803),
    .Y(_0714_));
 sg13g2_nand3_1 _0938_ (.B(\latch_mem.addr_write[1] ),
    .C(_0714_),
    .A(\latch_mem.addr_write[0] ),
    .Y(_0715_));
 sg13g2_nor2_1 _0939_ (.A(net794),
    .B(_0715_),
    .Y(\latch_mem.genblk1[55].sel_byte ));
 sg13g2_nand2_2 _0940_ (.Y(_0716_),
    .A(_0703_),
    .B(_0714_));
 sg13g2_nor2_1 _0941_ (.A(net795),
    .B(_0716_),
    .Y(\latch_mem.genblk1[54].sel_byte ));
 sg13g2_nand2_2 _0942_ (.Y(_0717_),
    .A(_0705_),
    .B(_0714_));
 sg13g2_nor2_1 _0943_ (.A(net794),
    .B(_0717_),
    .Y(\latch_mem.genblk1[53].sel_byte ));
 sg13g2_nand2_2 _0944_ (.Y(_0718_),
    .A(_0707_),
    .B(_0714_));
 sg13g2_nor2_1 _0945_ (.A(net795),
    .B(_0718_),
    .Y(\latch_mem.genblk1[52].sel_byte ));
 sg13g2_nor4_2 _0946_ (.A(_0660_),
    .B(_0661_),
    .C(net805),
    .Y(_0719_),
    .D(net804));
 sg13g2_nor2b_1 _0947_ (.A(net794),
    .B_N(_0719_),
    .Y(\latch_mem.genblk1[51].sel_byte ));
 sg13g2_nor4_2 _0948_ (.A(\latch_mem.addr_write[0] ),
    .B(_0661_),
    .C(net805),
    .Y(_0720_),
    .D(net803));
 sg13g2_nor2b_1 _0949_ (.A(net794),
    .B_N(_0720_),
    .Y(\latch_mem.genblk1[50].sel_byte ));
 sg13g2_nor4_2 _0950_ (.A(_0660_),
    .B(\latch_mem.addr_write[1] ),
    .C(net805),
    .Y(_0721_),
    .D(net804));
 sg13g2_nor2b_1 _0951_ (.A(net795),
    .B_N(_0721_),
    .Y(\latch_mem.genblk1[49].sel_byte ));
 sg13g2_nand2b_2 _0952_ (.Y(_0722_),
    .B(_0712_),
    .A_N(net803));
 sg13g2_nor2_1 _0953_ (.A(net795),
    .B(_0722_),
    .Y(\latch_mem.genblk1[48].sel_byte ));
 sg13g2_nor2b_1 _0954_ (.A(\latch_mem.addr_write[4] ),
    .B_N(\latch_mem.addr_write[5] ),
    .Y(_0723_));
 sg13g2_nand2b_1 _0955_ (.Y(_0724_),
    .B(\latch_mem.addr_write[5] ),
    .A_N(\latch_mem.addr_write[4] ));
 sg13g2_nor2_1 _0956_ (.A(_0701_),
    .B(net793),
    .Y(\latch_mem.genblk1[47].sel_byte ));
 sg13g2_nor2_1 _0957_ (.A(_0704_),
    .B(net792),
    .Y(\latch_mem.genblk1[46].sel_byte ));
 sg13g2_nor2_1 _0958_ (.A(_0706_),
    .B(net792),
    .Y(\latch_mem.genblk1[45].sel_byte ));
 sg13g2_nor2_1 _0959_ (.A(_0708_),
    .B(net793),
    .Y(\latch_mem.genblk1[44].sel_byte ));
 sg13g2_nor2_1 _0960_ (.A(_0709_),
    .B(net792),
    .Y(\latch_mem.genblk1[43].sel_byte ));
 sg13g2_nor2_1 _0961_ (.A(_0710_),
    .B(net792),
    .Y(\latch_mem.genblk1[42].sel_byte ));
 sg13g2_nor2_1 _0962_ (.A(_0711_),
    .B(net793),
    .Y(\latch_mem.genblk1[41].sel_byte ));
 sg13g2_nor2_1 _0963_ (.A(_0713_),
    .B(net792),
    .Y(\latch_mem.genblk1[40].sel_byte ));
 sg13g2_nor2_1 _0964_ (.A(_0715_),
    .B(net792),
    .Y(\latch_mem.genblk1[39].sel_byte ));
 sg13g2_nor2_1 _0965_ (.A(_0716_),
    .B(net792),
    .Y(\latch_mem.genblk1[38].sel_byte ));
 sg13g2_nor2_1 _0966_ (.A(_0717_),
    .B(net793),
    .Y(\latch_mem.genblk1[37].sel_byte ));
 sg13g2_nor2_1 _0967_ (.A(_0718_),
    .B(net792),
    .Y(\latch_mem.genblk1[36].sel_byte ));
 sg13g2_and2_1 _0968_ (.A(_0719_),
    .B(_0723_),
    .X(\latch_mem.genblk1[35].sel_byte ));
 sg13g2_and2_1 _0969_ (.A(_0720_),
    .B(_0723_),
    .X(\latch_mem.genblk1[34].sel_byte ));
 sg13g2_and2_1 _0970_ (.A(_0721_),
    .B(_0723_),
    .X(\latch_mem.genblk1[33].sel_byte ));
 sg13g2_nor2_1 _0971_ (.A(_0722_),
    .B(net793),
    .Y(\latch_mem.genblk1[32].sel_byte ));
 sg13g2_nor2b_1 _0972_ (.A(\latch_mem.addr_write[5] ),
    .B_N(\latch_mem.addr_write[4] ),
    .Y(_0725_));
 sg13g2_nand2b_1 _0973_ (.Y(_0726_),
    .B(\latch_mem.addr_write[4] ),
    .A_N(\latch_mem.addr_write[5] ));
 sg13g2_nor2_1 _0974_ (.A(_0701_),
    .B(net790),
    .Y(\latch_mem.genblk1[31].sel_byte ));
 sg13g2_nor2_1 _0975_ (.A(_0704_),
    .B(net791),
    .Y(\latch_mem.genblk1[30].sel_byte ));
 sg13g2_nor2_1 _0976_ (.A(_0706_),
    .B(net790),
    .Y(\latch_mem.genblk1[29].sel_byte ));
 sg13g2_nor2_1 _0977_ (.A(_0708_),
    .B(net791),
    .Y(\latch_mem.genblk1[28].sel_byte ));
 sg13g2_nor2_1 _0978_ (.A(_0709_),
    .B(net791),
    .Y(\latch_mem.genblk1[27].sel_byte ));
 sg13g2_nor2_1 _0979_ (.A(_0710_),
    .B(net790),
    .Y(\latch_mem.genblk1[26].sel_byte ));
 sg13g2_nor2_1 _0980_ (.A(_0711_),
    .B(net791),
    .Y(\latch_mem.genblk1[25].sel_byte ));
 sg13g2_nor2_1 _0981_ (.A(_0713_),
    .B(net790),
    .Y(\latch_mem.genblk1[24].sel_byte ));
 sg13g2_nor2_1 _0982_ (.A(_0715_),
    .B(net790),
    .Y(\latch_mem.genblk1[23].sel_byte ));
 sg13g2_nor2_1 _0983_ (.A(_0716_),
    .B(net790),
    .Y(\latch_mem.genblk1[22].sel_byte ));
 sg13g2_nor2_1 _0984_ (.A(_0717_),
    .B(net790),
    .Y(\latch_mem.genblk1[21].sel_byte ));
 sg13g2_nor2_1 _0985_ (.A(_0718_),
    .B(net790),
    .Y(\latch_mem.genblk1[20].sel_byte ));
 sg13g2_and2_1 _0986_ (.A(_0719_),
    .B(_0725_),
    .X(\latch_mem.genblk1[19].sel_byte ));
 sg13g2_and2_1 _0987_ (.A(_0720_),
    .B(_0725_),
    .X(\latch_mem.genblk1[18].sel_byte ));
 sg13g2_and2_1 _0988_ (.A(_0721_),
    .B(_0725_),
    .X(\latch_mem.genblk1[17].sel_byte ));
 sg13g2_nor2_1 _0989_ (.A(_0722_),
    .B(net791),
    .Y(\latch_mem.genblk1[16].sel_byte ));
 sg13g2_nor2_1 _0990_ (.A(\latch_mem.addr_write[4] ),
    .B(\latch_mem.addr_write[5] ),
    .Y(_0727_));
 sg13g2_or2_1 _0991_ (.X(_0728_),
    .B(\latch_mem.addr_write[5] ),
    .A(\latch_mem.addr_write[4] ));
 sg13g2_nor2_1 _0992_ (.A(_0701_),
    .B(net788),
    .Y(\latch_mem.genblk1[15].sel_byte ));
 sg13g2_nor2_1 _0993_ (.A(_0704_),
    .B(net789),
    .Y(\latch_mem.genblk1[14].sel_byte ));
 sg13g2_nor2_1 _0994_ (.A(_0706_),
    .B(net788),
    .Y(\latch_mem.genblk1[13].sel_byte ));
 sg13g2_nor2_1 _0995_ (.A(_0708_),
    .B(net788),
    .Y(\latch_mem.genblk1[12].sel_byte ));
 sg13g2_nor2_1 _0996_ (.A(_0709_),
    .B(net789),
    .Y(\latch_mem.genblk1[11].sel_byte ));
 sg13g2_nor2_1 _0997_ (.A(_0710_),
    .B(net789),
    .Y(\latch_mem.genblk1[10].sel_byte ));
 sg13g2_nor2_1 _0998_ (.A(_0711_),
    .B(net788),
    .Y(\latch_mem.genblk1[9].sel_byte ));
 sg13g2_nor2_1 _0999_ (.A(_0713_),
    .B(net788),
    .Y(\latch_mem.genblk1[8].sel_byte ));
 sg13g2_nor2_1 _1000_ (.A(_0715_),
    .B(net788),
    .Y(\latch_mem.genblk1[7].sel_byte ));
 sg13g2_nor2_1 _1001_ (.A(_0716_),
    .B(net788),
    .Y(\latch_mem.genblk1[6].sel_byte ));
 sg13g2_nor2_1 _1002_ (.A(_0717_),
    .B(net788),
    .Y(\latch_mem.genblk1[5].sel_byte ));
 sg13g2_nor2_1 _1003_ (.A(_0718_),
    .B(net789),
    .Y(\latch_mem.genblk1[4].sel_byte ));
 sg13g2_and2_1 _1004_ (.A(_0719_),
    .B(_0727_),
    .X(\latch_mem.genblk1[3].sel_byte ));
 sg13g2_and2_1 _1005_ (.A(_0720_),
    .B(_0727_),
    .X(\latch_mem.genblk1[2].sel_byte ));
 sg13g2_and2_1 _1006_ (.A(_0721_),
    .B(_0727_),
    .X(\latch_mem.genblk1[1].sel_byte ));
 sg13g2_nor2_1 _1007_ (.A(_0722_),
    .B(net789),
    .Y(\latch_mem.genblk1[0].sel_byte ));
 sg13g2_and2_2 _1008_ (.A(\latch_mem.wr_en_valid ),
    .B(\latch_mem.wr_en_ok ),
    .X(\latch_mem.wr_en ));
 sg13g2_nand2b_2 _1009_ (.Y(_0729_),
    .B(\latch_mem.addr_read[1] ),
    .A_N(\latch_mem.addr_read[0] ));
 sg13g2_nor3_1 _1010_ (.A(\latch_mem.addr_read[2] ),
    .B(\latch_mem.addr_read[3] ),
    .C(_0729_),
    .Y(_0730_));
 sg13g2_nor4_1 _1011_ (.A(\latch_mem.addr_read[2] ),
    .B(\latch_mem.addr_read[3] ),
    .C(\latch_mem.addr_read[1] ),
    .D(\latch_mem.addr_read[0] ),
    .Y(_0731_));
 sg13g2_nand2b_1 _1012_ (.Y(_0732_),
    .B(\latch_mem.addr_read[0] ),
    .A_N(\latch_mem.addr_read[1] ));
 sg13g2_nor3_1 _1013_ (.A(\latch_mem.addr_read[2] ),
    .B(\latch_mem.addr_read[3] ),
    .C(_0732_),
    .Y(_0733_));
 sg13g2_nand2_2 _1014_ (.Y(_0734_),
    .A(\latch_mem.addr_read[1] ),
    .B(\latch_mem.addr_read[0] ));
 sg13g2_nand2b_2 _1015_ (.Y(_0735_),
    .B(\latch_mem.addr_read[2] ),
    .A_N(\latch_mem.addr_read[3] ));
 sg13g2_nor2_2 _1016_ (.A(_0734_),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_nand2_2 _1017_ (.Y(_0737_),
    .A(\latch_mem.addr_read[2] ),
    .B(\latch_mem.addr_read[3] ));
 sg13g2_nor2_2 _1018_ (.A(_0734_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_nor3_2 _1019_ (.A(\latch_mem.addr_read[2] ),
    .B(\latch_mem.addr_read[3] ),
    .C(_0734_),
    .Y(_0739_));
 sg13g2_nand2b_2 _1020_ (.Y(_0740_),
    .B(\latch_mem.addr_read[3] ),
    .A_N(\latch_mem.addr_read[2] ));
 sg13g2_nor2_1 _1021_ (.A(_0732_),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_nor3_1 _1022_ (.A(\latch_mem.addr_read[1] ),
    .B(\latch_mem.addr_read[0] ),
    .C(_0735_),
    .Y(_0742_));
 sg13g2_nor3_1 _1023_ (.A(\latch_mem.addr_read[1] ),
    .B(\latch_mem.addr_read[0] ),
    .C(_0740_),
    .Y(_0743_));
 sg13g2_nor2_1 _1024_ (.A(_0729_),
    .B(_0735_),
    .Y(_0744_));
 sg13g2_a22oi_1 _1025_ (.Y(_0745_),
    .B1(net726),
    .B2(\latch_mem.RAM[54][0] ),
    .A2(net731),
    .A1(\latch_mem.RAM[56][0] ));
 sg13g2_nor2_1 _1026_ (.A(_0732_),
    .B(_0737_),
    .Y(_0746_));
 sg13g2_nor2_2 _1027_ (.A(_0729_),
    .B(_0737_),
    .Y(_0747_));
 sg13g2_nor3_1 _1028_ (.A(\latch_mem.addr_read[1] ),
    .B(\latch_mem.addr_read[0] ),
    .C(_0737_),
    .Y(_0748_));
 sg13g2_nor2_2 _1029_ (.A(_0729_),
    .B(_0740_),
    .Y(_0749_));
 sg13g2_nor2_1 _1030_ (.A(_0732_),
    .B(_0735_),
    .Y(_0750_));
 sg13g2_nor2_1 _1031_ (.A(_0734_),
    .B(_0740_),
    .Y(_0751_));
 sg13g2_a22oi_1 _1032_ (.Y(_0752_),
    .B1(net753),
    .B2(\latch_mem.RAM[63][0] ),
    .A2(net762),
    .A1(\latch_mem.RAM[49][0] ));
 sg13g2_a22oi_1 _1033_ (.Y(_0753_),
    .B1(net711),
    .B2(\latch_mem.RAM[60][0] ),
    .A2(net742),
    .A1(\latch_mem.RAM[57][0] ));
 sg13g2_a22oi_1 _1034_ (.Y(_0754_),
    .B1(net757),
    .B2(\latch_mem.RAM[55][0] ),
    .A2(net764),
    .A1(\latch_mem.RAM[50][0] ));
 sg13g2_a22oi_1 _1035_ (.Y(_0755_),
    .B1(net701),
    .B2(\latch_mem.RAM[53][0] ),
    .A2(net786),
    .A1(\latch_mem.RAM[48][0] ));
 sg13g2_nand4_1 _1036_ (.B(_0753_),
    .C(_0754_),
    .A(_0752_),
    .Y(_0756_),
    .D(_0755_));
 sg13g2_a22oi_1 _1037_ (.Y(_0757_),
    .B1(net707),
    .B2(\latch_mem.RAM[58][0] ),
    .A2(net736),
    .A1(\latch_mem.RAM[52][0] ));
 sg13g2_a22oi_1 _1038_ (.Y(_0758_),
    .B1(net721),
    .B2(\latch_mem.RAM[61][0] ),
    .A2(net747),
    .A1(\latch_mem.RAM[51][0] ));
 sg13g2_a22oi_1 _1039_ (.Y(_0759_),
    .B1(net696),
    .B2(\latch_mem.RAM[59][0] ),
    .A2(net716),
    .A1(\latch_mem.RAM[62][0] ));
 sg13g2_nand4_1 _1040_ (.B(_0757_),
    .C(_0758_),
    .A(_0745_),
    .Y(_0760_),
    .D(_0759_));
 sg13g2_or2_1 _1041_ (.X(\latch_mem.genblk2[3].selected_out[0] ),
    .B(_0760_),
    .A(_0756_));
 sg13g2_a22oi_1 _1042_ (.Y(_0761_),
    .B1(net696),
    .B2(\latch_mem.RAM[59][1] ),
    .A2(net761),
    .A1(\latch_mem.RAM[49][1] ));
 sg13g2_a22oi_1 _1043_ (.Y(_0762_),
    .B1(net721),
    .B2(\latch_mem.RAM[61][1] ),
    .A2(net752),
    .A1(\latch_mem.RAM[63][1] ));
 sg13g2_a22oi_1 _1044_ (.Y(_0763_),
    .B1(net711),
    .B2(\latch_mem.RAM[60][1] ),
    .A2(net766),
    .A1(\latch_mem.RAM[50][1] ));
 sg13g2_a22oi_1 _1045_ (.Y(_0764_),
    .B1(net701),
    .B2(\latch_mem.RAM[53][1] ),
    .A2(net747),
    .A1(\latch_mem.RAM[51][1] ));
 sg13g2_a22oi_1 _1046_ (.Y(_0765_),
    .B1(net716),
    .B2(\latch_mem.RAM[62][1] ),
    .A2(net736),
    .A1(\latch_mem.RAM[52][1] ));
 sg13g2_nand4_1 _1047_ (.B(_0763_),
    .C(_0764_),
    .A(_0762_),
    .Y(_0766_),
    .D(_0765_));
 sg13g2_a22oi_1 _1048_ (.Y(_0767_),
    .B1(net731),
    .B2(\latch_mem.RAM[56][1] ),
    .A2(net741),
    .A1(\latch_mem.RAM[57][1] ));
 sg13g2_a22oi_1 _1049_ (.Y(_0768_),
    .B1(net707),
    .B2(\latch_mem.RAM[58][1] ),
    .A2(net786),
    .A1(\latch_mem.RAM[48][1] ));
 sg13g2_a22oi_1 _1050_ (.Y(_0769_),
    .B1(net726),
    .B2(\latch_mem.RAM[54][1] ),
    .A2(_0736_),
    .A1(\latch_mem.RAM[55][1] ));
 sg13g2_nand4_1 _1051_ (.B(_0767_),
    .C(_0768_),
    .A(_0761_),
    .Y(_0770_),
    .D(_0769_));
 sg13g2_or2_1 _1052_ (.X(\latch_mem.genblk2[3].selected_out[1] ),
    .B(_0770_),
    .A(_0766_));
 sg13g2_a22oi_1 _1053_ (.Y(_0089_),
    .B1(net732),
    .B2(\latch_mem.RAM[56][2] ),
    .A2(net748),
    .A1(\latch_mem.RAM[51][2] ));
 sg13g2_a22oi_1 _1054_ (.Y(_0090_),
    .B1(net707),
    .B2(\latch_mem.RAM[58][2] ),
    .A2(net761),
    .A1(\latch_mem.RAM[49][2] ));
 sg13g2_a22oi_1 _1055_ (.Y(_0091_),
    .B1(net736),
    .B2(\latch_mem.RAM[52][2] ),
    .A2(net741),
    .A1(\latch_mem.RAM[57][2] ));
 sg13g2_a22oi_1 _1056_ (.Y(_0092_),
    .B1(net696),
    .B2(\latch_mem.RAM[59][2] ),
    .A2(net727),
    .A1(\latch_mem.RAM[54][2] ));
 sg13g2_a22oi_1 _1057_ (.Y(_0093_),
    .B1(net701),
    .B2(\latch_mem.RAM[53][2] ),
    .A2(net716),
    .A1(\latch_mem.RAM[62][2] ));
 sg13g2_a22oi_1 _1058_ (.Y(_0094_),
    .B1(net721),
    .B2(\latch_mem.RAM[61][2] ),
    .A2(net752),
    .A1(\latch_mem.RAM[63][2] ));
 sg13g2_nand4_1 _1059_ (.B(_0091_),
    .C(_0093_),
    .A(_0090_),
    .Y(_0095_),
    .D(_0094_));
 sg13g2_a22oi_1 _1060_ (.Y(_0096_),
    .B1(net786),
    .B2(\latch_mem.RAM[48][2] ),
    .A2(net766),
    .A1(\latch_mem.RAM[50][2] ));
 sg13g2_a22oi_1 _1061_ (.Y(_0097_),
    .B1(net711),
    .B2(\latch_mem.RAM[60][2] ),
    .A2(net757),
    .A1(\latch_mem.RAM[55][2] ));
 sg13g2_nand4_1 _1062_ (.B(_0092_),
    .C(_0096_),
    .A(_0089_),
    .Y(_0098_),
    .D(_0097_));
 sg13g2_or2_1 _1063_ (.X(\latch_mem.genblk2[3].selected_out[2] ),
    .B(_0098_),
    .A(_0095_));
 sg13g2_a22oi_1 _1064_ (.Y(_0099_),
    .B1(net716),
    .B2(\latch_mem.RAM[62][3] ),
    .A2(net786),
    .A1(\latch_mem.RAM[48][3] ));
 sg13g2_a22oi_1 _1065_ (.Y(_0100_),
    .B1(net707),
    .B2(\latch_mem.RAM[58][3] ),
    .A2(net736),
    .A1(\latch_mem.RAM[52][3] ));
 sg13g2_a22oi_1 _1066_ (.Y(_0101_),
    .B1(net753),
    .B2(\latch_mem.RAM[63][3] ),
    .A2(net766),
    .A1(\latch_mem.RAM[50][3] ));
 sg13g2_a22oi_1 _1067_ (.Y(_0102_),
    .B1(net742),
    .B2(\latch_mem.RAM[57][3] ),
    .A2(net757),
    .A1(\latch_mem.RAM[55][3] ));
 sg13g2_a22oi_1 _1068_ (.Y(_0103_),
    .B1(net731),
    .B2(\latch_mem.RAM[56][3] ),
    .A2(net747),
    .A1(\latch_mem.RAM[51][3] ));
 sg13g2_a22oi_1 _1069_ (.Y(_0104_),
    .B1(net711),
    .B2(\latch_mem.RAM[60][3] ),
    .A2(net721),
    .A1(\latch_mem.RAM[61][3] ));
 sg13g2_nand4_1 _1070_ (.B(_0100_),
    .C(_0103_),
    .A(_0099_),
    .Y(_0105_),
    .D(_0104_));
 sg13g2_a22oi_1 _1071_ (.Y(_0106_),
    .B1(net701),
    .B2(\latch_mem.RAM[53][3] ),
    .A2(net762),
    .A1(\latch_mem.RAM[49][3] ));
 sg13g2_a22oi_1 _1072_ (.Y(_0107_),
    .B1(net696),
    .B2(\latch_mem.RAM[59][3] ),
    .A2(net727),
    .A1(\latch_mem.RAM[54][3] ));
 sg13g2_nand4_1 _1073_ (.B(_0102_),
    .C(_0106_),
    .A(_0101_),
    .Y(_0108_),
    .D(_0107_));
 sg13g2_or2_1 _1074_ (.X(\latch_mem.genblk2[3].selected_out[3] ),
    .B(_0108_),
    .A(_0105_));
 sg13g2_a22oi_1 _1075_ (.Y(_0109_),
    .B1(net716),
    .B2(\latch_mem.RAM[62][4] ),
    .A2(net752),
    .A1(\latch_mem.RAM[63][4] ));
 sg13g2_a22oi_1 _1076_ (.Y(_0110_),
    .B1(net707),
    .B2(\latch_mem.RAM[58][4] ),
    .A2(net721),
    .A1(\latch_mem.RAM[61][4] ));
 sg13g2_a22oi_1 _1077_ (.Y(_0111_),
    .B1(net736),
    .B2(\latch_mem.RAM[52][4] ),
    .A2(net766),
    .A1(\latch_mem.RAM[50][4] ));
 sg13g2_a22oi_1 _1078_ (.Y(_0112_),
    .B1(net696),
    .B2(\latch_mem.RAM[59][4] ),
    .A2(net731),
    .A1(\latch_mem.RAM[56][4] ));
 sg13g2_nand4_1 _1079_ (.B(_0110_),
    .C(_0111_),
    .A(_0109_),
    .Y(_0113_),
    .D(_0112_));
 sg13g2_a22oi_1 _1080_ (.Y(_0114_),
    .B1(net742),
    .B2(\latch_mem.RAM[57][4] ),
    .A2(net762),
    .A1(\latch_mem.RAM[49][4] ));
 sg13g2_a22oi_1 _1081_ (.Y(_0115_),
    .B1(net701),
    .B2(\latch_mem.RAM[53][4] ),
    .A2(net757),
    .A1(\latch_mem.RAM[55][4] ));
 sg13g2_a22oi_1 _1082_ (.Y(_0116_),
    .B1(net727),
    .B2(\latch_mem.RAM[54][4] ),
    .A2(net786),
    .A1(\latch_mem.RAM[48][4] ));
 sg13g2_a22oi_1 _1083_ (.Y(_0117_),
    .B1(net711),
    .B2(\latch_mem.RAM[60][4] ),
    .A2(net748),
    .A1(\latch_mem.RAM[51][4] ));
 sg13g2_nand4_1 _1084_ (.B(_0115_),
    .C(_0116_),
    .A(_0114_),
    .Y(_0118_),
    .D(_0117_));
 sg13g2_or2_1 _1085_ (.X(\latch_mem.genblk2[3].selected_out[4] ),
    .B(_0118_),
    .A(_0113_));
 sg13g2_a22oi_1 _1086_ (.Y(_0119_),
    .B1(net716),
    .B2(\latch_mem.RAM[62][5] ),
    .A2(net747),
    .A1(\latch_mem.RAM[51][5] ));
 sg13g2_a22oi_1 _1087_ (.Y(_0120_),
    .B1(net707),
    .B2(\latch_mem.RAM[58][5] ),
    .A2(net726),
    .A1(\latch_mem.RAM[54][5] ));
 sg13g2_a22oi_1 _1088_ (.Y(_0121_),
    .B1(net711),
    .B2(\latch_mem.RAM[60][5] ),
    .A2(net732),
    .A1(\latch_mem.RAM[56][5] ));
 sg13g2_a22oi_1 _1089_ (.Y(_0122_),
    .B1(net721),
    .B2(\latch_mem.RAM[61][5] ),
    .A2(net741),
    .A1(\latch_mem.RAM[57][5] ));
 sg13g2_a22oi_1 _1090_ (.Y(_0123_),
    .B1(net696),
    .B2(\latch_mem.RAM[59][5] ),
    .A2(net786),
    .A1(\latch_mem.RAM[48][5] ));
 sg13g2_nand4_1 _1091_ (.B(_0120_),
    .C(_0122_),
    .A(_0119_),
    .Y(_0124_),
    .D(_0123_));
 sg13g2_a22oi_1 _1092_ (.Y(_0125_),
    .B1(net737),
    .B2(\latch_mem.RAM[52][5] ),
    .A2(net762),
    .A1(\latch_mem.RAM[49][5] ));
 sg13g2_a22oi_1 _1093_ (.Y(_0126_),
    .B1(net753),
    .B2(\latch_mem.RAM[63][5] ),
    .A2(net757),
    .A1(\latch_mem.RAM[55][5] ));
 sg13g2_a22oi_1 _1094_ (.Y(_0127_),
    .B1(net701),
    .B2(\latch_mem.RAM[53][5] ),
    .A2(net766),
    .A1(\latch_mem.RAM[50][5] ));
 sg13g2_nand4_1 _1095_ (.B(_0125_),
    .C(_0126_),
    .A(_0121_),
    .Y(_0128_),
    .D(_0127_));
 sg13g2_or2_1 _1096_ (.X(\latch_mem.genblk2[3].selected_out[5] ),
    .B(_0128_),
    .A(_0124_));
 sg13g2_a22oi_1 _1097_ (.Y(_0129_),
    .B1(net732),
    .B2(\latch_mem.RAM[56][6] ),
    .A2(net766),
    .A1(\latch_mem.RAM[50][6] ));
 sg13g2_a22oi_1 _1098_ (.Y(_0130_),
    .B1(net707),
    .B2(\latch_mem.RAM[58][6] ),
    .A2(net716),
    .A1(\latch_mem.RAM[62][6] ));
 sg13g2_a22oi_1 _1099_ (.Y(_0131_),
    .B1(net701),
    .B2(\latch_mem.RAM[53][6] ),
    .A2(net737),
    .A1(\latch_mem.RAM[52][6] ));
 sg13g2_a22oi_1 _1100_ (.Y(_0132_),
    .B1(net711),
    .B2(\latch_mem.RAM[60][6] ),
    .A2(net741),
    .A1(\latch_mem.RAM[57][6] ));
 sg13g2_a22oi_1 _1101_ (.Y(_0133_),
    .B1(net721),
    .B2(\latch_mem.RAM[61][6] ),
    .A2(net726),
    .A1(\latch_mem.RAM[54][6] ));
 sg13g2_a22oi_1 _1102_ (.Y(_0134_),
    .B1(net752),
    .B2(\latch_mem.RAM[63][6] ),
    .A2(net786),
    .A1(\latch_mem.RAM[48][6] ));
 sg13g2_a22oi_1 _1103_ (.Y(_0135_),
    .B1(net758),
    .B2(\latch_mem.RAM[55][6] ),
    .A2(net761),
    .A1(\latch_mem.RAM[49][6] ));
 sg13g2_nand4_1 _1104_ (.B(_0133_),
    .C(_0134_),
    .A(_0130_),
    .Y(_0136_),
    .D(_0135_));
 sg13g2_a22oi_1 _1105_ (.Y(_0137_),
    .B1(net696),
    .B2(\latch_mem.RAM[59][6] ),
    .A2(net747),
    .A1(\latch_mem.RAM[51][6] ));
 sg13g2_nand4_1 _1106_ (.B(_0131_),
    .C(_0132_),
    .A(_0129_),
    .Y(_0138_),
    .D(_0137_));
 sg13g2_or2_1 _1107_ (.X(\latch_mem.genblk2[3].selected_out[6] ),
    .B(_0138_),
    .A(_0136_));
 sg13g2_a22oi_1 _1108_ (.Y(_0139_),
    .B1(net718),
    .B2(\latch_mem.RAM[62][7] ),
    .A2(net721),
    .A1(\latch_mem.RAM[61][7] ));
 sg13g2_a22oi_1 _1109_ (.Y(_0140_),
    .B1(net732),
    .B2(\latch_mem.RAM[56][7] ),
    .A2(net766),
    .A1(\latch_mem.RAM[50][7] ));
 sg13g2_a22oi_1 _1110_ (.Y(_0141_),
    .B1(net701),
    .B2(\latch_mem.RAM[53][7] ),
    .A2(net786),
    .A1(\latch_mem.RAM[48][7] ));
 sg13g2_a22oi_1 _1111_ (.Y(_0142_),
    .B1(net737),
    .B2(\latch_mem.RAM[52][7] ),
    .A2(net762),
    .A1(\latch_mem.RAM[49][7] ));
 sg13g2_nand4_1 _1112_ (.B(_0140_),
    .C(_0141_),
    .A(_0139_),
    .Y(_0143_),
    .D(_0142_));
 sg13g2_a22oi_1 _1113_ (.Y(_0144_),
    .B1(net711),
    .B2(\latch_mem.RAM[60][7] ),
    .A2(net758),
    .A1(\latch_mem.RAM[55][7] ));
 sg13g2_a22oi_1 _1114_ (.Y(_0145_),
    .B1(net707),
    .B2(\latch_mem.RAM[58][7] ),
    .A2(net747),
    .A1(\latch_mem.RAM[51][7] ));
 sg13g2_a22oi_1 _1115_ (.Y(_0146_),
    .B1(net726),
    .B2(\latch_mem.RAM[54][7] ),
    .A2(net752),
    .A1(\latch_mem.RAM[63][7] ));
 sg13g2_a22oi_1 _1116_ (.Y(_0147_),
    .B1(net696),
    .B2(\latch_mem.RAM[59][7] ),
    .A2(net741),
    .A1(\latch_mem.RAM[57][7] ));
 sg13g2_nand4_1 _1117_ (.B(_0145_),
    .C(_0146_),
    .A(_0144_),
    .Y(_0148_),
    .D(_0147_));
 sg13g2_or2_1 _1118_ (.X(\latch_mem.genblk2[3].selected_out[7] ),
    .B(_0148_),
    .A(_0143_));
 sg13g2_a22oi_1 _1119_ (.Y(_0149_),
    .B1(net705),
    .B2(\latch_mem.RAM[42][0] ),
    .A2(net710),
    .A1(\latch_mem.RAM[44][0] ));
 sg13g2_a22oi_1 _1120_ (.Y(_0150_),
    .B1(net700),
    .B2(\latch_mem.RAM[37][0] ),
    .A2(net725),
    .A1(\latch_mem.RAM[38][0] ));
 sg13g2_a22oi_1 _1121_ (.Y(_0151_),
    .B1(net715),
    .B2(\latch_mem.RAM[46][0] ),
    .A2(net740),
    .A1(\latch_mem.RAM[41][0] ));
 sg13g2_a22oi_1 _1122_ (.Y(_0152_),
    .B1(net720),
    .B2(\latch_mem.RAM[45][0] ),
    .A2(net783),
    .A1(\latch_mem.RAM[32][0] ));
 sg13g2_nand4_1 _1123_ (.B(_0150_),
    .C(_0151_),
    .A(_0149_),
    .Y(_0153_),
    .D(_0152_));
 sg13g2_a22oi_1 _1124_ (.Y(_0154_),
    .B1(net695),
    .B2(\latch_mem.RAM[43][0] ),
    .A2(net756),
    .A1(\latch_mem.RAM[39][0] ));
 sg13g2_a22oi_1 _1125_ (.Y(_0155_),
    .B1(net730),
    .B2(\latch_mem.RAM[40][0] ),
    .A2(net768),
    .A1(\latch_mem.RAM[34][0] ));
 sg13g2_a22oi_1 _1126_ (.Y(_0156_),
    .B1(net735),
    .B2(\latch_mem.RAM[36][0] ),
    .A2(net751),
    .A1(\latch_mem.RAM[47][0] ));
 sg13g2_a22oi_1 _1127_ (.Y(_0157_),
    .B1(net746),
    .B2(\latch_mem.RAM[35][0] ),
    .A2(net760),
    .A1(\latch_mem.RAM[33][0] ));
 sg13g2_nand4_1 _1128_ (.B(_0155_),
    .C(_0156_),
    .A(_0154_),
    .Y(_0158_),
    .D(_0157_));
 sg13g2_or2_1 _1129_ (.X(\latch_mem.genblk2[2].selected_out[0] ),
    .B(_0158_),
    .A(_0153_));
 sg13g2_a22oi_1 _1130_ (.Y(_0159_),
    .B1(net720),
    .B2(\latch_mem.RAM[45][1] ),
    .A2(net745),
    .A1(\latch_mem.RAM[35][1] ));
 sg13g2_a22oi_1 _1131_ (.Y(_0160_),
    .B1(net760),
    .B2(\latch_mem.RAM[33][1] ),
    .A2(net768),
    .A1(\latch_mem.RAM[34][1] ));
 sg13g2_a22oi_1 _1132_ (.Y(_0161_),
    .B1(net700),
    .B2(\latch_mem.RAM[37][1] ),
    .A2(net755),
    .A1(\latch_mem.RAM[39][1] ));
 sg13g2_a22oi_1 _1133_ (.Y(_0162_),
    .B1(net729),
    .B2(\latch_mem.RAM[40][1] ),
    .A2(net783),
    .A1(\latch_mem.RAM[32][1] ));
 sg13g2_a22oi_1 _1134_ (.Y(_0163_),
    .B1(net735),
    .B2(\latch_mem.RAM[36][1] ),
    .A2(net750),
    .A1(\latch_mem.RAM[47][1] ));
 sg13g2_nand4_1 _1135_ (.B(_0161_),
    .C(_0162_),
    .A(_0160_),
    .Y(_0164_),
    .D(_0163_));
 sg13g2_a22oi_1 _1136_ (.Y(_0165_),
    .B1(net710),
    .B2(\latch_mem.RAM[44][1] ),
    .A2(net725),
    .A1(\latch_mem.RAM[38][1] ));
 sg13g2_a22oi_1 _1137_ (.Y(_0166_),
    .B1(net695),
    .B2(\latch_mem.RAM[43][1] ),
    .A2(net740),
    .A1(\latch_mem.RAM[41][1] ));
 sg13g2_a22oi_1 _1138_ (.Y(_0167_),
    .B1(net705),
    .B2(\latch_mem.RAM[42][1] ),
    .A2(net715),
    .A1(\latch_mem.RAM[46][1] ));
 sg13g2_nand4_1 _1139_ (.B(_0165_),
    .C(_0166_),
    .A(_0159_),
    .Y(_0168_),
    .D(_0167_));
 sg13g2_or2_1 _1140_ (.X(\latch_mem.genblk2[2].selected_out[1] ),
    .B(_0168_),
    .A(_0164_));
 sg13g2_a22oi_1 _1141_ (.Y(_0169_),
    .B1(net700),
    .B2(\latch_mem.RAM[37][2] ),
    .A2(net765),
    .A1(\latch_mem.RAM[34][2] ));
 sg13g2_a22oi_1 _1142_ (.Y(_0170_),
    .B1(net710),
    .B2(\latch_mem.RAM[44][2] ),
    .A2(net714),
    .A1(\latch_mem.RAM[46][2] ));
 sg13g2_a22oi_1 _1143_ (.Y(_0171_),
    .B1(net735),
    .B2(\latch_mem.RAM[36][2] ),
    .A2(net755),
    .A1(\latch_mem.RAM[39][2] ));
 sg13g2_a22oi_1 _1144_ (.Y(_0172_),
    .B1(net705),
    .B2(\latch_mem.RAM[42][2] ),
    .A2(net745),
    .A1(\latch_mem.RAM[35][2] ));
 sg13g2_a22oi_1 _1145_ (.Y(_0173_),
    .B1(net720),
    .B2(\latch_mem.RAM[45][2] ),
    .A2(net725),
    .A1(\latch_mem.RAM[38][2] ));
 sg13g2_nand4_1 _1146_ (.B(_0171_),
    .C(_0172_),
    .A(_0170_),
    .Y(_0174_),
    .D(_0173_));
 sg13g2_a22oi_1 _1147_ (.Y(_0175_),
    .B1(net695),
    .B2(\latch_mem.RAM[43][2] ),
    .A2(net760),
    .A1(\latch_mem.RAM[33][2] ));
 sg13g2_a22oi_1 _1148_ (.Y(_0176_),
    .B1(net740),
    .B2(\latch_mem.RAM[41][2] ),
    .A2(net751),
    .A1(\latch_mem.RAM[47][2] ));
 sg13g2_a22oi_1 _1149_ (.Y(_0177_),
    .B1(net730),
    .B2(\latch_mem.RAM[40][2] ),
    .A2(net783),
    .A1(\latch_mem.RAM[32][2] ));
 sg13g2_nand4_1 _1150_ (.B(_0175_),
    .C(_0176_),
    .A(_0169_),
    .Y(_0178_),
    .D(_0177_));
 sg13g2_or2_1 _1151_ (.X(\latch_mem.genblk2[2].selected_out[2] ),
    .B(_0178_),
    .A(_0174_));
 sg13g2_a22oi_1 _1152_ (.Y(_0179_),
    .B1(net720),
    .B2(\latch_mem.RAM[45][3] ),
    .A2(net759),
    .A1(\latch_mem.RAM[33][3] ));
 sg13g2_a22oi_1 _1153_ (.Y(_0180_),
    .B1(net704),
    .B2(\latch_mem.RAM[42][3] ),
    .A2(net710),
    .A1(\latch_mem.RAM[44][3] ));
 sg13g2_a22oi_1 _1154_ (.Y(_0181_),
    .B1(net695),
    .B2(\latch_mem.RAM[43][3] ),
    .A2(net730),
    .A1(\latch_mem.RAM[40][3] ));
 sg13g2_a22oi_1 _1155_ (.Y(_0182_),
    .B1(net725),
    .B2(\latch_mem.RAM[38][3] ),
    .A2(net734),
    .A1(\latch_mem.RAM[36][3] ));
 sg13g2_nand4_1 _1156_ (.B(_0180_),
    .C(_0181_),
    .A(_0179_),
    .Y(_0183_),
    .D(_0182_));
 sg13g2_a22oi_1 _1157_ (.Y(_0184_),
    .B1(net755),
    .B2(\latch_mem.RAM[39][3] ),
    .A2(net765),
    .A1(\latch_mem.RAM[34][3] ));
 sg13g2_a22oi_1 _1158_ (.Y(_0185_),
    .B1(net714),
    .B2(\latch_mem.RAM[46][3] ),
    .A2(net750),
    .A1(\latch_mem.RAM[47][3] ));
 sg13g2_a22oi_1 _1159_ (.Y(_0186_),
    .B1(net700),
    .B2(\latch_mem.RAM[37][3] ),
    .A2(net783),
    .A1(\latch_mem.RAM[32][3] ));
 sg13g2_a22oi_1 _1160_ (.Y(_0187_),
    .B1(net740),
    .B2(\latch_mem.RAM[41][3] ),
    .A2(net745),
    .A1(\latch_mem.RAM[35][3] ));
 sg13g2_nand4_1 _1161_ (.B(_0185_),
    .C(_0186_),
    .A(_0184_),
    .Y(_0188_),
    .D(_0187_));
 sg13g2_or2_1 _1162_ (.X(\latch_mem.genblk2[2].selected_out[3] ),
    .B(_0188_),
    .A(_0183_));
 sg13g2_a22oi_1 _1163_ (.Y(_0189_),
    .B1(net695),
    .B2(\latch_mem.RAM[43][4] ),
    .A2(net730),
    .A1(\latch_mem.RAM[40][4] ));
 sg13g2_a22oi_1 _1164_ (.Y(_0190_),
    .B1(net700),
    .B2(\latch_mem.RAM[37][4] ),
    .A2(net765),
    .A1(\latch_mem.RAM[34][4] ));
 sg13g2_a22oi_1 _1165_ (.Y(_0191_),
    .B1(net734),
    .B2(\latch_mem.RAM[36][4] ),
    .A2(net755),
    .A1(\latch_mem.RAM[39][4] ));
 sg13g2_a22oi_1 _1166_ (.Y(_0192_),
    .B1(net705),
    .B2(\latch_mem.RAM[42][4] ),
    .A2(net710),
    .A1(\latch_mem.RAM[44][4] ));
 sg13g2_a22oi_1 _1167_ (.Y(_0193_),
    .B1(net715),
    .B2(\latch_mem.RAM[46][4] ),
    .A2(net760),
    .A1(\latch_mem.RAM[33][4] ));
 sg13g2_a22oi_1 _1168_ (.Y(_0194_),
    .B1(net746),
    .B2(\latch_mem.RAM[35][4] ),
    .A2(net783),
    .A1(\latch_mem.RAM[32][4] ));
 sg13g2_nand4_1 _1169_ (.B(_0190_),
    .C(_0193_),
    .A(_0189_),
    .Y(_0195_),
    .D(_0194_));
 sg13g2_a22oi_1 _1170_ (.Y(_0196_),
    .B1(net739),
    .B2(\latch_mem.RAM[41][4] ),
    .A2(net750),
    .A1(\latch_mem.RAM[47][4] ));
 sg13g2_a22oi_1 _1171_ (.Y(_0197_),
    .B1(net720),
    .B2(\latch_mem.RAM[45][4] ),
    .A2(net725),
    .A1(\latch_mem.RAM[38][4] ));
 sg13g2_nand4_1 _1172_ (.B(_0192_),
    .C(_0196_),
    .A(_0191_),
    .Y(_0198_),
    .D(_0197_));
 sg13g2_or2_1 _1173_ (.X(\latch_mem.genblk2[2].selected_out[4] ),
    .B(_0198_),
    .A(_0195_));
 sg13g2_a22oi_1 _1174_ (.Y(_0199_),
    .B1(net714),
    .B2(\latch_mem.RAM[46][5] ),
    .A2(net759),
    .A1(\latch_mem.RAM[33][5] ));
 sg13g2_a22oi_1 _1175_ (.Y(_0200_),
    .B1(net734),
    .B2(\latch_mem.RAM[36][5] ),
    .A2(net739),
    .A1(\latch_mem.RAM[41][5] ));
 sg13g2_a22oi_1 _1176_ (.Y(_0201_),
    .B1(net704),
    .B2(\latch_mem.RAM[42][5] ),
    .A2(net745),
    .A1(\latch_mem.RAM[35][5] ));
 sg13g2_a22oi_1 _1177_ (.Y(_0202_),
    .B1(net720),
    .B2(\latch_mem.RAM[45][5] ),
    .A2(net754),
    .A1(\latch_mem.RAM[39][5] ));
 sg13g2_nand4_1 _1178_ (.B(_0200_),
    .C(_0201_),
    .A(_0199_),
    .Y(_0203_),
    .D(_0202_));
 sg13g2_a22oi_1 _1179_ (.Y(_0204_),
    .B1(net695),
    .B2(\latch_mem.RAM[43][5] ),
    .A2(net700),
    .A1(\latch_mem.RAM[37][5] ));
 sg13g2_a22oi_1 _1180_ (.Y(_0205_),
    .B1(net725),
    .B2(\latch_mem.RAM[38][5] ),
    .A2(net765),
    .A1(\latch_mem.RAM[34][5] ));
 sg13g2_a22oi_1 _1181_ (.Y(_0206_),
    .B1(net710),
    .B2(\latch_mem.RAM[44][5] ),
    .A2(net783),
    .A1(\latch_mem.RAM[32][5] ));
 sg13g2_a22oi_1 _1182_ (.Y(_0207_),
    .B1(net729),
    .B2(\latch_mem.RAM[40][5] ),
    .A2(net750),
    .A1(\latch_mem.RAM[47][5] ));
 sg13g2_nand4_1 _1183_ (.B(_0205_),
    .C(_0206_),
    .A(_0204_),
    .Y(_0208_),
    .D(_0207_));
 sg13g2_or2_1 _1184_ (.X(\latch_mem.genblk2[2].selected_out[5] ),
    .B(_0208_),
    .A(_0203_));
 sg13g2_a22oi_1 _1185_ (.Y(_0209_),
    .B1(net695),
    .B2(\latch_mem.RAM[43][6] ),
    .A2(net730),
    .A1(\latch_mem.RAM[40][6] ));
 sg13g2_a22oi_1 _1186_ (.Y(_0210_),
    .B1(net710),
    .B2(\latch_mem.RAM[44][6] ),
    .A2(net756),
    .A1(\latch_mem.RAM[39][6] ));
 sg13g2_a22oi_1 _1187_ (.Y(_0211_),
    .B1(net715),
    .B2(\latch_mem.RAM[46][6] ),
    .A2(net751),
    .A1(\latch_mem.RAM[47][6] ));
 sg13g2_a22oi_1 _1188_ (.Y(_0212_),
    .B1(net720),
    .B2(\latch_mem.RAM[45][6] ),
    .A2(net783),
    .A1(\latch_mem.RAM[32][6] ));
 sg13g2_a22oi_1 _1189_ (.Y(_0213_),
    .B1(net706),
    .B2(\latch_mem.RAM[42][6] ),
    .A2(net735),
    .A1(\latch_mem.RAM[36][6] ));
 sg13g2_a22oi_1 _1190_ (.Y(_0214_),
    .B1(net725),
    .B2(\latch_mem.RAM[38][6] ),
    .A2(net739),
    .A1(\latch_mem.RAM[41][6] ));
 sg13g2_nand4_1 _1191_ (.B(_0210_),
    .C(_0211_),
    .A(_0209_),
    .Y(_0215_),
    .D(_0213_));
 sg13g2_a22oi_1 _1192_ (.Y(_0216_),
    .B1(net745),
    .B2(\latch_mem.RAM[35][6] ),
    .A2(net765),
    .A1(\latch_mem.RAM[34][6] ));
 sg13g2_a22oi_1 _1193_ (.Y(_0217_),
    .B1(net700),
    .B2(\latch_mem.RAM[37][6] ),
    .A2(net760),
    .A1(\latch_mem.RAM[33][6] ));
 sg13g2_nand4_1 _1194_ (.B(_0214_),
    .C(_0216_),
    .A(_0212_),
    .Y(_0218_),
    .D(_0217_));
 sg13g2_or2_1 _1195_ (.X(\latch_mem.genblk2[2].selected_out[6] ),
    .B(_0218_),
    .A(_0215_));
 sg13g2_a22oi_1 _1196_ (.Y(_0219_),
    .B1(net706),
    .B2(\latch_mem.RAM[42][7] ),
    .A2(net735),
    .A1(\latch_mem.RAM[36][7] ));
 sg13g2_a22oi_1 _1197_ (.Y(_0220_),
    .B1(net739),
    .B2(\latch_mem.RAM[41][7] ),
    .A2(net783),
    .A1(\latch_mem.RAM[32][7] ));
 sg13g2_a22oi_1 _1198_ (.Y(_0221_),
    .B1(net724),
    .B2(\latch_mem.RAM[38][7] ),
    .A2(net754),
    .A1(\latch_mem.RAM[39][7] ));
 sg13g2_a22oi_1 _1199_ (.Y(_0222_),
    .B1(net720),
    .B2(\latch_mem.RAM[45][7] ),
    .A2(net750),
    .A1(\latch_mem.RAM[47][7] ));
 sg13g2_a22oi_1 _1200_ (.Y(_0223_),
    .B1(net700),
    .B2(\latch_mem.RAM[37][7] ),
    .A2(net744),
    .A1(\latch_mem.RAM[35][7] ));
 sg13g2_nand4_1 _1201_ (.B(_0221_),
    .C(_0222_),
    .A(_0220_),
    .Y(_0224_),
    .D(_0223_));
 sg13g2_a22oi_1 _1202_ (.Y(_0225_),
    .B1(net695),
    .B2(\latch_mem.RAM[43][7] ),
    .A2(net715),
    .A1(\latch_mem.RAM[46][7] ));
 sg13g2_a22oi_1 _1203_ (.Y(_0226_),
    .B1(net730),
    .B2(\latch_mem.RAM[40][7] ),
    .A2(net760),
    .A1(\latch_mem.RAM[33][7] ));
 sg13g2_a22oi_1 _1204_ (.Y(_0227_),
    .B1(net710),
    .B2(\latch_mem.RAM[44][7] ),
    .A2(net765),
    .A1(\latch_mem.RAM[34][7] ));
 sg13g2_nand4_1 _1205_ (.B(_0225_),
    .C(_0226_),
    .A(_0219_),
    .Y(_0228_),
    .D(_0227_));
 sg13g2_or2_1 _1206_ (.X(\latch_mem.genblk2[2].selected_out[7] ),
    .B(_0228_),
    .A(_0224_));
 sg13g2_a22oi_1 _1207_ (.Y(_0229_),
    .B1(net759),
    .B2(\latch_mem.RAM[17][0] ),
    .A2(net764),
    .A1(\latch_mem.RAM[18][0] ));
 sg13g2_a22oi_1 _1208_ (.Y(_0230_),
    .B1(net719),
    .B2(\latch_mem.RAM[29][0] ),
    .A2(net729),
    .A1(\latch_mem.RAM[24][0] ));
 sg13g2_a22oi_1 _1209_ (.Y(_0231_),
    .B1(net704),
    .B2(\latch_mem.RAM[26][0] ),
    .A2(net709),
    .A1(\latch_mem.RAM[28][0] ));
 sg13g2_a22oi_1 _1210_ (.Y(_0232_),
    .B1(net714),
    .B2(\latch_mem.RAM[30][0] ),
    .A2(net749),
    .A1(\latch_mem.RAM[31][0] ));
 sg13g2_nand4_1 _1211_ (.B(_0230_),
    .C(_0231_),
    .A(_0229_),
    .Y(_0233_),
    .D(_0232_));
 sg13g2_a22oi_1 _1212_ (.Y(_0234_),
    .B1(net724),
    .B2(\latch_mem.RAM[22][0] ),
    .A2(net754),
    .A1(\latch_mem.RAM[23][0] ));
 sg13g2_a22oi_1 _1213_ (.Y(_0235_),
    .B1(net694),
    .B2(\latch_mem.RAM[27][0] ),
    .A2(net734),
    .A1(\latch_mem.RAM[20][0] ));
 sg13g2_a22oi_1 _1214_ (.Y(_0236_),
    .B1(net699),
    .B2(\latch_mem.RAM[21][0] ),
    .A2(net744),
    .A1(\latch_mem.RAM[19][0] ));
 sg13g2_a22oi_1 _1215_ (.Y(_0237_),
    .B1(net739),
    .B2(\latch_mem.RAM[25][0] ),
    .A2(net782),
    .A1(\latch_mem.RAM[16][0] ));
 sg13g2_nand4_1 _1216_ (.B(_0235_),
    .C(_0236_),
    .A(_0234_),
    .Y(_0238_),
    .D(_0237_));
 sg13g2_or2_1 _1217_ (.X(\latch_mem.genblk2[1].selected_out[0] ),
    .B(_0238_),
    .A(_0233_));
 sg13g2_a22oi_1 _1218_ (.Y(_0239_),
    .B1(net734),
    .B2(\latch_mem.RAM[20][1] ),
    .A2(net744),
    .A1(\latch_mem.RAM[19][1] ));
 sg13g2_a22oi_1 _1219_ (.Y(_0240_),
    .B1(net719),
    .B2(\latch_mem.RAM[29][1] ),
    .A2(net764),
    .A1(\latch_mem.RAM[18][1] ));
 sg13g2_a22oi_1 _1220_ (.Y(_0241_),
    .B1(net728),
    .B2(\latch_mem.RAM[22][1] ),
    .A2(net740),
    .A1(\latch_mem.RAM[25][1] ));
 sg13g2_a22oi_1 _1221_ (.Y(_0242_),
    .B1(net694),
    .B2(\latch_mem.RAM[27][1] ),
    .A2(net782),
    .A1(\latch_mem.RAM[16][1] ));
 sg13g2_a22oi_1 _1222_ (.Y(_0243_),
    .B1(net706),
    .B2(\latch_mem.RAM[26][1] ),
    .A2(net709),
    .A1(\latch_mem.RAM[28][1] ));
 sg13g2_nand4_1 _1223_ (.B(_0241_),
    .C(_0242_),
    .A(_0240_),
    .Y(_0244_),
    .D(_0243_));
 sg13g2_a22oi_1 _1224_ (.Y(_0245_),
    .B1(net714),
    .B2(\latch_mem.RAM[30][1] ),
    .A2(net754),
    .A1(\latch_mem.RAM[23][1] ));
 sg13g2_a22oi_1 _1225_ (.Y(_0246_),
    .B1(net729),
    .B2(\latch_mem.RAM[24][1] ),
    .A2(net749),
    .A1(\latch_mem.RAM[31][1] ));
 sg13g2_a22oi_1 _1226_ (.Y(_0247_),
    .B1(net699),
    .B2(\latch_mem.RAM[21][1] ),
    .A2(net759),
    .A1(\latch_mem.RAM[17][1] ));
 sg13g2_nand4_1 _1227_ (.B(_0245_),
    .C(_0246_),
    .A(_0239_),
    .Y(_0248_),
    .D(_0247_));
 sg13g2_or2_1 _1228_ (.X(\latch_mem.genblk2[1].selected_out[1] ),
    .B(_0248_),
    .A(_0244_));
 sg13g2_a22oi_1 _1229_ (.Y(_0249_),
    .B1(net694),
    .B2(\latch_mem.RAM[27][2] ),
    .A2(net743),
    .A1(\latch_mem.RAM[25][2] ));
 sg13g2_a22oi_1 _1230_ (.Y(_0250_),
    .B1(net738),
    .B2(\latch_mem.RAM[20][2] ),
    .A2(net782),
    .A1(\latch_mem.RAM[16][2] ));
 sg13g2_a22oi_1 _1231_ (.Y(_0251_),
    .B1(net763),
    .B2(\latch_mem.RAM[17][2] ),
    .A2(net765),
    .A1(\latch_mem.RAM[18][2] ));
 sg13g2_a22oi_1 _1232_ (.Y(_0252_),
    .B1(net730),
    .B2(\latch_mem.RAM[24][2] ),
    .A2(net746),
    .A1(\latch_mem.RAM[19][2] ));
 sg13g2_nand4_1 _1233_ (.B(_0250_),
    .C(_0251_),
    .A(_0249_),
    .Y(_0253_),
    .D(_0252_));
 sg13g2_a22oi_1 _1234_ (.Y(_0254_),
    .B1(net699),
    .B2(\latch_mem.RAM[21][2] ),
    .A2(net749),
    .A1(\latch_mem.RAM[31][2] ));
 sg13g2_a22oi_1 _1235_ (.Y(_0255_),
    .B1(net709),
    .B2(\latch_mem.RAM[28][2] ),
    .A2(net754),
    .A1(\latch_mem.RAM[23][2] ));
 sg13g2_a22oi_1 _1236_ (.Y(_0256_),
    .B1(net704),
    .B2(\latch_mem.RAM[26][2] ),
    .A2(net719),
    .A1(\latch_mem.RAM[29][2] ));
 sg13g2_a22oi_1 _1237_ (.Y(_0257_),
    .B1(net714),
    .B2(\latch_mem.RAM[30][2] ),
    .A2(net724),
    .A1(\latch_mem.RAM[22][2] ));
 sg13g2_nand4_1 _1238_ (.B(_0255_),
    .C(_0256_),
    .A(_0254_),
    .Y(_0258_),
    .D(_0257_));
 sg13g2_or2_1 _1239_ (.X(\latch_mem.genblk2[1].selected_out[2] ),
    .B(_0258_),
    .A(_0253_));
 sg13g2_a22oi_1 _1240_ (.Y(_0259_),
    .B1(net714),
    .B2(\latch_mem.RAM[30][3] ),
    .A2(net759),
    .A1(\latch_mem.RAM[17][3] ));
 sg13g2_a22oi_1 _1241_ (.Y(_0260_),
    .B1(net754),
    .B2(\latch_mem.RAM[23][3] ),
    .A2(net764),
    .A1(\latch_mem.RAM[18][3] ));
 sg13g2_a22oi_1 _1242_ (.Y(_0261_),
    .B1(net719),
    .B2(\latch_mem.RAM[29][3] ),
    .A2(net734),
    .A1(\latch_mem.RAM[20][3] ));
 sg13g2_a22oi_1 _1243_ (.Y(_0262_),
    .B1(net699),
    .B2(\latch_mem.RAM[21][3] ),
    .A2(net709),
    .A1(\latch_mem.RAM[28][3] ));
 sg13g2_a22oi_1 _1244_ (.Y(_0263_),
    .B1(net724),
    .B2(\latch_mem.RAM[22][3] ),
    .A2(net739),
    .A1(\latch_mem.RAM[25][3] ));
 sg13g2_nand4_1 _1245_ (.B(_0261_),
    .C(_0262_),
    .A(_0259_),
    .Y(_0264_),
    .D(_0263_));
 sg13g2_a22oi_1 _1246_ (.Y(_0265_),
    .B1(net729),
    .B2(\latch_mem.RAM[24][3] ),
    .A2(net744),
    .A1(\latch_mem.RAM[19][3] ));
 sg13g2_a22oi_1 _1247_ (.Y(_0266_),
    .B1(net704),
    .B2(\latch_mem.RAM[26][3] ),
    .A2(net749),
    .A1(\latch_mem.RAM[31][3] ));
 sg13g2_a22oi_1 _1248_ (.Y(_0267_),
    .B1(net694),
    .B2(\latch_mem.RAM[27][3] ),
    .A2(net782),
    .A1(\latch_mem.RAM[16][3] ));
 sg13g2_nand4_1 _1249_ (.B(_0265_),
    .C(_0266_),
    .A(_0260_),
    .Y(_0268_),
    .D(_0267_));
 sg13g2_or2_1 _1250_ (.X(\latch_mem.genblk2[1].selected_out[3] ),
    .B(_0268_),
    .A(_0264_));
 sg13g2_a22oi_1 _1251_ (.Y(_0269_),
    .B1(net699),
    .B2(\latch_mem.RAM[21][4] ),
    .A2(net739),
    .A1(\latch_mem.RAM[25][4] ));
 sg13g2_a22oi_1 _1252_ (.Y(_0270_),
    .B1(net729),
    .B2(\latch_mem.RAM[24][4] ),
    .A2(net782),
    .A1(\latch_mem.RAM[16][4] ));
 sg13g2_a22oi_1 _1253_ (.Y(_0271_),
    .B1(net709),
    .B2(\latch_mem.RAM[28][4] ),
    .A2(net719),
    .A1(\latch_mem.RAM[29][4] ));
 sg13g2_a22oi_1 _1254_ (.Y(_0272_),
    .B1(net704),
    .B2(\latch_mem.RAM[26][4] ),
    .A2(net724),
    .A1(\latch_mem.RAM[22][4] ));
 sg13g2_nand4_1 _1255_ (.B(_0270_),
    .C(_0271_),
    .A(_0269_),
    .Y(_0273_),
    .D(_0272_));
 sg13g2_a22oi_1 _1256_ (.Y(_0274_),
    .B1(net734),
    .B2(\latch_mem.RAM[20][4] ),
    .A2(net754),
    .A1(\latch_mem.RAM[23][4] ));
 sg13g2_a22oi_1 _1257_ (.Y(_0275_),
    .B1(net744),
    .B2(\latch_mem.RAM[19][4] ),
    .A2(net759),
    .A1(\latch_mem.RAM[17][4] ));
 sg13g2_a22oi_1 _1258_ (.Y(_0276_),
    .B1(net714),
    .B2(\latch_mem.RAM[30][4] ),
    .A2(net749),
    .A1(\latch_mem.RAM[31][4] ));
 sg13g2_a22oi_1 _1259_ (.Y(_0277_),
    .B1(net694),
    .B2(\latch_mem.RAM[27][4] ),
    .A2(net764),
    .A1(\latch_mem.RAM[18][4] ));
 sg13g2_nand4_1 _1260_ (.B(_0275_),
    .C(_0276_),
    .A(_0274_),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_or2_1 _1261_ (.X(\latch_mem.genblk2[1].selected_out[4] ),
    .B(_0278_),
    .A(_0273_));
 sg13g2_a22oi_1 _1262_ (.Y(_0279_),
    .B1(net709),
    .B2(\latch_mem.RAM[28][5] ),
    .A2(net719),
    .A1(\latch_mem.RAM[29][5] ));
 sg13g2_a22oi_1 _1263_ (.Y(_0280_),
    .B1(net694),
    .B2(\latch_mem.RAM[27][5] ),
    .A2(net733),
    .A1(\latch_mem.RAM[24][5] ));
 sg13g2_a22oi_1 _1264_ (.Y(_0281_),
    .B1(_0747_),
    .B2(\latch_mem.RAM[30][5] ),
    .A2(net764),
    .A1(\latch_mem.RAM[18][5] ));
 sg13g2_a22oi_1 _1265_ (.Y(_0282_),
    .B1(net704),
    .B2(\latch_mem.RAM[26][5] ),
    .A2(net724),
    .A1(\latch_mem.RAM[22][5] ));
 sg13g2_a22oi_1 _1266_ (.Y(_0283_),
    .B1(net734),
    .B2(\latch_mem.RAM[20][5] ),
    .A2(net759),
    .A1(\latch_mem.RAM[17][5] ));
 sg13g2_a22oi_1 _1267_ (.Y(_0284_),
    .B1(net699),
    .B2(\latch_mem.RAM[21][5] ),
    .A2(net756),
    .A1(\latch_mem.RAM[23][5] ));
 sg13g2_nand4_1 _1268_ (.B(_0281_),
    .C(_0283_),
    .A(_0280_),
    .Y(_0285_),
    .D(_0284_));
 sg13g2_a22oi_1 _1269_ (.Y(_0286_),
    .B1(net739),
    .B2(\latch_mem.RAM[25][5] ),
    .A2(net782),
    .A1(\latch_mem.RAM[16][5] ));
 sg13g2_a22oi_1 _1270_ (.Y(_0287_),
    .B1(net744),
    .B2(\latch_mem.RAM[19][5] ),
    .A2(net749),
    .A1(\latch_mem.RAM[31][5] ));
 sg13g2_nand4_1 _1271_ (.B(_0282_),
    .C(_0286_),
    .A(_0279_),
    .Y(_0288_),
    .D(_0287_));
 sg13g2_or2_1 _1272_ (.X(\latch_mem.genblk2[1].selected_out[5] ),
    .B(_0288_),
    .A(_0285_));
 sg13g2_a22oi_1 _1273_ (.Y(_0289_),
    .B1(net719),
    .B2(\latch_mem.RAM[29][6] ),
    .A2(net782),
    .A1(\latch_mem.RAM[16][6] ));
 sg13g2_a22oi_1 _1274_ (.Y(_0290_),
    .B1(net699),
    .B2(\latch_mem.RAM[21][6] ),
    .A2(net704),
    .A1(\latch_mem.RAM[26][6] ));
 sg13g2_a22oi_1 _1275_ (.Y(_0291_),
    .B1(net744),
    .B2(\latch_mem.RAM[19][6] ),
    .A2(net754),
    .A1(\latch_mem.RAM[23][6] ));
 sg13g2_a22oi_1 _1276_ (.Y(_0292_),
    .B1(net749),
    .B2(\latch_mem.RAM[31][6] ),
    .A2(net759),
    .A1(\latch_mem.RAM[17][6] ));
 sg13g2_a22oi_1 _1277_ (.Y(_0293_),
    .B1(net724),
    .B2(\latch_mem.RAM[22][6] ),
    .A2(net729),
    .A1(\latch_mem.RAM[24][6] ));
 sg13g2_nand4_1 _1278_ (.B(_0291_),
    .C(_0292_),
    .A(_0290_),
    .Y(_0294_),
    .D(_0293_));
 sg13g2_a22oi_1 _1279_ (.Y(_0295_),
    .B1(net740),
    .B2(\latch_mem.RAM[25][6] ),
    .A2(net764),
    .A1(\latch_mem.RAM[18][6] ));
 sg13g2_a22oi_1 _1280_ (.Y(_0296_),
    .B1(net694),
    .B2(\latch_mem.RAM[27][6] ),
    .A2(net715),
    .A1(\latch_mem.RAM[30][6] ));
 sg13g2_a22oi_1 _1281_ (.Y(_0297_),
    .B1(net709),
    .B2(\latch_mem.RAM[28][6] ),
    .A2(net735),
    .A1(\latch_mem.RAM[20][6] ));
 sg13g2_nand4_1 _1282_ (.B(_0295_),
    .C(_0296_),
    .A(_0289_),
    .Y(_0298_),
    .D(_0297_));
 sg13g2_or2_1 _1283_ (.X(\latch_mem.genblk2[1].selected_out[6] ),
    .B(_0298_),
    .A(_0294_));
 sg13g2_a22oi_1 _1284_ (.Y(_0299_),
    .B1(net744),
    .B2(\latch_mem.RAM[19][7] ),
    .A2(net749),
    .A1(\latch_mem.RAM[31][7] ));
 sg13g2_a22oi_1 _1285_ (.Y(_0300_),
    .B1(net706),
    .B2(\latch_mem.RAM[26][7] ),
    .A2(net735),
    .A1(\latch_mem.RAM[20][7] ));
 sg13g2_a22oi_1 _1286_ (.Y(_0301_),
    .B1(net756),
    .B2(\latch_mem.RAM[23][7] ),
    .A2(net760),
    .A1(\latch_mem.RAM[17][7] ));
 sg13g2_a22oi_1 _1287_ (.Y(_0302_),
    .B1(net782),
    .B2(\latch_mem.RAM[16][7] ),
    .A2(net764),
    .A1(\latch_mem.RAM[18][7] ));
 sg13g2_a22oi_1 _1288_ (.Y(_0303_),
    .B1(net715),
    .B2(\latch_mem.RAM[30][7] ),
    .A2(net740),
    .A1(\latch_mem.RAM[25][7] ));
 sg13g2_nand4_1 _1289_ (.B(_0301_),
    .C(_0302_),
    .A(_0300_),
    .Y(_0304_),
    .D(_0303_));
 sg13g2_a22oi_1 _1290_ (.Y(_0305_),
    .B1(net699),
    .B2(\latch_mem.RAM[21][7] ),
    .A2(net719),
    .A1(\latch_mem.RAM[29][7] ));
 sg13g2_a22oi_1 _1291_ (.Y(_0306_),
    .B1(net694),
    .B2(\latch_mem.RAM[27][7] ),
    .A2(net729),
    .A1(\latch_mem.RAM[24][7] ));
 sg13g2_a22oi_1 _1292_ (.Y(_0307_),
    .B1(net709),
    .B2(\latch_mem.RAM[28][7] ),
    .A2(net724),
    .A1(\latch_mem.RAM[22][7] ));
 sg13g2_nand4_1 _1293_ (.B(_0305_),
    .C(_0306_),
    .A(_0299_),
    .Y(_0308_),
    .D(_0307_));
 sg13g2_or2_1 _1294_ (.X(\latch_mem.genblk2[1].selected_out[7] ),
    .B(_0308_),
    .A(_0304_));
 sg13g2_a21oi_1 _1295_ (.A1(\latch_mem.RAM[8][0] ),
    .A2(net732),
    .Y(_0309_),
    .B1(net785));
 sg13g2_a22oi_1 _1296_ (.Y(_0310_),
    .B1(net702),
    .B2(\latch_mem.RAM[5][0] ),
    .A2(net722),
    .A1(\latch_mem.RAM[13][0] ));
 sg13g2_a22oi_1 _1297_ (.Y(_0311_),
    .B1(net712),
    .B2(\latch_mem.RAM[12][0] ),
    .A2(net767),
    .A1(\latch_mem.RAM[2][0] ));
 sg13g2_nand3_1 _1298_ (.B(_0310_),
    .C(_0311_),
    .A(_0309_),
    .Y(_0312_));
 sg13g2_a221oi_1 _1299_ (.B2(\latch_mem.RAM[6][0] ),
    .C1(_0312_),
    .B1(net727),
    .A1(\latch_mem.RAM[9][0] ),
    .Y(_0313_),
    .A2(net742));
 sg13g2_a22oi_1 _1300_ (.Y(_0314_),
    .B1(net697),
    .B2(\latch_mem.RAM[11][0] ),
    .A2(net737),
    .A1(\latch_mem.RAM[4][0] ));
 sg13g2_a22oi_1 _1301_ (.Y(_0315_),
    .B1(net758),
    .B2(\latch_mem.RAM[7][0] ),
    .A2(net763),
    .A1(\latch_mem.RAM[1][0] ));
 sg13g2_a22oi_1 _1302_ (.Y(_0316_),
    .B1(net708),
    .B2(\latch_mem.RAM[10][0] ),
    .A2(net717),
    .A1(\latch_mem.RAM[14][0] ));
 sg13g2_nand3_1 _1303_ (.B(_0315_),
    .C(_0316_),
    .A(_0314_),
    .Y(_0317_));
 sg13g2_a221oi_1 _1304_ (.B2(\latch_mem.RAM[3][0] ),
    .C1(_0317_),
    .B1(net748),
    .A1(\latch_mem.RAM[15][0] ),
    .Y(_0318_),
    .A2(net753));
 sg13g2_a22oi_1 _1305_ (.Y(\latch_mem.genblk2[0].selected_out[0] ),
    .B1(_0313_),
    .B2(_0318_),
    .A2(net785),
    .A1(_0664_));
 sg13g2_a22oi_1 _1306_ (.Y(_0319_),
    .B1(net712),
    .B2(\latch_mem.RAM[12][1] ),
    .A2(net767),
    .A1(\latch_mem.RAM[2][1] ));
 sg13g2_a21oi_1 _1307_ (.A1(\latch_mem.RAM[15][1] ),
    .A2(net753),
    .Y(_0320_),
    .B1(net785));
 sg13g2_a22oi_1 _1308_ (.Y(_0321_),
    .B1(net722),
    .B2(\latch_mem.RAM[13][1] ),
    .A2(net758),
    .A1(\latch_mem.RAM[7][1] ));
 sg13g2_nand3_1 _1309_ (.B(_0320_),
    .C(_0321_),
    .A(_0319_),
    .Y(_0322_));
 sg13g2_a221oi_1 _1310_ (.B2(\latch_mem.RAM[5][1] ),
    .C1(_0322_),
    .B1(net702),
    .A1(\latch_mem.RAM[3][1] ),
    .Y(_0323_),
    .A2(net748));
 sg13g2_a22oi_1 _1311_ (.Y(_0324_),
    .B1(net708),
    .B2(\latch_mem.RAM[10][1] ),
    .A2(net717),
    .A1(\latch_mem.RAM[14][1] ));
 sg13g2_a22oi_1 _1312_ (.Y(_0325_),
    .B1(net733),
    .B2(\latch_mem.RAM[8][1] ),
    .A2(net737),
    .A1(\latch_mem.RAM[4][1] ));
 sg13g2_a22oi_1 _1313_ (.Y(_0326_),
    .B1(net727),
    .B2(\latch_mem.RAM[6][1] ),
    .A2(net762),
    .A1(\latch_mem.RAM[1][1] ));
 sg13g2_nand3_1 _1314_ (.B(_0325_),
    .C(_0326_),
    .A(_0324_),
    .Y(_0327_));
 sg13g2_a221oi_1 _1315_ (.B2(\latch_mem.RAM[11][1] ),
    .C1(_0327_),
    .B1(net697),
    .A1(\latch_mem.RAM[9][1] ),
    .Y(_0328_),
    .A2(net743));
 sg13g2_a22oi_1 _1316_ (.Y(\latch_mem.genblk2[0].selected_out[1] ),
    .B1(_0323_),
    .B2(_0328_),
    .A2(net785),
    .A1(_0665_));
 sg13g2_a21oi_1 _1317_ (.A1(\latch_mem.RAM[9][2] ),
    .A2(net741),
    .Y(_0329_),
    .B1(net784));
 sg13g2_a22oi_1 _1318_ (.Y(_0330_),
    .B1(net722),
    .B2(\latch_mem.RAM[13][2] ),
    .A2(_0738_),
    .A1(\latch_mem.RAM[15][2] ));
 sg13g2_a22oi_1 _1319_ (.Y(_0331_),
    .B1(net748),
    .B2(\latch_mem.RAM[3][2] ),
    .A2(net762),
    .A1(\latch_mem.RAM[1][2] ));
 sg13g2_a22oi_1 _1320_ (.Y(_0332_),
    .B1(net717),
    .B2(\latch_mem.RAM[14][2] ),
    .A2(net758),
    .A1(\latch_mem.RAM[7][2] ));
 sg13g2_nand3_1 _1321_ (.B(_0331_),
    .C(_0332_),
    .A(_0329_),
    .Y(_0333_));
 sg13g2_a221oi_1 _1322_ (.B2(\latch_mem.RAM[6][2] ),
    .C1(_0333_),
    .B1(net728),
    .A1(\latch_mem.RAM[2][2] ),
    .Y(_0334_),
    .A2(net767));
 sg13g2_a22oi_1 _1323_ (.Y(_0335_),
    .B1(net708),
    .B2(\latch_mem.RAM[10][2] ),
    .A2(net731),
    .A1(\latch_mem.RAM[8][2] ));
 sg13g2_a22oi_1 _1324_ (.Y(_0336_),
    .B1(net697),
    .B2(\latch_mem.RAM[11][2] ),
    .A2(net712),
    .A1(\latch_mem.RAM[12][2] ));
 sg13g2_nand3_1 _1325_ (.B(_0335_),
    .C(_0336_),
    .A(_0330_),
    .Y(_0337_));
 sg13g2_a221oi_1 _1326_ (.B2(\latch_mem.RAM[5][2] ),
    .C1(_0337_),
    .B1(net702),
    .A1(\latch_mem.RAM[4][2] ),
    .Y(_0338_),
    .A2(net738));
 sg13g2_a22oi_1 _1327_ (.Y(\latch_mem.genblk2[0].selected_out[2] ),
    .B1(_0334_),
    .B2(_0338_),
    .A2(net784),
    .A1(_0666_));
 sg13g2_a22oi_1 _1328_ (.Y(_0339_),
    .B1(net722),
    .B2(\latch_mem.RAM[13][3] ),
    .A2(net748),
    .A1(\latch_mem.RAM[3][3] ));
 sg13g2_a22oi_1 _1329_ (.Y(_0340_),
    .B1(net718),
    .B2(\latch_mem.RAM[14][3] ),
    .A2(net767),
    .A1(\latch_mem.RAM[2][3] ));
 sg13g2_a21oi_1 _1330_ (.A1(\latch_mem.RAM[9][3] ),
    .A2(net742),
    .Y(_0341_),
    .B1(net785));
 sg13g2_nand3_1 _1331_ (.B(_0340_),
    .C(_0341_),
    .A(_0339_),
    .Y(_0342_));
 sg13g2_a221oi_1 _1332_ (.B2(\latch_mem.RAM[5][3] ),
    .C1(_0342_),
    .B1(net702),
    .A1(\latch_mem.RAM[7][3] ),
    .Y(_0343_),
    .A2(net757));
 sg13g2_a22oi_1 _1333_ (.Y(_0344_),
    .B1(net712),
    .B2(\latch_mem.RAM[12][3] ),
    .A2(net752),
    .A1(\latch_mem.RAM[15][3] ));
 sg13g2_a22oi_1 _1334_ (.Y(_0345_),
    .B1(net708),
    .B2(\latch_mem.RAM[10][3] ),
    .A2(net731),
    .A1(\latch_mem.RAM[8][3] ));
 sg13g2_a22oi_1 _1335_ (.Y(_0346_),
    .B1(net697),
    .B2(\latch_mem.RAM[11][3] ),
    .A2(net761),
    .A1(\latch_mem.RAM[1][3] ));
 sg13g2_nand3_1 _1336_ (.B(_0345_),
    .C(_0346_),
    .A(_0344_),
    .Y(_0347_));
 sg13g2_a221oi_1 _1337_ (.B2(\latch_mem.RAM[6][3] ),
    .C1(_0347_),
    .B1(net726),
    .A1(\latch_mem.RAM[4][3] ),
    .Y(_0348_),
    .A2(net736));
 sg13g2_a22oi_1 _1338_ (.Y(\latch_mem.genblk2[0].selected_out[3] ),
    .B1(_0343_),
    .B2(_0348_),
    .A2(net785),
    .A1(_0667_));
 sg13g2_a22oi_1 _1339_ (.Y(_0349_),
    .B1(net712),
    .B2(\latch_mem.RAM[12][4] ),
    .A2(net731),
    .A1(\latch_mem.RAM[8][4] ));
 sg13g2_a21oi_1 _1340_ (.A1(\latch_mem.RAM[7][4] ),
    .A2(net758),
    .Y(_0350_),
    .B1(net784));
 sg13g2_a22oi_1 _1341_ (.Y(_0351_),
    .B1(net702),
    .B2(\latch_mem.RAM[5][4] ),
    .A2(net761),
    .A1(\latch_mem.RAM[1][4] ));
 sg13g2_nand3_1 _1342_ (.B(_0350_),
    .C(_0351_),
    .A(_0349_),
    .Y(_0352_));
 sg13g2_a221oi_1 _1343_ (.B2(\latch_mem.RAM[11][4] ),
    .C1(_0352_),
    .B1(net697),
    .A1(\latch_mem.RAM[4][4] ),
    .Y(_0353_),
    .A2(net736));
 sg13g2_a22oi_1 _1344_ (.Y(_0354_),
    .B1(net717),
    .B2(\latch_mem.RAM[14][4] ),
    .A2(_0739_),
    .A1(\latch_mem.RAM[3][4] ));
 sg13g2_a22oi_1 _1345_ (.Y(_0355_),
    .B1(net752),
    .B2(\latch_mem.RAM[15][4] ),
    .A2(net767),
    .A1(\latch_mem.RAM[2][4] ));
 sg13g2_a22oi_1 _1346_ (.Y(_0356_),
    .B1(net722),
    .B2(\latch_mem.RAM[13][4] ),
    .A2(net741),
    .A1(\latch_mem.RAM[9][4] ));
 sg13g2_nand3_1 _1347_ (.B(_0355_),
    .C(_0356_),
    .A(_0354_),
    .Y(_0357_));
 sg13g2_a221oi_1 _1348_ (.B2(\latch_mem.RAM[10][4] ),
    .C1(_0357_),
    .B1(net708),
    .A1(\latch_mem.RAM[6][4] ),
    .Y(_0358_),
    .A2(net726));
 sg13g2_a22oi_1 _1349_ (.Y(\latch_mem.genblk2[0].selected_out[4] ),
    .B1(_0353_),
    .B2(_0358_),
    .A2(net784),
    .A1(_0668_));
 sg13g2_a21oi_1 _1350_ (.A1(\latch_mem.RAM[3][5] ),
    .A2(net747),
    .Y(_0359_),
    .B1(net784));
 sg13g2_a22oi_1 _1351_ (.Y(_0360_),
    .B1(net697),
    .B2(\latch_mem.RAM[11][5] ),
    .A2(net717),
    .A1(\latch_mem.RAM[14][5] ));
 sg13g2_a22oi_1 _1352_ (.Y(_0361_),
    .B1(net731),
    .B2(\latch_mem.RAM[8][5] ),
    .A2(net741),
    .A1(\latch_mem.RAM[9][5] ));
 sg13g2_nand3_1 _1353_ (.B(_0360_),
    .C(_0361_),
    .A(_0359_),
    .Y(_0362_));
 sg13g2_a221oi_1 _1354_ (.B2(\latch_mem.RAM[10][5] ),
    .C1(_0362_),
    .B1(net708),
    .A1(\latch_mem.RAM[1][5] ),
    .Y(_0363_),
    .A2(net761));
 sg13g2_a22oi_1 _1355_ (.Y(_0364_),
    .B1(net727),
    .B2(\latch_mem.RAM[6][5] ),
    .A2(net753),
    .A1(\latch_mem.RAM[15][5] ));
 sg13g2_a22oi_1 _1356_ (.Y(_0365_),
    .B1(net712),
    .B2(\latch_mem.RAM[12][5] ),
    .A2(net722),
    .A1(\latch_mem.RAM[13][5] ));
 sg13g2_a22oi_1 _1357_ (.Y(_0366_),
    .B1(net757),
    .B2(\latch_mem.RAM[7][5] ),
    .A2(net767),
    .A1(\latch_mem.RAM[2][5] ));
 sg13g2_nand3_1 _1358_ (.B(_0365_),
    .C(_0366_),
    .A(_0364_),
    .Y(_0367_));
 sg13g2_a221oi_1 _1359_ (.B2(\latch_mem.RAM[5][5] ),
    .C1(_0367_),
    .B1(net702),
    .A1(\latch_mem.RAM[4][5] ),
    .Y(_0368_),
    .A2(net737));
 sg13g2_a22oi_1 _1360_ (.Y(\latch_mem.genblk2[0].selected_out[5] ),
    .B1(_0363_),
    .B2(_0368_),
    .A2(net784),
    .A1(_0669_));
 sg13g2_a22oi_1 _1361_ (.Y(_0369_),
    .B1(net708),
    .B2(\latch_mem.RAM[10][6] ),
    .A2(net758),
    .A1(\latch_mem.RAM[7][6] ));
 sg13g2_a21oi_1 _1362_ (.A1(\latch_mem.RAM[1][6] ),
    .A2(net761),
    .Y(_0370_),
    .B1(net784));
 sg13g2_a22oi_1 _1363_ (.Y(_0371_),
    .B1(net697),
    .B2(\latch_mem.RAM[11][6] ),
    .A2(net747),
    .A1(\latch_mem.RAM[3][6] ));
 sg13g2_nand3_1 _1364_ (.B(_0370_),
    .C(_0371_),
    .A(_0369_),
    .Y(_0372_));
 sg13g2_a221oi_1 _1365_ (.B2(\latch_mem.RAM[13][6] ),
    .C1(_0372_),
    .B1(net722),
    .A1(\latch_mem.RAM[6][6] ),
    .Y(_0373_),
    .A2(net726));
 sg13g2_a22oi_1 _1366_ (.Y(_0374_),
    .B1(net737),
    .B2(\latch_mem.RAM[4][6] ),
    .A2(net767),
    .A1(\latch_mem.RAM[2][6] ));
 sg13g2_a22oi_1 _1367_ (.Y(_0375_),
    .B1(net702),
    .B2(\latch_mem.RAM[5][6] ),
    .A2(net752),
    .A1(\latch_mem.RAM[15][6] ));
 sg13g2_a22oi_1 _1368_ (.Y(_0376_),
    .B1(net718),
    .B2(\latch_mem.RAM[14][6] ),
    .A2(net742),
    .A1(\latch_mem.RAM[9][6] ));
 sg13g2_nand3_1 _1369_ (.B(_0375_),
    .C(_0376_),
    .A(_0374_),
    .Y(_0377_));
 sg13g2_a221oi_1 _1370_ (.B2(\latch_mem.RAM[12][6] ),
    .C1(_0377_),
    .B1(net712),
    .A1(\latch_mem.RAM[8][6] ),
    .Y(_0378_),
    .A2(net732));
 sg13g2_a22oi_1 _1371_ (.Y(\latch_mem.genblk2[0].selected_out[6] ),
    .B1(_0373_),
    .B2(_0378_),
    .A2(net787),
    .A1(_0670_));
 sg13g2_a22oi_1 _1372_ (.Y(_0379_),
    .B1(net697),
    .B2(\latch_mem.RAM[11][7] ),
    .A2(net708),
    .A1(\latch_mem.RAM[10][7] ));
 sg13g2_a21oi_1 _1373_ (.A1(\latch_mem.RAM[12][7] ),
    .A2(net712),
    .Y(_0380_),
    .B1(net784));
 sg13g2_a22oi_1 _1374_ (.Y(_0381_),
    .B1(net736),
    .B2(\latch_mem.RAM[4][7] ),
    .A2(net766),
    .A1(\latch_mem.RAM[2][7] ));
 sg13g2_nand3_1 _1375_ (.B(_0380_),
    .C(_0381_),
    .A(_0379_),
    .Y(_0382_));
 sg13g2_a221oi_1 _1376_ (.B2(\latch_mem.RAM[14][7] ),
    .C1(_0382_),
    .B1(net716),
    .A1(\latch_mem.RAM[1][7] ),
    .Y(_0383_),
    .A2(net761));
 sg13g2_a22oi_1 _1377_ (.Y(_0384_),
    .B1(net753),
    .B2(\latch_mem.RAM[15][7] ),
    .A2(net757),
    .A1(\latch_mem.RAM[7][7] ));
 sg13g2_a22oi_1 _1378_ (.Y(_0385_),
    .B1(net722),
    .B2(\latch_mem.RAM[13][7] ),
    .A2(net727),
    .A1(\latch_mem.RAM[6][7] ));
 sg13g2_a22oi_1 _1379_ (.Y(_0386_),
    .B1(net702),
    .B2(\latch_mem.RAM[5][7] ),
    .A2(net742),
    .A1(\latch_mem.RAM[9][7] ));
 sg13g2_nand3_1 _1380_ (.B(_0385_),
    .C(_0386_),
    .A(_0384_),
    .Y(_0387_));
 sg13g2_a221oi_1 _1381_ (.B2(\latch_mem.RAM[8][7] ),
    .C1(_0387_),
    .B1(net732),
    .A1(\latch_mem.RAM[3][7] ),
    .Y(_0388_),
    .A2(net748));
 sg13g2_a22oi_1 _1382_ (.Y(\latch_mem.genblk2[0].selected_out[7] ),
    .B1(_0383_),
    .B2(_0388_),
    .A2(net785),
    .A1(_0671_));
 sg13g2_and2_1 _1383_ (.A(net897),
    .B(net4),
    .X(_0023_));
 sg13g2_nand2b_1 _1384_ (.Y(_0389_),
    .B(\latch_mem.wr_en_in ),
    .A_N(\latch_mem.wr_en_next ));
 sg13g2_mux2_1 _1385_ (.A0(net138),
    .A1(net889),
    .S(net781),
    .X(_0024_));
 sg13g2_mux2_1 _1386_ (.A0(net121),
    .A1(net880),
    .S(net780),
    .X(_0025_));
 sg13g2_mux2_1 _1387_ (.A0(net111),
    .A1(net869),
    .S(net780),
    .X(_0026_));
 sg13g2_mux2_1 _1388_ (.A0(net124),
    .A1(net859),
    .S(net780),
    .X(_0027_));
 sg13g2_mux2_1 _1389_ (.A0(net120),
    .A1(net847),
    .S(net781),
    .X(_0028_));
 sg13g2_mux2_1 _1390_ (.A0(net147),
    .A1(net837),
    .S(net781),
    .X(_0029_));
 sg13g2_mux2_1 _1391_ (.A0(net113),
    .A1(net828),
    .S(net781),
    .X(_0030_));
 sg13g2_mux2_1 _1392_ (.A0(net108),
    .A1(net818),
    .S(net781),
    .X(_0031_));
 sg13g2_nor4_2 _1393_ (.A(_0651_),
    .B(history_buffer_empty_state),
    .C(_0659_),
    .Y(_0390_),
    .D(net143));
 sg13g2_and2_1 _1394_ (.A(net896),
    .B(history_buffer_empty_state),
    .X(_0391_));
 sg13g2_nand2_1 _1395_ (.Y(_0392_),
    .A(net896),
    .B(history_buffer_empty_state));
 sg13g2_nor2b_1 _1396_ (.A(\history_buffer_index[0] ),
    .B_N(\history_buffer_index[1] ),
    .Y(_0393_));
 sg13g2_nand2b_1 _1397_ (.Y(_0394_),
    .B(_0393_),
    .A_N(_0018_));
 sg13g2_a21o_1 _1398_ (.A2(_0394_),
    .A1(_0391_),
    .B1(net144),
    .X(_0032_));
 sg13g2_a21oi_1 _1399_ (.A1(_0642_),
    .A2(\history_buffer_index[0] ),
    .Y(_0395_),
    .B1(\history_buffer_index[1] ));
 sg13g2_o21ai_1 _1400_ (.B1(_0395_),
    .Y(_0396_),
    .A1(\history_buffer[1] ),
    .A2(\history_buffer_index[0] ));
 sg13g2_and2_1 _1401_ (.A(\history_buffer_index[0] ),
    .B(net135),
    .X(_0397_));
 sg13g2_a221oi_1 _1402_ (.B2(\history_buffer[4] ),
    .C1(net140),
    .B1(_0397_),
    .A1(\history_buffer[3] ),
    .Y(_0398_),
    .A2(_0393_));
 sg13g2_nand2_1 _1403_ (.Y(_0399_),
    .A(_0396_),
    .B(_0398_));
 sg13g2_mux2_1 _1404_ (.A0(_0639_),
    .A1(_0638_),
    .S(\history_buffer_index[0] ),
    .X(_0400_));
 sg13g2_o21ai_1 _1405_ (.B1(net140),
    .Y(_0401_),
    .A1(\history_buffer_index[1] ),
    .A2(_0400_));
 sg13g2_a21oi_1 _1406_ (.A1(net161),
    .A2(_0393_),
    .Y(_0402_),
    .B1(_0401_));
 sg13g2_nor2_1 _1407_ (.A(_0392_),
    .B(net162),
    .Y(_0403_));
 sg13g2_a22oi_1 _1408_ (.Y(_0404_),
    .B1(_0399_),
    .B2(net163),
    .A2(net144),
    .A1(net154));
 sg13g2_inv_1 _1409_ (.Y(_0033_),
    .A(net164));
 sg13g2_nand2b_1 _1410_ (.Y(_0405_),
    .B(\substate[2] ),
    .A_N(\substate[0] ));
 sg13g2_and2_1 _1411_ (.A(\substate[1] ),
    .B(_0405_),
    .X(_0406_));
 sg13g2_nor2b_1 _1412_ (.A(\substate[0] ),
    .B_N(net796),
    .Y(_0407_));
 sg13g2_nor4_2 _1413_ (.A(\substate[0] ),
    .B(net806),
    .C(_0674_),
    .Y(_0408_),
    .D(_0406_));
 sg13g2_o21ai_1 _1414_ (.B1(_0012_),
    .Y(_0409_),
    .A1(uo_out[6]),
    .A2(net807));
 sg13g2_a21oi_1 _1415_ (.A1(_0673_),
    .A2(_0678_),
    .Y(_0410_),
    .B1(_0409_));
 sg13g2_nor2_1 _1416_ (.A(_0011_),
    .B(_0674_),
    .Y(_0411_));
 sg13g2_nor3_1 _1417_ (.A(net806),
    .B(net103),
    .C(_0674_),
    .Y(_0412_));
 sg13g2_a21oi_1 _1418_ (.A1(net806),
    .A2(net171),
    .Y(_0413_),
    .B1(_0412_));
 sg13g2_or3_1 _1419_ (.A(_0408_),
    .B(_0410_),
    .C(_0413_),
    .X(_0414_));
 sg13g2_o21ai_1 _1420_ (.B1(net146),
    .Y(_0415_),
    .A1(_0408_),
    .A2(_0410_));
 sg13g2_nand3_1 _1421_ (.B(_0414_),
    .C(_0415_),
    .A(net897),
    .Y(_0034_));
 sg13g2_and3_1 _1422_ (.X(_0416_),
    .A(net802),
    .B(_0686_),
    .C(_0694_));
 sg13g2_nand3_1 _1423_ (.B(_0686_),
    .C(_0694_),
    .A(net802),
    .Y(_0417_));
 sg13g2_nand3_1 _1424_ (.B(_0012_),
    .C(_0416_),
    .A(net896),
    .Y(_0418_));
 sg13g2_mux2_1 _1425_ (.A0(net109),
    .A1(prediction),
    .S(_0418_),
    .X(_0035_));
 sg13g2_o21ai_1 _1426_ (.B1(net116),
    .Y(_0419_),
    .A1(net808),
    .A2(_0677_));
 sg13g2_o21ai_1 _1427_ (.B1(_0419_),
    .Y(_0036_),
    .A1(_0677_),
    .A2(_0417_));
 sg13g2_nor4_2 _1428_ (.A(\sum[1] ),
    .B(\abs_sum[0] ),
    .C(\sum[2] ),
    .Y(_0420_),
    .D(\sum[3] ));
 sg13g2_nand3_1 _1429_ (.B(\sum[5] ),
    .C(\sum[6] ),
    .A(\sum[7] ),
    .Y(_0421_));
 sg13g2_or4_1 _1430_ (.A(_0657_),
    .B(_0016_),
    .C(_0420_),
    .D(_0421_),
    .X(_0422_));
 sg13g2_a21oi_1 _1431_ (.A1(\sum[9] ),
    .A2(_0422_),
    .Y(_0423_),
    .B1(net5));
 sg13g2_nand3_1 _1432_ (.B(_0016_),
    .C(_0420_),
    .A(_0656_),
    .Y(_0424_));
 sg13g2_nand2_1 _1433_ (.Y(_0425_),
    .A(\sum[9] ),
    .B(_0424_));
 sg13g2_a21oi_1 _1434_ (.A1(_0015_),
    .A2(_0658_),
    .Y(_0426_),
    .B1(\sum[9] ));
 sg13g2_nor4_1 _1435_ (.A(\sum[5] ),
    .B(\sum[4] ),
    .C(\sum[6] ),
    .D(_0426_),
    .Y(_0427_));
 sg13g2_a221oi_1 _1436_ (.B2(_0427_),
    .C1(_0423_),
    .B1(_0425_),
    .A1(net5),
    .Y(_0428_),
    .A2(\sum[9] ));
 sg13g2_nor2_1 _1437_ (.A(_0417_),
    .B(_0428_),
    .Y(_0429_));
 sg13g2_a21oi_2 _1438_ (.B1(_0687_),
    .Y(_0430_),
    .A2(_0694_),
    .A1(net802));
 sg13g2_nand2_1 _1439_ (.Y(_0431_),
    .A(_0696_),
    .B(_0430_));
 sg13g2_o21ai_1 _1440_ (.B1(net807),
    .Y(_0432_),
    .A1(_0695_),
    .A2(_0407_));
 sg13g2_nand3_1 _1441_ (.B(_0696_),
    .C(_0411_),
    .A(net185),
    .Y(_0433_));
 sg13g2_nand3_1 _1442_ (.B(_0432_),
    .C(_0433_),
    .A(_0431_),
    .Y(_0434_));
 sg13g2_nand2_1 _1443_ (.Y(_0435_),
    .A(\substate[0] ),
    .B(_0673_));
 sg13g2_o21ai_1 _1444_ (.B1(_0685_),
    .Y(_0436_),
    .A1(_0696_),
    .A2(_0435_));
 sg13g2_nor3_1 _1445_ (.A(_0429_),
    .B(_0434_),
    .C(_0436_),
    .Y(_0437_));
 sg13g2_nor2_1 _1446_ (.A(net122),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_a21oi_1 _1447_ (.A1(_0650_),
    .A2(_0437_),
    .Y(_0037_),
    .B1(_0438_));
 sg13g2_and3_1 _1448_ (.X(_0439_),
    .A(\latch_mem.addr_in[2] ),
    .B(\latch_mem.addr_in[1] ),
    .C(\latch_mem.addr_in[0] ));
 sg13g2_and2_1 _1449_ (.A(\latch_mem.addr_in[3] ),
    .B(_0439_),
    .X(_0440_));
 sg13g2_nor2b_1 _1450_ (.A(_0004_),
    .B_N(_0440_),
    .Y(_0441_));
 sg13g2_nor2_1 _1451_ (.A(net117),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_nor2_1 _1452_ (.A(_0681_),
    .B(net118),
    .Y(_0038_));
 sg13g2_nand2b_1 _1453_ (.Y(_0443_),
    .B(_0672_),
    .A_N(new_data_avail_posedge));
 sg13g2_nand2_1 _1454_ (.Y(_0444_),
    .A(net184),
    .B(_0443_));
 sg13g2_nor2_1 _1455_ (.A(_0434_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_nand2_1 _1456_ (.Y(_0446_),
    .A(net808),
    .B(_0445_));
 sg13g2_o21ai_1 _1457_ (.B1(net896),
    .Y(_0447_),
    .A1(net807),
    .A2(_0445_));
 sg13g2_nor2b_1 _1458_ (.A(_0447_),
    .B_N(_0446_),
    .Y(_0039_));
 sg13g2_nor2b_1 _1459_ (.A(net802),
    .B_N(_0412_),
    .Y(_0448_));
 sg13g2_o21ai_1 _1460_ (.B1(net899),
    .Y(_0449_),
    .A1(net138),
    .A2(net691));
 sg13g2_a21oi_1 _1461_ (.A1(\latch_mem.uo_out[0] ),
    .A2(net691),
    .Y(_0040_),
    .B1(_0449_));
 sg13g2_mux4_1 _1462_ (.S0(_0019_),
    .A0(\history_buffer[4] ),
    .A1(\history_buffer[0] ),
    .A2(\history_buffer[6] ),
    .A3(\history_buffer[2] ),
    .S1(net799),
    .X(_0450_));
 sg13g2_nand2_1 _1463_ (.Y(_0451_),
    .A(net797),
    .B(_0450_));
 sg13g2_nor2_1 _1464_ (.A(net797),
    .B(_0691_),
    .Y(_0452_));
 sg13g2_nand2_1 _1465_ (.Y(_0453_),
    .A(\history_buffer[5] ),
    .B(net799));
 sg13g2_nand2_1 _1466_ (.Y(_0454_),
    .A(\history_buffer[3] ),
    .B(_0654_));
 sg13g2_mux4_1 _1467_ (.S0(net799),
    .A0(\history_buffer[3] ),
    .A1(\history_buffer[5] ),
    .A2(\history_buffer[7] ),
    .A3(\history_buffer[1] ),
    .S1(_0019_),
    .X(_0455_));
 sg13g2_nand3_1 _1468_ (.B(_0692_),
    .C(_0455_),
    .A(_0653_),
    .Y(_0456_));
 sg13g2_and3_1 _1469_ (.X(_0457_),
    .A(_0696_),
    .B(_0451_),
    .C(_0456_));
 sg13g2_xnor2_1 _1470_ (.Y(_0458_),
    .A(\latch_mem.uo_out[0] ),
    .B(\latch_mem.uo_out[1] ));
 sg13g2_xnor2_1 _1471_ (.Y(_0459_),
    .A(_0645_),
    .B(_0458_));
 sg13g2_xnor2_1 _1472_ (.Y(_0460_),
    .A(_0457_),
    .B(_0459_));
 sg13g2_o21ai_1 _1473_ (.B1(net895),
    .Y(_0461_),
    .A1(net121),
    .A2(_0448_));
 sg13g2_a21oi_1 _1474_ (.A1(net691),
    .A2(_0460_),
    .Y(_0041_),
    .B1(_0461_));
 sg13g2_a22oi_1 _1475_ (.Y(_0462_),
    .B1(_0451_),
    .B2(_0456_),
    .A2(_0694_),
    .A1(net801));
 sg13g2_xnor2_1 _1476_ (.Y(_0463_),
    .A(net5),
    .B(_0462_));
 sg13g2_nand2_1 _1477_ (.Y(_0464_),
    .A(_0458_),
    .B(_0463_));
 sg13g2_nor3_2 _1478_ (.A(\latch_mem.uo_out[0] ),
    .B(\latch_mem.uo_out[1] ),
    .C(\latch_mem.uo_out[2] ),
    .Y(_0465_));
 sg13g2_o21ai_1 _1479_ (.B1(\latch_mem.uo_out[2] ),
    .Y(_0466_),
    .A1(\latch_mem.uo_out[0] ),
    .A2(\latch_mem.uo_out[1] ));
 sg13g2_nand2b_1 _1480_ (.Y(_0467_),
    .B(_0466_),
    .A_N(_0465_));
 sg13g2_nand2_1 _1481_ (.Y(_0468_),
    .A(_0695_),
    .B(_0458_));
 sg13g2_xnor2_1 _1482_ (.Y(_0469_),
    .A(_0467_),
    .B(_0468_));
 sg13g2_o21ai_1 _1483_ (.B1(net691),
    .Y(_0470_),
    .A1(_0464_),
    .A2(_0469_));
 sg13g2_a21oi_1 _1484_ (.A1(_0464_),
    .A2(_0469_),
    .Y(_0471_),
    .B1(_0470_));
 sg13g2_o21ai_1 _1485_ (.B1(net899),
    .Y(_0472_),
    .A1(net111),
    .A2(net691));
 sg13g2_nor2_1 _1486_ (.A(_0471_),
    .B(_0472_),
    .Y(_0042_));
 sg13g2_a22oi_1 _1487_ (.Y(_0473_),
    .B1(_0696_),
    .B2(_0463_),
    .A2(_0693_),
    .A1(net5));
 sg13g2_nand3_1 _1488_ (.B(\latch_mem.uo_out[1] ),
    .C(\latch_mem.uo_out[2] ),
    .A(\latch_mem.uo_out[0] ),
    .Y(_0474_));
 sg13g2_nor2_1 _1489_ (.A(_0663_),
    .B(_0474_),
    .Y(_0475_));
 sg13g2_and2_1 _1490_ (.A(_0663_),
    .B(_0474_),
    .X(_0476_));
 sg13g2_nor3_1 _1491_ (.A(_0473_),
    .B(_0475_),
    .C(_0476_),
    .Y(_0477_));
 sg13g2_and2_1 _1492_ (.A(_0663_),
    .B(_0465_),
    .X(_0478_));
 sg13g2_xnor2_1 _1493_ (.Y(_0479_),
    .A(_0663_),
    .B(_0465_));
 sg13g2_nand2_1 _1494_ (.Y(_0480_),
    .A(_0645_),
    .B(_0693_));
 sg13g2_o21ai_1 _1495_ (.B1(_0480_),
    .Y(_0481_),
    .A1(_0695_),
    .A2(_0463_));
 sg13g2_a21oi_1 _1496_ (.A1(_0479_),
    .A2(_0481_),
    .Y(_0482_),
    .B1(_0477_));
 sg13g2_o21ai_1 _1497_ (.B1(net899),
    .Y(_0483_),
    .A1(net124),
    .A2(net691));
 sg13g2_a21oi_1 _1498_ (.A1(net691),
    .A2(_0482_),
    .Y(_0043_),
    .B1(_0483_));
 sg13g2_mux2_2 _1499_ (.A0(net5),
    .A1(_0463_),
    .S(_0696_),
    .X(_0484_));
 sg13g2_mux2_1 _1500_ (.A0(_0478_),
    .A1(_0475_),
    .S(_0484_),
    .X(_0485_));
 sg13g2_xnor2_1 _1501_ (.Y(_0486_),
    .A(\latch_mem.uo_out[4] ),
    .B(_0485_));
 sg13g2_o21ai_1 _1502_ (.B1(net899),
    .Y(_0487_),
    .A1(net120),
    .A2(net690));
 sg13g2_a21oi_1 _1503_ (.A1(net690),
    .A2(_0486_),
    .Y(_0044_),
    .B1(_0487_));
 sg13g2_and2_1 _1504_ (.A(\latch_mem.uo_out[4] ),
    .B(_0475_),
    .X(_0488_));
 sg13g2_nor2b_1 _1505_ (.A(\latch_mem.uo_out[4] ),
    .B_N(_0478_),
    .Y(_0489_));
 sg13g2_mux2_1 _1506_ (.A0(_0489_),
    .A1(_0488_),
    .S(_0484_),
    .X(_0490_));
 sg13g2_xnor2_1 _1507_ (.Y(_0491_),
    .A(\latch_mem.uo_out[5] ),
    .B(_0490_));
 sg13g2_o21ai_1 _1508_ (.B1(net899),
    .Y(_0492_),
    .A1(net147),
    .A2(net690));
 sg13g2_a21oi_1 _1509_ (.A1(net690),
    .A2(_0491_),
    .Y(_0045_),
    .B1(_0492_));
 sg13g2_nand2_1 _1510_ (.Y(_0493_),
    .A(\latch_mem.uo_out[5] ),
    .B(_0488_));
 sg13g2_nand2b_1 _1511_ (.Y(_0494_),
    .B(_0489_),
    .A_N(\latch_mem.uo_out[5] ));
 sg13g2_mux2_1 _1512_ (.A0(_0494_),
    .A1(_0493_),
    .S(_0484_),
    .X(_0495_));
 sg13g2_xor2_1 _1513_ (.B(_0495_),
    .A(\latch_mem.uo_out[6] ),
    .X(_0496_));
 sg13g2_o21ai_1 _1514_ (.B1(net899),
    .Y(_0497_),
    .A1(net113),
    .A2(net690));
 sg13g2_a21oi_1 _1515_ (.A1(net690),
    .A2(_0496_),
    .Y(_0046_),
    .B1(_0497_));
 sg13g2_xor2_1 _1516_ (.B(_0484_),
    .A(\latch_mem.uo_out[6] ),
    .X(_0498_));
 sg13g2_nor2_1 _1517_ (.A(_0495_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_xnor2_1 _1518_ (.Y(_0500_),
    .A(\latch_mem.uo_out[7] ),
    .B(_0499_));
 sg13g2_o21ai_1 _1519_ (.B1(net899),
    .Y(_0501_),
    .A1(net108),
    .A2(net690));
 sg13g2_a21oi_1 _1520_ (.A1(net690),
    .A2(_0500_),
    .Y(_0047_),
    .B1(_0501_));
 sg13g2_o21ai_1 _1521_ (.B1(net897),
    .Y(_0048_),
    .A1(_0652_),
    .A2(_0441_));
 sg13g2_a21oi_1 _1522_ (.A1(_0416_),
    .A2(_0428_),
    .Y(_0502_),
    .B1(_0684_));
 sg13g2_nand2b_1 _1523_ (.Y(_0503_),
    .B(_0012_),
    .A_N(_0502_));
 sg13g2_a21oi_1 _1524_ (.A1(_0435_),
    .A2(_0443_),
    .Y(_0504_),
    .B1(net806));
 sg13g2_a21oi_1 _1525_ (.A1(\latch_mem.wr_en_in ),
    .A2(net806),
    .Y(_0505_),
    .B1(_0504_));
 sg13g2_nand3b_1 _1526_ (.B(_0503_),
    .C(_0505_),
    .Y(_0506_),
    .A_N(_0408_));
 sg13g2_nor2b_1 _1527_ (.A(net123),
    .B_N(net687),
    .Y(_0507_));
 sg13g2_nor2_1 _1528_ (.A(\latch_mem.addr_in[0] ),
    .B(net806),
    .Y(_0508_));
 sg13g2_a221oi_1 _1529_ (.B2(_0508_),
    .C1(net687),
    .B1(_0430_),
    .A1(net127),
    .Y(_0509_),
    .A2(_0675_));
 sg13g2_nor3_1 _1530_ (.A(_0651_),
    .B(_0507_),
    .C(net128),
    .Y(_0049_));
 sg13g2_a21oi_2 _1531_ (.B1(net167),
    .Y(_0510_),
    .A2(_0417_),
    .A1(net808));
 sg13g2_xnor2_1 _1532_ (.Y(_0511_),
    .A(net169),
    .B(net177));
 sg13g2_nor2_1 _1533_ (.A(_0510_),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_o21ai_1 _1534_ (.B1(net898),
    .Y(_0513_),
    .A1(net686),
    .A2(_0512_));
 sg13g2_a21oi_1 _1535_ (.A1(_0649_),
    .A2(net686),
    .Y(_0050_),
    .B1(_0513_));
 sg13g2_a21oi_1 _1536_ (.A1(net169),
    .A2(\latch_mem.addr_in[0] ),
    .Y(_0514_),
    .B1(net102));
 sg13g2_nor3_1 _1537_ (.A(_0439_),
    .B(_0510_),
    .C(net170),
    .Y(_0515_));
 sg13g2_nor2_1 _1538_ (.A(net686),
    .B(_0515_),
    .Y(_0516_));
 sg13g2_nor2b_1 _1539_ (.A(net102),
    .B_N(net686),
    .Y(_0517_));
 sg13g2_nor3_1 _1540_ (.A(_0651_),
    .B(_0516_),
    .C(_0517_),
    .Y(_0051_));
 sg13g2_nor2_1 _1541_ (.A(net101),
    .B(_0439_),
    .Y(_0518_));
 sg13g2_or3_1 _1542_ (.A(_0440_),
    .B(_0510_),
    .C(_0518_),
    .X(_0519_));
 sg13g2_a21oi_1 _1543_ (.A1(net1),
    .A2(_0510_),
    .Y(_0520_),
    .B1(net686));
 sg13g2_a221oi_1 _1544_ (.B2(_0520_),
    .C1(_0651_),
    .B1(_0519_),
    .A1(_0648_),
    .Y(_0052_),
    .A2(net687));
 sg13g2_xnor2_1 _1545_ (.Y(_0521_),
    .A(net180),
    .B(_0440_));
 sg13g2_nand2_1 _1546_ (.Y(_0522_),
    .A(net2),
    .B(_0510_));
 sg13g2_o21ai_1 _1547_ (.B1(_0522_),
    .Y(_0523_),
    .A1(_0510_),
    .A2(_0521_));
 sg13g2_o21ai_1 _1548_ (.B1(net898),
    .Y(_0524_),
    .A1(net687),
    .A2(_0523_));
 sg13g2_a21oi_1 _1549_ (.A1(_0647_),
    .A2(net686),
    .Y(_0053_),
    .B1(_0524_));
 sg13g2_a21oi_1 _1550_ (.A1(\latch_mem.addr_in[4] ),
    .A2(_0440_),
    .Y(_0525_),
    .B1(\latch_mem.addr_in[5] ));
 sg13g2_nor2_1 _1551_ (.A(_0441_),
    .B(_0525_),
    .Y(_0526_));
 sg13g2_mux2_1 _1552_ (.A0(_0526_),
    .A1(net3),
    .S(_0510_),
    .X(_0527_));
 sg13g2_o21ai_1 _1553_ (.B1(net897),
    .Y(_0528_),
    .A1(net686),
    .A2(_0527_));
 sg13g2_a21oi_1 _1554_ (.A1(_0646_),
    .A2(net686),
    .Y(_0054_),
    .B1(_0528_));
 sg13g2_o21ai_1 _1555_ (.B1(net895),
    .Y(_0529_),
    .A1(net809),
    .A2(net154));
 sg13g2_a21oi_1 _1556_ (.A1(net810),
    .A2(_0645_),
    .Y(_0055_),
    .B1(_0529_));
 sg13g2_o21ai_1 _1557_ (.B1(net895),
    .Y(_0530_),
    .A1(net809),
    .A2(\history_buffer[1] ));
 sg13g2_a21oi_1 _1558_ (.A1(net809),
    .A2(_0644_),
    .Y(_0056_),
    .B1(_0530_));
 sg13g2_o21ai_1 _1559_ (.B1(net895),
    .Y(_0531_),
    .A1(net809),
    .A2(net151));
 sg13g2_a21oi_1 _1560_ (.A1(net809),
    .A2(_0643_),
    .Y(_0057_),
    .B1(_0531_));
 sg13g2_o21ai_1 _1561_ (.B1(net895),
    .Y(_0532_),
    .A1(net810),
    .A2(net148));
 sg13g2_a21oi_1 _1562_ (.A1(net810),
    .A2(_0642_),
    .Y(_0058_),
    .B1(_0532_));
 sg13g2_o21ai_1 _1563_ (.B1(net895),
    .Y(_0533_),
    .A1(net810),
    .A2(\history_buffer[4] ));
 sg13g2_a21oi_1 _1564_ (.A1(net809),
    .A2(_0641_),
    .Y(_0059_),
    .B1(_0533_));
 sg13g2_o21ai_1 _1565_ (.B1(net895),
    .Y(_0534_),
    .A1(net809),
    .A2(net156));
 sg13g2_a21oi_1 _1566_ (.A1(net809),
    .A2(_0640_),
    .Y(_0060_),
    .B1(_0534_));
 sg13g2_o21ai_1 _1567_ (.B1(net896),
    .Y(_0535_),
    .A1(net133),
    .A2(net811));
 sg13g2_a21oi_1 _1568_ (.A1(net811),
    .A2(_0639_),
    .Y(_0061_),
    .B1(_0535_));
 sg13g2_o21ai_1 _1569_ (.B1(net896),
    .Y(_0536_),
    .A1(\history_buffer[7] ),
    .A2(net811));
 sg13g2_a21oi_1 _1570_ (.A1(_0638_),
    .A2(net811),
    .Y(_0062_),
    .B1(_0536_));
 sg13g2_nand3_1 _1571_ (.B(_0453_),
    .C(_0454_),
    .A(net800),
    .Y(_0537_));
 sg13g2_nor3_1 _1572_ (.A(\history_buffer[1] ),
    .B(_0654_),
    .C(net800),
    .Y(_0538_));
 sg13g2_nor3_1 _1573_ (.A(_0653_),
    .B(net801),
    .C(_0538_),
    .Y(_0539_));
 sg13g2_mux2_1 _1574_ (.A0(_0644_),
    .A1(_0640_),
    .S(net800),
    .X(_0540_));
 sg13g2_a22oi_1 _1575_ (.Y(_0541_),
    .B1(_0540_),
    .B2(net799),
    .A2(_0690_),
    .A1(_0642_));
 sg13g2_a22oi_1 _1576_ (.Y(_0542_),
    .B1(_0541_),
    .B2(_0452_),
    .A2(_0539_),
    .A1(_0537_));
 sg13g2_nand2b_1 _1577_ (.Y(_0543_),
    .B(\history_buffer[6] ),
    .A_N(net799));
 sg13g2_o21ai_1 _1578_ (.B1(net801),
    .Y(_0544_),
    .A1(\cnt[2] ),
    .A2(_0543_));
 sg13g2_nand4_1 _1579_ (.B(_0012_),
    .C(_0686_),
    .A(net895),
    .Y(_0545_),
    .D(_0544_));
 sg13g2_nor2_1 _1580_ (.A(_0542_),
    .B(_0545_),
    .Y(_0546_));
 sg13g2_inv_1 _1581_ (.Y(_0547_),
    .A(_0546_));
 sg13g2_nand2_1 _1582_ (.Y(_0548_),
    .A(\latch_mem.uo_out[0] ),
    .B(net689));
 sg13g2_nor2_1 _1583_ (.A(_0653_),
    .B(_0692_),
    .Y(_0549_));
 sg13g2_nand2_1 _1584_ (.Y(_0550_),
    .A(net797),
    .B(_0691_));
 sg13g2_o21ai_1 _1585_ (.B1(net150),
    .Y(_0551_),
    .A1(net688),
    .A2(net692));
 sg13g2_xor2_1 _1586_ (.B(_0551_),
    .A(_0548_),
    .X(_0063_));
 sg13g2_nand2_1 _1587_ (.Y(_0552_),
    .A(\abs_sum[0] ),
    .B(\latch_mem.uo_out[0] ));
 sg13g2_nand2_1 _1588_ (.Y(_0553_),
    .A(\sum[1] ),
    .B(\latch_mem.uo_out[1] ));
 sg13g2_xnor2_1 _1589_ (.Y(_0554_),
    .A(\sum[1] ),
    .B(\latch_mem.uo_out[1] ));
 sg13g2_xnor2_1 _1590_ (.Y(_0555_),
    .A(_0552_),
    .B(_0554_));
 sg13g2_nand2_1 _1591_ (.Y(_0556_),
    .A(net692),
    .B(_0555_));
 sg13g2_o21ai_1 _1592_ (.B1(_0556_),
    .Y(_0557_),
    .A1(\latch_mem.uo_out[1] ),
    .A2(net692));
 sg13g2_nor2_1 _1593_ (.A(net158),
    .B(net689),
    .Y(_0558_));
 sg13g2_a21oi_1 _1594_ (.A1(net689),
    .A2(_0557_),
    .Y(_0064_),
    .B1(_0558_));
 sg13g2_and2_1 _1595_ (.A(\sum[2] ),
    .B(\latch_mem.uo_out[2] ),
    .X(_0559_));
 sg13g2_xor2_1 _1596_ (.B(\latch_mem.uo_out[2] ),
    .A(\sum[2] ),
    .X(_0560_));
 sg13g2_o21ai_1 _1597_ (.B1(_0553_),
    .Y(_0561_),
    .A1(_0552_),
    .A2(_0554_));
 sg13g2_xnor2_1 _1598_ (.Y(_0562_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_nand2_1 _1599_ (.Y(_0563_),
    .A(net692),
    .B(_0562_));
 sg13g2_o21ai_1 _1600_ (.B1(_0563_),
    .Y(_0564_),
    .A1(\latch_mem.uo_out[2] ),
    .A2(net692));
 sg13g2_nor2_1 _1601_ (.A(net168),
    .B(net689),
    .Y(_0565_));
 sg13g2_a21oi_1 _1602_ (.A1(net689),
    .A2(_0564_),
    .Y(_0065_),
    .B1(_0565_));
 sg13g2_a21oi_1 _1603_ (.A1(_0560_),
    .A2(_0561_),
    .Y(_0566_),
    .B1(_0559_));
 sg13g2_nand2_1 _1604_ (.Y(_0567_),
    .A(\sum[3] ),
    .B(\latch_mem.uo_out[3] ));
 sg13g2_xnor2_1 _1605_ (.Y(_0568_),
    .A(\sum[3] ),
    .B(\latch_mem.uo_out[3] ));
 sg13g2_xnor2_1 _1606_ (.Y(_0569_),
    .A(_0566_),
    .B(_0568_));
 sg13g2_o21ai_1 _1607_ (.B1(net689),
    .Y(_0570_),
    .A1(\latch_mem.uo_out[3] ),
    .A2(net692));
 sg13g2_a21oi_1 _1608_ (.A1(net692),
    .A2(_0569_),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_a21o_1 _1609_ (.A2(net688),
    .A1(net165),
    .B1(_0571_),
    .X(_0066_));
 sg13g2_o21ai_1 _1610_ (.B1(_0567_),
    .Y(_0572_),
    .A1(_0566_),
    .A2(_0568_));
 sg13g2_and2_1 _1611_ (.A(\sum[4] ),
    .B(\latch_mem.uo_out[4] ),
    .X(_0573_));
 sg13g2_xor2_1 _1612_ (.B(\latch_mem.uo_out[4] ),
    .A(\sum[4] ),
    .X(_0574_));
 sg13g2_a21oi_1 _1613_ (.A1(\latch_mem.uo_out[4] ),
    .A2(_0549_),
    .Y(_0575_),
    .B1(_0547_));
 sg13g2_o21ai_1 _1614_ (.B1(net693),
    .Y(_0576_),
    .A1(_0572_),
    .A2(_0574_));
 sg13g2_a21o_1 _1615_ (.A2(_0574_),
    .A1(_0572_),
    .B1(_0576_),
    .X(_0577_));
 sg13g2_a22oi_1 _1616_ (.Y(_0067_),
    .B1(_0575_),
    .B2(_0577_),
    .A2(net688),
    .A1(_0657_));
 sg13g2_nand2_1 _1617_ (.Y(_0578_),
    .A(\sum[5] ),
    .B(\latch_mem.uo_out[5] ));
 sg13g2_xor2_1 _1618_ (.B(\latch_mem.uo_out[5] ),
    .A(\sum[5] ),
    .X(_0579_));
 sg13g2_a21oi_1 _1619_ (.A1(_0572_),
    .A2(_0574_),
    .Y(_0580_),
    .B1(_0573_));
 sg13g2_xor2_1 _1620_ (.B(_0580_),
    .A(_0579_),
    .X(_0581_));
 sg13g2_o21ai_1 _1621_ (.B1(net689),
    .Y(_0582_),
    .A1(\latch_mem.uo_out[5] ),
    .A2(net693));
 sg13g2_a21oi_1 _1622_ (.A1(net692),
    .A2(_0581_),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_a21o_1 _1623_ (.A2(net688),
    .A1(net174),
    .B1(_0583_),
    .X(_0068_));
 sg13g2_nand2_1 _1624_ (.Y(_0584_),
    .A(\sum[6] ),
    .B(\latch_mem.uo_out[6] ));
 sg13g2_nor2_1 _1625_ (.A(\sum[6] ),
    .B(\latch_mem.uo_out[6] ),
    .Y(_0585_));
 sg13g2_xnor2_1 _1626_ (.Y(_0586_),
    .A(\sum[6] ),
    .B(\latch_mem.uo_out[6] ));
 sg13g2_and2_1 _1627_ (.A(_0574_),
    .B(_0579_),
    .X(_0587_));
 sg13g2_o21ai_1 _1628_ (.B1(_0573_),
    .Y(_0588_),
    .A1(\sum[5] ),
    .A2(\latch_mem.uo_out[5] ));
 sg13g2_nand2_1 _1629_ (.Y(_0589_),
    .A(_0578_),
    .B(_0588_));
 sg13g2_a21oi_2 _1630_ (.B1(_0589_),
    .Y(_0590_),
    .A2(_0587_),
    .A1(_0572_));
 sg13g2_xnor2_1 _1631_ (.Y(_0591_),
    .A(_0586_),
    .B(_0590_));
 sg13g2_nor2_1 _1632_ (.A(\latch_mem.uo_out[6] ),
    .B(net693),
    .Y(_0592_));
 sg13g2_a21oi_1 _1633_ (.A1(net693),
    .A2(_0591_),
    .Y(_0593_),
    .B1(_0592_));
 sg13g2_mux2_1 _1634_ (.A0(net175),
    .A1(_0593_),
    .S(net689),
    .X(_0069_));
 sg13g2_a21oi_2 _1635_ (.B1(net688),
    .Y(_0594_),
    .A2(_0549_),
    .A1(\latch_mem.uo_out[7] ));
 sg13g2_nor2_1 _1636_ (.A(\sum[7] ),
    .B(\latch_mem.uo_out[7] ),
    .Y(_0595_));
 sg13g2_nand2_1 _1637_ (.Y(_0596_),
    .A(\sum[7] ),
    .B(\latch_mem.uo_out[7] ));
 sg13g2_nand2b_1 _1638_ (.Y(_0597_),
    .B(_0596_),
    .A_N(_0595_));
 sg13g2_o21ai_1 _1639_ (.B1(_0584_),
    .Y(_0598_),
    .A1(_0585_),
    .A2(_0590_));
 sg13g2_xnor2_1 _1640_ (.Y(_0599_),
    .A(_0597_),
    .B(_0598_));
 sg13g2_nand2_1 _1641_ (.Y(_0600_),
    .A(net693),
    .B(_0599_));
 sg13g2_a22oi_1 _1642_ (.Y(_0070_),
    .B1(_0594_),
    .B2(_0600_),
    .A2(net688),
    .A1(_0656_));
 sg13g2_nand2_1 _1643_ (.Y(_0601_),
    .A(net153),
    .B(\latch_mem.uo_out[7] ));
 sg13g2_xnor2_1 _1644_ (.Y(_0602_),
    .A(net153),
    .B(\latch_mem.uo_out[7] ));
 sg13g2_o21ai_1 _1645_ (.B1(_0596_),
    .Y(_0603_),
    .A1(_0584_),
    .A2(_0595_));
 sg13g2_or2_1 _1646_ (.X(_0604_),
    .B(_0603_),
    .A(_0589_));
 sg13g2_a21oi_1 _1647_ (.A1(_0572_),
    .A2(_0587_),
    .Y(_0605_),
    .B1(_0604_));
 sg13g2_a21o_1 _1648_ (.A2(_0596_),
    .A1(_0585_),
    .B1(_0595_),
    .X(_0606_));
 sg13g2_or3_1 _1649_ (.A(_0602_),
    .B(_0605_),
    .C(_0606_),
    .X(_0607_));
 sg13g2_o21ai_1 _1650_ (.B1(_0602_),
    .Y(_0608_),
    .A1(_0605_),
    .A2(_0606_));
 sg13g2_nand3_1 _1651_ (.B(_0607_),
    .C(_0608_),
    .A(net693),
    .Y(_0609_));
 sg13g2_a22oi_1 _1652_ (.Y(_0071_),
    .B1(_0594_),
    .B2(_0609_),
    .A2(net688),
    .A1(_0658_));
 sg13g2_xnor2_1 _1653_ (.Y(_0610_),
    .A(\sum[9] ),
    .B(\latch_mem.uo_out[7] ));
 sg13g2_nand3_1 _1654_ (.B(_0607_),
    .C(_0610_),
    .A(_0601_),
    .Y(_0611_));
 sg13g2_a21o_1 _1655_ (.A2(_0607_),
    .A1(_0601_),
    .B1(_0610_),
    .X(_0612_));
 sg13g2_nand3_1 _1656_ (.B(_0611_),
    .C(_0612_),
    .A(net693),
    .Y(_0613_));
 sg13g2_a22oi_1 _1657_ (.Y(_0072_),
    .B1(_0594_),
    .B2(_0613_),
    .A2(net688),
    .A1(_0655_));
 sg13g2_and2_1 _1658_ (.A(net99),
    .B(_0391_),
    .X(_0073_));
 sg13g2_nor2_1 _1659_ (.A(\history_buffer_index[0] ),
    .B(net135),
    .Y(_0614_));
 sg13g2_nor3_1 _1660_ (.A(_0392_),
    .B(_0397_),
    .C(net136),
    .Y(_0074_));
 sg13g2_xnor2_1 _1661_ (.Y(_0615_),
    .A(net140),
    .B(_0397_));
 sg13g2_nor2_1 _1662_ (.A(_0392_),
    .B(net141),
    .Y(_0075_));
 sg13g2_nor2_2 _1663_ (.A(net123),
    .B(net779),
    .Y(_0616_));
 sg13g2_a21oi_1 _1664_ (.A1(_0660_),
    .A2(net781),
    .Y(_0076_),
    .B1(_0616_));
 sg13g2_nor2_2 _1665_ (.A(net107),
    .B(net779),
    .Y(_0617_));
 sg13g2_a21oi_1 _1666_ (.A1(_0661_),
    .A2(net781),
    .Y(_0077_),
    .B1(_0617_));
 sg13g2_nor2_2 _1667_ (.A(net102),
    .B(net779),
    .Y(_0618_));
 sg13g2_a21oi_1 _1668_ (.A1(_0662_),
    .A2(net781),
    .Y(_0078_),
    .B1(_0618_));
 sg13g2_nand2_1 _1669_ (.Y(_0619_),
    .A(net166),
    .B(net779));
 sg13g2_o21ai_1 _1670_ (.B1(_0619_),
    .Y(_0079_),
    .A1(_0648_),
    .A2(net779));
 sg13g2_nand2_1 _1671_ (.Y(_0620_),
    .A(net181),
    .B(net780));
 sg13g2_o21ai_1 _1672_ (.B1(_0620_),
    .Y(_0080_),
    .A1(_0647_),
    .A2(net779));
 sg13g2_nand2_1 _1673_ (.Y(_0621_),
    .A(net178),
    .B(net780));
 sg13g2_o21ai_1 _1674_ (.B1(_0621_),
    .Y(_0081_),
    .A1(_0646_),
    .A2(net779));
 sg13g2_nor2_1 _1675_ (.A(_0651_),
    .B(net779),
    .Y(_0082_));
 sg13g2_and2_1 _1676_ (.A(net898),
    .B(net112),
    .X(_0083_));
 sg13g2_nor2b_1 _1677_ (.A(\substate[1] ),
    .B_N(_0407_),
    .Y(_0622_));
 sg13g2_o21ai_1 _1678_ (.B1(_0685_),
    .Y(_0623_),
    .A1(_0674_),
    .A2(_0405_));
 sg13g2_or3_2 _1679_ (.A(_0411_),
    .B(_0622_),
    .C(_0623_),
    .X(_0624_));
 sg13g2_nor3_2 _1680_ (.A(_0650_),
    .B(_0416_),
    .C(_0624_),
    .Y(_0625_));
 sg13g2_nand2_1 _1681_ (.Y(_0626_),
    .A(net176),
    .B(net798));
 sg13g2_nor2_1 _1682_ (.A(net188),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_xnor2_1 _1683_ (.Y(_0628_),
    .A(net173),
    .B(_0627_));
 sg13g2_a22oi_1 _1684_ (.Y(_0629_),
    .B1(_0625_),
    .B2(_0628_),
    .A2(_0624_),
    .A1(net801));
 sg13g2_inv_1 _1685_ (.Y(_0084_),
    .A(_0629_));
 sg13g2_xor2_1 _1686_ (.B(_0626_),
    .A(net179),
    .X(_0630_));
 sg13g2_a22oi_1 _1687_ (.Y(_0631_),
    .B1(_0625_),
    .B2(_0630_),
    .A2(_0624_),
    .A1(net800));
 sg13g2_inv_1 _1688_ (.Y(_0085_),
    .A(_0631_));
 sg13g2_xor2_1 _1689_ (.B(net798),
    .A(net176),
    .X(_0632_));
 sg13g2_a22oi_1 _1690_ (.Y(_0633_),
    .B1(_0625_),
    .B2(_0632_),
    .A2(_0624_),
    .A1(net798));
 sg13g2_inv_1 _1691_ (.Y(_0086_),
    .A(_0633_));
 sg13g2_a21oi_1 _1692_ (.A1(net807),
    .A2(_0417_),
    .Y(_0634_),
    .B1(_0651_));
 sg13g2_nor3_1 _1693_ (.A(net797),
    .B(_0624_),
    .C(_0634_),
    .Y(_0635_));
 sg13g2_a21o_1 _1694_ (.A2(_0624_),
    .A1(net797),
    .B1(_0635_),
    .X(_0087_));
 sg13g2_nand2_1 _1695_ (.Y(_0636_),
    .A(net796),
    .B(_0446_));
 sg13g2_nand3b_1 _1696_ (.B(_0445_),
    .C(_0686_),
    .Y(_0637_),
    .A_N(_0428_));
 sg13g2_a21oi_1 _1697_ (.A1(_0636_),
    .A2(_0637_),
    .Y(_0088_),
    .B1(_0651_));
 sg13g2_inv_1 _1698_ (.Y(_0638_),
    .A(net133));
 sg13g2_inv_1 _1699_ (.Y(_0639_),
    .A(net156));
 sg13g2_inv_1 _1700_ (.Y(_0640_),
    .A(net159));
 sg13g2_inv_1 _1701_ (.Y(_0641_),
    .A(net148));
 sg13g2_inv_1 _1702_ (.Y(_0642_),
    .A(net151));
 sg13g2_inv_1 _1703_ (.Y(_0643_),
    .A(\history_buffer[1] ));
 sg13g2_inv_1 _1704_ (.Y(_0644_),
    .A(net154));
 sg13g2_inv_1 _1705_ (.Y(_0645_),
    .A(net5));
 sg13g2_inv_1 _1706_ (.Y(_0646_),
    .A(net132));
 sg13g2_inv_1 _1707_ (.Y(_0647_),
    .A(net130));
 sg13g2_inv_1 _1708_ (.Y(_0648_),
    .A(net101));
 sg13g2_inv_1 _1709_ (.Y(_0649_),
    .A(net107));
 sg13g2_inv_1 _1710_ (.Y(_0650_),
    .A(net807));
 sg13g2_inv_2 _1711_ (.Y(_0651_),
    .A(net897));
 sg13g2_inv_1 _1712_ (.Y(_0652_),
    .A(net806));
 sg13g2_inv_1 _1713_ (.Y(_0653_),
    .A(net797));
 sg13g2_inv_1 _1714_ (.Y(_0654_),
    .A(net799));
 sg13g2_inv_1 _1715_ (.Y(_0655_),
    .A(net172));
 sg13g2_inv_1 _1716_ (.Y(_0656_),
    .A(net157));
 sg13g2_inv_1 _1717_ (.Y(_0657_),
    .A(net160));
 sg13g2_inv_1 _1718_ (.Y(_0658_),
    .A(net153));
 sg13g2_inv_1 _1719_ (.Y(_0659_),
    .A(net6));
 sg13g2_inv_1 _1720_ (.Y(_0660_),
    .A(net186));
 sg13g2_inv_2 _1721_ (.Y(_0661_),
    .A(net182));
 sg13g2_inv_2 _1722_ (.Y(_0662_),
    .A(net805));
 sg13g2_inv_1 _1723_ (.Y(_0663_),
    .A(\latch_mem.uo_out[3] ));
 sg13g2_inv_1 _1724_ (.Y(_0664_),
    .A(\latch_mem.RAM[0][0] ));
 sg13g2_inv_1 _1725_ (.Y(_0665_),
    .A(\latch_mem.RAM[0][1] ));
 sg13g2_inv_1 _1726_ (.Y(_0666_),
    .A(\latch_mem.RAM[0][2] ));
 sg13g2_inv_1 _1727_ (.Y(_0667_),
    .A(\latch_mem.RAM[0][3] ));
 sg13g2_inv_1 _1728_ (.Y(_0668_),
    .A(\latch_mem.RAM[0][4] ));
 sg13g2_inv_1 _1729_ (.Y(_0669_),
    .A(\latch_mem.RAM[0][5] ));
 sg13g2_inv_1 _1730_ (.Y(_0670_),
    .A(\latch_mem.RAM[0][6] ));
 sg13g2_inv_1 _1731_ (.Y(_0671_),
    .A(\latch_mem.RAM[0][7] ));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_nand2_1 _1733_ (.Y(_0004_),
    .A(net132),
    .B(net130));
 sg13g2_nor2_1 _1734_ (.A(net796),
    .B(net808),
    .Y(_0672_));
 sg13g2_and2_1 _1735_ (.A(net796),
    .B(net808),
    .X(_0673_));
 sg13g2_nand2_2 _1736_ (.Y(_0674_),
    .A(net796),
    .B(net807));
 sg13g2_nand2_1 _1737_ (.Y(_0675_),
    .A(_0652_),
    .B(_0674_));
 sg13g2_o21ai_1 _1738_ (.B1(net897),
    .Y(_0676_),
    .A1(_0672_),
    .A2(_0675_));
 sg13g2_nand2_2 _1739_ (.Y(_0677_),
    .A(net897),
    .B(_0652_));
 sg13g2_nand2_1 _1740_ (.Y(_0678_),
    .A(\substate[0] ),
    .B(net801));
 sg13g2_a21oi_1 _1741_ (.A1(\substate[3] ),
    .A2(_0673_),
    .Y(_0679_),
    .B1(_0672_));
 sg13g2_a21oi_1 _1742_ (.A1(_0678_),
    .A2(_0679_),
    .Y(_0680_),
    .B1(_0677_));
 sg13g2_nand2_1 _1743_ (.Y(_0681_),
    .A(net897),
    .B(net806));
 sg13g2_a21oi_1 _1744_ (.A1(\substate[0] ),
    .A2(_0676_),
    .Y(_0682_),
    .B1(_0680_));
 sg13g2_o21ai_1 _1745_ (.B1(_0682_),
    .Y(_0000_),
    .A1(net103),
    .A2(_0681_));
 sg13g2_nor2b_1 _1746_ (.A(new_data_avail_prev),
    .B_N(net4),
    .Y(new_data_avail_posedge));
 sg13g2_nor2_1 _1747_ (.A(_0674_),
    .B(_0677_),
    .Y(_0683_));
 sg13g2_nor2b_1 _1748_ (.A(net807),
    .B_N(net796),
    .Y(_0684_));
 sg13g2_nor2_1 _1749_ (.A(_0677_),
    .B(_0684_),
    .Y(_0685_));
 sg13g2_nor2_2 _1750_ (.A(net796),
    .B(_0650_),
    .Y(_0686_));
 sg13g2_nand2b_1 _1751_ (.Y(_0687_),
    .B(net807),
    .A_N(net796));
 sg13g2_nand2_1 _1752_ (.Y(_0688_),
    .A(_0685_),
    .B(_0687_));
 sg13g2_a22oi_1 _1753_ (.Y(_0689_),
    .B1(_0688_),
    .B2(net105),
    .A2(_0683_),
    .A1(\substate[1] ));
 sg13g2_inv_1 _1754_ (.Y(_0003_),
    .A(net106));
 sg13g2_nor2_1 _1755_ (.A(net798),
    .B(net801),
    .Y(_0690_));
 sg13g2_nor3_2 _1756_ (.A(net798),
    .B(net801),
    .C(net800),
    .Y(_0691_));
 sg13g2_or3_1 _1757_ (.A(net798),
    .B(net801),
    .C(net800),
    .X(_0692_));
 sg13g2_nor3_1 _1758_ (.A(net797),
    .B(net798),
    .C(net800),
    .Y(_0693_));
 sg13g2_or3_2 _1759_ (.A(net797),
    .B(net798),
    .C(net800),
    .X(_0694_));
 sg13g2_nor2_2 _1760_ (.A(net802),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_nand2_2 _1761_ (.Y(_0696_),
    .A(_0653_),
    .B(_0691_));
 sg13g2_nor2_1 _1762_ (.A(_0017_),
    .B(_0695_),
    .Y(_0697_));
 sg13g2_nor2b_1 _1763_ (.A(_0697_),
    .B_N(_0683_),
    .Y(_0698_));
 sg13g2_a22oi_1 _1764_ (.Y(_0699_),
    .B1(_0698_),
    .B2(\substate[0] ),
    .A2(_0688_),
    .A1(net125));
 sg13g2_inv_1 _1765_ (.Y(_0002_),
    .A(net126));
 sg13g2_a22oi_1 _1766_ (.Y(_0700_),
    .B1(_0688_),
    .B2(net114),
    .A2(_0683_),
    .A1(\substate[2] ));
 sg13g2_inv_1 _1767_ (.Y(_0001_),
    .A(net115));
 sg13g2_nand2_1 _1768_ (.Y(_0007_),
    .A(net132),
    .B(_0647_));
 sg13g2_nand2_1 _1769_ (.Y(_0006_),
    .A(_0646_),
    .B(net130));
 sg13g2_nand2_1 _1770_ (.Y(_0005_),
    .A(_0646_),
    .B(_0647_));
 sg13g2_nand4_1 _1771_ (.B(\latch_mem.addr_write[1] ),
    .C(net805),
    .A(\latch_mem.addr_write[0] ),
    .Y(_0701_),
    .D(net803));
 sg13g2_dfrbp_1 _1772_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net14),
    .D(net104),
    .Q_N(_0011_),
    .Q(\substate[0] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net15),
    .D(_0001_),
    .Q_N(_0827_),
    .Q(\substate[1] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net26),
    .D(_0002_),
    .Q_N(_0828_),
    .Q(\substate[2] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net13),
    .D(_0003_),
    .Q_N(_0826_),
    .Q(\substate[3] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net92),
    .D(_0023_),
    .Q_N(_0825_),
    .Q(new_data_avail_prev));
 sg13g2_dfrbp_1 _1777_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net91),
    .D(_0024_),
    .Q_N(_0824_),
    .Q(\latch_mem.data_to_write[0] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net90),
    .D(_0025_),
    .Q_N(_0823_),
    .Q(\latch_mem.data_to_write[1] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net89),
    .D(_0026_),
    .Q_N(_0822_),
    .Q(\latch_mem.data_to_write[2] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net88),
    .D(_0027_),
    .Q_N(_0821_),
    .Q(\latch_mem.data_to_write[3] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net87),
    .D(_0028_),
    .Q_N(_0820_),
    .Q(\latch_mem.data_to_write[4] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net86),
    .D(_0029_),
    .Q_N(_0819_),
    .Q(\latch_mem.data_to_write[5] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net85),
    .D(_0030_),
    .Q_N(_0818_),
    .Q(\latch_mem.data_to_write[6] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net84),
    .D(_0031_),
    .Q_N(_0817_),
    .Q(\latch_mem.data_to_write[7] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net70),
    .D(net145),
    .Q_N(_0829_),
    .Q(history_buffer_empty_state));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net83),
    .D(net6),
    .Q_N(_0816_),
    .Q(history_buffer_request_prev));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net82),
    .D(_0033_),
    .Q_N(_0815_),
    .Q(history_buffer_output));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net81),
    .D(_0034_),
    .Q_N(_0010_),
    .Q(\latch_mem.wr_en_in ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net79),
    .D(net110),
    .Q_N(_0814_),
    .Q(prediction));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net74),
    .D(_0036_),
    .Q_N(_0813_),
    .Q(pred_ready));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net69),
    .D(_0037_),
    .Q_N(_0812_),
    .Q(training_done));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net68),
    .D(net119),
    .Q_N(_0811_),
    .Q(mem_reset_done));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net66),
    .D(_0039_),
    .Q_N(_0810_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net64),
    .D(_0040_),
    .Q_N(_0809_),
    .Q(\latch_mem.uio_in[0] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net62),
    .D(_0041_),
    .Q_N(_0808_),
    .Q(\latch_mem.uio_in[1] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net60),
    .D(_0042_),
    .Q_N(_0807_),
    .Q(\latch_mem.uio_in[2] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net58),
    .D(_0043_),
    .Q_N(_0806_),
    .Q(\latch_mem.uio_in[3] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net56),
    .D(_0044_),
    .Q_N(_0805_),
    .Q(\latch_mem.uio_in[4] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net54),
    .D(_0045_),
    .Q_N(_0804_),
    .Q(\latch_mem.uio_in[5] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net52),
    .D(_0046_),
    .Q_N(_0803_),
    .Q(\latch_mem.uio_in[6] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net50),
    .D(_0047_),
    .Q_N(_0802_),
    .Q(\latch_mem.uio_in[7] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net48),
    .D(_0048_),
    .Q_N(_0012_),
    .Q(state_rst_memory));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net47),
    .D(_0049_),
    .Q_N(_0009_),
    .Q(\latch_mem.addr_in[0] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net45),
    .D(_0050_),
    .Q_N(_0801_),
    .Q(\latch_mem.addr_in[1] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net43),
    .D(_0051_),
    .Q_N(_0800_),
    .Q(\latch_mem.addr_in[2] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net41),
    .D(_0052_),
    .Q_N(_0799_),
    .Q(\latch_mem.addr_in[3] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net39),
    .D(_0053_),
    .Q_N(_0798_),
    .Q(\latch_mem.addr_in[4] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net37),
    .D(_0054_),
    .Q_N(_0797_),
    .Q(\latch_mem.addr_in[5] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net35),
    .D(_0055_),
    .Q_N(_0796_),
    .Q(\history_buffer[0] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net33),
    .D(net155),
    .Q_N(_0795_),
    .Q(\history_buffer[1] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net31),
    .D(net152),
    .Q_N(_0794_),
    .Q(\history_buffer[2] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net29),
    .D(_0058_),
    .Q_N(_0793_),
    .Q(\history_buffer[3] ));
 sg13g2_dfrbp_1 _1813_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net27),
    .D(net149),
    .Q_N(_0792_),
    .Q(\history_buffer[4] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net24),
    .D(_0060_),
    .Q_N(_0791_),
    .Q(\history_buffer[5] ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net22),
    .D(_0061_),
    .Q_N(_0790_),
    .Q(\history_buffer[6] ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net20),
    .D(net134),
    .Q_N(_0789_),
    .Q(\history_buffer[7] ));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net18),
    .D(_0063_),
    .Q_N(_0788_),
    .Q(\abs_sum[0] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net17),
    .D(_0064_),
    .Q_N(_0787_),
    .Q(\sum[1] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net16),
    .D(_0065_),
    .Q_N(_0013_),
    .Q(\sum[2] ));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net80),
    .D(_0066_),
    .Q_N(_0014_),
    .Q(\sum[3] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net67),
    .D(_0067_),
    .Q_N(_0786_),
    .Q(\sum[4] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net65),
    .D(_0068_),
    .Q_N(_0785_),
    .Q(\sum[5] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net63),
    .D(_0069_),
    .Q_N(_0784_),
    .Q(\sum[6] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net61),
    .D(_0070_),
    .Q_N(_0015_),
    .Q(\sum[7] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net59),
    .D(_0071_),
    .Q_N(_0016_),
    .Q(\sum[8] ));
 sg13g2_dfrbp_1 _1826_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net57),
    .D(_0072_),
    .Q_N(_0021_),
    .Q(\sum[9] ));
 sg13g2_dfrbp_1 _1827_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net55),
    .D(net100),
    .Q_N(_0020_),
    .Q(\history_buffer_index[0] ));
 sg13g2_dfrbp_1 _1828_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net53),
    .D(net137),
    .Q_N(_0783_),
    .Q(\history_buffer_index[1] ));
 sg13g2_dfrbp_1 _1829_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net71),
    .D(net142),
    .Q_N(_0018_),
    .Q(\history_buffer_index[2] ));
 sg13g2_dlhq_1 _1830_ (.D(net886),
    .GATE(\latch_mem.genblk1[17].wr_en_this_byte ),
    .Q(\latch_mem.RAM[17][0] ));
 sg13g2_dlhq_1 _1831_ (.D(net874),
    .GATE(\latch_mem.genblk1[17].wr_en_this_byte ),
    .Q(\latch_mem.RAM[17][1] ));
 sg13g2_dlhq_1 _1832_ (.D(net865),
    .GATE(\latch_mem.genblk1[17].wr_en_this_byte ),
    .Q(\latch_mem.RAM[17][2] ));
 sg13g2_dlhq_1 _1833_ (.D(net854),
    .GATE(\latch_mem.genblk1[17].wr_en_this_byte ),
    .Q(\latch_mem.RAM[17][3] ));
 sg13g2_dlhq_1 _1834_ (.D(net843),
    .GATE(\latch_mem.genblk1[17].wr_en_this_byte ),
    .Q(\latch_mem.RAM[17][4] ));
 sg13g2_dlhq_1 _1835_ (.D(net833),
    .GATE(\latch_mem.genblk1[17].wr_en_this_byte ),
    .Q(\latch_mem.RAM[17][5] ));
 sg13g2_dlhq_1 _1836_ (.D(net822),
    .GATE(\latch_mem.genblk1[17].wr_en_this_byte ),
    .Q(\latch_mem.RAM[17][6] ));
 sg13g2_dlhq_1 _1837_ (.D(net814),
    .GATE(\latch_mem.genblk1[17].wr_en_this_byte ),
    .Q(\latch_mem.RAM[17][7] ));
 sg13g2_dlhq_1 _1838_ (.D(net889),
    .GATE(\latch_mem.genblk1[52].wr_en_this_byte ),
    .Q(\latch_mem.RAM[52][0] ));
 sg13g2_dlhq_1 _1839_ (.D(net880),
    .GATE(\latch_mem.genblk1[52].wr_en_this_byte ),
    .Q(\latch_mem.RAM[52][1] ));
 sg13g2_dlhq_1 _1840_ (.D(net869),
    .GATE(\latch_mem.genblk1[52].wr_en_this_byte ),
    .Q(\latch_mem.RAM[52][2] ));
 sg13g2_dlhq_1 _1841_ (.D(net859),
    .GATE(\latch_mem.genblk1[52].wr_en_this_byte ),
    .Q(\latch_mem.RAM[52][3] ));
 sg13g2_dlhq_1 _1842_ (.D(net848),
    .GATE(\latch_mem.genblk1[52].wr_en_this_byte ),
    .Q(\latch_mem.RAM[52][4] ));
 sg13g2_dlhq_1 _1843_ (.D(net837),
    .GATE(\latch_mem.genblk1[52].wr_en_this_byte ),
    .Q(\latch_mem.RAM[52][5] ));
 sg13g2_dlhq_1 _1844_ (.D(net827),
    .GATE(\latch_mem.genblk1[52].wr_en_this_byte ),
    .Q(\latch_mem.RAM[52][6] ));
 sg13g2_dlhq_1 _1845_ (.D(net818),
    .GATE(\latch_mem.genblk1[52].wr_en_this_byte ),
    .Q(\latch_mem.RAM[52][7] ));
 sg13g2_dlhq_1 _1846_ (.D(net888),
    .GATE(\latch_mem.genblk1[35].wr_en_this_byte ),
    .Q(\latch_mem.RAM[35][0] ));
 sg13g2_dlhq_1 _1847_ (.D(net876),
    .GATE(\latch_mem.genblk1[35].wr_en_this_byte ),
    .Q(\latch_mem.RAM[35][1] ));
 sg13g2_dlhq_1 _1848_ (.D(net866),
    .GATE(\latch_mem.genblk1[35].wr_en_this_byte ),
    .Q(\latch_mem.RAM[35][2] ));
 sg13g2_dlhq_1 _1849_ (.D(net857),
    .GATE(\latch_mem.genblk1[35].wr_en_this_byte ),
    .Q(\latch_mem.RAM[35][3] ));
 sg13g2_dlhq_1 _1850_ (.D(net845),
    .GATE(\latch_mem.genblk1[35].wr_en_this_byte ),
    .Q(\latch_mem.RAM[35][4] ));
 sg13g2_dlhq_1 _1851_ (.D(net834),
    .GATE(\latch_mem.genblk1[35].wr_en_this_byte ),
    .Q(\latch_mem.RAM[35][5] ));
 sg13g2_dlhq_1 _1852_ (.D(net824),
    .GATE(\latch_mem.genblk1[35].wr_en_this_byte ),
    .Q(\latch_mem.RAM[35][6] ));
 sg13g2_dlhq_1 _1853_ (.D(net813),
    .GATE(\latch_mem.genblk1[35].wr_en_this_byte ),
    .Q(\latch_mem.RAM[35][7] ));
 sg13g2_dlhq_1 _1854_ (.D(net884),
    .GATE(\latch_mem.genblk1[28].wr_en_this_byte ),
    .Q(\latch_mem.RAM[28][0] ));
 sg13g2_dlhq_1 _1855_ (.D(net875),
    .GATE(\latch_mem.genblk1[28].wr_en_this_byte ),
    .Q(\latch_mem.RAM[28][1] ));
 sg13g2_dlhq_1 _1856_ (.D(net864),
    .GATE(\latch_mem.genblk1[28].wr_en_this_byte ),
    .Q(\latch_mem.RAM[28][2] ));
 sg13g2_dlhq_1 _1857_ (.D(net852),
    .GATE(\latch_mem.genblk1[28].wr_en_this_byte ),
    .Q(\latch_mem.RAM[28][3] ));
 sg13g2_dlhq_1 _1858_ (.D(net842),
    .GATE(\latch_mem.genblk1[28].wr_en_this_byte ),
    .Q(\latch_mem.RAM[28][4] ));
 sg13g2_dlhq_1 _1859_ (.D(net832),
    .GATE(\latch_mem.genblk1[28].wr_en_this_byte ),
    .Q(\latch_mem.RAM[28][5] ));
 sg13g2_dlhq_1 _1860_ (.D(net823),
    .GATE(\latch_mem.genblk1[28].wr_en_this_byte ),
    .Q(\latch_mem.RAM[28][6] ));
 sg13g2_dlhq_1 _1861_ (.D(net812),
    .GATE(\latch_mem.genblk1[28].wr_en_this_byte ),
    .Q(\latch_mem.RAM[28][7] ));
 sg13g2_dlhq_1 _1862_ (.D(net890),
    .GATE(\latch_mem.genblk1[53].wr_en_this_byte ),
    .Q(\latch_mem.RAM[53][0] ));
 sg13g2_dlhq_1 _1863_ (.D(net880),
    .GATE(\latch_mem.genblk1[53].wr_en_this_byte ),
    .Q(\latch_mem.RAM[53][1] ));
 sg13g2_dlhq_1 _1864_ (.D(net869),
    .GATE(\latch_mem.genblk1[53].wr_en_this_byte ),
    .Q(\latch_mem.RAM[53][2] ));
 sg13g2_dlhq_1 _1865_ (.D(net860),
    .GATE(\latch_mem.genblk1[53].wr_en_this_byte ),
    .Q(\latch_mem.RAM[53][3] ));
 sg13g2_dlhq_1 _1866_ (.D(net848),
    .GATE(\latch_mem.genblk1[53].wr_en_this_byte ),
    .Q(\latch_mem.RAM[53][4] ));
 sg13g2_dlhq_1 _1867_ (.D(net838),
    .GATE(\latch_mem.genblk1[53].wr_en_this_byte ),
    .Q(\latch_mem.RAM[53][5] ));
 sg13g2_dlhq_1 _1868_ (.D(net827),
    .GATE(\latch_mem.genblk1[53].wr_en_this_byte ),
    .Q(\latch_mem.RAM[53][6] ));
 sg13g2_dlhq_1 _1869_ (.D(net818),
    .GATE(\latch_mem.genblk1[53].wr_en_this_byte ),
    .Q(\latch_mem.RAM[53][7] ));
 sg13g2_dlhq_1 _1870_ (.D(net885),
    .GATE(\latch_mem.genblk1[16].wr_en_this_byte ),
    .Q(\latch_mem.RAM[16][0] ));
 sg13g2_dlhq_1 _1871_ (.D(net875),
    .GATE(\latch_mem.genblk1[16].wr_en_this_byte ),
    .Q(\latch_mem.RAM[16][1] ));
 sg13g2_dlhq_1 _1872_ (.D(net865),
    .GATE(\latch_mem.genblk1[16].wr_en_this_byte ),
    .Q(\latch_mem.RAM[16][2] ));
 sg13g2_dlhq_1 _1873_ (.D(net852),
    .GATE(\latch_mem.genblk1[16].wr_en_this_byte ),
    .Q(\latch_mem.RAM[16][3] ));
 sg13g2_dlhq_1 _1874_ (.D(net842),
    .GATE(\latch_mem.genblk1[16].wr_en_this_byte ),
    .Q(\latch_mem.RAM[16][4] ));
 sg13g2_dlhq_1 _1875_ (.D(net832),
    .GATE(\latch_mem.genblk1[16].wr_en_this_byte ),
    .Q(\latch_mem.RAM[16][5] ));
 sg13g2_dlhq_1 _1876_ (.D(net823),
    .GATE(\latch_mem.genblk1[16].wr_en_this_byte ),
    .Q(\latch_mem.RAM[16][6] ));
 sg13g2_dlhq_1 _1877_ (.D(net814),
    .GATE(\latch_mem.genblk1[16].wr_en_this_byte ),
    .Q(\latch_mem.RAM[16][7] ));
 sg13g2_dlhq_1 _1878_ (.D(net887),
    .GATE(\latch_mem.genblk1[41].wr_en_this_byte ),
    .Q(\latch_mem.RAM[41][0] ));
 sg13g2_dlhq_1 _1879_ (.D(net876),
    .GATE(\latch_mem.genblk1[41].wr_en_this_byte ),
    .Q(\latch_mem.RAM[41][1] ));
 sg13g2_dlhq_1 _1880_ (.D(net867),
    .GATE(\latch_mem.genblk1[41].wr_en_this_byte ),
    .Q(\latch_mem.RAM[41][2] ));
 sg13g2_dlhq_1 _1881_ (.D(net857),
    .GATE(\latch_mem.genblk1[41].wr_en_this_byte ),
    .Q(\latch_mem.RAM[41][3] ));
 sg13g2_dlhq_1 _1882_ (.D(net844),
    .GATE(\latch_mem.genblk1[41].wr_en_this_byte ),
    .Q(\latch_mem.RAM[41][4] ));
 sg13g2_dlhq_1 _1883_ (.D(net834),
    .GATE(\latch_mem.genblk1[41].wr_en_this_byte ),
    .Q(\latch_mem.RAM[41][5] ));
 sg13g2_dlhq_1 _1884_ (.D(net824),
    .GATE(\latch_mem.genblk1[41].wr_en_this_byte ),
    .Q(\latch_mem.RAM[41][6] ));
 sg13g2_dlhq_1 _1885_ (.D(net813),
    .GATE(\latch_mem.genblk1[41].wr_en_this_byte ),
    .Q(\latch_mem.RAM[41][7] ));
 sg13g2_dlhq_1 _1886_ (.D(net889),
    .GATE(\latch_mem.genblk1[54].wr_en_this_byte ),
    .Q(\latch_mem.RAM[54][0] ));
 sg13g2_dlhq_1 _1887_ (.D(net879),
    .GATE(\latch_mem.genblk1[54].wr_en_this_byte ),
    .Q(\latch_mem.RAM[54][1] ));
 sg13g2_dlhq_1 _1888_ (.D(net870),
    .GATE(\latch_mem.genblk1[54].wr_en_this_byte ),
    .Q(\latch_mem.RAM[54][2] ));
 sg13g2_dlhq_1 _1889_ (.D(net860),
    .GATE(\latch_mem.genblk1[54].wr_en_this_byte ),
    .Q(\latch_mem.RAM[54][3] ));
 sg13g2_dlhq_1 _1890_ (.D(net847),
    .GATE(\latch_mem.genblk1[54].wr_en_this_byte ),
    .Q(\latch_mem.RAM[54][4] ));
 sg13g2_dlhq_1 _1891_ (.D(net838),
    .GATE(\latch_mem.genblk1[54].wr_en_this_byte ),
    .Q(\latch_mem.RAM[54][5] ));
 sg13g2_dlhq_1 _1892_ (.D(net827),
    .GATE(\latch_mem.genblk1[54].wr_en_this_byte ),
    .Q(\latch_mem.RAM[54][6] ));
 sg13g2_dlhq_1 _1893_ (.D(net819),
    .GATE(\latch_mem.genblk1[54].wr_en_this_byte ),
    .Q(\latch_mem.RAM[54][7] ));
 sg13g2_dlhq_1 _1894_ (.D(net884),
    .GATE(\latch_mem.genblk1[24].wr_en_this_byte ),
    .Q(\latch_mem.RAM[24][0] ));
 sg13g2_dlhq_1 _1895_ (.D(net874),
    .GATE(\latch_mem.genblk1[24].wr_en_this_byte ),
    .Q(\latch_mem.RAM[24][1] ));
 sg13g2_dlhq_1 _1896_ (.D(net865),
    .GATE(\latch_mem.genblk1[24].wr_en_this_byte ),
    .Q(\latch_mem.RAM[24][2] ));
 sg13g2_dlhq_1 _1897_ (.D(net853),
    .GATE(\latch_mem.genblk1[24].wr_en_this_byte ),
    .Q(\latch_mem.RAM[24][3] ));
 sg13g2_dlhq_1 _1898_ (.D(net842),
    .GATE(\latch_mem.genblk1[24].wr_en_this_byte ),
    .Q(\latch_mem.RAM[24][4] ));
 sg13g2_dlhq_1 _1899_ (.D(net833),
    .GATE(\latch_mem.genblk1[24].wr_en_this_byte ),
    .Q(\latch_mem.RAM[24][5] ));
 sg13g2_dlhq_1 _1900_ (.D(net822),
    .GATE(\latch_mem.genblk1[24].wr_en_this_byte ),
    .Q(\latch_mem.RAM[24][6] ));
 sg13g2_dlhq_1 _1901_ (.D(net812),
    .GATE(\latch_mem.genblk1[24].wr_en_this_byte ),
    .Q(\latch_mem.RAM[24][7] ));
 sg13g2_dlhq_1 _1902_ (.D(net892),
    .GATE(\latch_mem.genblk1[15].wr_en_this_byte ),
    .Q(\latch_mem.RAM[15][0] ));
 sg13g2_dlhq_1 _1903_ (.D(net882),
    .GATE(\latch_mem.genblk1[15].wr_en_this_byte ),
    .Q(\latch_mem.RAM[15][1] ));
 sg13g2_dlhq_1 _1904_ (.D(net872),
    .GATE(\latch_mem.genblk1[15].wr_en_this_byte ),
    .Q(\latch_mem.RAM[15][2] ));
 sg13g2_dlhq_1 _1905_ (.D(net862),
    .GATE(\latch_mem.genblk1[15].wr_en_this_byte ),
    .Q(\latch_mem.RAM[15][3] ));
 sg13g2_dlhq_1 _1906_ (.D(net850),
    .GATE(\latch_mem.genblk1[15].wr_en_this_byte ),
    .Q(\latch_mem.RAM[15][4] ));
 sg13g2_dlhq_1 _1907_ (.D(net840),
    .GATE(\latch_mem.genblk1[15].wr_en_this_byte ),
    .Q(\latch_mem.RAM[15][5] ));
 sg13g2_dlhq_1 _1908_ (.D(net830),
    .GATE(\latch_mem.genblk1[15].wr_en_this_byte ),
    .Q(\latch_mem.RAM[15][6] ));
 sg13g2_dlhq_1 _1909_ (.D(net817),
    .GATE(\latch_mem.genblk1[15].wr_en_this_byte ),
    .Q(\latch_mem.RAM[15][7] ));
 sg13g2_dlhq_1 _1910_ (.D(net890),
    .GATE(\latch_mem.genblk1[55].wr_en_this_byte ),
    .Q(\latch_mem.RAM[55][0] ));
 sg13g2_dlhq_1 _1911_ (.D(net879),
    .GATE(\latch_mem.genblk1[55].wr_en_this_byte ),
    .Q(\latch_mem.RAM[55][1] ));
 sg13g2_dlhq_1 _1912_ (.D(net870),
    .GATE(\latch_mem.genblk1[55].wr_en_this_byte ),
    .Q(\latch_mem.RAM[55][2] ));
 sg13g2_dlhq_1 _1913_ (.D(net855),
    .GATE(\latch_mem.genblk1[55].wr_en_this_byte ),
    .Q(\latch_mem.RAM[55][3] ));
 sg13g2_dlhq_1 _1914_ (.D(net847),
    .GATE(\latch_mem.genblk1[55].wr_en_this_byte ),
    .Q(\latch_mem.RAM[55][4] ));
 sg13g2_dlhq_1 _1915_ (.D(net837),
    .GATE(\latch_mem.genblk1[55].wr_en_this_byte ),
    .Q(\latch_mem.RAM[55][5] ));
 sg13g2_dlhq_1 _1916_ (.D(net828),
    .GATE(\latch_mem.genblk1[55].wr_en_this_byte ),
    .Q(\latch_mem.RAM[55][6] ));
 sg13g2_dlhq_1 _1917_ (.D(net819),
    .GATE(\latch_mem.genblk1[55].wr_en_this_byte ),
    .Q(\latch_mem.RAM[55][7] ));
 sg13g2_dlhq_1 _1918_ (.D(net888),
    .GATE(\latch_mem.genblk1[33].wr_en_this_byte ),
    .Q(\latch_mem.RAM[33][0] ));
 sg13g2_dlhq_1 _1919_ (.D(net877),
    .GATE(\latch_mem.genblk1[33].wr_en_this_byte ),
    .Q(\latch_mem.RAM[33][1] ));
 sg13g2_dlhq_1 _1920_ (.D(net867),
    .GATE(\latch_mem.genblk1[33].wr_en_this_byte ),
    .Q(\latch_mem.RAM[33][2] ));
 sg13g2_dlhq_1 _1921_ (.D(net856),
    .GATE(\latch_mem.genblk1[33].wr_en_this_byte ),
    .Q(\latch_mem.RAM[33][3] ));
 sg13g2_dlhq_1 _1922_ (.D(net845),
    .GATE(\latch_mem.genblk1[33].wr_en_this_byte ),
    .Q(\latch_mem.RAM[33][4] ));
 sg13g2_dlhq_1 _1923_ (.D(net834),
    .GATE(\latch_mem.genblk1[33].wr_en_this_byte ),
    .Q(\latch_mem.RAM[33][5] ));
 sg13g2_dlhq_1 _1924_ (.D(net824),
    .GATE(\latch_mem.genblk1[33].wr_en_this_byte ),
    .Q(\latch_mem.RAM[33][6] ));
 sg13g2_dlhq_1 _1925_ (.D(net815),
    .GATE(\latch_mem.genblk1[33].wr_en_this_byte ),
    .Q(\latch_mem.RAM[33][7] ));
 sg13g2_dlhq_1 _1926_ (.D(net887),
    .GATE(\latch_mem.genblk1[42].wr_en_this_byte ),
    .Q(\latch_mem.RAM[42][0] ));
 sg13g2_dlhq_1 _1927_ (.D(net876),
    .GATE(\latch_mem.genblk1[42].wr_en_this_byte ),
    .Q(\latch_mem.RAM[42][1] ));
 sg13g2_dlhq_1 _1928_ (.D(net866),
    .GATE(\latch_mem.genblk1[42].wr_en_this_byte ),
    .Q(\latch_mem.RAM[42][2] ));
 sg13g2_dlhq_1 _1929_ (.D(net856),
    .GATE(\latch_mem.genblk1[42].wr_en_this_byte ),
    .Q(\latch_mem.RAM[42][3] ));
 sg13g2_dlhq_1 _1930_ (.D(net844),
    .GATE(\latch_mem.genblk1[42].wr_en_this_byte ),
    .Q(\latch_mem.RAM[42][4] ));
 sg13g2_dlhq_1 _1931_ (.D(net834),
    .GATE(\latch_mem.genblk1[42].wr_en_this_byte ),
    .Q(\latch_mem.RAM[42][5] ));
 sg13g2_dlhq_1 _1932_ (.D(net825),
    .GATE(\latch_mem.genblk1[42].wr_en_this_byte ),
    .Q(\latch_mem.RAM[42][6] ));
 sg13g2_dlhq_1 _1933_ (.D(net815),
    .GATE(\latch_mem.genblk1[42].wr_en_this_byte ),
    .Q(\latch_mem.RAM[42][7] ));
 sg13g2_dlhq_1 _1934_ (.D(net889),
    .GATE(\latch_mem.genblk1[56].wr_en_this_byte ),
    .Q(\latch_mem.RAM[56][0] ));
 sg13g2_dlhq_1 _1935_ (.D(net879),
    .GATE(\latch_mem.genblk1[56].wr_en_this_byte ),
    .Q(\latch_mem.RAM[56][1] ));
 sg13g2_dlhq_1 _1936_ (.D(net870),
    .GATE(\latch_mem.genblk1[56].wr_en_this_byte ),
    .Q(\latch_mem.RAM[56][2] ));
 sg13g2_dlhq_1 _1937_ (.D(net859),
    .GATE(\latch_mem.genblk1[56].wr_en_this_byte ),
    .Q(\latch_mem.RAM[56][3] ));
 sg13g2_dlhq_1 _1938_ (.D(net848),
    .GATE(\latch_mem.genblk1[56].wr_en_this_byte ),
    .Q(\latch_mem.RAM[56][4] ));
 sg13g2_dlhq_1 _1939_ (.D(net837),
    .GATE(\latch_mem.genblk1[56].wr_en_this_byte ),
    .Q(\latch_mem.RAM[56][5] ));
 sg13g2_dlhq_1 _1940_ (.D(net828),
    .GATE(\latch_mem.genblk1[56].wr_en_this_byte ),
    .Q(\latch_mem.RAM[56][6] ));
 sg13g2_dlhq_1 _1941_ (.D(net818),
    .GATE(\latch_mem.genblk1[56].wr_en_this_byte ),
    .Q(\latch_mem.RAM[56][7] ));
 sg13g2_dlhq_1 _1942_ (.D(net892),
    .GATE(\latch_mem.genblk1[14].wr_en_this_byte ),
    .Q(\latch_mem.RAM[14][0] ));
 sg13g2_dlhq_1 _1943_ (.D(net881),
    .GATE(\latch_mem.genblk1[14].wr_en_this_byte ),
    .Q(\latch_mem.RAM[14][1] ));
 sg13g2_dlhq_1 _1944_ (.D(net872),
    .GATE(\latch_mem.genblk1[14].wr_en_this_byte ),
    .Q(\latch_mem.RAM[14][2] ));
 sg13g2_dlhq_1 _1945_ (.D(net861),
    .GATE(\latch_mem.genblk1[14].wr_en_this_byte ),
    .Q(\latch_mem.RAM[14][3] ));
 sg13g2_dlhq_1 _1946_ (.D(net849),
    .GATE(\latch_mem.genblk1[14].wr_en_this_byte ),
    .Q(\latch_mem.RAM[14][4] ));
 sg13g2_dlhq_1 _1947_ (.D(net840),
    .GATE(\latch_mem.genblk1[14].wr_en_this_byte ),
    .Q(\latch_mem.RAM[14][5] ));
 sg13g2_dlhq_1 _1948_ (.D(net830),
    .GATE(\latch_mem.genblk1[14].wr_en_this_byte ),
    .Q(\latch_mem.RAM[14][6] ));
 sg13g2_dlhq_1 _1949_ (.D(net820),
    .GATE(\latch_mem.genblk1[14].wr_en_this_byte ),
    .Q(\latch_mem.RAM[14][7] ));
 sg13g2_dlhq_1 _1950_ (.D(net888),
    .GATE(\latch_mem.genblk1[36].wr_en_this_byte ),
    .Q(\latch_mem.RAM[36][0] ));
 sg13g2_dlhq_1 _1951_ (.D(net877),
    .GATE(\latch_mem.genblk1[36].wr_en_this_byte ),
    .Q(\latch_mem.RAM[36][1] ));
 sg13g2_dlhq_1 _1952_ (.D(net866),
    .GATE(\latch_mem.genblk1[36].wr_en_this_byte ),
    .Q(\latch_mem.RAM[36][2] ));
 sg13g2_dlhq_1 _1953_ (.D(net856),
    .GATE(\latch_mem.genblk1[36].wr_en_this_byte ),
    .Q(\latch_mem.RAM[36][3] ));
 sg13g2_dlhq_1 _1954_ (.D(net844),
    .GATE(\latch_mem.genblk1[36].wr_en_this_byte ),
    .Q(\latch_mem.RAM[36][4] ));
 sg13g2_dlhq_1 _1955_ (.D(net834),
    .GATE(\latch_mem.genblk1[36].wr_en_this_byte ),
    .Q(\latch_mem.RAM[36][5] ));
 sg13g2_dlhq_1 _1956_ (.D(net825),
    .GATE(\latch_mem.genblk1[36].wr_en_this_byte ),
    .Q(\latch_mem.RAM[36][6] ));
 sg13g2_dlhq_1 _1957_ (.D(net815),
    .GATE(\latch_mem.genblk1[36].wr_en_this_byte ),
    .Q(\latch_mem.RAM[36][7] ));
 sg13g2_dlhq_1 _1958_ (.D(net890),
    .GATE(\latch_mem.genblk1[57].wr_en_this_byte ),
    .Q(\latch_mem.RAM[57][0] ));
 sg13g2_dlhq_1 _1959_ (.D(net879),
    .GATE(\latch_mem.genblk1[57].wr_en_this_byte ),
    .Q(\latch_mem.RAM[57][1] ));
 sg13g2_dlhq_1 _1960_ (.D(net873),
    .GATE(\latch_mem.genblk1[57].wr_en_this_byte ),
    .Q(\latch_mem.RAM[57][2] ));
 sg13g2_dlhq_1 _1961_ (.D(net855),
    .GATE(\latch_mem.genblk1[57].wr_en_this_byte ),
    .Q(\latch_mem.RAM[57][3] ));
 sg13g2_dlhq_1 _1962_ (.D(net847),
    .GATE(\latch_mem.genblk1[57].wr_en_this_byte ),
    .Q(\latch_mem.RAM[57][4] ));
 sg13g2_dlhq_1 _1963_ (.D(net841),
    .GATE(\latch_mem.genblk1[57].wr_en_this_byte ),
    .Q(\latch_mem.RAM[57][5] ));
 sg13g2_dlhq_1 _1964_ (.D(net828),
    .GATE(\latch_mem.genblk1[57].wr_en_this_byte ),
    .Q(\latch_mem.RAM[57][6] ));
 sg13g2_dlhq_1 _1965_ (.D(net819),
    .GATE(\latch_mem.genblk1[57].wr_en_this_byte ),
    .Q(\latch_mem.RAM[57][7] ));
 sg13g2_dlhq_1 _1966_ (.D(net884),
    .GATE(\latch_mem.genblk1[23].wr_en_this_byte ),
    .Q(\latch_mem.RAM[23][0] ));
 sg13g2_dlhq_1 _1967_ (.D(net874),
    .GATE(\latch_mem.genblk1[23].wr_en_this_byte ),
    .Q(\latch_mem.RAM[23][1] ));
 sg13g2_dlhq_1 _1968_ (.D(net864),
    .GATE(\latch_mem.genblk1[23].wr_en_this_byte ),
    .Q(\latch_mem.RAM[23][2] ));
 sg13g2_dlhq_1 _1969_ (.D(net854),
    .GATE(\latch_mem.genblk1[23].wr_en_this_byte ),
    .Q(\latch_mem.RAM[23][3] ));
 sg13g2_dlhq_1 _1970_ (.D(net843),
    .GATE(\latch_mem.genblk1[23].wr_en_this_byte ),
    .Q(\latch_mem.RAM[23][4] ));
 sg13g2_dlhq_1 _1971_ (.D(net836),
    .GATE(\latch_mem.genblk1[23].wr_en_this_byte ),
    .Q(\latch_mem.RAM[23][5] ));
 sg13g2_dlhq_1 _1972_ (.D(net822),
    .GATE(\latch_mem.genblk1[23].wr_en_this_byte ),
    .Q(\latch_mem.RAM[23][6] ));
 sg13g2_dlhq_1 _1973_ (.D(net814),
    .GATE(\latch_mem.genblk1[23].wr_en_this_byte ),
    .Q(\latch_mem.RAM[23][7] ));
 sg13g2_dlhq_1 _1974_ (.D(net891),
    .GATE(\latch_mem.genblk1[13].wr_en_this_byte ),
    .Q(\latch_mem.RAM[13][0] ));
 sg13g2_dlhq_1 _1975_ (.D(net882),
    .GATE(\latch_mem.genblk1[13].wr_en_this_byte ),
    .Q(\latch_mem.RAM[13][1] ));
 sg13g2_dlhq_1 _1976_ (.D(net871),
    .GATE(\latch_mem.genblk1[13].wr_en_this_byte ),
    .Q(\latch_mem.RAM[13][2] ));
 sg13g2_dlhq_1 _1977_ (.D(net858),
    .GATE(\latch_mem.genblk1[13].wr_en_this_byte ),
    .Q(\latch_mem.RAM[13][3] ));
 sg13g2_dlhq_1 _1978_ (.D(net850),
    .GATE(\latch_mem.genblk1[13].wr_en_this_byte ),
    .Q(\latch_mem.RAM[13][4] ));
 sg13g2_dlhq_1 _1979_ (.D(net839),
    .GATE(\latch_mem.genblk1[13].wr_en_this_byte ),
    .Q(\latch_mem.RAM[13][5] ));
 sg13g2_dlhq_1 _1980_ (.D(net829),
    .GATE(\latch_mem.genblk1[13].wr_en_this_byte ),
    .Q(\latch_mem.RAM[13][6] ));
 sg13g2_dlhq_1 _1981_ (.D(net817),
    .GATE(\latch_mem.genblk1[13].wr_en_this_byte ),
    .Q(\latch_mem.RAM[13][7] ));
 sg13g2_dlhq_1 _1982_ (.D(net889),
    .GATE(\latch_mem.genblk1[58].wr_en_this_byte ),
    .Q(\latch_mem.RAM[58][0] ));
 sg13g2_dlhq_1 _1983_ (.D(net879),
    .GATE(\latch_mem.genblk1[58].wr_en_this_byte ),
    .Q(\latch_mem.RAM[58][1] ));
 sg13g2_dlhq_1 _1984_ (.D(net869),
    .GATE(\latch_mem.genblk1[58].wr_en_this_byte ),
    .Q(\latch_mem.RAM[58][2] ));
 sg13g2_dlhq_1 _1985_ (.D(net859),
    .GATE(\latch_mem.genblk1[58].wr_en_this_byte ),
    .Q(\latch_mem.RAM[58][3] ));
 sg13g2_dlhq_1 _1986_ (.D(net848),
    .GATE(\latch_mem.genblk1[58].wr_en_this_byte ),
    .Q(\latch_mem.RAM[58][4] ));
 sg13g2_dlhq_1 _1987_ (.D(net838),
    .GATE(\latch_mem.genblk1[58].wr_en_this_byte ),
    .Q(\latch_mem.RAM[58][5] ));
 sg13g2_dlhq_1 _1988_ (.D(net827),
    .GATE(\latch_mem.genblk1[58].wr_en_this_byte ),
    .Q(\latch_mem.RAM[58][6] ));
 sg13g2_dlhq_1 _1989_ (.D(net819),
    .GATE(\latch_mem.genblk1[58].wr_en_this_byte ),
    .Q(\latch_mem.RAM[58][7] ));
 sg13g2_dlhq_1 _1990_ (.D(net888),
    .GATE(\latch_mem.genblk1[43].wr_en_this_byte ),
    .Q(\latch_mem.RAM[43][0] ));
 sg13g2_dlhq_1 _1991_ (.D(net876),
    .GATE(\latch_mem.genblk1[43].wr_en_this_byte ),
    .Q(\latch_mem.RAM[43][1] ));
 sg13g2_dlhq_1 _1992_ (.D(net867),
    .GATE(\latch_mem.genblk1[43].wr_en_this_byte ),
    .Q(\latch_mem.RAM[43][2] ));
 sg13g2_dlhq_1 _1993_ (.D(net856),
    .GATE(\latch_mem.genblk1[43].wr_en_this_byte ),
    .Q(\latch_mem.RAM[43][3] ));
 sg13g2_dlhq_1 _1994_ (.D(net845),
    .GATE(\latch_mem.genblk1[43].wr_en_this_byte ),
    .Q(\latch_mem.RAM[43][4] ));
 sg13g2_dlhq_1 _1995_ (.D(net835),
    .GATE(\latch_mem.genblk1[43].wr_en_this_byte ),
    .Q(\latch_mem.RAM[43][5] ));
 sg13g2_dlhq_1 _1996_ (.D(net825),
    .GATE(\latch_mem.genblk1[43].wr_en_this_byte ),
    .Q(\latch_mem.RAM[43][6] ));
 sg13g2_dlhq_1 _1997_ (.D(net815),
    .GATE(\latch_mem.genblk1[43].wr_en_this_byte ),
    .Q(\latch_mem.RAM[43][7] ));
 sg13g2_dlhq_1 _1998_ (.D(net887),
    .GATE(\latch_mem.genblk1[32].wr_en_this_byte ),
    .Q(\latch_mem.RAM[32][0] ));
 sg13g2_dlhq_1 _1999_ (.D(net877),
    .GATE(\latch_mem.genblk1[32].wr_en_this_byte ),
    .Q(\latch_mem.RAM[32][1] ));
 sg13g2_dlhq_1 _2000_ (.D(net867),
    .GATE(\latch_mem.genblk1[32].wr_en_this_byte ),
    .Q(\latch_mem.RAM[32][2] ));
 sg13g2_dlhq_1 _2001_ (.D(net857),
    .GATE(\latch_mem.genblk1[32].wr_en_this_byte ),
    .Q(\latch_mem.RAM[32][3] ));
 sg13g2_dlhq_1 _2002_ (.D(net845),
    .GATE(\latch_mem.genblk1[32].wr_en_this_byte ),
    .Q(\latch_mem.RAM[32][4] ));
 sg13g2_dlhq_1 _2003_ (.D(net835),
    .GATE(\latch_mem.genblk1[32].wr_en_this_byte ),
    .Q(\latch_mem.RAM[32][5] ));
 sg13g2_dlhq_1 _2004_ (.D(net824),
    .GATE(\latch_mem.genblk1[32].wr_en_this_byte ),
    .Q(\latch_mem.RAM[32][6] ));
 sg13g2_dlhq_1 _2005_ (.D(net813),
    .GATE(\latch_mem.genblk1[32].wr_en_this_byte ),
    .Q(\latch_mem.RAM[32][7] ));
 sg13g2_dlhq_1 _2006_ (.D(net893),
    .GATE(\latch_mem.genblk1[59].wr_en_this_byte ),
    .Q(\latch_mem.RAM[59][0] ));
 sg13g2_dlhq_1 _2007_ (.D(net879),
    .GATE(\latch_mem.genblk1[59].wr_en_this_byte ),
    .Q(\latch_mem.RAM[59][1] ));
 sg13g2_dlhq_1 _2008_ (.D(net870),
    .GATE(\latch_mem.genblk1[59].wr_en_this_byte ),
    .Q(\latch_mem.RAM[59][2] ));
 sg13g2_dlhq_1 _2009_ (.D(net860),
    .GATE(\latch_mem.genblk1[59].wr_en_this_byte ),
    .Q(\latch_mem.RAM[59][3] ));
 sg13g2_dlhq_1 _2010_ (.D(net848),
    .GATE(\latch_mem.genblk1[59].wr_en_this_byte ),
    .Q(\latch_mem.RAM[59][4] ));
 sg13g2_dlhq_1 _2011_ (.D(net838),
    .GATE(\latch_mem.genblk1[59].wr_en_this_byte ),
    .Q(\latch_mem.RAM[59][5] ));
 sg13g2_dlhq_1 _2012_ (.D(net828),
    .GATE(\latch_mem.genblk1[59].wr_en_this_byte ),
    .Q(\latch_mem.RAM[59][6] ));
 sg13g2_dlhq_1 _2013_ (.D(net819),
    .GATE(\latch_mem.genblk1[59].wr_en_this_byte ),
    .Q(\latch_mem.RAM[59][7] ));
 sg13g2_dlhq_1 _2014_ (.D(net891),
    .GATE(\latch_mem.genblk1[12].wr_en_this_byte ),
    .Q(\latch_mem.RAM[12][0] ));
 sg13g2_dlhq_1 _2015_ (.D(net882),
    .GATE(\latch_mem.genblk1[12].wr_en_this_byte ),
    .Q(\latch_mem.RAM[12][1] ));
 sg13g2_dlhq_1 _2016_ (.D(net871),
    .GATE(\latch_mem.genblk1[12].wr_en_this_byte ),
    .Q(\latch_mem.RAM[12][2] ));
 sg13g2_dlhq_1 _2017_ (.D(net862),
    .GATE(\latch_mem.genblk1[12].wr_en_this_byte ),
    .Q(\latch_mem.RAM[12][3] ));
 sg13g2_dlhq_1 _2018_ (.D(net849),
    .GATE(\latch_mem.genblk1[12].wr_en_this_byte ),
    .Q(\latch_mem.RAM[12][4] ));
 sg13g2_dlhq_1 _2019_ (.D(net839),
    .GATE(\latch_mem.genblk1[12].wr_en_this_byte ),
    .Q(\latch_mem.RAM[12][5] ));
 sg13g2_dlhq_1 _2020_ (.D(net830),
    .GATE(\latch_mem.genblk1[12].wr_en_this_byte ),
    .Q(\latch_mem.RAM[12][6] ));
 sg13g2_dlhq_1 _2021_ (.D(net820),
    .GATE(\latch_mem.genblk1[12].wr_en_this_byte ),
    .Q(\latch_mem.RAM[12][7] ));
 sg13g2_dlhq_1 _2022_ (.D(net885),
    .GATE(\latch_mem.genblk1[27].wr_en_this_byte ),
    .Q(\latch_mem.RAM[27][0] ));
 sg13g2_dlhq_1 _2023_ (.D(net875),
    .GATE(\latch_mem.genblk1[27].wr_en_this_byte ),
    .Q(\latch_mem.RAM[27][1] ));
 sg13g2_dlhq_1 _2024_ (.D(net865),
    .GATE(\latch_mem.genblk1[27].wr_en_this_byte ),
    .Q(\latch_mem.RAM[27][2] ));
 sg13g2_dlhq_1 _2025_ (.D(net852),
    .GATE(\latch_mem.genblk1[27].wr_en_this_byte ),
    .Q(\latch_mem.RAM[27][3] ));
 sg13g2_dlhq_1 _2026_ (.D(net843),
    .GATE(\latch_mem.genblk1[27].wr_en_this_byte ),
    .Q(\latch_mem.RAM[27][4] ));
 sg13g2_dlhq_1 _2027_ (.D(net833),
    .GATE(\latch_mem.genblk1[27].wr_en_this_byte ),
    .Q(\latch_mem.RAM[27][5] ));
 sg13g2_dlhq_1 _2028_ (.D(net823),
    .GATE(\latch_mem.genblk1[27].wr_en_this_byte ),
    .Q(\latch_mem.RAM[27][6] ));
 sg13g2_dlhq_1 _2029_ (.D(net812),
    .GATE(\latch_mem.genblk1[27].wr_en_this_byte ),
    .Q(\latch_mem.RAM[27][7] ));
 sg13g2_dlhq_1 _2030_ (.D(net890),
    .GATE(\latch_mem.genblk1[60].wr_en_this_byte ),
    .Q(\latch_mem.RAM[60][0] ));
 sg13g2_dlhq_1 _2031_ (.D(net883),
    .GATE(\latch_mem.genblk1[60].wr_en_this_byte ),
    .Q(\latch_mem.RAM[60][1] ));
 sg13g2_dlhq_1 _2032_ (.D(net870),
    .GATE(\latch_mem.genblk1[60].wr_en_this_byte ),
    .Q(\latch_mem.RAM[60][2] ));
 sg13g2_dlhq_1 _2033_ (.D(net859),
    .GATE(\latch_mem.genblk1[60].wr_en_this_byte ),
    .Q(\latch_mem.RAM[60][3] ));
 sg13g2_dlhq_1 _2034_ (.D(net847),
    .GATE(\latch_mem.genblk1[60].wr_en_this_byte ),
    .Q(\latch_mem.RAM[60][4] ));
 sg13g2_dlhq_1 _2035_ (.D(net837),
    .GATE(\latch_mem.genblk1[60].wr_en_this_byte ),
    .Q(\latch_mem.RAM[60][5] ));
 sg13g2_dlhq_1 _2036_ (.D(net828),
    .GATE(\latch_mem.genblk1[60].wr_en_this_byte ),
    .Q(\latch_mem.RAM[60][6] ));
 sg13g2_dlhq_1 _2037_ (.D(net819),
    .GATE(\latch_mem.genblk1[60].wr_en_this_byte ),
    .Q(\latch_mem.RAM[60][7] ));
 sg13g2_dlhq_1 _2038_ (.D(net887),
    .GATE(\latch_mem.genblk1[44].wr_en_this_byte ),
    .Q(\latch_mem.RAM[44][0] ));
 sg13g2_dlhq_1 _2039_ (.D(net876),
    .GATE(\latch_mem.genblk1[44].wr_en_this_byte ),
    .Q(\latch_mem.RAM[44][1] ));
 sg13g2_dlhq_1 _2040_ (.D(net866),
    .GATE(\latch_mem.genblk1[44].wr_en_this_byte ),
    .Q(\latch_mem.RAM[44][2] ));
 sg13g2_dlhq_1 _2041_ (.D(net856),
    .GATE(\latch_mem.genblk1[44].wr_en_this_byte ),
    .Q(\latch_mem.RAM[44][3] ));
 sg13g2_dlhq_1 _2042_ (.D(net844),
    .GATE(\latch_mem.genblk1[44].wr_en_this_byte ),
    .Q(\latch_mem.RAM[44][4] ));
 sg13g2_dlhq_1 _2043_ (.D(net835),
    .GATE(\latch_mem.genblk1[44].wr_en_this_byte ),
    .Q(\latch_mem.RAM[44][5] ));
 sg13g2_dlhq_1 _2044_ (.D(net825),
    .GATE(\latch_mem.genblk1[44].wr_en_this_byte ),
    .Q(\latch_mem.RAM[44][6] ));
 sg13g2_dlhq_1 _2045_ (.D(net815),
    .GATE(\latch_mem.genblk1[44].wr_en_this_byte ),
    .Q(\latch_mem.RAM[44][7] ));
 sg13g2_dlhq_1 _2046_ (.D(net892),
    .GATE(\latch_mem.genblk1[11].wr_en_this_byte ),
    .Q(\latch_mem.RAM[11][0] ));
 sg13g2_dlhq_1 _2047_ (.D(net881),
    .GATE(\latch_mem.genblk1[11].wr_en_this_byte ),
    .Q(\latch_mem.RAM[11][1] ));
 sg13g2_dlhq_1 _2048_ (.D(net872),
    .GATE(\latch_mem.genblk1[11].wr_en_this_byte ),
    .Q(\latch_mem.RAM[11][2] ));
 sg13g2_dlhq_1 _2049_ (.D(net862),
    .GATE(\latch_mem.genblk1[11].wr_en_this_byte ),
    .Q(\latch_mem.RAM[11][3] ));
 sg13g2_dlhq_1 _2050_ (.D(net851),
    .GATE(\latch_mem.genblk1[11].wr_en_this_byte ),
    .Q(\latch_mem.RAM[11][4] ));
 sg13g2_dlhq_1 _2051_ (.D(net841),
    .GATE(\latch_mem.genblk1[11].wr_en_this_byte ),
    .Q(\latch_mem.RAM[11][5] ));
 sg13g2_dlhq_1 _2052_ (.D(net829),
    .GATE(\latch_mem.genblk1[11].wr_en_this_byte ),
    .Q(\latch_mem.RAM[11][6] ));
 sg13g2_dlhq_1 _2053_ (.D(net820),
    .GATE(\latch_mem.genblk1[11].wr_en_this_byte ),
    .Q(\latch_mem.RAM[11][7] ));
 sg13g2_dlhq_1 _2054_ (.D(net889),
    .GATE(\latch_mem.genblk1[61].wr_en_this_byte ),
    .Q(\latch_mem.RAM[61][0] ));
 sg13g2_dlhq_1 _2055_ (.D(net881),
    .GATE(\latch_mem.genblk1[61].wr_en_this_byte ),
    .Q(\latch_mem.RAM[61][1] ));
 sg13g2_dlhq_1 _2056_ (.D(net869),
    .GATE(\latch_mem.genblk1[61].wr_en_this_byte ),
    .Q(\latch_mem.RAM[61][2] ));
 sg13g2_dlhq_1 _2057_ (.D(net859),
    .GATE(\latch_mem.genblk1[61].wr_en_this_byte ),
    .Q(\latch_mem.RAM[61][3] ));
 sg13g2_dlhq_1 _2058_ (.D(net851),
    .GATE(\latch_mem.genblk1[61].wr_en_this_byte ),
    .Q(\latch_mem.RAM[61][4] ));
 sg13g2_dlhq_1 _2059_ (.D(net838),
    .GATE(\latch_mem.genblk1[61].wr_en_this_byte ),
    .Q(\latch_mem.RAM[61][5] ));
 sg13g2_dlhq_1 _2060_ (.D(net827),
    .GATE(\latch_mem.genblk1[61].wr_en_this_byte ),
    .Q(\latch_mem.RAM[61][6] ));
 sg13g2_dlhq_1 _2061_ (.D(net821),
    .GATE(\latch_mem.genblk1[61].wr_en_this_byte ),
    .Q(\latch_mem.RAM[61][7] ));
 sg13g2_dlhq_1 _2062_ (.D(net884),
    .GATE(\latch_mem.genblk1[22].wr_en_this_byte ),
    .Q(\latch_mem.RAM[22][0] ));
 sg13g2_dlhq_1 _2063_ (.D(net875),
    .GATE(\latch_mem.genblk1[22].wr_en_this_byte ),
    .Q(\latch_mem.RAM[22][1] ));
 sg13g2_dlhq_1 _2064_ (.D(net864),
    .GATE(\latch_mem.genblk1[22].wr_en_this_byte ),
    .Q(\latch_mem.RAM[22][2] ));
 sg13g2_dlhq_1 _2065_ (.D(net852),
    .GATE(\latch_mem.genblk1[22].wr_en_this_byte ),
    .Q(\latch_mem.RAM[22][3] ));
 sg13g2_dlhq_1 _2066_ (.D(net842),
    .GATE(\latch_mem.genblk1[22].wr_en_this_byte ),
    .Q(\latch_mem.RAM[22][4] ));
 sg13g2_dlhq_1 _2067_ (.D(net832),
    .GATE(\latch_mem.genblk1[22].wr_en_this_byte ),
    .Q(\latch_mem.RAM[22][5] ));
 sg13g2_dlhq_1 _2068_ (.D(net822),
    .GATE(\latch_mem.genblk1[22].wr_en_this_byte ),
    .Q(\latch_mem.RAM[22][6] ));
 sg13g2_dlhq_1 _2069_ (.D(net812),
    .GATE(\latch_mem.genblk1[22].wr_en_this_byte ),
    .Q(\latch_mem.RAM[22][7] ));
 sg13g2_dlhq_1 _2070_ (.D(net887),
    .GATE(\latch_mem.genblk1[37].wr_en_this_byte ),
    .Q(\latch_mem.RAM[37][0] ));
 sg13g2_dlhq_1 _2071_ (.D(net877),
    .GATE(\latch_mem.genblk1[37].wr_en_this_byte ),
    .Q(\latch_mem.RAM[37][1] ));
 sg13g2_dlhq_1 _2072_ (.D(net867),
    .GATE(\latch_mem.genblk1[37].wr_en_this_byte ),
    .Q(\latch_mem.RAM[37][2] ));
 sg13g2_dlhq_1 _2073_ (.D(net857),
    .GATE(\latch_mem.genblk1[37].wr_en_this_byte ),
    .Q(\latch_mem.RAM[37][3] ));
 sg13g2_dlhq_1 _2074_ (.D(net845),
    .GATE(\latch_mem.genblk1[37].wr_en_this_byte ),
    .Q(\latch_mem.RAM[37][4] ));
 sg13g2_dlhq_1 _2075_ (.D(net836),
    .GATE(\latch_mem.genblk1[37].wr_en_this_byte ),
    .Q(\latch_mem.RAM[37][5] ));
 sg13g2_dlhq_1 _2076_ (.D(net824),
    .GATE(\latch_mem.genblk1[37].wr_en_this_byte ),
    .Q(\latch_mem.RAM[37][6] ));
 sg13g2_dlhq_1 _2077_ (.D(net813),
    .GATE(\latch_mem.genblk1[37].wr_en_this_byte ),
    .Q(\latch_mem.RAM[37][7] ));
 sg13g2_dlhq_1 _2078_ (.D(net889),
    .GATE(\latch_mem.genblk1[62].wr_en_this_byte ),
    .Q(\latch_mem.RAM[62][0] ));
 sg13g2_dlhq_1 _2079_ (.D(net880),
    .GATE(\latch_mem.genblk1[62].wr_en_this_byte ),
    .Q(\latch_mem.RAM[62][1] ));
 sg13g2_dlhq_1 _2080_ (.D(net869),
    .GATE(\latch_mem.genblk1[62].wr_en_this_byte ),
    .Q(\latch_mem.RAM[62][2] ));
 sg13g2_dlhq_1 _2081_ (.D(net859),
    .GATE(\latch_mem.genblk1[62].wr_en_this_byte ),
    .Q(\latch_mem.RAM[62][3] ));
 sg13g2_dlhq_1 _2082_ (.D(net851),
    .GATE(\latch_mem.genblk1[62].wr_en_this_byte ),
    .Q(\latch_mem.RAM[62][4] ));
 sg13g2_dlhq_1 _2083_ (.D(net838),
    .GATE(\latch_mem.genblk1[62].wr_en_this_byte ),
    .Q(\latch_mem.RAM[62][5] ));
 sg13g2_dlhq_1 _2084_ (.D(net827),
    .GATE(\latch_mem.genblk1[62].wr_en_this_byte ),
    .Q(\latch_mem.RAM[62][6] ));
 sg13g2_dlhq_1 _2085_ (.D(net821),
    .GATE(\latch_mem.genblk1[62].wr_en_this_byte ),
    .Q(\latch_mem.RAM[62][7] ));
 sg13g2_dlhq_1 _2086_ (.D(net892),
    .GATE(\latch_mem.genblk1[10].wr_en_this_byte ),
    .Q(\latch_mem.RAM[10][0] ));
 sg13g2_dlhq_1 _2087_ (.D(net883),
    .GATE(\latch_mem.genblk1[10].wr_en_this_byte ),
    .Q(\latch_mem.RAM[10][1] ));
 sg13g2_dlhq_1 _2088_ (.D(net873),
    .GATE(\latch_mem.genblk1[10].wr_en_this_byte ),
    .Q(\latch_mem.RAM[10][2] ));
 sg13g2_dlhq_1 _2089_ (.D(net862),
    .GATE(\latch_mem.genblk1[10].wr_en_this_byte ),
    .Q(\latch_mem.RAM[10][3] ));
 sg13g2_dlhq_1 _2090_ (.D(net849),
    .GATE(\latch_mem.genblk1[10].wr_en_this_byte ),
    .Q(\latch_mem.RAM[10][4] ));
 sg13g2_dlhq_1 _2091_ (.D(net840),
    .GATE(\latch_mem.genblk1[10].wr_en_this_byte ),
    .Q(\latch_mem.RAM[10][5] ));
 sg13g2_dlhq_1 _2092_ (.D(net829),
    .GATE(\latch_mem.genblk1[10].wr_en_this_byte ),
    .Q(\latch_mem.RAM[10][6] ));
 sg13g2_dlhq_1 _2093_ (.D(net820),
    .GATE(\latch_mem.genblk1[10].wr_en_this_byte ),
    .Q(\latch_mem.RAM[10][7] ));
 sg13g2_dlhq_1 _2094_ (.D(net887),
    .GATE(\latch_mem.genblk1[45].wr_en_this_byte ),
    .Q(\latch_mem.RAM[45][0] ));
 sg13g2_dlhq_1 _2095_ (.D(net876),
    .GATE(\latch_mem.genblk1[45].wr_en_this_byte ),
    .Q(\latch_mem.RAM[45][1] ));
 sg13g2_dlhq_1 _2096_ (.D(net866),
    .GATE(\latch_mem.genblk1[45].wr_en_this_byte ),
    .Q(\latch_mem.RAM[45][2] ));
 sg13g2_dlhq_1 _2097_ (.D(net856),
    .GATE(\latch_mem.genblk1[45].wr_en_this_byte ),
    .Q(\latch_mem.RAM[45][3] ));
 sg13g2_dlhq_1 _2098_ (.D(net844),
    .GATE(\latch_mem.genblk1[45].wr_en_this_byte ),
    .Q(\latch_mem.RAM[45][4] ));
 sg13g2_dlhq_1 _2099_ (.D(net834),
    .GATE(\latch_mem.genblk1[45].wr_en_this_byte ),
    .Q(\latch_mem.RAM[45][5] ));
 sg13g2_dlhq_1 _2100_ (.D(net824),
    .GATE(\latch_mem.genblk1[45].wr_en_this_byte ),
    .Q(\latch_mem.RAM[45][6] ));
 sg13g2_dlhq_1 _2101_ (.D(net813),
    .GATE(\latch_mem.genblk1[45].wr_en_this_byte ),
    .Q(\latch_mem.RAM[45][7] ));
 sg13g2_dlhq_1 _2102_ (.D(net890),
    .GATE(\latch_mem.genblk1[63].wr_en_this_byte ),
    .Q(\latch_mem.RAM[63][0] ));
 sg13g2_dlhq_1 _2103_ (.D(net880),
    .GATE(\latch_mem.genblk1[63].wr_en_this_byte ),
    .Q(\latch_mem.RAM[63][1] ));
 sg13g2_dlhq_1 _2104_ (.D(net869),
    .GATE(\latch_mem.genblk1[63].wr_en_this_byte ),
    .Q(\latch_mem.RAM[63][2] ));
 sg13g2_dlhq_1 _2105_ (.D(net855),
    .GATE(\latch_mem.genblk1[63].wr_en_this_byte ),
    .Q(\latch_mem.RAM[63][3] ));
 sg13g2_dlhq_1 _2106_ (.D(net851),
    .GATE(\latch_mem.genblk1[63].wr_en_this_byte ),
    .Q(\latch_mem.RAM[63][4] ));
 sg13g2_dlhq_1 _2107_ (.D(net837),
    .GATE(\latch_mem.genblk1[63].wr_en_this_byte ),
    .Q(\latch_mem.RAM[63][5] ));
 sg13g2_dlhq_1 _2108_ (.D(net827),
    .GATE(\latch_mem.genblk1[63].wr_en_this_byte ),
    .Q(\latch_mem.RAM[63][6] ));
 sg13g2_dlhq_1 _2109_ (.D(net819),
    .GATE(\latch_mem.genblk1[63].wr_en_this_byte ),
    .Q(\latch_mem.RAM[63][7] ));
 sg13g2_dlhq_1 _2110_ (.D(net884),
    .GATE(\latch_mem.genblk1[29].wr_en_this_byte ),
    .Q(\latch_mem.RAM[29][0] ));
 sg13g2_dlhq_1 _2111_ (.D(net875),
    .GATE(\latch_mem.genblk1[29].wr_en_this_byte ),
    .Q(\latch_mem.RAM[29][1] ));
 sg13g2_dlhq_1 _2112_ (.D(net864),
    .GATE(\latch_mem.genblk1[29].wr_en_this_byte ),
    .Q(\latch_mem.RAM[29][2] ));
 sg13g2_dlhq_1 _2113_ (.D(net852),
    .GATE(\latch_mem.genblk1[29].wr_en_this_byte ),
    .Q(\latch_mem.RAM[29][3] ));
 sg13g2_dlhq_1 _2114_ (.D(net842),
    .GATE(\latch_mem.genblk1[29].wr_en_this_byte ),
    .Q(\latch_mem.RAM[29][4] ));
 sg13g2_dlhq_1 _2115_ (.D(net832),
    .GATE(\latch_mem.genblk1[29].wr_en_this_byte ),
    .Q(\latch_mem.RAM[29][5] ));
 sg13g2_dlhq_1 _2116_ (.D(net823),
    .GATE(\latch_mem.genblk1[29].wr_en_this_byte ),
    .Q(\latch_mem.RAM[29][6] ));
 sg13g2_dlhq_1 _2117_ (.D(net812),
    .GATE(\latch_mem.genblk1[29].wr_en_this_byte ),
    .Q(\latch_mem.RAM[29][7] ));
 sg13g2_dlhq_1 _2118_ (.D(net891),
    .GATE(\latch_mem.genblk1[9].wr_en_this_byte ),
    .Q(\latch_mem.RAM[9][0] ));
 sg13g2_dlhq_1 _2119_ (.D(net881),
    .GATE(\latch_mem.genblk1[9].wr_en_this_byte ),
    .Q(\latch_mem.RAM[9][1] ));
 sg13g2_dlhq_1 _2120_ (.D(net872),
    .GATE(\latch_mem.genblk1[9].wr_en_this_byte ),
    .Q(\latch_mem.RAM[9][2] ));
 sg13g2_dlhq_1 _2121_ (.D(net861),
    .GATE(\latch_mem.genblk1[9].wr_en_this_byte ),
    .Q(\latch_mem.RAM[9][3] ));
 sg13g2_dlhq_1 _2122_ (.D(net850),
    .GATE(\latch_mem.genblk1[9].wr_en_this_byte ),
    .Q(\latch_mem.RAM[9][4] ));
 sg13g2_dlhq_1 _2123_ (.D(net840),
    .GATE(\latch_mem.genblk1[9].wr_en_this_byte ),
    .Q(\latch_mem.RAM[9][5] ));
 sg13g2_dlhq_1 _2124_ (.D(net830),
    .GATE(\latch_mem.genblk1[9].wr_en_this_byte ),
    .Q(\latch_mem.RAM[9][6] ));
 sg13g2_dlhq_1 _2125_ (.D(net817),
    .GATE(\latch_mem.genblk1[9].wr_en_this_byte ),
    .Q(\latch_mem.RAM[9][7] ));
 sg13g2_dlhq_1 _2126_ (.D(net884),
    .GATE(\latch_mem.genblk1[21].wr_en_this_byte ),
    .Q(\latch_mem.RAM[21][0] ));
 sg13g2_dlhq_1 _2127_ (.D(net874),
    .GATE(\latch_mem.genblk1[21].wr_en_this_byte ),
    .Q(\latch_mem.RAM[21][1] ));
 sg13g2_dlhq_1 _2128_ (.D(net864),
    .GATE(\latch_mem.genblk1[21].wr_en_this_byte ),
    .Q(\latch_mem.RAM[21][2] ));
 sg13g2_dlhq_1 _2129_ (.D(net852),
    .GATE(\latch_mem.genblk1[21].wr_en_this_byte ),
    .Q(\latch_mem.RAM[21][3] ));
 sg13g2_dlhq_1 _2130_ (.D(net842),
    .GATE(\latch_mem.genblk1[21].wr_en_this_byte ),
    .Q(\latch_mem.RAM[21][4] ));
 sg13g2_dlhq_1 _2131_ (.D(net833),
    .GATE(\latch_mem.genblk1[21].wr_en_this_byte ),
    .Q(\latch_mem.RAM[21][5] ));
 sg13g2_dlhq_1 _2132_ (.D(net822),
    .GATE(\latch_mem.genblk1[21].wr_en_this_byte ),
    .Q(\latch_mem.RAM[21][6] ));
 sg13g2_dlhq_1 _2133_ (.D(net812),
    .GATE(\latch_mem.genblk1[21].wr_en_this_byte ),
    .Q(\latch_mem.RAM[21][7] ));
 sg13g2_dlhq_1 _2134_ (.D(net887),
    .GATE(\latch_mem.genblk1[46].wr_en_this_byte ),
    .Q(\latch_mem.RAM[46][0] ));
 sg13g2_dlhq_1 _2135_ (.D(net876),
    .GATE(\latch_mem.genblk1[46].wr_en_this_byte ),
    .Q(\latch_mem.RAM[46][1] ));
 sg13g2_dlhq_1 _2136_ (.D(net866),
    .GATE(\latch_mem.genblk1[46].wr_en_this_byte ),
    .Q(\latch_mem.RAM[46][2] ));
 sg13g2_dlhq_1 _2137_ (.D(net857),
    .GATE(\latch_mem.genblk1[46].wr_en_this_byte ),
    .Q(\latch_mem.RAM[46][3] ));
 sg13g2_dlhq_1 _2138_ (.D(net845),
    .GATE(\latch_mem.genblk1[46].wr_en_this_byte ),
    .Q(\latch_mem.RAM[46][4] ));
 sg13g2_dlhq_1 _2139_ (.D(net834),
    .GATE(\latch_mem.genblk1[46].wr_en_this_byte ),
    .Q(\latch_mem.RAM[46][5] ));
 sg13g2_dlhq_1 _2140_ (.D(net825),
    .GATE(\latch_mem.genblk1[46].wr_en_this_byte ),
    .Q(\latch_mem.RAM[46][6] ));
 sg13g2_dlhq_1 _2141_ (.D(net815),
    .GATE(\latch_mem.genblk1[46].wr_en_this_byte ),
    .Q(\latch_mem.RAM[46][7] ));
 sg13g2_dlhq_1 _2142_ (.D(net891),
    .GATE(\latch_mem.genblk1[8].wr_en_this_byte ),
    .Q(\latch_mem.RAM[8][0] ));
 sg13g2_dlhq_1 _2143_ (.D(net881),
    .GATE(\latch_mem.genblk1[8].wr_en_this_byte ),
    .Q(\latch_mem.RAM[8][1] ));
 sg13g2_dlhq_1 _2144_ (.D(net871),
    .GATE(\latch_mem.genblk1[8].wr_en_this_byte ),
    .Q(\latch_mem.RAM[8][2] ));
 sg13g2_dlhq_1 _2145_ (.D(net861),
    .GATE(\latch_mem.genblk1[8].wr_en_this_byte ),
    .Q(\latch_mem.RAM[8][3] ));
 sg13g2_dlhq_1 _2146_ (.D(net849),
    .GATE(\latch_mem.genblk1[8].wr_en_this_byte ),
    .Q(\latch_mem.RAM[8][4] ));
 sg13g2_dlhq_1 _2147_ (.D(net840),
    .GATE(\latch_mem.genblk1[8].wr_en_this_byte ),
    .Q(\latch_mem.RAM[8][5] ));
 sg13g2_dlhq_1 _2148_ (.D(net830),
    .GATE(\latch_mem.genblk1[8].wr_en_this_byte ),
    .Q(\latch_mem.RAM[8][6] ));
 sg13g2_dlhq_1 _2149_ (.D(net817),
    .GATE(\latch_mem.genblk1[8].wr_en_this_byte ),
    .Q(\latch_mem.RAM[8][7] ));
 sg13g2_dlhq_1 _2150_ (.D(net888),
    .GATE(\latch_mem.genblk1[34].wr_en_this_byte ),
    .Q(\latch_mem.RAM[34][0] ));
 sg13g2_dlhq_1 _2151_ (.D(net877),
    .GATE(\latch_mem.genblk1[34].wr_en_this_byte ),
    .Q(\latch_mem.RAM[34][1] ));
 sg13g2_dlhq_1 _2152_ (.D(net867),
    .GATE(\latch_mem.genblk1[34].wr_en_this_byte ),
    .Q(\latch_mem.RAM[34][2] ));
 sg13g2_dlhq_1 _2153_ (.D(net857),
    .GATE(\latch_mem.genblk1[34].wr_en_this_byte ),
    .Q(\latch_mem.RAM[34][3] ));
 sg13g2_dlhq_1 _2154_ (.D(net845),
    .GATE(\latch_mem.genblk1[34].wr_en_this_byte ),
    .Q(\latch_mem.RAM[34][4] ));
 sg13g2_dlhq_1 _2155_ (.D(net835),
    .GATE(\latch_mem.genblk1[34].wr_en_this_byte ),
    .Q(\latch_mem.RAM[34][5] ));
 sg13g2_dlhq_1 _2156_ (.D(net824),
    .GATE(\latch_mem.genblk1[34].wr_en_this_byte ),
    .Q(\latch_mem.RAM[34][6] ));
 sg13g2_dlhq_1 _2157_ (.D(net815),
    .GATE(\latch_mem.genblk1[34].wr_en_this_byte ),
    .Q(\latch_mem.RAM[34][7] ));
 sg13g2_dlhq_1 _2158_ (.D(net887),
    .GATE(\latch_mem.genblk1[38].wr_en_this_byte ),
    .Q(\latch_mem.RAM[38][0] ));
 sg13g2_dlhq_1 _2159_ (.D(net876),
    .GATE(\latch_mem.genblk1[38].wr_en_this_byte ),
    .Q(\latch_mem.RAM[38][1] ));
 sg13g2_dlhq_1 _2160_ (.D(net866),
    .GATE(\latch_mem.genblk1[38].wr_en_this_byte ),
    .Q(\latch_mem.RAM[38][2] ));
 sg13g2_dlhq_1 _2161_ (.D(net856),
    .GATE(\latch_mem.genblk1[38].wr_en_this_byte ),
    .Q(\latch_mem.RAM[38][3] ));
 sg13g2_dlhq_1 _2162_ (.D(net844),
    .GATE(\latch_mem.genblk1[38].wr_en_this_byte ),
    .Q(\latch_mem.RAM[38][4] ));
 sg13g2_dlhq_1 _2163_ (.D(net835),
    .GATE(\latch_mem.genblk1[38].wr_en_this_byte ),
    .Q(\latch_mem.RAM[38][5] ));
 sg13g2_dlhq_1 _2164_ (.D(net824),
    .GATE(\latch_mem.genblk1[38].wr_en_this_byte ),
    .Q(\latch_mem.RAM[38][6] ));
 sg13g2_dlhq_1 _2165_ (.D(net813),
    .GATE(\latch_mem.genblk1[38].wr_en_this_byte ),
    .Q(\latch_mem.RAM[38][7] ));
 sg13g2_dlhq_1 _2166_ (.D(net892),
    .GATE(\latch_mem.genblk1[7].wr_en_this_byte ),
    .Q(\latch_mem.RAM[7][0] ));
 sg13g2_dlhq_1 _2167_ (.D(net882),
    .GATE(\latch_mem.genblk1[7].wr_en_this_byte ),
    .Q(\latch_mem.RAM[7][1] ));
 sg13g2_dlhq_1 _2168_ (.D(net872),
    .GATE(\latch_mem.genblk1[7].wr_en_this_byte ),
    .Q(\latch_mem.RAM[7][2] ));
 sg13g2_dlhq_1 _2169_ (.D(net861),
    .GATE(\latch_mem.genblk1[7].wr_en_this_byte ),
    .Q(\latch_mem.RAM[7][3] ));
 sg13g2_dlhq_1 _2170_ (.D(net849),
    .GATE(\latch_mem.genblk1[7].wr_en_this_byte ),
    .Q(\latch_mem.RAM[7][4] ));
 sg13g2_dlhq_1 _2171_ (.D(net839),
    .GATE(\latch_mem.genblk1[7].wr_en_this_byte ),
    .Q(\latch_mem.RAM[7][5] ));
 sg13g2_dlhq_1 _2172_ (.D(net829),
    .GATE(\latch_mem.genblk1[7].wr_en_this_byte ),
    .Q(\latch_mem.RAM[7][6] ));
 sg13g2_dlhq_1 _2173_ (.D(net817),
    .GATE(\latch_mem.genblk1[7].wr_en_this_byte ),
    .Q(\latch_mem.RAM[7][7] ));
 sg13g2_dlhq_1 _2174_ (.D(net888),
    .GATE(\latch_mem.genblk1[47].wr_en_this_byte ),
    .Q(\latch_mem.RAM[47][0] ));
 sg13g2_dlhq_1 _2175_ (.D(net877),
    .GATE(\latch_mem.genblk1[47].wr_en_this_byte ),
    .Q(\latch_mem.RAM[47][1] ));
 sg13g2_dlhq_1 _2176_ (.D(net867),
    .GATE(\latch_mem.genblk1[47].wr_en_this_byte ),
    .Q(\latch_mem.RAM[47][2] ));
 sg13g2_dlhq_1 _2177_ (.D(net857),
    .GATE(\latch_mem.genblk1[47].wr_en_this_byte ),
    .Q(\latch_mem.RAM[47][3] ));
 sg13g2_dlhq_1 _2178_ (.D(net844),
    .GATE(\latch_mem.genblk1[47].wr_en_this_byte ),
    .Q(\latch_mem.RAM[47][4] ));
 sg13g2_dlhq_1 _2179_ (.D(net835),
    .GATE(\latch_mem.genblk1[47].wr_en_this_byte ),
    .Q(\latch_mem.RAM[47][5] ));
 sg13g2_dlhq_1 _2180_ (.D(net825),
    .GATE(\latch_mem.genblk1[47].wr_en_this_byte ),
    .Q(\latch_mem.RAM[47][6] ));
 sg13g2_dlhq_1 _2181_ (.D(net813),
    .GATE(\latch_mem.genblk1[47].wr_en_this_byte ),
    .Q(\latch_mem.RAM[47][7] ));
 sg13g2_dlhq_1 _2182_ (.D(net885),
    .GATE(\latch_mem.genblk1[20].wr_en_this_byte ),
    .Q(\latch_mem.RAM[20][0] ));
 sg13g2_dlhq_1 _2183_ (.D(net874),
    .GATE(\latch_mem.genblk1[20].wr_en_this_byte ),
    .Q(\latch_mem.RAM[20][1] ));
 sg13g2_dlhq_1 _2184_ (.D(net865),
    .GATE(\latch_mem.genblk1[20].wr_en_this_byte ),
    .Q(\latch_mem.RAM[20][2] ));
 sg13g2_dlhq_1 _2185_ (.D(net852),
    .GATE(\latch_mem.genblk1[20].wr_en_this_byte ),
    .Q(\latch_mem.RAM[20][3] ));
 sg13g2_dlhq_1 _2186_ (.D(net843),
    .GATE(\latch_mem.genblk1[20].wr_en_this_byte ),
    .Q(\latch_mem.RAM[20][4] ));
 sg13g2_dlhq_1 _2187_ (.D(net833),
    .GATE(\latch_mem.genblk1[20].wr_en_this_byte ),
    .Q(\latch_mem.RAM[20][5] ));
 sg13g2_dlhq_1 _2188_ (.D(net823),
    .GATE(\latch_mem.genblk1[20].wr_en_this_byte ),
    .Q(\latch_mem.RAM[20][6] ));
 sg13g2_dlhq_1 _2189_ (.D(net814),
    .GATE(\latch_mem.genblk1[20].wr_en_this_byte ),
    .Q(\latch_mem.RAM[20][7] ));
 sg13g2_dlhq_1 _2190_ (.D(net891),
    .GATE(\latch_mem.genblk1[6].wr_en_this_byte ),
    .Q(\latch_mem.RAM[6][0] ));
 sg13g2_dlhq_1 _2191_ (.D(net881),
    .GATE(\latch_mem.genblk1[6].wr_en_this_byte ),
    .Q(\latch_mem.RAM[6][1] ));
 sg13g2_dlhq_1 _2192_ (.D(net871),
    .GATE(\latch_mem.genblk1[6].wr_en_this_byte ),
    .Q(\latch_mem.RAM[6][2] ));
 sg13g2_dlhq_1 _2193_ (.D(net862),
    .GATE(\latch_mem.genblk1[6].wr_en_this_byte ),
    .Q(\latch_mem.RAM[6][3] ));
 sg13g2_dlhq_1 _2194_ (.D(net849),
    .GATE(\latch_mem.genblk1[6].wr_en_this_byte ),
    .Q(\latch_mem.RAM[6][4] ));
 sg13g2_dlhq_1 _2195_ (.D(net839),
    .GATE(\latch_mem.genblk1[6].wr_en_this_byte ),
    .Q(\latch_mem.RAM[6][5] ));
 sg13g2_dlhq_1 _2196_ (.D(net829),
    .GATE(\latch_mem.genblk1[6].wr_en_this_byte ),
    .Q(\latch_mem.RAM[6][6] ));
 sg13g2_dlhq_1 _2197_ (.D(net817),
    .GATE(\latch_mem.genblk1[6].wr_en_this_byte ),
    .Q(\latch_mem.RAM[6][7] ));
 sg13g2_dlhq_1 _2198_ (.D(net884),
    .GATE(\latch_mem.genblk1[26].wr_en_this_byte ),
    .Q(\latch_mem.RAM[26][0] ));
 sg13g2_dlhq_1 _2199_ (.D(net875),
    .GATE(\latch_mem.genblk1[26].wr_en_this_byte ),
    .Q(\latch_mem.RAM[26][1] ));
 sg13g2_dlhq_1 _2200_ (.D(net864),
    .GATE(\latch_mem.genblk1[26].wr_en_this_byte ),
    .Q(\latch_mem.RAM[26][2] ));
 sg13g2_dlhq_1 _2201_ (.D(net853),
    .GATE(\latch_mem.genblk1[26].wr_en_this_byte ),
    .Q(\latch_mem.RAM[26][3] ));
 sg13g2_dlhq_1 _2202_ (.D(net842),
    .GATE(\latch_mem.genblk1[26].wr_en_this_byte ),
    .Q(\latch_mem.RAM[26][4] ));
 sg13g2_dlhq_1 _2203_ (.D(net832),
    .GATE(\latch_mem.genblk1[26].wr_en_this_byte ),
    .Q(\latch_mem.RAM[26][5] ));
 sg13g2_dlhq_1 _2204_ (.D(net822),
    .GATE(\latch_mem.genblk1[26].wr_en_this_byte ),
    .Q(\latch_mem.RAM[26][6] ));
 sg13g2_dlhq_1 _2205_ (.D(net814),
    .GATE(\latch_mem.genblk1[26].wr_en_this_byte ),
    .Q(\latch_mem.RAM[26][7] ));
 sg13g2_dlhq_1 _2206_ (.D(net890),
    .GATE(\latch_mem.genblk1[48].wr_en_this_byte ),
    .Q(\latch_mem.RAM[48][0] ));
 sg13g2_dlhq_1 _2207_ (.D(net879),
    .GATE(\latch_mem.genblk1[48].wr_en_this_byte ),
    .Q(\latch_mem.RAM[48][1] ));
 sg13g2_dlhq_1 _2208_ (.D(net870),
    .GATE(\latch_mem.genblk1[48].wr_en_this_byte ),
    .Q(\latch_mem.RAM[48][2] ));
 sg13g2_dlhq_1 _2209_ (.D(net860),
    .GATE(\latch_mem.genblk1[48].wr_en_this_byte ),
    .Q(\latch_mem.RAM[48][3] ));
 sg13g2_dlhq_1 _2210_ (.D(net847),
    .GATE(\latch_mem.genblk1[48].wr_en_this_byte ),
    .Q(\latch_mem.RAM[48][4] ));
 sg13g2_dlhq_1 _2211_ (.D(net841),
    .GATE(\latch_mem.genblk1[48].wr_en_this_byte ),
    .Q(\latch_mem.RAM[48][5] ));
 sg13g2_dlhq_1 _2212_ (.D(net831),
    .GATE(\latch_mem.genblk1[48].wr_en_this_byte ),
    .Q(\latch_mem.RAM[48][6] ));
 sg13g2_dlhq_1 _2213_ (.D(net818),
    .GATE(\latch_mem.genblk1[48].wr_en_this_byte ),
    .Q(\latch_mem.RAM[48][7] ));
 sg13g2_dlhq_1 _2214_ (.D(net891),
    .GATE(\latch_mem.genblk1[5].wr_en_this_byte ),
    .Q(\latch_mem.RAM[5][0] ));
 sg13g2_dlhq_1 _2215_ (.D(net882),
    .GATE(\latch_mem.genblk1[5].wr_en_this_byte ),
    .Q(\latch_mem.RAM[5][1] ));
 sg13g2_dlhq_1 _2216_ (.D(net871),
    .GATE(\latch_mem.genblk1[5].wr_en_this_byte ),
    .Q(\latch_mem.RAM[5][2] ));
 sg13g2_dlhq_1 _2217_ (.D(net861),
    .GATE(\latch_mem.genblk1[5].wr_en_this_byte ),
    .Q(\latch_mem.RAM[5][3] ));
 sg13g2_dlhq_1 _2218_ (.D(net850),
    .GATE(\latch_mem.genblk1[5].wr_en_this_byte ),
    .Q(\latch_mem.RAM[5][4] ));
 sg13g2_dlhq_1 _2219_ (.D(net839),
    .GATE(\latch_mem.genblk1[5].wr_en_this_byte ),
    .Q(\latch_mem.RAM[5][5] ));
 sg13g2_dlhq_1 _2220_ (.D(net830),
    .GATE(\latch_mem.genblk1[5].wr_en_this_byte ),
    .Q(\latch_mem.RAM[5][6] ));
 sg13g2_dlhq_1 _2221_ (.D(net817),
    .GATE(\latch_mem.genblk1[5].wr_en_this_byte ),
    .Q(\latch_mem.RAM[5][7] ));
 sg13g2_dlhq_1 _2222_ (.D(net886),
    .GATE(\latch_mem.genblk1[30].wr_en_this_byte ),
    .Q(\latch_mem.RAM[30][0] ));
 sg13g2_dlhq_1 _2223_ (.D(net874),
    .GATE(\latch_mem.genblk1[30].wr_en_this_byte ),
    .Q(\latch_mem.RAM[30][1] ));
 sg13g2_dlhq_1 _2224_ (.D(net864),
    .GATE(\latch_mem.genblk1[30].wr_en_this_byte ),
    .Q(\latch_mem.RAM[30][2] ));
 sg13g2_dlhq_1 _2225_ (.D(net854),
    .GATE(\latch_mem.genblk1[30].wr_en_this_byte ),
    .Q(\latch_mem.RAM[30][3] ));
 sg13g2_dlhq_1 _2226_ (.D(net843),
    .GATE(\latch_mem.genblk1[30].wr_en_this_byte ),
    .Q(\latch_mem.RAM[30][4] ));
 sg13g2_dlhq_1 _2227_ (.D(net833),
    .GATE(\latch_mem.genblk1[30].wr_en_this_byte ),
    .Q(\latch_mem.RAM[30][5] ));
 sg13g2_dlhq_1 _2228_ (.D(net823),
    .GATE(\latch_mem.genblk1[30].wr_en_this_byte ),
    .Q(\latch_mem.RAM[30][6] ));
 sg13g2_dlhq_1 _2229_ (.D(net814),
    .GATE(\latch_mem.genblk1[30].wr_en_this_byte ),
    .Q(\latch_mem.RAM[30][7] ));
 sg13g2_dlhq_1 _2230_ (.D(net884),
    .GATE(\latch_mem.genblk1[19].wr_en_this_byte ),
    .Q(\latch_mem.RAM[19][0] ));
 sg13g2_dlhq_1 _2231_ (.D(net874),
    .GATE(\latch_mem.genblk1[19].wr_en_this_byte ),
    .Q(\latch_mem.RAM[19][1] ));
 sg13g2_dlhq_1 _2232_ (.D(net865),
    .GATE(\latch_mem.genblk1[19].wr_en_this_byte ),
    .Q(\latch_mem.RAM[19][2] ));
 sg13g2_dlhq_1 _2233_ (.D(net853),
    .GATE(\latch_mem.genblk1[19].wr_en_this_byte ),
    .Q(\latch_mem.RAM[19][3] ));
 sg13g2_dlhq_1 _2234_ (.D(net843),
    .GATE(\latch_mem.genblk1[19].wr_en_this_byte ),
    .Q(\latch_mem.RAM[19][4] ));
 sg13g2_dlhq_1 _2235_ (.D(net832),
    .GATE(\latch_mem.genblk1[19].wr_en_this_byte ),
    .Q(\latch_mem.RAM[19][5] ));
 sg13g2_dlhq_1 _2236_ (.D(net822),
    .GATE(\latch_mem.genblk1[19].wr_en_this_byte ),
    .Q(\latch_mem.RAM[19][6] ));
 sg13g2_dlhq_1 _2237_ (.D(net812),
    .GATE(\latch_mem.genblk1[19].wr_en_this_byte ),
    .Q(\latch_mem.RAM[19][7] ));
 sg13g2_dlhq_1 _2238_ (.D(net892),
    .GATE(\latch_mem.genblk1[4].wr_en_this_byte ),
    .Q(\latch_mem.RAM[4][0] ));
 sg13g2_dlhq_1 _2239_ (.D(net881),
    .GATE(\latch_mem.genblk1[4].wr_en_this_byte ),
    .Q(\latch_mem.RAM[4][1] ));
 sg13g2_dlhq_1 _2240_ (.D(net871),
    .GATE(\latch_mem.genblk1[4].wr_en_this_byte ),
    .Q(\latch_mem.RAM[4][2] ));
 sg13g2_dlhq_1 _2241_ (.D(net862),
    .GATE(\latch_mem.genblk1[4].wr_en_this_byte ),
    .Q(\latch_mem.RAM[4][3] ));
 sg13g2_dlhq_1 _2242_ (.D(net849),
    .GATE(\latch_mem.genblk1[4].wr_en_this_byte ),
    .Q(\latch_mem.RAM[4][4] ));
 sg13g2_dlhq_1 _2243_ (.D(net839),
    .GATE(\latch_mem.genblk1[4].wr_en_this_byte ),
    .Q(\latch_mem.RAM[4][5] ));
 sg13g2_dlhq_1 _2244_ (.D(net830),
    .GATE(\latch_mem.genblk1[4].wr_en_this_byte ),
    .Q(\latch_mem.RAM[4][6] ));
 sg13g2_dlhq_1 _2245_ (.D(net820),
    .GATE(\latch_mem.genblk1[4].wr_en_this_byte ),
    .Q(\latch_mem.RAM[4][7] ));
 sg13g2_dlhq_1 _2246_ (.D(net890),
    .GATE(\latch_mem.genblk1[49].wr_en_this_byte ),
    .Q(\latch_mem.RAM[49][0] ));
 sg13g2_dlhq_1 _2247_ (.D(net879),
    .GATE(\latch_mem.genblk1[49].wr_en_this_byte ),
    .Q(\latch_mem.RAM[49][1] ));
 sg13g2_dlhq_1 _2248_ (.D(net869),
    .GATE(\latch_mem.genblk1[49].wr_en_this_byte ),
    .Q(\latch_mem.RAM[49][2] ));
 sg13g2_dlhq_1 _2249_ (.D(net860),
    .GATE(\latch_mem.genblk1[49].wr_en_this_byte ),
    .Q(\latch_mem.RAM[49][3] ));
 sg13g2_dlhq_1 _2250_ (.D(net847),
    .GATE(\latch_mem.genblk1[49].wr_en_this_byte ),
    .Q(\latch_mem.RAM[49][4] ));
 sg13g2_dlhq_1 _2251_ (.D(net837),
    .GATE(\latch_mem.genblk1[49].wr_en_this_byte ),
    .Q(\latch_mem.RAM[49][5] ));
 sg13g2_dlhq_1 _2252_ (.D(net828),
    .GATE(\latch_mem.genblk1[49].wr_en_this_byte ),
    .Q(\latch_mem.RAM[49][6] ));
 sg13g2_dlhq_1 _2253_ (.D(net818),
    .GATE(\latch_mem.genblk1[49].wr_en_this_byte ),
    .Q(\latch_mem.RAM[49][7] ));
 sg13g2_dlhq_1 _2254_ (.D(net888),
    .GATE(\latch_mem.genblk1[39].wr_en_this_byte ),
    .Q(\latch_mem.RAM[39][0] ));
 sg13g2_dlhq_1 _2255_ (.D(net877),
    .GATE(\latch_mem.genblk1[39].wr_en_this_byte ),
    .Q(\latch_mem.RAM[39][1] ));
 sg13g2_dlhq_1 _2256_ (.D(net866),
    .GATE(\latch_mem.genblk1[39].wr_en_this_byte ),
    .Q(\latch_mem.RAM[39][2] ));
 sg13g2_dlhq_1 _2257_ (.D(net857),
    .GATE(\latch_mem.genblk1[39].wr_en_this_byte ),
    .Q(\latch_mem.RAM[39][3] ));
 sg13g2_dlhq_1 _2258_ (.D(net844),
    .GATE(\latch_mem.genblk1[39].wr_en_this_byte ),
    .Q(\latch_mem.RAM[39][4] ));
 sg13g2_dlhq_1 _2259_ (.D(net834),
    .GATE(\latch_mem.genblk1[39].wr_en_this_byte ),
    .Q(\latch_mem.RAM[39][5] ));
 sg13g2_dlhq_1 _2260_ (.D(net825),
    .GATE(\latch_mem.genblk1[39].wr_en_this_byte ),
    .Q(\latch_mem.RAM[39][6] ));
 sg13g2_dlhq_1 _2261_ (.D(net813),
    .GATE(\latch_mem.genblk1[39].wr_en_this_byte ),
    .Q(\latch_mem.RAM[39][7] ));
 sg13g2_dlhq_1 _2262_ (.D(net892),
    .GATE(\latch_mem.genblk1[3].wr_en_this_byte ),
    .Q(\latch_mem.RAM[3][0] ));
 sg13g2_dlhq_1 _2263_ (.D(net882),
    .GATE(\latch_mem.genblk1[3].wr_en_this_byte ),
    .Q(\latch_mem.RAM[3][1] ));
 sg13g2_dlhq_1 _2264_ (.D(net872),
    .GATE(\latch_mem.genblk1[3].wr_en_this_byte ),
    .Q(\latch_mem.RAM[3][2] ));
 sg13g2_dlhq_1 _2265_ (.D(net861),
    .GATE(\latch_mem.genblk1[3].wr_en_this_byte ),
    .Q(\latch_mem.RAM[3][3] ));
 sg13g2_dlhq_1 _2266_ (.D(net849),
    .GATE(\latch_mem.genblk1[3].wr_en_this_byte ),
    .Q(\latch_mem.RAM[3][4] ));
 sg13g2_dlhq_1 _2267_ (.D(net840),
    .GATE(\latch_mem.genblk1[3].wr_en_this_byte ),
    .Q(\latch_mem.RAM[3][5] ));
 sg13g2_dlhq_1 _2268_ (.D(net829),
    .GATE(\latch_mem.genblk1[3].wr_en_this_byte ),
    .Q(\latch_mem.RAM[3][6] ));
 sg13g2_dlhq_1 _2269_ (.D(net817),
    .GATE(\latch_mem.genblk1[3].wr_en_this_byte ),
    .Q(\latch_mem.RAM[3][7] ));
 sg13g2_dlhq_1 _2270_ (.D(net886),
    .GATE(\latch_mem.genblk1[31].wr_en_this_byte ),
    .Q(\latch_mem.RAM[31][0] ));
 sg13g2_dlhq_1 _2271_ (.D(net874),
    .GATE(\latch_mem.genblk1[31].wr_en_this_byte ),
    .Q(\latch_mem.RAM[31][1] ));
 sg13g2_dlhq_1 _2272_ (.D(net864),
    .GATE(\latch_mem.genblk1[31].wr_en_this_byte ),
    .Q(\latch_mem.RAM[31][2] ));
 sg13g2_dlhq_1 _2273_ (.D(net853),
    .GATE(\latch_mem.genblk1[31].wr_en_this_byte ),
    .Q(\latch_mem.RAM[31][3] ));
 sg13g2_dlhq_1 _2274_ (.D(net843),
    .GATE(\latch_mem.genblk1[31].wr_en_this_byte ),
    .Q(\latch_mem.RAM[31][4] ));
 sg13g2_dlhq_1 _2275_ (.D(net832),
    .GATE(\latch_mem.genblk1[31].wr_en_this_byte ),
    .Q(\latch_mem.RAM[31][5] ));
 sg13g2_dlhq_1 _2276_ (.D(net822),
    .GATE(\latch_mem.genblk1[31].wr_en_this_byte ),
    .Q(\latch_mem.RAM[31][6] ));
 sg13g2_dlhq_1 _2277_ (.D(net812),
    .GATE(\latch_mem.genblk1[31].wr_en_this_byte ),
    .Q(\latch_mem.RAM[31][7] ));
 sg13g2_dlhq_1 _2278_ (.D(net890),
    .GATE(\latch_mem.genblk1[50].wr_en_this_byte ),
    .Q(\latch_mem.RAM[50][0] ));
 sg13g2_dlhq_1 _2279_ (.D(net880),
    .GATE(\latch_mem.genblk1[50].wr_en_this_byte ),
    .Q(\latch_mem.RAM[50][1] ));
 sg13g2_dlhq_1 _2280_ (.D(net870),
    .GATE(\latch_mem.genblk1[50].wr_en_this_byte ),
    .Q(\latch_mem.RAM[50][2] ));
 sg13g2_dlhq_1 _2281_ (.D(net855),
    .GATE(\latch_mem.genblk1[50].wr_en_this_byte ),
    .Q(\latch_mem.RAM[50][3] ));
 sg13g2_dlhq_1 _2282_ (.D(net848),
    .GATE(\latch_mem.genblk1[50].wr_en_this_byte ),
    .Q(\latch_mem.RAM[50][4] ));
 sg13g2_dlhq_1 _2283_ (.D(net837),
    .GATE(\latch_mem.genblk1[50].wr_en_this_byte ),
    .Q(\latch_mem.RAM[50][5] ));
 sg13g2_dlhq_1 _2284_ (.D(net827),
    .GATE(\latch_mem.genblk1[50].wr_en_this_byte ),
    .Q(\latch_mem.RAM[50][6] ));
 sg13g2_dlhq_1 _2285_ (.D(net818),
    .GATE(\latch_mem.genblk1[50].wr_en_this_byte ),
    .Q(\latch_mem.RAM[50][7] ));
 sg13g2_dlhq_1 _2286_ (.D(net891),
    .GATE(\latch_mem.genblk1[2].wr_en_this_byte ),
    .Q(\latch_mem.RAM[2][0] ));
 sg13g2_dlhq_1 _2287_ (.D(net882),
    .GATE(\latch_mem.genblk1[2].wr_en_this_byte ),
    .Q(\latch_mem.RAM[2][1] ));
 sg13g2_dlhq_1 _2288_ (.D(net871),
    .GATE(\latch_mem.genblk1[2].wr_en_this_byte ),
    .Q(\latch_mem.RAM[2][2] ));
 sg13g2_dlhq_1 _2289_ (.D(net861),
    .GATE(\latch_mem.genblk1[2].wr_en_this_byte ),
    .Q(\latch_mem.RAM[2][3] ));
 sg13g2_dlhq_1 _2290_ (.D(net850),
    .GATE(\latch_mem.genblk1[2].wr_en_this_byte ),
    .Q(\latch_mem.RAM[2][4] ));
 sg13g2_dlhq_1 _2291_ (.D(net839),
    .GATE(\latch_mem.genblk1[2].wr_en_this_byte ),
    .Q(\latch_mem.RAM[2][5] ));
 sg13g2_dlhq_1 _2292_ (.D(net830),
    .GATE(\latch_mem.genblk1[2].wr_en_this_byte ),
    .Q(\latch_mem.RAM[2][6] ));
 sg13g2_dlhq_1 _2293_ (.D(net820),
    .GATE(\latch_mem.genblk1[2].wr_en_this_byte ),
    .Q(\latch_mem.RAM[2][7] ));
 sg13g2_dlhq_1 _2294_ (.D(net886),
    .GATE(\latch_mem.genblk1[18].wr_en_this_byte ),
    .Q(\latch_mem.RAM[18][0] ));
 sg13g2_dlhq_1 _2295_ (.D(net875),
    .GATE(\latch_mem.genblk1[18].wr_en_this_byte ),
    .Q(\latch_mem.RAM[18][1] ));
 sg13g2_dlhq_1 _2296_ (.D(net865),
    .GATE(\latch_mem.genblk1[18].wr_en_this_byte ),
    .Q(\latch_mem.RAM[18][2] ));
 sg13g2_dlhq_1 _2297_ (.D(net853),
    .GATE(\latch_mem.genblk1[18].wr_en_this_byte ),
    .Q(\latch_mem.RAM[18][3] ));
 sg13g2_dlhq_1 _2298_ (.D(net843),
    .GATE(\latch_mem.genblk1[18].wr_en_this_byte ),
    .Q(\latch_mem.RAM[18][4] ));
 sg13g2_dlhq_1 _2299_ (.D(net833),
    .GATE(\latch_mem.genblk1[18].wr_en_this_byte ),
    .Q(\latch_mem.RAM[18][5] ));
 sg13g2_dlhq_1 _2300_ (.D(net823),
    .GATE(\latch_mem.genblk1[18].wr_en_this_byte ),
    .Q(\latch_mem.RAM[18][6] ));
 sg13g2_dlhq_1 _2301_ (.D(net814),
    .GATE(\latch_mem.genblk1[18].wr_en_this_byte ),
    .Q(\latch_mem.RAM[18][7] ));
 sg13g2_dlhq_1 _2302_ (.D(net885),
    .GATE(\latch_mem.genblk1[25].wr_en_this_byte ),
    .Q(\latch_mem.RAM[25][0] ));
 sg13g2_dlhq_1 _2303_ (.D(net875),
    .GATE(\latch_mem.genblk1[25].wr_en_this_byte ),
    .Q(\latch_mem.RAM[25][1] ));
 sg13g2_dlhq_1 _2304_ (.D(net865),
    .GATE(\latch_mem.genblk1[25].wr_en_this_byte ),
    .Q(\latch_mem.RAM[25][2] ));
 sg13g2_dlhq_1 _2305_ (.D(net852),
    .GATE(\latch_mem.genblk1[25].wr_en_this_byte ),
    .Q(\latch_mem.RAM[25][3] ));
 sg13g2_dlhq_1 _2306_ (.D(net842),
    .GATE(\latch_mem.genblk1[25].wr_en_this_byte ),
    .Q(\latch_mem.RAM[25][4] ));
 sg13g2_dlhq_1 _2307_ (.D(net832),
    .GATE(\latch_mem.genblk1[25].wr_en_this_byte ),
    .Q(\latch_mem.RAM[25][5] ));
 sg13g2_dlhq_1 _2308_ (.D(net823),
    .GATE(\latch_mem.genblk1[25].wr_en_this_byte ),
    .Q(\latch_mem.RAM[25][6] ));
 sg13g2_dlhq_1 _2309_ (.D(net814),
    .GATE(\latch_mem.genblk1[25].wr_en_this_byte ),
    .Q(\latch_mem.RAM[25][7] ));
 sg13g2_dlhq_1 _2310_ (.D(net892),
    .GATE(\latch_mem.genblk1[1].wr_en_this_byte ),
    .Q(\latch_mem.RAM[1][0] ));
 sg13g2_dlhq_1 _2311_ (.D(net881),
    .GATE(\latch_mem.genblk1[1].wr_en_this_byte ),
    .Q(\latch_mem.RAM[1][1] ));
 sg13g2_dlhq_1 _2312_ (.D(net872),
    .GATE(\latch_mem.genblk1[1].wr_en_this_byte ),
    .Q(\latch_mem.RAM[1][2] ));
 sg13g2_dlhq_1 _2313_ (.D(net862),
    .GATE(\latch_mem.genblk1[1].wr_en_this_byte ),
    .Q(\latch_mem.RAM[1][3] ));
 sg13g2_dlhq_1 _2314_ (.D(net850),
    .GATE(\latch_mem.genblk1[1].wr_en_this_byte ),
    .Q(\latch_mem.RAM[1][4] ));
 sg13g2_dlhq_1 _2315_ (.D(net840),
    .GATE(\latch_mem.genblk1[1].wr_en_this_byte ),
    .Q(\latch_mem.RAM[1][5] ));
 sg13g2_dlhq_1 _2316_ (.D(net829),
    .GATE(\latch_mem.genblk1[1].wr_en_this_byte ),
    .Q(\latch_mem.RAM[1][6] ));
 sg13g2_dlhq_1 _2317_ (.D(net820),
    .GATE(\latch_mem.genblk1[1].wr_en_this_byte ),
    .Q(\latch_mem.RAM[1][7] ));
 sg13g2_dlhq_1 _2318_ (.D(net889),
    .GATE(\latch_mem.genblk1[51].wr_en_this_byte ),
    .Q(\latch_mem.RAM[51][0] ));
 sg13g2_dlhq_1 _2319_ (.D(net880),
    .GATE(\latch_mem.genblk1[51].wr_en_this_byte ),
    .Q(\latch_mem.RAM[51][1] ));
 sg13g2_dlhq_1 _2320_ (.D(net870),
    .GATE(\latch_mem.genblk1[51].wr_en_this_byte ),
    .Q(\latch_mem.RAM[51][2] ));
 sg13g2_dlhq_1 _2321_ (.D(net859),
    .GATE(\latch_mem.genblk1[51].wr_en_this_byte ),
    .Q(\latch_mem.RAM[51][3] ));
 sg13g2_dlhq_1 _2322_ (.D(net847),
    .GATE(\latch_mem.genblk1[51].wr_en_this_byte ),
    .Q(\latch_mem.RAM[51][4] ));
 sg13g2_dlhq_1 _2323_ (.D(net838),
    .GATE(\latch_mem.genblk1[51].wr_en_this_byte ),
    .Q(\latch_mem.RAM[51][5] ));
 sg13g2_dlhq_1 _2324_ (.D(net828),
    .GATE(\latch_mem.genblk1[51].wr_en_this_byte ),
    .Q(\latch_mem.RAM[51][6] ));
 sg13g2_dlhq_1 _2325_ (.D(net819),
    .GATE(\latch_mem.genblk1[51].wr_en_this_byte ),
    .Q(\latch_mem.RAM[51][7] ));
 sg13g2_dlhq_1 _2326_ (.D(net888),
    .GATE(\latch_mem.genblk1[40].wr_en_this_byte ),
    .Q(\latch_mem.RAM[40][0] ));
 sg13g2_dlhq_1 _2327_ (.D(net877),
    .GATE(\latch_mem.genblk1[40].wr_en_this_byte ),
    .Q(\latch_mem.RAM[40][1] ));
 sg13g2_dlhq_1 _2328_ (.D(net867),
    .GATE(\latch_mem.genblk1[40].wr_en_this_byte ),
    .Q(\latch_mem.RAM[40][2] ));
 sg13g2_dlhq_1 _2329_ (.D(net856),
    .GATE(\latch_mem.genblk1[40].wr_en_this_byte ),
    .Q(\latch_mem.RAM[40][3] ));
 sg13g2_dlhq_1 _2330_ (.D(net845),
    .GATE(\latch_mem.genblk1[40].wr_en_this_byte ),
    .Q(\latch_mem.RAM[40][4] ));
 sg13g2_dlhq_1 _2331_ (.D(net835),
    .GATE(\latch_mem.genblk1[40].wr_en_this_byte ),
    .Q(\latch_mem.RAM[40][5] ));
 sg13g2_dlhq_1 _2332_ (.D(net825),
    .GATE(\latch_mem.genblk1[40].wr_en_this_byte ),
    .Q(\latch_mem.RAM[40][6] ));
 sg13g2_dlhq_1 _2333_ (.D(net815),
    .GATE(\latch_mem.genblk1[40].wr_en_this_byte ),
    .Q(\latch_mem.RAM[40][7] ));
 sg13g2_dlhq_1 _2334_ (.D(net891),
    .GATE(\latch_mem.genblk1[0].wr_en_this_byte ),
    .Q(\latch_mem.RAM[0][0] ));
 sg13g2_dlhq_1 _2335_ (.D(net882),
    .GATE(\latch_mem.genblk1[0].wr_en_this_byte ),
    .Q(\latch_mem.RAM[0][1] ));
 sg13g2_dlhq_1 _2336_ (.D(net871),
    .GATE(\latch_mem.genblk1[0].wr_en_this_byte ),
    .Q(\latch_mem.RAM[0][2] ));
 sg13g2_dlhq_1 _2337_ (.D(net861),
    .GATE(\latch_mem.genblk1[0].wr_en_this_byte ),
    .Q(\latch_mem.RAM[0][3] ));
 sg13g2_dlhq_1 _2338_ (.D(net850),
    .GATE(\latch_mem.genblk1[0].wr_en_this_byte ),
    .Q(\latch_mem.RAM[0][4] ));
 sg13g2_dlhq_1 _2339_ (.D(net839),
    .GATE(\latch_mem.genblk1[0].wr_en_this_byte ),
    .Q(\latch_mem.RAM[0][5] ));
 sg13g2_dlhq_1 _2340_ (.D(net829),
    .GATE(\latch_mem.genblk1[0].wr_en_this_byte ),
    .Q(\latch_mem.RAM[0][6] ));
 sg13g2_dlhq_1 _2341_ (.D(net821),
    .GATE(\latch_mem.genblk1[0].wr_en_this_byte ),
    .Q(\latch_mem.RAM[0][7] ));
 sg13g2_dfrbp_1 _2342_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net72),
    .D(_0004_),
    .Q_N(_0830_),
    .Q(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_dfrbp_1 _2343_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net73),
    .D(_0007_),
    .Q_N(_0831_),
    .Q(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_dfrbp_1 _2344_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net75),
    .D(net131),
    .Q_N(_0832_),
    .Q(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_dfrbp_1 _2345_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net51),
    .D(_0005_),
    .Q_N(_0782_),
    .Q(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_dfrbp_1 _2346_ (.CLK(net98),
    .RESET_B(net76),
    .D(_0008_),
    .Q_N(_0833_),
    .Q(\latch_mem.wr_en_ok ));
 sg13g2_dfrbp_1 _2347_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net77),
    .D(net123),
    .Q_N(_0834_),
    .Q(\latch_mem.addr_read[0] ));
 sg13g2_dfrbp_1 _2348_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net78),
    .D(net107),
    .Q_N(_0835_),
    .Q(\latch_mem.addr_read[1] ));
 sg13g2_dfrbp_1 _2349_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net23),
    .D(net102),
    .Q_N(_0836_),
    .Q(\latch_mem.addr_read[2] ));
 sg13g2_dfrbp_1 _2350_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net49),
    .D(net101),
    .Q_N(_0781_),
    .Q(\latch_mem.addr_read[3] ));
 sg13g2_dfrbp_1 _2351_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net46),
    .D(_0076_),
    .Q_N(_0780_),
    .Q(\latch_mem.addr_write[0] ));
 sg13g2_dfrbp_1 _2352_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net44),
    .D(_0077_),
    .Q_N(_0779_),
    .Q(\latch_mem.addr_write[1] ));
 sg13g2_dfrbp_1 _2353_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net42),
    .D(_0078_),
    .Q_N(_0778_),
    .Q(\latch_mem.addr_write[2] ));
 sg13g2_dfrbp_1 _2354_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net40),
    .D(_0079_),
    .Q_N(_0777_),
    .Q(\latch_mem.addr_write[3] ));
 sg13g2_dfrbp_1 _2355_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net38),
    .D(_0080_),
    .Q_N(_0776_),
    .Q(\latch_mem.addr_write[4] ));
 sg13g2_dfrbp_1 _2356_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net36),
    .D(_0081_),
    .Q_N(_0775_),
    .Q(\latch_mem.addr_write[5] ));
 sg13g2_dfrbp_1 _2357_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net34),
    .D(_0082_),
    .Q_N(_0774_),
    .Q(\latch_mem.wr_en_next ));
 sg13g2_dfrbp_1 _2358_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net32),
    .D(_0083_),
    .Q_N(_0008_),
    .Q(\latch_mem.wr_en_valid ));
 sg13g2_dfrbp_1 _2359_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net30),
    .D(_0084_),
    .Q_N(_0017_),
    .Q(\cnt[3] ));
 sg13g2_dfrbp_1 _2360_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net25),
    .D(_0085_),
    .Q_N(_0019_),
    .Q(\cnt[2] ));
 sg13g2_dfrbp_1 _2361_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net21),
    .D(_0086_),
    .Q_N(_0773_),
    .Q(\cnt[1] ));
 sg13g2_dfrbp_1 _2362_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net28),
    .D(_0087_),
    .Q_N(_0772_),
    .Q(\cnt[0] ));
 sg13g2_dfrbp_1 _2363_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net19),
    .D(_0088_),
    .Q_N(_0771_),
    .Q(uo_out[6]));
 sg13g2_tiehi _1772__14 (.L_HI(net14));
 sg13g2_tiehi _1773__15 (.L_HI(net15));
 sg13g2_tiehi _1819__16 (.L_HI(net16));
 sg13g2_tiehi _1818__17 (.L_HI(net17));
 sg13g2_tiehi _1817__18 (.L_HI(net18));
 sg13g2_tiehi _2363__19 (.L_HI(net19));
 sg13g2_tiehi _1816__20 (.L_HI(net20));
 sg13g2_tiehi _2361__21 (.L_HI(net21));
 sg13g2_tiehi _1815__22 (.L_HI(net22));
 sg13g2_tiehi _2349__23 (.L_HI(net23));
 sg13g2_tiehi _1814__24 (.L_HI(net24));
 sg13g2_tiehi _2360__25 (.L_HI(net25));
 sg13g2_tiehi _1774__26 (.L_HI(net26));
 sg13g2_tiehi _1813__27 (.L_HI(net27));
 sg13g2_tiehi _2362__28 (.L_HI(net28));
 sg13g2_tiehi _1812__29 (.L_HI(net29));
 sg13g2_tiehi _2359__30 (.L_HI(net30));
 sg13g2_tiehi _1811__31 (.L_HI(net31));
 sg13g2_tiehi _2358__32 (.L_HI(net32));
 sg13g2_tiehi _1810__33 (.L_HI(net33));
 sg13g2_tiehi _2357__34 (.L_HI(net34));
 sg13g2_tiehi _1809__35 (.L_HI(net35));
 sg13g2_tiehi _2356__36 (.L_HI(net36));
 sg13g2_tiehi _1808__37 (.L_HI(net37));
 sg13g2_tiehi _2355__38 (.L_HI(net38));
 sg13g2_tiehi _1807__39 (.L_HI(net39));
 sg13g2_tiehi _2354__40 (.L_HI(net40));
 sg13g2_tiehi _1806__41 (.L_HI(net41));
 sg13g2_tiehi _2353__42 (.L_HI(net42));
 sg13g2_tiehi _1805__43 (.L_HI(net43));
 sg13g2_tiehi _2352__44 (.L_HI(net44));
 sg13g2_tiehi _1804__45 (.L_HI(net45));
 sg13g2_tiehi _2351__46 (.L_HI(net46));
 sg13g2_tiehi _1803__47 (.L_HI(net47));
 sg13g2_tiehi _1802__48 (.L_HI(net48));
 sg13g2_tiehi _2350__49 (.L_HI(net49));
 sg13g2_tiehi _1801__50 (.L_HI(net50));
 sg13g2_tiehi _2345__51 (.L_HI(net51));
 sg13g2_tiehi _1800__52 (.L_HI(net52));
 sg13g2_tiehi _1828__53 (.L_HI(net53));
 sg13g2_tiehi _1799__54 (.L_HI(net54));
 sg13g2_tiehi _1827__55 (.L_HI(net55));
 sg13g2_tiehi _1798__56 (.L_HI(net56));
 sg13g2_tiehi _1826__57 (.L_HI(net57));
 sg13g2_tiehi _1797__58 (.L_HI(net58));
 sg13g2_tiehi _1825__59 (.L_HI(net59));
 sg13g2_tiehi _1796__60 (.L_HI(net60));
 sg13g2_tiehi _1824__61 (.L_HI(net61));
 sg13g2_tiehi _1795__62 (.L_HI(net62));
 sg13g2_tiehi _1823__63 (.L_HI(net63));
 sg13g2_tiehi _1794__64 (.L_HI(net64));
 sg13g2_tiehi _1822__65 (.L_HI(net65));
 sg13g2_tiehi _1793__66 (.L_HI(net66));
 sg13g2_tiehi _1821__67 (.L_HI(net67));
 sg13g2_tiehi _1792__68 (.L_HI(net68));
 sg13g2_tiehi _1791__69 (.L_HI(net69));
 sg13g2_tiehi _1785__70 (.L_HI(net70));
 sg13g2_tiehi _1829__71 (.L_HI(net71));
 sg13g2_tiehi _2342__72 (.L_HI(net72));
 sg13g2_tiehi _2343__73 (.L_HI(net73));
 sg13g2_tiehi _1790__74 (.L_HI(net74));
 sg13g2_tiehi _2344__75 (.L_HI(net75));
 sg13g2_tiehi _2346__76 (.L_HI(net76));
 sg13g2_tiehi _2347__77 (.L_HI(net77));
 sg13g2_tiehi _2348__78 (.L_HI(net78));
 sg13g2_tiehi _1789__79 (.L_HI(net79));
 sg13g2_tiehi _1820__80 (.L_HI(net80));
 sg13g2_tiehi _1788__81 (.L_HI(net81));
 sg13g2_tiehi _1787__82 (.L_HI(net82));
 sg13g2_tiehi _1786__83 (.L_HI(net83));
 sg13g2_tiehi _1784__84 (.L_HI(net84));
 sg13g2_tiehi _1783__85 (.L_HI(net85));
 sg13g2_tiehi _1782__86 (.L_HI(net86));
 sg13g2_tiehi _1781__87 (.L_HI(net87));
 sg13g2_tiehi _1780__88 (.L_HI(net88));
 sg13g2_tiehi _1779__89 (.L_HI(net89));
 sg13g2_tiehi _1778__90 (.L_HI(net90));
 sg13g2_tiehi _1777__91 (.L_HI(net91));
 sg13g2_tiehi _1776__92 (.L_HI(net92));
 sg13g2_tiehi tt_um_branch_pred_93 (.L_HI(net93));
 sg13g2_tiehi tt_um_branch_pred_94 (.L_HI(net94));
 sg13g2_tiehi tt_um_branch_pred_95 (.L_HI(net95));
 sg13g2_tiehi tt_um_branch_pred_96 (.L_HI(net96));
 sg13g2_tiehi tt_um_branch_pred_97 (.L_HI(net97));
 sg13g2_inv_1 _1732__1 (.Y(net98),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_branch_pred_8 (.L_LO(net8));
 sg13g2_tielo tt_um_branch_pred_9 (.L_LO(net9));
 sg13g2_tielo tt_um_branch_pred_10 (.L_LO(net10));
 sg13g2_tielo tt_um_branch_pred_11 (.L_LO(net11));
 sg13g2_tielo tt_um_branch_pred_12 (.L_LO(net12));
 sg13g2_tiehi _1775__13 (.L_HI(net13));
 sg13g2_buf_1 _2455_ (.A(net1),
    .X(uio_out[2]));
 sg13g2_buf_1 _2456_ (.A(net2),
    .X(uio_out[3]));
 sg13g2_buf_1 _2457_ (.A(net3),
    .X(uio_out[4]));
 sg13g2_buf_1 _2458_ (.A(\latch_mem.wr_en_in ),
    .X(uio_out[5]));
 sg13g2_buf_2 _2459_ (.A(history_buffer_output),
    .X(uio_out[6]));
 sg13g2_buf_1 _2460_ (.A(pred_ready),
    .X(uo_out[0]));
 sg13g2_buf_2 _2461_ (.A(prediction),
    .X(uo_out[1]));
 sg13g2_buf_2 _2462_ (.A(training_done),
    .X(uo_out[2]));
 sg13g2_buf_1 _2463_ (.A(mem_reset_done),
    .X(uo_out[3]));
 sg13g2_buf_1 _2464_ (.A(new_data_avail_posedge),
    .X(uo_out[4]));
 sg13g2_buf_1 _2465_ (.A(state_rst_memory),
    .X(uo_out[7]));
 sg13g2_and2_2 \latch_mem.genblk1[0].lm_gate  (.A(net777),
    .B(\latch_mem.genblk1[0].sel_byte ),
    .X(\latch_mem.genblk1[0].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[10].lm_gate  (.A(net778),
    .B(\latch_mem.genblk1[10].sel_byte ),
    .X(\latch_mem.genblk1[10].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[11].lm_gate  (.A(net778),
    .B(\latch_mem.genblk1[11].sel_byte ),
    .X(\latch_mem.genblk1[11].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[12].lm_gate  (.A(net775),
    .B(\latch_mem.genblk1[12].sel_byte ),
    .X(\latch_mem.genblk1[12].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[13].lm_gate  (.A(net777),
    .B(\latch_mem.genblk1[13].sel_byte ),
    .X(\latch_mem.genblk1[13].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[14].lm_gate  (.A(net777),
    .B(\latch_mem.genblk1[14].sel_byte ),
    .X(\latch_mem.genblk1[14].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[15].lm_gate  (.A(net775),
    .B(\latch_mem.genblk1[15].sel_byte ),
    .X(\latch_mem.genblk1[15].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[16].lm_gate  (.A(net770),
    .B(\latch_mem.genblk1[16].sel_byte ),
    .X(\latch_mem.genblk1[16].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[17].lm_gate  (.A(net769),
    .B(\latch_mem.genblk1[17].sel_byte ),
    .X(\latch_mem.genblk1[17].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[18].lm_gate  (.A(net769),
    .B(\latch_mem.genblk1[18].sel_byte ),
    .X(\latch_mem.genblk1[18].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[19].lm_gate  (.A(net769),
    .B(\latch_mem.genblk1[19].sel_byte ),
    .X(\latch_mem.genblk1[19].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[1].lm_gate  (.A(net777),
    .B(\latch_mem.genblk1[1].sel_byte ),
    .X(\latch_mem.genblk1[1].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[20].lm_gate  (.A(net769),
    .B(\latch_mem.genblk1[20].sel_byte ),
    .X(\latch_mem.genblk1[20].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[21].lm_gate  (.A(net769),
    .B(\latch_mem.genblk1[21].sel_byte ),
    .X(\latch_mem.genblk1[21].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[22].lm_gate  (.A(net770),
    .B(\latch_mem.genblk1[22].sel_byte ),
    .X(\latch_mem.genblk1[22].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[23].lm_gate  (.A(net769),
    .B(\latch_mem.genblk1[23].sel_byte ),
    .X(\latch_mem.genblk1[23].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[24].lm_gate  (.A(net769),
    .B(\latch_mem.genblk1[24].sel_byte ),
    .X(\latch_mem.genblk1[24].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[25].lm_gate  (.A(net770),
    .B(\latch_mem.genblk1[25].sel_byte ),
    .X(\latch_mem.genblk1[25].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[26].lm_gate  (.A(net770),
    .B(\latch_mem.genblk1[26].sel_byte ),
    .X(\latch_mem.genblk1[26].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[27].lm_gate  (.A(net770),
    .B(\latch_mem.genblk1[27].sel_byte ),
    .X(\latch_mem.genblk1[27].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[28].lm_gate  (.A(net770),
    .B(\latch_mem.genblk1[28].sel_byte ),
    .X(\latch_mem.genblk1[28].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[29].lm_gate  (.A(net770),
    .B(\latch_mem.genblk1[29].sel_byte ),
    .X(\latch_mem.genblk1[29].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[2].lm_gate  (.A(net775),
    .B(\latch_mem.genblk1[2].sel_byte ),
    .X(\latch_mem.genblk1[2].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[30].lm_gate  (.A(net771),
    .B(\latch_mem.genblk1[30].sel_byte ),
    .X(\latch_mem.genblk1[30].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[31].lm_gate  (.A(net769),
    .B(\latch_mem.genblk1[31].sel_byte ),
    .X(\latch_mem.genblk1[31].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[32].lm_gate  (.A(net774),
    .B(\latch_mem.genblk1[32].sel_byte ),
    .X(\latch_mem.genblk1[32].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[33].lm_gate  (.A(net774),
    .B(\latch_mem.genblk1[33].sel_byte ),
    .X(\latch_mem.genblk1[33].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[34].lm_gate  (.A(net774),
    .B(\latch_mem.genblk1[34].sel_byte ),
    .X(\latch_mem.genblk1[34].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[35].lm_gate  (.A(net773),
    .B(\latch_mem.genblk1[35].sel_byte ),
    .X(\latch_mem.genblk1[35].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[36].lm_gate  (.A(net773),
    .B(\latch_mem.genblk1[36].sel_byte ),
    .X(\latch_mem.genblk1[36].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[37].lm_gate  (.A(net774),
    .B(\latch_mem.genblk1[37].sel_byte ),
    .X(\latch_mem.genblk1[37].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[38].lm_gate  (.A(net772),
    .B(\latch_mem.genblk1[38].sel_byte ),
    .X(\latch_mem.genblk1[38].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[39].lm_gate  (.A(net772),
    .B(\latch_mem.genblk1[39].sel_byte ),
    .X(\latch_mem.genblk1[39].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[3].lm_gate  (.A(net777),
    .B(\latch_mem.genblk1[3].sel_byte ),
    .X(\latch_mem.genblk1[3].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[40].lm_gate  (.A(net773),
    .B(\latch_mem.genblk1[40].sel_byte ),
    .X(\latch_mem.genblk1[40].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[41].lm_gate  (.A(net772),
    .B(\latch_mem.genblk1[41].sel_byte ),
    .X(\latch_mem.genblk1[41].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[42].lm_gate  (.A(net772),
    .B(\latch_mem.genblk1[42].sel_byte ),
    .X(\latch_mem.genblk1[42].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[43].lm_gate  (.A(net772),
    .B(\latch_mem.genblk1[43].sel_byte ),
    .X(\latch_mem.genblk1[43].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[44].lm_gate  (.A(net773),
    .B(\latch_mem.genblk1[44].sel_byte ),
    .X(\latch_mem.genblk1[44].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[45].lm_gate  (.A(net772),
    .B(\latch_mem.genblk1[45].sel_byte ),
    .X(\latch_mem.genblk1[45].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[46].lm_gate  (.A(net772),
    .B(\latch_mem.genblk1[46].sel_byte ),
    .X(\latch_mem.genblk1[46].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[47].lm_gate  (.A(net772),
    .B(\latch_mem.genblk1[47].sel_byte ),
    .X(\latch_mem.genblk1[47].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[48].lm_gate  (.A(net776),
    .B(\latch_mem.genblk1[48].sel_byte ),
    .X(\latch_mem.genblk1[48].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[49].lm_gate  (.A(net776),
    .B(\latch_mem.genblk1[49].sel_byte ),
    .X(\latch_mem.genblk1[49].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[4].lm_gate  (.A(net777),
    .B(\latch_mem.genblk1[4].sel_byte ),
    .X(\latch_mem.genblk1[4].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[50].lm_gate  (.A(net771),
    .B(\latch_mem.genblk1[50].sel_byte ),
    .X(\latch_mem.genblk1[50].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[51].lm_gate  (.A(net776),
    .B(\latch_mem.genblk1[51].sel_byte ),
    .X(\latch_mem.genblk1[51].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[52].lm_gate  (.A(net776),
    .B(\latch_mem.genblk1[52].sel_byte ),
    .X(\latch_mem.genblk1[52].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[53].lm_gate  (.A(net771),
    .B(\latch_mem.genblk1[53].sel_byte ),
    .X(\latch_mem.genblk1[53].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[54].lm_gate  (.A(net776),
    .B(\latch_mem.genblk1[54].sel_byte ),
    .X(\latch_mem.genblk1[54].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[55].lm_gate  (.A(net771),
    .B(\latch_mem.genblk1[55].sel_byte ),
    .X(\latch_mem.genblk1[55].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[56].lm_gate  (.A(net776),
    .B(\latch_mem.genblk1[56].sel_byte ),
    .X(\latch_mem.genblk1[56].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[57].lm_gate  (.A(net771),
    .B(\latch_mem.genblk1[57].sel_byte ),
    .X(\latch_mem.genblk1[57].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[58].lm_gate  (.A(net778),
    .B(\latch_mem.genblk1[58].sel_byte ),
    .X(\latch_mem.genblk1[58].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[59].lm_gate  (.A(net778),
    .B(\latch_mem.genblk1[59].sel_byte ),
    .X(\latch_mem.genblk1[59].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[5].lm_gate  (.A(net775),
    .B(\latch_mem.genblk1[5].sel_byte ),
    .X(\latch_mem.genblk1[5].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[60].lm_gate  (.A(net771),
    .B(\latch_mem.genblk1[60].sel_byte ),
    .X(\latch_mem.genblk1[60].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[61].lm_gate  (.A(net776),
    .B(\latch_mem.genblk1[61].sel_byte ),
    .X(\latch_mem.genblk1[61].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[62].lm_gate  (.A(net776),
    .B(\latch_mem.genblk1[62].sel_byte ),
    .X(\latch_mem.genblk1[62].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[63].lm_gate  (.A(net771),
    .B(\latch_mem.genblk1[63].sel_byte ),
    .X(\latch_mem.genblk1[63].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[6].lm_gate  (.A(net777),
    .B(\latch_mem.genblk1[6].sel_byte ),
    .X(\latch_mem.genblk1[6].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[7].lm_gate  (.A(net775),
    .B(\latch_mem.genblk1[7].sel_byte ),
    .X(\latch_mem.genblk1[7].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[8].lm_gate  (.A(net777),
    .B(\latch_mem.genblk1[8].sel_byte ),
    .X(\latch_mem.genblk1[8].wr_en_this_byte ));
 sg13g2_and2_2 \latch_mem.genblk1[9].lm_gate  (.A(net775),
    .B(\latch_mem.genblk1[9].sel_byte ),
    .X(\latch_mem.genblk1[9].wr_en_this_byte ));
 sg13g2_ebufn_8 \latch_mem.genblk2[0].lm_dt_out_buf[0]  (.Z(\latch_mem.combined_out[0] ),
    .A(\latch_mem.genblk2[0].selected_out[0] ),
    .TE_B(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[0].lm_dt_out_buf[1]  (.Z(\latch_mem.combined_out[1] ),
    .A(\latch_mem.genblk2[0].selected_out[1] ),
    .TE_B(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[0].lm_dt_out_buf[2]  (.Z(\latch_mem.combined_out[2] ),
    .A(\latch_mem.genblk2[0].selected_out[2] ),
    .TE_B(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[0].lm_dt_out_buf[3]  (.Z(\latch_mem.combined_out[3] ),
    .A(\latch_mem.genblk2[0].selected_out[3] ),
    .TE_B(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[0].lm_dt_out_buf[4]  (.Z(\latch_mem.combined_out[4] ),
    .A(\latch_mem.genblk2[0].selected_out[4] ),
    .TE_B(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[0].lm_dt_out_buf[5]  (.Z(\latch_mem.combined_out[5] ),
    .A(\latch_mem.genblk2[0].selected_out[5] ),
    .TE_B(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[0].lm_dt_out_buf[6]  (.Z(\latch_mem.combined_out[6] ),
    .A(\latch_mem.genblk2[0].selected_out[6] ),
    .TE_B(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[0].lm_dt_out_buf[7]  (.Z(\latch_mem.combined_out[7] ),
    .A(\latch_mem.genblk2[0].selected_out[7] ),
    .TE_B(\latch_mem.genblk2[0].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[1].lm_dt_out_buf[0]  (.Z(\latch_mem.combined_out[0] ),
    .A(\latch_mem.genblk2[1].selected_out[0] ),
    .TE_B(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[1].lm_dt_out_buf[1]  (.Z(\latch_mem.combined_out[1] ),
    .A(\latch_mem.genblk2[1].selected_out[1] ),
    .TE_B(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[1].lm_dt_out_buf[2]  (.Z(\latch_mem.combined_out[2] ),
    .A(\latch_mem.genblk2[1].selected_out[2] ),
    .TE_B(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[1].lm_dt_out_buf[3]  (.Z(\latch_mem.combined_out[3] ),
    .A(\latch_mem.genblk2[1].selected_out[3] ),
    .TE_B(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[1].lm_dt_out_buf[4]  (.Z(\latch_mem.combined_out[4] ),
    .A(\latch_mem.genblk2[1].selected_out[4] ),
    .TE_B(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[1].lm_dt_out_buf[5]  (.Z(\latch_mem.combined_out[5] ),
    .A(\latch_mem.genblk2[1].selected_out[5] ),
    .TE_B(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[1].lm_dt_out_buf[6]  (.Z(\latch_mem.combined_out[6] ),
    .A(\latch_mem.genblk2[1].selected_out[6] ),
    .TE_B(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[1].lm_dt_out_buf[7]  (.Z(\latch_mem.combined_out[7] ),
    .A(\latch_mem.genblk2[1].selected_out[7] ),
    .TE_B(\latch_mem.genblk2[1].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[2].lm_dt_out_buf[0]  (.Z(\latch_mem.combined_out[0] ),
    .A(\latch_mem.genblk2[2].selected_out[0] ),
    .TE_B(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[2].lm_dt_out_buf[1]  (.Z(\latch_mem.combined_out[1] ),
    .A(\latch_mem.genblk2[2].selected_out[1] ),
    .TE_B(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[2].lm_dt_out_buf[2]  (.Z(\latch_mem.combined_out[2] ),
    .A(\latch_mem.genblk2[2].selected_out[2] ),
    .TE_B(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[2].lm_dt_out_buf[3]  (.Z(\latch_mem.combined_out[3] ),
    .A(\latch_mem.genblk2[2].selected_out[3] ),
    .TE_B(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[2].lm_dt_out_buf[4]  (.Z(\latch_mem.combined_out[4] ),
    .A(\latch_mem.genblk2[2].selected_out[4] ),
    .TE_B(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[2].lm_dt_out_buf[5]  (.Z(\latch_mem.combined_out[5] ),
    .A(\latch_mem.genblk2[2].selected_out[5] ),
    .TE_B(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[2].lm_dt_out_buf[6]  (.Z(\latch_mem.combined_out[6] ),
    .A(\latch_mem.genblk2[2].selected_out[6] ),
    .TE_B(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[2].lm_dt_out_buf[7]  (.Z(\latch_mem.combined_out[7] ),
    .A(\latch_mem.genblk2[2].selected_out[7] ),
    .TE_B(\latch_mem.genblk2[2].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[3].lm_dt_out_buf[0]  (.Z(\latch_mem.combined_out[0] ),
    .A(\latch_mem.genblk2[3].selected_out[0] ),
    .TE_B(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[3].lm_dt_out_buf[1]  (.Z(\latch_mem.combined_out[1] ),
    .A(\latch_mem.genblk2[3].selected_out[1] ),
    .TE_B(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[3].lm_dt_out_buf[2]  (.Z(\latch_mem.combined_out[2] ),
    .A(\latch_mem.genblk2[3].selected_out[2] ),
    .TE_B(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[3].lm_dt_out_buf[3]  (.Z(\latch_mem.combined_out[3] ),
    .A(\latch_mem.genblk2[3].selected_out[3] ),
    .TE_B(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[3].lm_dt_out_buf[4]  (.Z(\latch_mem.combined_out[4] ),
    .A(\latch_mem.genblk2[3].selected_out[4] ),
    .TE_B(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[3].lm_dt_out_buf[5]  (.Z(\latch_mem.combined_out[5] ),
    .A(\latch_mem.genblk2[3].selected_out[5] ),
    .TE_B(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[3].lm_dt_out_buf[6]  (.Z(\latch_mem.combined_out[6] ),
    .A(\latch_mem.genblk2[3].selected_out[6] ),
    .TE_B(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_ebufn_8 \latch_mem.genblk2[3].lm_dt_out_buf[7]  (.Z(\latch_mem.combined_out[7] ),
    .A(\latch_mem.genblk2[3].selected_out[7] ),
    .TE_B(\latch_mem.genblk2[3].partition_sel_n ));
 sg13g2_buf_4 \latch_mem.lm_dt_final_buf[0]  (.X(\latch_mem.uo_out[0] ),
    .A(\latch_mem.combined_out[0] ));
 sg13g2_buf_4 \latch_mem.lm_dt_final_buf[1]  (.X(\latch_mem.uo_out[1] ),
    .A(\latch_mem.combined_out[1] ));
 sg13g2_buf_2 \latch_mem.lm_dt_final_buf[2]  (.A(\latch_mem.combined_out[2] ),
    .X(\latch_mem.uo_out[2] ));
 sg13g2_buf_2 \latch_mem.lm_dt_final_buf[3]  (.A(\latch_mem.combined_out[3] ),
    .X(\latch_mem.uo_out[3] ));
 sg13g2_buf_2 \latch_mem.lm_dt_final_buf[4]  (.A(\latch_mem.combined_out[4] ),
    .X(\latch_mem.uo_out[4] ));
 sg13g2_buf_2 \latch_mem.lm_dt_final_buf[5]  (.A(\latch_mem.combined_out[5] ),
    .X(\latch_mem.uo_out[5] ));
 sg13g2_buf_2 \latch_mem.lm_dt_final_buf[6]  (.A(\latch_mem.combined_out[6] ),
    .X(\latch_mem.uo_out[6] ));
 sg13g2_buf_4 \latch_mem.lm_dt_final_buf[7]  (.X(\latch_mem.uo_out[7] ),
    .A(\latch_mem.combined_out[7] ));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_1 fanout687 (.A(_0506_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_0547_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_0546_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_0448_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_0550_),
    .X(net693));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(net698));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(net698));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(net698));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(net698));
 sg13g2_buf_2 fanout698 (.A(_0751_),
    .X(net698));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(net703));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(net703));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(net703));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(net703));
 sg13g2_buf_2 fanout703 (.A(_0750_),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(net706));
 sg13g2_buf_2 fanout705 (.A(net706),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(_0749_));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(_0749_));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(_0749_));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(net713));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(net713));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(net713));
 sg13g2_buf_4 fanout712 (.X(net712),
    .A(net713));
 sg13g2_buf_2 fanout713 (.A(_0748_),
    .X(net713));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(net715));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(_0747_));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(net718));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_0747_),
    .X(net718));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(net723));
 sg13g2_buf_4 fanout720 (.X(net720),
    .A(net723));
 sg13g2_buf_4 fanout721 (.X(net721),
    .A(net723));
 sg13g2_buf_4 fanout722 (.X(net722),
    .A(net723));
 sg13g2_buf_2 fanout723 (.A(_0746_),
    .X(net723));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(net728));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(net728));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(net727));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(net728));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(_0744_));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net730));
 sg13g2_buf_4 fanout730 (.X(net730),
    .A(net733));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(net732));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(net733));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(_0743_));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(net735));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(net738));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(net737));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net738));
 sg13g2_buf_4 fanout738 (.X(net738),
    .A(_0742_));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(net740));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net743));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net742));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(net743));
 sg13g2_buf_2 fanout743 (.A(_0741_),
    .X(net743));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(net746));
 sg13g2_buf_2 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_0739_),
    .X(net746));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(net748));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(_0739_));
 sg13g2_buf_4 fanout749 (.X(net749),
    .A(net751));
 sg13g2_buf_2 fanout750 (.A(net751),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_0738_),
    .X(net751));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(net753));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(_0738_));
 sg13g2_buf_4 fanout754 (.X(net754),
    .A(net756));
 sg13g2_buf_2 fanout755 (.A(net756),
    .X(net755));
 sg13g2_buf_4 fanout756 (.X(net756),
    .A(_0736_));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(net758));
 sg13g2_buf_4 fanout758 (.X(net758),
    .A(_0736_));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(net760));
 sg13g2_buf_4 fanout760 (.X(net760),
    .A(net763));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(net762));
 sg13g2_buf_4 fanout762 (.X(net762),
    .A(net763));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(_0733_));
 sg13g2_buf_4 fanout764 (.X(net764),
    .A(net765));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(net768));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(net768));
 sg13g2_buf_4 fanout767 (.X(net767),
    .A(net768));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(_0730_));
 sg13g2_buf_2 fanout769 (.A(net770),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(\latch_mem.wr_en ),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(net774),
    .X(net772));
 sg13g2_buf_1 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_1 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(\latch_mem.wr_en ),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(net778),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(\latch_mem.wr_en ),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(net780));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(_0389_));
 sg13g2_buf_4 fanout781 (.X(net781),
    .A(_0389_));
 sg13g2_buf_4 fanout782 (.X(net782),
    .A(net787));
 sg13g2_buf_4 fanout783 (.X(net783),
    .A(net787));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(net785));
 sg13g2_buf_2 fanout785 (.A(net787),
    .X(net785));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(net787));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(_0731_));
 sg13g2_buf_2 fanout788 (.A(_0728_),
    .X(net788));
 sg13g2_buf_1 fanout789 (.A(_0728_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_0726_),
    .X(net790));
 sg13g2_buf_1 fanout791 (.A(_0726_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_1 fanout793 (.A(_0724_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_0702_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(uo_out[6]),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(net176),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(net799),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(\cnt[1] ),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(net139),
    .X(net800));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(net129));
 sg13g2_buf_2 fanout802 (.A(net129),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(\latch_mem.addr_write[3] ),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(net183),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(net187),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(uo_out[5]),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net810),
    .X(net809));
 sg13g2_buf_1 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_1 fanout811 (.A(net122),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(net816),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(net816),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(net816),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(\latch_mem.data_to_write[7] ));
 sg13g2_buf_2 fanout817 (.A(net818),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net821),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(net821),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(\latch_mem.data_to_write[7] ));
 sg13g2_buf_2 fanout822 (.A(net826),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net826),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(net826),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(\latch_mem.data_to_write[6] ));
 sg13g2_buf_2 fanout827 (.A(net831),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(net831),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(net831),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(net831),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(\latch_mem.data_to_write[6] ),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net836),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(net835),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(net836),
    .X(net835));
 sg13g2_buf_1 fanout836 (.A(\latch_mem.data_to_write[5] ),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(net838),
    .X(net837));
 sg13g2_buf_4 fanout838 (.X(net838),
    .A(net841));
 sg13g2_buf_2 fanout839 (.A(net840),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(\latch_mem.data_to_write[5] ));
 sg13g2_buf_2 fanout842 (.A(net846),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net846),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net846),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(\latch_mem.data_to_write[4] ),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(net848),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(\latch_mem.data_to_write[4] ),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(\latch_mem.data_to_write[4] ),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_1 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_1 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(net858),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(net858),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(net858),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(net863),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net863),
    .X(net860));
 sg13g2_buf_4 fanout861 (.X(net861),
    .A(net863));
 sg13g2_buf_2 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(\latch_mem.data_to_write[3] ));
 sg13g2_buf_2 fanout864 (.A(net868),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(net868),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net868),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net868),
    .X(net867));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(\latch_mem.data_to_write[2] ));
 sg13g2_buf_2 fanout869 (.A(net873),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(net873),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(net872),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(\latch_mem.data_to_write[2] ),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net878),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net878),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net878),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(\latch_mem.data_to_write[1] ),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(net880),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(net883),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net883),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(net883),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(\latch_mem.data_to_write[1] ),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(net886),
    .X(net884));
 sg13g2_buf_1 fanout885 (.A(net886),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(net894),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net894),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net894),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net893),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net893),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(net893),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(net893),
    .X(net892));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net894));
 sg13g2_buf_4 fanout894 (.X(net894),
    .A(\latch_mem.data_to_write[0] ));
 sg13g2_buf_2 fanout895 (.A(rst_n),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(rst_n),
    .X(net896));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(net898));
 sg13g2_buf_1 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(rst_n),
    .X(net899));
 sg13g2_buf_2 input1 (.A(ui_in[2]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_4 input5 (.X(net5),
    .A(uio_in[1]));
 sg13g2_buf_2 input6 (.A(uio_in[7]),
    .X(net6));
 sg13g2_tielo tt_um_branch_pred_7 (.L_LO(net7));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(delaynet_1_clk));
 sg13g2_buf_2 delaybuf_1_clk (.A(delaynet_1_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0020_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0073_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold3 (.A(\latch_mem.addr_in[3] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold4 (.A(\latch_mem.addr_in[2] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0011_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0000_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold7 (.A(\substate[3] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0689_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold9 (.A(\latch_mem.addr_in[1] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold10 (.A(\latch_mem.uio_in[7] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0021_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0035_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold13 (.A(\latch_mem.uio_in[2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold14 (.A(\latch_mem.wr_en_next ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold15 (.A(\latch_mem.uio_in[6] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold16 (.A(\substate[1] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0700_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold18 (.A(pred_ready),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold19 (.A(mem_reset_done),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0442_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0038_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold22 (.A(\latch_mem.uio_in[4] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold23 (.A(\latch_mem.uio_in[1] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold24 (.A(training_done),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold25 (.A(\latch_mem.addr_in[0] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold26 (.A(\latch_mem.uio_in[3] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold27 (.A(\substate[2] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0699_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0009_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0509_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cnt[3] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold32 (.A(\latch_mem.addr_in[4] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0006_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold34 (.A(\latch_mem.addr_in[5] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold35 (.A(\history_buffer[6] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0062_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold37 (.A(\history_buffer_index[1] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0614_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0074_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold40 (.A(\latch_mem.uio_in[0] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cnt[2] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold42 (.A(\history_buffer_index[2] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0615_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0075_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold45 (.A(history_buffer_request_prev),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0390_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0032_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold48 (.A(\latch_mem.wr_en_in ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold49 (.A(\latch_mem.uio_in[5] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold50 (.A(\history_buffer[3] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0059_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold52 (.A(\abs_sum[0] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold53 (.A(\history_buffer[2] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0057_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold55 (.A(\sum[8] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold56 (.A(\history_buffer[0] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0056_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold58 (.A(\history_buffer[5] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold59 (.A(\sum[7] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold60 (.A(\sum[1] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold61 (.A(\history_buffer[4] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold62 (.A(\sum[4] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold63 (.A(\history_buffer[7] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0402_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0403_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0404_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold67 (.A(\sum[3] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold68 (.A(\latch_mem.addr_write[3] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold69 (.A(state_rst_memory),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold70 (.A(\sum[2] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold71 (.A(\latch_mem.addr_in[1] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0514_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0010_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold74 (.A(\sum[9] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0017_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold76 (.A(\sum[5] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold77 (.A(\sum[6] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cnt[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold79 (.A(\latch_mem.addr_in[0] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold80 (.A(\latch_mem.addr_write[5] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0019_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold82 (.A(\latch_mem.addr_in[4] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold83 (.A(\latch_mem.addr_write[4] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold84 (.A(\latch_mem.addr_write[1] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold85 (.A(\latch_mem.addr_write[2] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0012_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0017_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold88 (.A(\latch_mem.addr_write[0] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold89 (.A(state_rst_memory),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0019_),
    .X(net188));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_fill_2 FILLER_0_175 ();
 sg13g2_fill_1 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_195 ();
 sg13g2_decap_8 FILLER_0_202 ();
 sg13g2_decap_8 FILLER_0_209 ();
 sg13g2_decap_8 FILLER_0_216 ();
 sg13g2_decap_8 FILLER_0_223 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_decap_8 FILLER_0_237 ();
 sg13g2_decap_8 FILLER_0_244 ();
 sg13g2_decap_8 FILLER_0_251 ();
 sg13g2_decap_8 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_272 ();
 sg13g2_decap_8 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_321 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_4 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_fill_1 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_227 ();
 sg13g2_fill_1 FILLER_1_234 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_4 FILLER_1_294 ();
 sg13g2_fill_2 FILLER_1_298 ();
 sg13g2_fill_1 FILLER_1_306 ();
 sg13g2_fill_2 FILLER_1_324 ();
 sg13g2_fill_2 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_fill_2 FILLER_2_235 ();
 sg13g2_fill_1 FILLER_2_237 ();
 sg13g2_decap_8 FILLER_2_255 ();
 sg13g2_decap_8 FILLER_2_262 ();
 sg13g2_decap_8 FILLER_2_269 ();
 sg13g2_decap_8 FILLER_2_276 ();
 sg13g2_decap_8 FILLER_2_283 ();
 sg13g2_fill_1 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_fill_1 FILLER_3_216 ();
 sg13g2_fill_1 FILLER_3_234 ();
 sg13g2_decap_4 FILLER_3_252 ();
 sg13g2_fill_1 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_fill_1 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_4 FILLER_4_168 ();
 sg13g2_decap_4 FILLER_4_183 ();
 sg13g2_decap_4 FILLER_4_222 ();
 sg13g2_fill_1 FILLER_4_226 ();
 sg13g2_decap_4 FILLER_4_233 ();
 sg13g2_fill_2 FILLER_4_254 ();
 sg13g2_fill_1 FILLER_4_313 ();
 sg13g2_fill_2 FILLER_4_332 ();
 sg13g2_decap_4 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_4 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_197 ();
 sg13g2_fill_2 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_212 ();
 sg13g2_fill_2 FILLER_5_219 ();
 sg13g2_decap_8 FILLER_5_227 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_decap_8 FILLER_5_241 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_fill_1 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_4 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_fill_2 FILLER_6_154 ();
 sg13g2_fill_2 FILLER_6_213 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_251 ();
 sg13g2_decap_8 FILLER_6_258 ();
 sg13g2_decap_8 FILLER_6_265 ();
 sg13g2_decap_8 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_fill_2 FILLER_6_304 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_1 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_fill_2 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_154 ();
 sg13g2_fill_1 FILLER_7_173 ();
 sg13g2_fill_2 FILLER_7_180 ();
 sg13g2_decap_8 FILLER_7_188 ();
 sg13g2_fill_2 FILLER_7_195 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_fill_2 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_265 ();
 sg13g2_fill_2 FILLER_7_272 ();
 sg13g2_fill_2 FILLER_7_305 ();
 sg13g2_fill_2 FILLER_7_324 ();
 sg13g2_fill_1 FILLER_7_326 ();
 sg13g2_fill_2 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_154 ();
 sg13g2_decap_4 FILLER_8_195 ();
 sg13g2_fill_2 FILLER_8_199 ();
 sg13g2_decap_8 FILLER_8_218 ();
 sg13g2_fill_2 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_233 ();
 sg13g2_decap_4 FILLER_8_281 ();
 sg13g2_fill_1 FILLER_8_285 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_fill_1 FILLER_9_195 ();
 sg13g2_fill_1 FILLER_9_200 ();
 sg13g2_fill_1 FILLER_9_236 ();
 sg13g2_decap_4 FILLER_9_254 ();
 sg13g2_fill_2 FILLER_9_258 ();
 sg13g2_decap_4 FILLER_9_317 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_fill_2 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_4 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_178 ();
 sg13g2_decap_4 FILLER_10_185 ();
 sg13g2_fill_1 FILLER_10_189 ();
 sg13g2_fill_2 FILLER_10_207 ();
 sg13g2_fill_1 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_4 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_285 ();
 sg13g2_decap_4 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_fill_2 FILLER_10_333 ();
 sg13g2_fill_1 FILLER_10_335 ();
 sg13g2_decap_4 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_190 ();
 sg13g2_fill_1 FILLER_11_208 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_250 ();
 sg13g2_fill_1 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_fill_2 FILLER_11_287 ();
 sg13g2_decap_4 FILLER_11_294 ();
 sg13g2_fill_1 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_316 ();
 sg13g2_fill_1 FILLER_11_350 ();
 sg13g2_fill_2 FILLER_11_368 ();
 sg13g2_fill_1 FILLER_11_370 ();
 sg13g2_decap_4 FILLER_11_376 ();
 sg13g2_fill_1 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_4 FILLER_12_133 ();
 sg13g2_fill_1 FILLER_12_137 ();
 sg13g2_fill_2 FILLER_12_172 ();
 sg13g2_fill_1 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_205 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_274 ();
 sg13g2_fill_1 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_325 ();
 sg13g2_fill_2 FILLER_12_350 ();
 sg13g2_decap_4 FILLER_12_358 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_fill_1 FILLER_12_375 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_191 ();
 sg13g2_decap_8 FILLER_13_209 ();
 sg13g2_decap_8 FILLER_13_216 ();
 sg13g2_decap_4 FILLER_13_223 ();
 sg13g2_decap_4 FILLER_13_249 ();
 sg13g2_decap_4 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_308 ();
 sg13g2_decap_4 FILLER_13_332 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_decap_4 FILLER_13_354 ();
 sg13g2_fill_1 FILLER_13_358 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_4 FILLER_14_171 ();
 sg13g2_fill_1 FILLER_14_175 ();
 sg13g2_decap_4 FILLER_14_182 ();
 sg13g2_fill_2 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_223 ();
 sg13g2_decap_4 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_decap_4 FILLER_14_269 ();
 sg13g2_decap_4 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_290 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_387 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_4 FILLER_15_154 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_183 ();
 sg13g2_decap_8 FILLER_15_190 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_236 ();
 sg13g2_decap_4 FILLER_15_243 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_fill_2 FILLER_15_260 ();
 sg13g2_decap_4 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_decap_4 FILLER_15_379 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_4 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_202 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_4 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_4 FILLER_16_346 ();
 sg13g2_fill_1 FILLER_16_350 ();
 sg13g2_decap_4 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_4 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_decap_4 FILLER_18_183 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_decap_4 FILLER_18_237 ();
 sg13g2_fill_2 FILLER_18_258 ();
 sg13g2_decap_4 FILLER_18_302 ();
 sg13g2_fill_2 FILLER_18_306 ();
 sg13g2_decap_4 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_368 ();
 sg13g2_decap_4 FILLER_18_374 ();
 sg13g2_fill_1 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_158 ();
 sg13g2_decap_4 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_224 ();
 sg13g2_decap_4 FILLER_19_238 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_fill_2 FILLER_19_327 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_decap_4 FILLER_19_364 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_4 FILLER_20_171 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_243 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_fill_1 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_244 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_4 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_fill_2 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_4 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_387 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_fill_2 FILLER_22_179 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_decap_4 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_250 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_fill_2 FILLER_22_284 ();
 sg13g2_fill_1 FILLER_22_286 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_317 ();
 sg13g2_decap_4 FILLER_22_324 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_decap_4 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_4 FILLER_22_370 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_decap_4 FILLER_22_392 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_4 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_170 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_192 ();
 sg13g2_decap_4 FILLER_23_200 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_decap_8 FILLER_23_216 ();
 sg13g2_decap_4 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_decap_4 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_decap_4 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_decap_8 FILLER_24_185 ();
 sg13g2_decap_8 FILLER_24_192 ();
 sg13g2_decap_8 FILLER_24_199 ();
 sg13g2_decap_4 FILLER_24_206 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_218 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_293 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_238 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_decap_4 FILLER_25_278 ();
 sg13g2_decap_8 FILLER_25_306 ();
 sg13g2_decap_4 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_4 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_151 ();
 sg13g2_decap_4 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_decap_8 FILLER_26_215 ();
 sg13g2_decap_8 FILLER_26_222 ();
 sg13g2_decap_8 FILLER_26_229 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_decap_4 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_decap_4 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_fill_2 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_2 FILLER_27_151 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_283 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_27_313 ();
 sg13g2_decap_8 FILLER_27_320 ();
 sg13g2_decap_8 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_334 ();
 sg13g2_decap_8 FILLER_27_341 ();
 sg13g2_fill_2 FILLER_27_348 ();
 sg13g2_fill_2 FILLER_27_373 ();
 sg13g2_fill_1 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_fill_2 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_fill_2 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_decap_4 FILLER_28_339 ();
 sg13g2_fill_2 FILLER_28_343 ();
 sg13g2_fill_2 FILLER_28_384 ();
 sg13g2_fill_1 FILLER_28_386 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_decap_4 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_decap_4 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_182 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_249 ();
 sg13g2_fill_2 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_276 ();
 sg13g2_fill_2 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_298 ();
 sg13g2_decap_4 FILLER_30_305 ();
 sg13g2_decap_4 FILLER_30_332 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_283 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_decap_4 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_363 ();
 sg13g2_fill_1 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_decap_4 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_376 ();
 sg13g2_decap_4 FILLER_32_382 ();
 sg13g2_fill_2 FILLER_32_386 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_132 ();
 sg13g2_decap_8 FILLER_33_139 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_4 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_286 ();
 sg13g2_fill_1 FILLER_33_288 ();
 sg13g2_decap_4 FILLER_33_334 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_386 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_137 ();
 sg13g2_fill_2 FILLER_34_142 ();
 sg13g2_decap_8 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_decap_4 FILLER_34_162 ();
 sg13g2_decap_8 FILLER_34_216 ();
 sg13g2_decap_8 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_251 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_290 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_309 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_4 FILLER_35_70 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_decap_4 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_decap_4 FILLER_35_191 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_decap_4 FILLER_35_327 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_fill_2 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_95 ();
 sg13g2_fill_2 FILLER_36_123 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_188 ();
 sg13g2_decap_4 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_decap_4 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_298 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_fill_2 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_decap_4 FILLER_36_340 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_4 FILLER_37_185 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_290 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_306 ();
 sg13g2_decap_8 FILLER_37_313 ();
 sg13g2_decap_8 FILLER_37_320 ();
 sg13g2_decap_8 FILLER_37_327 ();
 sg13g2_decap_4 FILLER_37_334 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_fill_2 FILLER_37_374 ();
 sg13g2_fill_1 FILLER_37_376 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_74 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_fill_2 FILLER_38_111 ();
 sg13g2_fill_1 FILLER_38_113 ();
 sg13g2_decap_8 FILLER_38_159 ();
 sg13g2_decap_4 FILLER_38_166 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_4 FILLER_38_186 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_2 FILLER_38_238 ();
 sg13g2_fill_1 FILLER_38_240 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_331 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_342 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_decap_8 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_370 ();
 sg13g2_decap_4 FILLER_38_377 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_fill_1 FILLER_39_70 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_fill_2 FILLER_39_108 ();
 sg13g2_fill_2 FILLER_39_131 ();
 sg13g2_decap_8 FILLER_39_164 ();
 sg13g2_fill_2 FILLER_39_171 ();
 sg13g2_fill_1 FILLER_39_173 ();
 sg13g2_decap_8 FILLER_39_191 ();
 sg13g2_decap_4 FILLER_39_198 ();
 sg13g2_fill_2 FILLER_39_202 ();
 sg13g2_decap_8 FILLER_39_226 ();
 sg13g2_decap_4 FILLER_39_233 ();
 sg13g2_fill_1 FILLER_39_258 ();
 sg13g2_fill_2 FILLER_39_264 ();
 sg13g2_fill_1 FILLER_39_266 ();
 sg13g2_decap_4 FILLER_39_277 ();
 sg13g2_fill_1 FILLER_39_281 ();
 sg13g2_fill_2 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_fill_2 FILLER_39_406 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_fill_1 FILLER_40_107 ();
 sg13g2_decap_4 FILLER_40_165 ();
 sg13g2_fill_1 FILLER_40_174 ();
 sg13g2_decap_4 FILLER_40_198 ();
 sg13g2_fill_2 FILLER_40_208 ();
 sg13g2_decap_8 FILLER_40_233 ();
 sg13g2_fill_2 FILLER_40_240 ();
 sg13g2_fill_1 FILLER_40_242 ();
 sg13g2_decap_8 FILLER_40_277 ();
 sg13g2_fill_2 FILLER_40_284 ();
 sg13g2_decap_8 FILLER_40_302 ();
 sg13g2_fill_2 FILLER_40_309 ();
 sg13g2_fill_1 FILLER_40_311 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_4 FILLER_41_56 ();
 sg13g2_fill_1 FILLER_41_82 ();
 sg13g2_fill_2 FILLER_41_99 ();
 sg13g2_fill_1 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_128 ();
 sg13g2_decap_8 FILLER_41_229 ();
 sg13g2_decap_4 FILLER_41_236 ();
 sg13g2_decap_4 FILLER_41_271 ();
 sg13g2_fill_2 FILLER_41_275 ();
 sg13g2_fill_2 FILLER_41_281 ();
 sg13g2_fill_2 FILLER_41_302 ();
 sg13g2_decap_4 FILLER_41_351 ();
 sg13g2_decap_8 FILLER_41_389 ();
 sg13g2_decap_8 FILLER_41_396 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_fill_2 FILLER_42_56 ();
 sg13g2_fill_1 FILLER_42_58 ();
 sg13g2_fill_1 FILLER_42_102 ();
 sg13g2_decap_4 FILLER_42_132 ();
 sg13g2_decap_4 FILLER_42_148 ();
 sg13g2_fill_1 FILLER_42_152 ();
 sg13g2_fill_2 FILLER_42_167 ();
 sg13g2_fill_1 FILLER_42_169 ();
 sg13g2_fill_1 FILLER_42_254 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_fill_2 FILLER_42_266 ();
 sg13g2_fill_2 FILLER_42_276 ();
 sg13g2_fill_1 FILLER_42_283 ();
 sg13g2_decap_8 FILLER_42_317 ();
 sg13g2_fill_2 FILLER_42_324 ();
 sg13g2_fill_2 FILLER_42_337 ();
 sg13g2_decap_8 FILLER_42_395 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_4 FILLER_43_49 ();
 sg13g2_fill_1 FILLER_43_53 ();
 sg13g2_decap_8 FILLER_43_58 ();
 sg13g2_decap_4 FILLER_43_65 ();
 sg13g2_fill_1 FILLER_43_69 ();
 sg13g2_fill_2 FILLER_43_74 ();
 sg13g2_fill_1 FILLER_43_76 ();
 sg13g2_fill_2 FILLER_43_95 ();
 sg13g2_fill_2 FILLER_43_109 ();
 sg13g2_decap_8 FILLER_43_120 ();
 sg13g2_decap_4 FILLER_43_127 ();
 sg13g2_decap_8 FILLER_43_141 ();
 sg13g2_decap_4 FILLER_43_148 ();
 sg13g2_fill_2 FILLER_43_152 ();
 sg13g2_fill_1 FILLER_43_194 ();
 sg13g2_fill_2 FILLER_43_201 ();
 sg13g2_fill_1 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_fill_1 FILLER_43_217 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_4 FILLER_43_238 ();
 sg13g2_fill_2 FILLER_43_257 ();
 sg13g2_fill_1 FILLER_43_259 ();
 sg13g2_decap_4 FILLER_43_269 ();
 sg13g2_fill_2 FILLER_43_273 ();
 sg13g2_fill_2 FILLER_43_285 ();
 sg13g2_decap_8 FILLER_43_326 ();
 sg13g2_decap_8 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_340 ();
 sg13g2_decap_8 FILLER_43_347 ();
 sg13g2_decap_4 FILLER_43_354 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_decap_4 FILLER_43_365 ();
 sg13g2_fill_2 FILLER_43_374 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_4 FILLER_44_35 ();
 sg13g2_fill_1 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_114 ();
 sg13g2_decap_4 FILLER_44_121 ();
 sg13g2_fill_1 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_131 ();
 sg13g2_decap_4 FILLER_44_137 ();
 sg13g2_decap_8 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_201 ();
 sg13g2_decap_8 FILLER_44_208 ();
 sg13g2_decap_8 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_decap_8 FILLER_44_229 ();
 sg13g2_decap_4 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_240 ();
 sg13g2_fill_2 FILLER_44_277 ();
 sg13g2_fill_1 FILLER_44_279 ();
 sg13g2_decap_4 FILLER_44_301 ();
 sg13g2_fill_1 FILLER_44_305 ();
 sg13g2_fill_1 FILLER_44_323 ();
 sg13g2_decap_4 FILLER_44_341 ();
 sg13g2_fill_1 FILLER_44_345 ();
 sg13g2_decap_8 FILLER_44_351 ();
 sg13g2_decap_8 FILLER_44_358 ();
 sg13g2_fill_2 FILLER_44_365 ();
 sg13g2_decap_8 FILLER_44_372 ();
 sg13g2_decap_8 FILLER_44_379 ();
 sg13g2_fill_1 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_395 ();
 sg13g2_decap_8 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_69 ();
 sg13g2_decap_4 FILLER_45_80 ();
 sg13g2_fill_2 FILLER_45_84 ();
 sg13g2_fill_1 FILLER_45_95 ();
 sg13g2_decap_4 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_109 ();
 sg13g2_fill_1 FILLER_45_114 ();
 sg13g2_fill_2 FILLER_45_178 ();
 sg13g2_fill_1 FILLER_45_180 ();
 sg13g2_decap_4 FILLER_45_198 ();
 sg13g2_fill_2 FILLER_45_227 ();
 sg13g2_decap_8 FILLER_45_241 ();
 sg13g2_decap_8 FILLER_45_248 ();
 sg13g2_fill_2 FILLER_45_255 ();
 sg13g2_fill_1 FILLER_45_257 ();
 sg13g2_fill_2 FILLER_45_272 ();
 sg13g2_fill_1 FILLER_45_274 ();
 sg13g2_fill_2 FILLER_45_295 ();
 sg13g2_fill_1 FILLER_45_297 ();
 sg13g2_decap_8 FILLER_45_307 ();
 sg13g2_fill_2 FILLER_45_314 ();
 sg13g2_decap_8 FILLER_45_358 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_4 FILLER_45_378 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_fill_2 FILLER_46_21 ();
 sg13g2_fill_1 FILLER_46_23 ();
 sg13g2_fill_2 FILLER_46_76 ();
 sg13g2_decap_4 FILLER_46_84 ();
 sg13g2_fill_1 FILLER_46_108 ();
 sg13g2_decap_4 FILLER_46_167 ();
 sg13g2_fill_2 FILLER_46_211 ();
 sg13g2_fill_1 FILLER_46_213 ();
 sg13g2_fill_2 FILLER_46_231 ();
 sg13g2_fill_1 FILLER_46_233 ();
 sg13g2_fill_2 FILLER_46_279 ();
 sg13g2_fill_1 FILLER_46_281 ();
 sg13g2_fill_2 FILLER_46_292 ();
 sg13g2_fill_1 FILLER_46_294 ();
 sg13g2_fill_2 FILLER_46_311 ();
 sg13g2_fill_1 FILLER_46_319 ();
 sg13g2_decap_8 FILLER_46_325 ();
 sg13g2_decap_4 FILLER_46_332 ();
 sg13g2_fill_1 FILLER_46_336 ();
 sg13g2_decap_4 FILLER_46_343 ();
 sg13g2_decap_4 FILLER_46_372 ();
 sg13g2_fill_1 FILLER_46_376 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_4 FILLER_47_21 ();
 sg13g2_fill_1 FILLER_47_41 ();
 sg13g2_decap_4 FILLER_47_110 ();
 sg13g2_fill_2 FILLER_47_132 ();
 sg13g2_fill_2 FILLER_47_139 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_fill_2 FILLER_47_161 ();
 sg13g2_fill_1 FILLER_47_163 ();
 sg13g2_fill_2 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_194 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_fill_1 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_369 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_decap_8 FILLER_47_383 ();
 sg13g2_decap_8 FILLER_47_390 ();
 sg13g2_decap_8 FILLER_47_397 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_fill_1 FILLER_48_69 ();
 sg13g2_fill_1 FILLER_48_79 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_fill_1 FILLER_48_123 ();
 sg13g2_decap_8 FILLER_48_146 ();
 sg13g2_fill_2 FILLER_48_153 ();
 sg13g2_fill_1 FILLER_48_155 ();
 sg13g2_decap_8 FILLER_48_173 ();
 sg13g2_decap_8 FILLER_48_180 ();
 sg13g2_decap_8 FILLER_48_187 ();
 sg13g2_decap_4 FILLER_48_194 ();
 sg13g2_fill_1 FILLER_48_198 ();
 sg13g2_decap_4 FILLER_48_254 ();
 sg13g2_fill_2 FILLER_48_258 ();
 sg13g2_fill_2 FILLER_48_271 ();
 sg13g2_decap_8 FILLER_48_281 ();
 sg13g2_fill_2 FILLER_48_288 ();
 sg13g2_decap_8 FILLER_48_302 ();
 sg13g2_fill_1 FILLER_48_309 ();
 sg13g2_fill_2 FILLER_48_321 ();
 sg13g2_fill_1 FILLER_48_323 ();
 sg13g2_fill_1 FILLER_48_366 ();
 sg13g2_decap_8 FILLER_48_384 ();
 sg13g2_decap_8 FILLER_48_391 ();
 sg13g2_decap_8 FILLER_48_398 ();
 sg13g2_decap_4 FILLER_48_405 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_4 FILLER_49_14 ();
 sg13g2_fill_1 FILLER_49_18 ();
 sg13g2_fill_1 FILLER_49_54 ();
 sg13g2_fill_1 FILLER_49_89 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_fill_1 FILLER_49_97 ();
 sg13g2_decap_8 FILLER_49_107 ();
 sg13g2_fill_1 FILLER_49_127 ();
 sg13g2_fill_2 FILLER_49_188 ();
 sg13g2_decap_4 FILLER_49_196 ();
 sg13g2_fill_1 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_209 ();
 sg13g2_decap_8 FILLER_49_216 ();
 sg13g2_decap_8 FILLER_49_223 ();
 sg13g2_decap_8 FILLER_49_230 ();
 sg13g2_fill_1 FILLER_49_237 ();
 sg13g2_decap_8 FILLER_49_244 ();
 sg13g2_decap_8 FILLER_49_251 ();
 sg13g2_decap_8 FILLER_49_258 ();
 sg13g2_fill_2 FILLER_49_265 ();
 sg13g2_fill_1 FILLER_49_267 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_333 ();
 sg13g2_decap_4 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_384 ();
 sg13g2_decap_8 FILLER_49_391 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_21 ();
 sg13g2_fill_1 FILLER_50_25 ();
 sg13g2_fill_1 FILLER_50_88 ();
 sg13g2_decap_8 FILLER_50_97 ();
 sg13g2_decap_4 FILLER_50_104 ();
 sg13g2_fill_2 FILLER_50_108 ();
 sg13g2_fill_1 FILLER_50_115 ();
 sg13g2_fill_2 FILLER_50_126 ();
 sg13g2_decap_4 FILLER_50_169 ();
 sg13g2_fill_1 FILLER_50_173 ();
 sg13g2_decap_8 FILLER_50_203 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_4 FILLER_50_217 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_decap_4 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_252 ();
 sg13g2_decap_4 FILLER_50_262 ();
 sg13g2_decap_8 FILLER_50_274 ();
 sg13g2_fill_1 FILLER_50_281 ();
 sg13g2_fill_2 FILLER_50_305 ();
 sg13g2_decap_8 FILLER_50_341 ();
 sg13g2_fill_2 FILLER_50_365 ();
 sg13g2_fill_1 FILLER_50_367 ();
 sg13g2_decap_8 FILLER_50_390 ();
 sg13g2_decap_8 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_404 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_4 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_39 ();
 sg13g2_fill_2 FILLER_51_95 ();
 sg13g2_fill_2 FILLER_51_120 ();
 sg13g2_fill_2 FILLER_51_136 ();
 sg13g2_decap_4 FILLER_51_178 ();
 sg13g2_fill_2 FILLER_51_233 ();
 sg13g2_fill_1 FILLER_51_235 ();
 sg13g2_fill_2 FILLER_51_275 ();
 sg13g2_fill_2 FILLER_51_311 ();
 sg13g2_decap_8 FILLER_51_380 ();
 sg13g2_decap_8 FILLER_51_387 ();
 sg13g2_decap_8 FILLER_51_394 ();
 sg13g2_decap_8 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_28 ();
 sg13g2_fill_1 FILLER_52_44 ();
 sg13g2_fill_1 FILLER_52_50 ();
 sg13g2_fill_1 FILLER_52_55 ();
 sg13g2_fill_1 FILLER_52_92 ();
 sg13g2_fill_1 FILLER_52_103 ();
 sg13g2_decap_8 FILLER_52_132 ();
 sg13g2_decap_8 FILLER_52_139 ();
 sg13g2_decap_4 FILLER_52_146 ();
 sg13g2_fill_2 FILLER_52_150 ();
 sg13g2_fill_2 FILLER_52_173 ();
 sg13g2_fill_1 FILLER_52_175 ();
 sg13g2_fill_2 FILLER_52_204 ();
 sg13g2_fill_2 FILLER_52_229 ();
 sg13g2_fill_1 FILLER_52_231 ();
 sg13g2_fill_2 FILLER_52_263 ();
 sg13g2_fill_2 FILLER_52_275 ();
 sg13g2_fill_1 FILLER_52_277 ();
 sg13g2_decap_8 FILLER_52_335 ();
 sg13g2_decap_8 FILLER_52_342 ();
 sg13g2_decap_4 FILLER_52_349 ();
 sg13g2_fill_1 FILLER_52_353 ();
 sg13g2_decap_4 FILLER_52_362 ();
 sg13g2_fill_1 FILLER_52_366 ();
 sg13g2_decap_4 FILLER_52_375 ();
 sg13g2_decap_4 FILLER_52_404 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_50 ();
 sg13g2_fill_2 FILLER_53_81 ();
 sg13g2_fill_1 FILLER_53_88 ();
 sg13g2_decap_8 FILLER_53_116 ();
 sg13g2_decap_8 FILLER_53_123 ();
 sg13g2_fill_2 FILLER_53_130 ();
 sg13g2_fill_1 FILLER_53_132 ();
 sg13g2_fill_1 FILLER_53_138 ();
 sg13g2_fill_2 FILLER_53_143 ();
 sg13g2_decap_4 FILLER_53_154 ();
 sg13g2_decap_4 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_191 ();
 sg13g2_decap_8 FILLER_53_198 ();
 sg13g2_fill_2 FILLER_53_205 ();
 sg13g2_fill_1 FILLER_53_207 ();
 sg13g2_decap_8 FILLER_53_225 ();
 sg13g2_decap_8 FILLER_53_237 ();
 sg13g2_decap_4 FILLER_53_244 ();
 sg13g2_fill_1 FILLER_53_258 ();
 sg13g2_fill_2 FILLER_53_285 ();
 sg13g2_fill_1 FILLER_53_287 ();
 sg13g2_fill_2 FILLER_53_313 ();
 sg13g2_fill_2 FILLER_53_323 ();
 sg13g2_fill_2 FILLER_53_333 ();
 sg13g2_fill_1 FILLER_53_335 ();
 sg13g2_fill_2 FILLER_53_353 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_4 FILLER_53_403 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_4 ();
 sg13g2_fill_1 FILLER_54_32 ();
 sg13g2_fill_2 FILLER_54_41 ();
 sg13g2_fill_1 FILLER_54_43 ();
 sg13g2_fill_2 FILLER_54_54 ();
 sg13g2_fill_2 FILLER_54_80 ();
 sg13g2_fill_2 FILLER_54_86 ();
 sg13g2_fill_1 FILLER_54_88 ();
 sg13g2_decap_8 FILLER_54_102 ();
 sg13g2_fill_1 FILLER_54_109 ();
 sg13g2_decap_4 FILLER_54_123 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_fill_2 FILLER_54_178 ();
 sg13g2_fill_2 FILLER_54_203 ();
 sg13g2_fill_1 FILLER_54_205 ();
 sg13g2_decap_8 FILLER_54_229 ();
 sg13g2_fill_2 FILLER_54_236 ();
 sg13g2_fill_1 FILLER_54_238 ();
 sg13g2_decap_4 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_248 ();
 sg13g2_fill_2 FILLER_54_257 ();
 sg13g2_decap_4 FILLER_54_291 ();
 sg13g2_fill_2 FILLER_54_295 ();
 sg13g2_decap_8 FILLER_54_310 ();
 sg13g2_decap_8 FILLER_54_317 ();
 sg13g2_decap_8 FILLER_54_324 ();
 sg13g2_fill_2 FILLER_54_331 ();
 sg13g2_fill_2 FILLER_54_358 ();
 sg13g2_decap_8 FILLER_54_377 ();
 sg13g2_decap_8 FILLER_54_384 ();
 sg13g2_decap_8 FILLER_54_391 ();
 sg13g2_decap_8 FILLER_54_398 ();
 sg13g2_decap_4 FILLER_54_405 ();
 sg13g2_fill_2 FILLER_55_39 ();
 sg13g2_fill_1 FILLER_55_41 ();
 sg13g2_fill_2 FILLER_55_81 ();
 sg13g2_fill_1 FILLER_55_83 ();
 sg13g2_fill_2 FILLER_55_92 ();
 sg13g2_fill_1 FILLER_55_94 ();
 sg13g2_fill_1 FILLER_55_100 ();
 sg13g2_fill_2 FILLER_55_109 ();
 sg13g2_decap_4 FILLER_55_176 ();
 sg13g2_fill_1 FILLER_55_180 ();
 sg13g2_fill_1 FILLER_55_198 ();
 sg13g2_fill_2 FILLER_55_224 ();
 sg13g2_fill_1 FILLER_55_256 ();
 sg13g2_decap_8 FILLER_55_293 ();
 sg13g2_decap_4 FILLER_55_300 ();
 sg13g2_fill_2 FILLER_55_332 ();
 sg13g2_fill_2 FILLER_55_351 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_2 FILLER_56_42 ();
 sg13g2_fill_1 FILLER_56_117 ();
 sg13g2_fill_1 FILLER_56_205 ();
 sg13g2_decap_4 FILLER_56_211 ();
 sg13g2_decap_8 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_252 ();
 sg13g2_decap_8 FILLER_56_259 ();
 sg13g2_fill_1 FILLER_56_266 ();
 sg13g2_fill_2 FILLER_56_288 ();
 sg13g2_fill_1 FILLER_56_290 ();
 sg13g2_fill_2 FILLER_56_325 ();
 sg13g2_decap_8 FILLER_56_344 ();
 sg13g2_decap_8 FILLER_56_351 ();
 sg13g2_fill_1 FILLER_56_358 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_2 FILLER_57_23 ();
 sg13g2_fill_2 FILLER_57_48 ();
 sg13g2_fill_1 FILLER_57_68 ();
 sg13g2_fill_1 FILLER_57_107 ();
 sg13g2_fill_2 FILLER_57_138 ();
 sg13g2_fill_2 FILLER_57_166 ();
 sg13g2_fill_2 FILLER_57_173 ();
 sg13g2_decap_8 FILLER_57_192 ();
 sg13g2_decap_8 FILLER_57_199 ();
 sg13g2_decap_8 FILLER_57_206 ();
 sg13g2_decap_8 FILLER_57_213 ();
 sg13g2_decap_8 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_227 ();
 sg13g2_fill_2 FILLER_57_234 ();
 sg13g2_fill_1 FILLER_57_236 ();
 sg13g2_decap_8 FILLER_57_254 ();
 sg13g2_fill_2 FILLER_57_261 ();
 sg13g2_fill_1 FILLER_57_263 ();
 sg13g2_decap_8 FILLER_57_277 ();
 sg13g2_decap_4 FILLER_57_284 ();
 sg13g2_fill_2 FILLER_57_288 ();
 sg13g2_decap_8 FILLER_57_347 ();
 sg13g2_decap_8 FILLER_57_354 ();
 sg13g2_fill_1 FILLER_57_361 ();
 sg13g2_decap_4 FILLER_57_368 ();
 sg13g2_decap_8 FILLER_57_394 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_2 ();
 sg13g2_fill_2 FILLER_58_56 ();
 sg13g2_fill_2 FILLER_58_81 ();
 sg13g2_fill_1 FILLER_58_83 ();
 sg13g2_fill_2 FILLER_58_97 ();
 sg13g2_fill_1 FILLER_58_99 ();
 sg13g2_fill_1 FILLER_58_118 ();
 sg13g2_fill_1 FILLER_58_164 ();
 sg13g2_decap_8 FILLER_58_170 ();
 sg13g2_decap_8 FILLER_58_177 ();
 sg13g2_decap_8 FILLER_58_184 ();
 sg13g2_decap_8 FILLER_58_191 ();
 sg13g2_decap_8 FILLER_58_215 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_fill_2 FILLER_58_263 ();
 sg13g2_fill_2 FILLER_58_302 ();
 sg13g2_fill_1 FILLER_58_304 ();
 sg13g2_decap_4 FILLER_58_313 ();
 sg13g2_fill_2 FILLER_58_317 ();
 sg13g2_fill_1 FILLER_58_336 ();
 sg13g2_fill_1 FILLER_58_348 ();
 sg13g2_decap_4 FILLER_58_366 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_23 ();
 sg13g2_fill_1 FILLER_59_25 ();
 sg13g2_fill_1 FILLER_59_47 ();
 sg13g2_fill_2 FILLER_59_83 ();
 sg13g2_fill_2 FILLER_59_111 ();
 sg13g2_decap_8 FILLER_59_122 ();
 sg13g2_decap_4 FILLER_59_129 ();
 sg13g2_decap_8 FILLER_59_142 ();
 sg13g2_fill_2 FILLER_59_149 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_fill_1 FILLER_59_194 ();
 sg13g2_decap_4 FILLER_59_218 ();
 sg13g2_decap_4 FILLER_59_262 ();
 sg13g2_fill_1 FILLER_59_266 ();
 sg13g2_decap_4 FILLER_59_275 ();
 sg13g2_fill_1 FILLER_59_279 ();
 sg13g2_decap_8 FILLER_59_297 ();
 sg13g2_decap_8 FILLER_59_304 ();
 sg13g2_fill_1 FILLER_59_311 ();
 sg13g2_fill_1 FILLER_59_368 ();
 sg13g2_fill_1 FILLER_59_375 ();
 sg13g2_decap_8 FILLER_59_384 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_405 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_fill_2 FILLER_60_53 ();
 sg13g2_decap_4 FILLER_60_96 ();
 sg13g2_decap_8 FILLER_60_131 ();
 sg13g2_fill_2 FILLER_60_164 ();
 sg13g2_fill_1 FILLER_60_166 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_4 FILLER_60_224 ();
 sg13g2_fill_1 FILLER_60_228 ();
 sg13g2_decap_8 FILLER_60_234 ();
 sg13g2_fill_2 FILLER_60_241 ();
 sg13g2_decap_4 FILLER_60_266 ();
 sg13g2_fill_1 FILLER_60_270 ();
 sg13g2_fill_2 FILLER_60_280 ();
 sg13g2_decap_4 FILLER_60_290 ();
 sg13g2_decap_8 FILLER_60_311 ();
 sg13g2_decap_8 FILLER_60_318 ();
 sg13g2_decap_8 FILLER_60_325 ();
 sg13g2_fill_2 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_340 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_decap_8 FILLER_60_372 ();
 sg13g2_decap_8 FILLER_60_379 ();
 sg13g2_decap_8 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_393 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_11 ();
 sg13g2_fill_1 FILLER_61_64 ();
 sg13g2_fill_2 FILLER_61_108 ();
 sg13g2_fill_1 FILLER_61_110 ();
 sg13g2_fill_1 FILLER_61_156 ();
 sg13g2_fill_2 FILLER_61_179 ();
 sg13g2_fill_2 FILLER_61_187 ();
 sg13g2_fill_2 FILLER_61_223 ();
 sg13g2_fill_1 FILLER_61_225 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_fill_2 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_253 ();
 sg13g2_decap_4 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_271 ();
 sg13g2_fill_2 FILLER_61_281 ();
 sg13g2_fill_1 FILLER_61_283 ();
 sg13g2_fill_1 FILLER_61_318 ();
 sg13g2_decap_4 FILLER_61_329 ();
 sg13g2_fill_2 FILLER_61_333 ();
 sg13g2_fill_2 FILLER_61_352 ();
 sg13g2_decap_8 FILLER_61_379 ();
 sg13g2_decap_8 FILLER_61_386 ();
 sg13g2_decap_8 FILLER_61_393 ();
 sg13g2_decap_8 FILLER_61_400 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_14 ();
 sg13g2_fill_1 FILLER_62_16 ();
 sg13g2_fill_2 FILLER_62_112 ();
 sg13g2_fill_1 FILLER_62_114 ();
 sg13g2_fill_2 FILLER_62_120 ();
 sg13g2_fill_1 FILLER_62_122 ();
 sg13g2_fill_2 FILLER_62_158 ();
 sg13g2_fill_1 FILLER_62_160 ();
 sg13g2_decap_4 FILLER_62_183 ();
 sg13g2_fill_1 FILLER_62_187 ();
 sg13g2_decap_8 FILLER_62_194 ();
 sg13g2_decap_8 FILLER_62_201 ();
 sg13g2_decap_4 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_212 ();
 sg13g2_decap_8 FILLER_62_237 ();
 sg13g2_fill_1 FILLER_62_244 ();
 sg13g2_decap_4 FILLER_62_268 ();
 sg13g2_fill_2 FILLER_62_272 ();
 sg13g2_fill_1 FILLER_62_299 ();
 sg13g2_fill_1 FILLER_62_351 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_1 FILLER_63_39 ();
 sg13g2_fill_2 FILLER_63_53 ();
 sg13g2_fill_2 FILLER_63_59 ();
 sg13g2_fill_2 FILLER_63_65 ();
 sg13g2_fill_1 FILLER_63_71 ();
 sg13g2_fill_1 FILLER_63_129 ();
 sg13g2_decap_4 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_267 ();
 sg13g2_decap_4 FILLER_63_293 ();
 sg13g2_fill_1 FILLER_63_297 ();
 sg13g2_fill_2 FILLER_63_315 ();
 sg13g2_fill_1 FILLER_63_317 ();
 sg13g2_decap_4 FILLER_63_335 ();
 sg13g2_fill_2 FILLER_63_362 ();
 sg13g2_fill_1 FILLER_63_364 ();
 sg13g2_decap_4 FILLER_63_404 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_21 ();
 sg13g2_fill_1 FILLER_64_61 ();
 sg13g2_fill_2 FILLER_64_85 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_fill_1 FILLER_64_140 ();
 sg13g2_decap_4 FILLER_64_149 ();
 sg13g2_fill_1 FILLER_64_153 ();
 sg13g2_decap_4 FILLER_64_171 ();
 sg13g2_fill_1 FILLER_64_175 ();
 sg13g2_fill_2 FILLER_64_205 ();
 sg13g2_decap_8 FILLER_64_285 ();
 sg13g2_fill_2 FILLER_64_292 ();
 sg13g2_fill_1 FILLER_64_294 ();
 sg13g2_fill_2 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_313 ();
 sg13g2_decap_4 FILLER_64_320 ();
 sg13g2_fill_1 FILLER_64_324 ();
 sg13g2_fill_1 FILLER_64_348 ();
 sg13g2_decap_8 FILLER_64_355 ();
 sg13g2_decap_4 FILLER_64_362 ();
 sg13g2_decap_8 FILLER_64_389 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_4 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_70 ();
 sg13g2_fill_2 FILLER_65_91 ();
 sg13g2_fill_1 FILLER_65_93 ();
 sg13g2_fill_2 FILLER_65_99 ();
 sg13g2_fill_1 FILLER_65_110 ();
 sg13g2_decap_8 FILLER_65_115 ();
 sg13g2_decap_8 FILLER_65_122 ();
 sg13g2_fill_2 FILLER_65_129 ();
 sg13g2_fill_1 FILLER_65_131 ();
 sg13g2_decap_4 FILLER_65_149 ();
 sg13g2_fill_2 FILLER_65_153 ();
 sg13g2_fill_2 FILLER_65_172 ();
 sg13g2_fill_1 FILLER_65_174 ();
 sg13g2_decap_8 FILLER_65_181 ();
 sg13g2_decap_8 FILLER_65_188 ();
 sg13g2_fill_2 FILLER_65_195 ();
 sg13g2_fill_1 FILLER_65_197 ();
 sg13g2_decap_4 FILLER_65_204 ();
 sg13g2_fill_2 FILLER_65_208 ();
 sg13g2_fill_2 FILLER_65_227 ();
 sg13g2_fill_1 FILLER_65_229 ();
 sg13g2_decap_4 FILLER_65_242 ();
 sg13g2_fill_1 FILLER_65_246 ();
 sg13g2_decap_8 FILLER_65_253 ();
 sg13g2_decap_8 FILLER_65_260 ();
 sg13g2_fill_2 FILLER_65_267 ();
 sg13g2_fill_1 FILLER_65_269 ();
 sg13g2_fill_2 FILLER_65_295 ();
 sg13g2_decap_4 FILLER_65_324 ();
 sg13g2_fill_2 FILLER_65_328 ();
 sg13g2_decap_4 FILLER_65_336 ();
 sg13g2_decap_4 FILLER_65_345 ();
 sg13g2_fill_2 FILLER_65_349 ();
 sg13g2_decap_8 FILLER_65_368 ();
 sg13g2_decap_8 FILLER_65_375 ();
 sg13g2_decap_8 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_396 ();
 sg13g2_decap_4 FILLER_65_403 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_4 FILLER_66_35 ();
 sg13g2_fill_2 FILLER_66_39 ();
 sg13g2_decap_8 FILLER_66_104 ();
 sg13g2_decap_8 FILLER_66_111 ();
 sg13g2_fill_2 FILLER_66_118 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_decap_8 FILLER_66_125 ();
 sg13g2_fill_2 FILLER_66_132 ();
 sg13g2_fill_1 FILLER_66_134 ();
 sg13g2_fill_2 FILLER_66_147 ();
 sg13g2_fill_1 FILLER_66_149 ();
 sg13g2_decap_8 FILLER_66_172 ();
 sg13g2_decap_8 FILLER_66_179 ();
 sg13g2_decap_8 FILLER_66_186 ();
 sg13g2_decap_8 FILLER_66_193 ();
 sg13g2_fill_2 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_202 ();
 sg13g2_decap_8 FILLER_66_208 ();
 sg13g2_decap_8 FILLER_66_215 ();
 sg13g2_fill_2 FILLER_66_222 ();
 sg13g2_decap_8 FILLER_66_230 ();
 sg13g2_decap_8 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_244 ();
 sg13g2_fill_2 FILLER_66_251 ();
 sg13g2_fill_1 FILLER_66_253 ();
 sg13g2_decap_4 FILLER_66_316 ();
 sg13g2_fill_2 FILLER_66_337 ();
 sg13g2_fill_2 FILLER_66_365 ();
 sg13g2_decap_8 FILLER_66_384 ();
 sg13g2_decap_8 FILLER_66_391 ();
 sg13g2_decap_8 FILLER_66_398 ();
 sg13g2_decap_4 FILLER_66_405 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_fill_2 FILLER_67_42 ();
 sg13g2_fill_1 FILLER_67_44 ();
 sg13g2_fill_2 FILLER_67_49 ();
 sg13g2_fill_1 FILLER_67_51 ();
 sg13g2_fill_2 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_58 ();
 sg13g2_fill_1 FILLER_67_90 ();
 sg13g2_fill_1 FILLER_67_96 ();
 sg13g2_decap_4 FILLER_67_153 ();
 sg13g2_fill_2 FILLER_67_157 ();
 sg13g2_fill_2 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_230 ();
 sg13g2_fill_1 FILLER_67_232 ();
 sg13g2_fill_1 FILLER_67_250 ();
 sg13g2_decap_8 FILLER_67_274 ();
 sg13g2_decap_8 FILLER_67_281 ();
 sg13g2_decap_4 FILLER_67_288 ();
 sg13g2_fill_1 FILLER_67_292 ();
 sg13g2_fill_2 FILLER_67_316 ();
 sg13g2_fill_1 FILLER_67_318 ();
 sg13g2_decap_4 FILLER_67_361 ();
 sg13g2_fill_2 FILLER_67_365 ();
 sg13g2_decap_8 FILLER_67_390 ();
 sg13g2_decap_8 FILLER_67_397 ();
 sg13g2_decap_4 FILLER_67_404 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_4 FILLER_68_35 ();
 sg13g2_fill_2 FILLER_68_39 ();
 sg13g2_decap_8 FILLER_68_44 ();
 sg13g2_decap_8 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_74 ();
 sg13g2_fill_2 FILLER_68_83 ();
 sg13g2_fill_1 FILLER_68_90 ();
 sg13g2_decap_4 FILLER_68_153 ();
 sg13g2_decap_4 FILLER_68_203 ();
 sg13g2_decap_4 FILLER_68_224 ();
 sg13g2_fill_1 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_246 ();
 sg13g2_fill_2 FILLER_68_271 ();
 sg13g2_fill_1 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_290 ();
 sg13g2_decap_8 FILLER_68_297 ();
 sg13g2_decap_8 FILLER_68_331 ();
 sg13g2_decap_8 FILLER_68_338 ();
 sg13g2_decap_8 FILLER_68_345 ();
 sg13g2_decap_8 FILLER_68_374 ();
 sg13g2_decap_8 FILLER_68_381 ();
 sg13g2_decap_8 FILLER_68_388 ();
 sg13g2_decap_8 FILLER_68_395 ();
 sg13g2_decap_8 FILLER_68_402 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_4 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_32 ();
 sg13g2_fill_2 FILLER_69_69 ();
 sg13g2_fill_1 FILLER_69_71 ();
 sg13g2_fill_1 FILLER_69_197 ();
 sg13g2_decap_4 FILLER_69_221 ();
 sg13g2_decap_8 FILLER_69_276 ();
 sg13g2_fill_1 FILLER_69_289 ();
 sg13g2_fill_2 FILLER_69_324 ();
 sg13g2_fill_1 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_380 ();
 sg13g2_decap_8 FILLER_69_387 ();
 sg13g2_decap_8 FILLER_69_394 ();
 sg13g2_decap_8 FILLER_69_401 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_fill_1 FILLER_70_35 ();
 sg13g2_fill_2 FILLER_70_82 ();
 sg13g2_fill_1 FILLER_70_96 ();
 sg13g2_fill_1 FILLER_70_106 ();
 sg13g2_fill_2 FILLER_70_146 ();
 sg13g2_fill_2 FILLER_70_169 ();
 sg13g2_decap_8 FILLER_70_188 ();
 sg13g2_fill_1 FILLER_70_195 ();
 sg13g2_decap_8 FILLER_70_213 ();
 sg13g2_decap_8 FILLER_70_220 ();
 sg13g2_decap_8 FILLER_70_250 ();
 sg13g2_decap_8 FILLER_70_257 ();
 sg13g2_decap_8 FILLER_70_264 ();
 sg13g2_fill_1 FILLER_70_271 ();
 sg13g2_fill_2 FILLER_70_289 ();
 sg13g2_fill_1 FILLER_70_291 ();
 sg13g2_fill_2 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_325 ();
 sg13g2_decap_4 FILLER_70_332 ();
 sg13g2_fill_1 FILLER_70_336 ();
 sg13g2_fill_2 FILLER_70_354 ();
 sg13g2_decap_8 FILLER_70_373 ();
 sg13g2_decap_8 FILLER_70_380 ();
 sg13g2_decap_8 FILLER_70_387 ();
 sg13g2_decap_8 FILLER_70_394 ();
 sg13g2_decap_8 FILLER_70_401 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_4 FILLER_71_28 ();
 sg13g2_fill_2 FILLER_71_32 ();
 sg13g2_fill_1 FILLER_71_96 ();
 sg13g2_fill_1 FILLER_71_110 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_4 FILLER_71_154 ();
 sg13g2_fill_1 FILLER_71_158 ();
 sg13g2_decap_8 FILLER_71_199 ();
 sg13g2_decap_8 FILLER_71_206 ();
 sg13g2_fill_2 FILLER_71_213 ();
 sg13g2_fill_1 FILLER_71_215 ();
 sg13g2_decap_8 FILLER_71_233 ();
 sg13g2_decap_8 FILLER_71_240 ();
 sg13g2_decap_4 FILLER_71_247 ();
 sg13g2_fill_2 FILLER_71_251 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_fill_2 FILLER_71_266 ();
 sg13g2_fill_1 FILLER_71_268 ();
 sg13g2_decap_8 FILLER_71_291 ();
 sg13g2_decap_8 FILLER_71_298 ();
 sg13g2_fill_1 FILLER_71_310 ();
 sg13g2_fill_2 FILLER_71_316 ();
 sg13g2_fill_1 FILLER_71_318 ();
 sg13g2_decap_8 FILLER_71_341 ();
 sg13g2_decap_8 FILLER_71_348 ();
 sg13g2_decap_8 FILLER_71_355 ();
 sg13g2_decap_8 FILLER_71_362 ();
 sg13g2_decap_8 FILLER_71_369 ();
 sg13g2_decap_8 FILLER_71_376 ();
 sg13g2_decap_8 FILLER_71_383 ();
 sg13g2_decap_8 FILLER_71_390 ();
 sg13g2_decap_8 FILLER_71_397 ();
 sg13g2_decap_4 FILLER_71_404 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_35 ();
 sg13g2_fill_2 FILLER_72_85 ();
 sg13g2_decap_4 FILLER_72_154 ();
 sg13g2_fill_1 FILLER_72_158 ();
 sg13g2_fill_2 FILLER_72_176 ();
 sg13g2_fill_1 FILLER_72_178 ();
 sg13g2_decap_8 FILLER_72_191 ();
 sg13g2_decap_8 FILLER_72_198 ();
 sg13g2_fill_1 FILLER_72_240 ();
 sg13g2_fill_2 FILLER_72_270 ();
 sg13g2_fill_1 FILLER_72_272 ();
 sg13g2_decap_4 FILLER_72_281 ();
 sg13g2_fill_2 FILLER_72_285 ();
 sg13g2_fill_2 FILLER_72_309 ();
 sg13g2_fill_1 FILLER_72_311 ();
 sg13g2_fill_2 FILLER_72_341 ();
 sg13g2_fill_2 FILLER_72_360 ();
 sg13g2_decap_8 FILLER_72_379 ();
 sg13g2_decap_8 FILLER_72_386 ();
 sg13g2_decap_8 FILLER_72_393 ();
 sg13g2_decap_8 FILLER_72_400 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_fill_2 FILLER_73_119 ();
 sg13g2_fill_1 FILLER_73_121 ();
 sg13g2_fill_1 FILLER_73_228 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_fill_2 FILLER_73_287 ();
 sg13g2_fill_1 FILLER_73_289 ();
 sg13g2_decap_4 FILLER_73_295 ();
 sg13g2_fill_1 FILLER_73_299 ();
 sg13g2_decap_4 FILLER_73_317 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_4 FILLER_73_350 ();
 sg13g2_fill_2 FILLER_73_354 ();
 sg13g2_fill_1 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_386 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_4 FILLER_74_42 ();
 sg13g2_fill_1 FILLER_74_46 ();
 sg13g2_fill_1 FILLER_74_114 ();
 sg13g2_fill_1 FILLER_74_182 ();
 sg13g2_decap_4 FILLER_74_268 ();
 sg13g2_fill_2 FILLER_74_272 ();
 sg13g2_decap_8 FILLER_74_299 ();
 sg13g2_decap_4 FILLER_74_306 ();
 sg13g2_decap_8 FILLER_74_316 ();
 sg13g2_fill_2 FILLER_74_323 ();
 sg13g2_fill_1 FILLER_74_325 ();
 sg13g2_fill_1 FILLER_74_332 ();
 sg13g2_fill_2 FILLER_74_338 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_4 FILLER_75_42 ();
 sg13g2_fill_2 FILLER_75_72 ();
 sg13g2_fill_1 FILLER_75_114 ();
 sg13g2_fill_1 FILLER_75_120 ();
 sg13g2_fill_2 FILLER_75_148 ();
 sg13g2_decap_8 FILLER_75_163 ();
 sg13g2_decap_4 FILLER_75_170 ();
 sg13g2_fill_1 FILLER_75_174 ();
 sg13g2_fill_2 FILLER_75_198 ();
 sg13g2_decap_8 FILLER_75_229 ();
 sg13g2_decap_8 FILLER_75_236 ();
 sg13g2_decap_8 FILLER_75_243 ();
 sg13g2_fill_1 FILLER_75_250 ();
 sg13g2_fill_2 FILLER_75_291 ();
 sg13g2_decap_4 FILLER_75_350 ();
 sg13g2_fill_1 FILLER_75_354 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_4 FILLER_76_49 ();
 sg13g2_fill_1 FILLER_76_53 ();
 sg13g2_fill_2 FILLER_76_75 ();
 sg13g2_fill_1 FILLER_76_77 ();
 sg13g2_fill_2 FILLER_76_97 ();
 sg13g2_fill_1 FILLER_76_99 ();
 sg13g2_fill_1 FILLER_76_117 ();
 sg13g2_decap_8 FILLER_76_162 ();
 sg13g2_decap_8 FILLER_76_230 ();
 sg13g2_decap_8 FILLER_76_237 ();
 sg13g2_decap_4 FILLER_76_244 ();
 sg13g2_decap_8 FILLER_76_265 ();
 sg13g2_decap_4 FILLER_76_272 ();
 sg13g2_fill_2 FILLER_76_276 ();
 sg13g2_fill_2 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_297 ();
 sg13g2_decap_8 FILLER_76_366 ();
 sg13g2_decap_8 FILLER_76_373 ();
 sg13g2_decap_8 FILLER_76_380 ();
 sg13g2_decap_8 FILLER_76_387 ();
 sg13g2_decap_8 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_4 FILLER_77_56 ();
 sg13g2_fill_2 FILLER_77_60 ();
 sg13g2_fill_1 FILLER_77_111 ();
 sg13g2_fill_1 FILLER_77_146 ();
 sg13g2_fill_1 FILLER_77_157 ();
 sg13g2_fill_1 FILLER_77_205 ();
 sg13g2_fill_1 FILLER_77_223 ();
 sg13g2_decap_4 FILLER_77_250 ();
 sg13g2_fill_1 FILLER_77_254 ();
 sg13g2_decap_8 FILLER_77_272 ();
 sg13g2_fill_2 FILLER_77_279 ();
 sg13g2_fill_2 FILLER_77_298 ();
 sg13g2_fill_1 FILLER_77_300 ();
 sg13g2_decap_8 FILLER_77_318 ();
 sg13g2_decap_4 FILLER_77_325 ();
 sg13g2_fill_1 FILLER_77_346 ();
 sg13g2_decap_8 FILLER_77_353 ();
 sg13g2_decap_8 FILLER_77_360 ();
 sg13g2_decap_8 FILLER_77_367 ();
 sg13g2_decap_8 FILLER_77_374 ();
 sg13g2_decap_8 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_388 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_4 FILLER_78_63 ();
 sg13g2_fill_2 FILLER_78_67 ();
 sg13g2_fill_2 FILLER_78_108 ();
 sg13g2_fill_1 FILLER_78_120 ();
 sg13g2_fill_1 FILLER_78_139 ();
 sg13g2_decap_4 FILLER_78_183 ();
 sg13g2_fill_1 FILLER_78_204 ();
 sg13g2_fill_2 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_302 ();
 sg13g2_decap_8 FILLER_78_309 ();
 sg13g2_decap_8 FILLER_78_316 ();
 sg13g2_decap_8 FILLER_78_323 ();
 sg13g2_fill_1 FILLER_78_330 ();
 sg13g2_decap_8 FILLER_78_348 ();
 sg13g2_decap_8 FILLER_78_355 ();
 sg13g2_decap_8 FILLER_78_362 ();
 sg13g2_decap_8 FILLER_78_369 ();
 sg13g2_decap_8 FILLER_78_376 ();
 sg13g2_decap_8 FILLER_78_383 ();
 sg13g2_decap_8 FILLER_78_390 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_4 FILLER_79_63 ();
 sg13g2_fill_1 FILLER_79_67 ();
 sg13g2_fill_2 FILLER_79_102 ();
 sg13g2_fill_1 FILLER_79_104 ();
 sg13g2_fill_2 FILLER_79_183 ();
 sg13g2_fill_1 FILLER_79_202 ();
 sg13g2_decap_4 FILLER_79_254 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_338 ();
 sg13g2_decap_8 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_4 FILLER_80_49 ();
 sg13g2_fill_2 FILLER_80_53 ();
 sg13g2_fill_2 FILLER_80_84 ();
 sg13g2_fill_1 FILLER_80_86 ();
 sg13g2_fill_1 FILLER_80_99 ();
 sg13g2_fill_2 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_167 ();
 sg13g2_fill_1 FILLER_80_176 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_213 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_227 ();
 sg13g2_fill_1 FILLER_80_234 ();
 sg13g2_decap_4 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_decap_8 FILLER_80_253 ();
 sg13g2_decap_4 FILLER_80_260 ();
 sg13g2_fill_2 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_321 ();
 sg13g2_decap_8 FILLER_80_328 ();
 sg13g2_fill_1 FILLER_80_335 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_decap_8 FILLER_80_357 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_8 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_385 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net93;
 assign uio_oe[3] = net94;
 assign uio_oe[4] = net95;
 assign uio_oe[5] = net96;
 assign uio_oe[6] = net97;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[7] = net12;
endmodule

module tt_um_wokwi_group_3 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire net240;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net12 ;
 wire \proj_10.net13 ;
 wire \proj_10.net9 ;
 wire \proj_12.net10 ;
 wire \proj_12.net11 ;
 wire \proj_12.net12 ;
 wire \proj_12.net13 ;
 wire \proj_12.net18 ;
 wire \proj_12.net19 ;
 wire \proj_12.net20 ;
 wire \proj_12.net21 ;
 wire \proj_12.net22 ;
 wire \proj_12.net23 ;
 wire \proj_12.net24 ;
 wire \proj_12.net25 ;
 wire \proj_12.net26 ;
 wire \proj_12.net27 ;
 wire \proj_12.net28 ;
 wire \proj_12.net29 ;
 wire \proj_12.net9 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net7 ;
 wire \proj_13.net8 ;
 wire \proj_14.net100 ;
 wire \proj_14.net101 ;
 wire \proj_14.net102 ;
 wire \proj_14.net104 ;
 wire \proj_14.net105 ;
 wire \proj_14.net106 ;
 wire \proj_14.net108 ;
 wire \proj_14.net11 ;
 wire \proj_14.net110 ;
 wire \proj_14.net111 ;
 wire \proj_14.net112 ;
 wire \proj_14.net114 ;
 wire \proj_14.net115 ;
 wire \proj_14.net116 ;
 wire \proj_14.net117 ;
 wire \proj_14.net119 ;
 wire \proj_14.net12 ;
 wire \proj_14.net120 ;
 wire \proj_14.net121 ;
 wire \proj_14.net122 ;
 wire \proj_14.net124 ;
 wire \proj_14.net125 ;
 wire \proj_14.net126 ;
 wire \proj_14.net127 ;
 wire \proj_14.net129 ;
 wire \proj_14.net13 ;
 wire \proj_14.net130 ;
 wire \proj_14.net131 ;
 wire \proj_14.net132 ;
 wire \proj_14.net133 ;
 wire \proj_14.net135 ;
 wire \proj_14.net136 ;
 wire \proj_14.net137 ;
 wire \proj_14.net138 ;
 wire \proj_14.net14 ;
 wire \proj_14.net140 ;
 wire \proj_14.net141 ;
 wire \proj_14.net142 ;
 wire \proj_14.net143 ;
 wire \proj_14.net145 ;
 wire \proj_14.net146 ;
 wire \proj_14.net147 ;
 wire \proj_14.net148 ;
 wire \proj_14.net15 ;
 wire \proj_14.net150 ;
 wire \proj_14.net151 ;
 wire \proj_14.net152 ;
 wire \proj_14.net153 ;
 wire \proj_14.net155 ;
 wire \proj_14.net156 ;
 wire \proj_14.net157 ;
 wire \proj_14.net158 ;
 wire \proj_14.net16 ;
 wire \proj_14.net160 ;
 wire \proj_14.net161 ;
 wire \proj_14.net162 ;
 wire \proj_14.net163 ;
 wire \proj_14.net165 ;
 wire \proj_14.net166 ;
 wire \proj_14.net167 ;
 wire \proj_14.net168 ;
 wire \proj_14.net17 ;
 wire \proj_14.net170 ;
 wire \proj_14.net171 ;
 wire \proj_14.net172 ;
 wire \proj_14.net173 ;
 wire \proj_14.net175 ;
 wire \proj_14.net176 ;
 wire \proj_14.net177 ;
 wire \proj_14.net178 ;
 wire \proj_14.net180 ;
 wire \proj_14.net181 ;
 wire \proj_14.net182 ;
 wire \proj_14.net183 ;
 wire \proj_14.net184 ;
 wire \proj_14.net185 ;
 wire \proj_14.net186 ;
 wire \proj_14.net187 ;
 wire \proj_14.net188 ;
 wire \proj_14.net189 ;
 wire \proj_14.net190 ;
 wire \proj_14.net191 ;
 wire \proj_14.net192 ;
 wire \proj_14.net193 ;
 wire \proj_14.net194 ;
 wire \proj_14.net195 ;
 wire \proj_14.net196 ;
 wire \proj_14.net197 ;
 wire \proj_14.net198 ;
 wire \proj_14.net199 ;
 wire \proj_14.net200 ;
 wire \proj_14.net201 ;
 wire \proj_14.net202 ;
 wire \proj_14.net203 ;
 wire \proj_14.net204 ;
 wire \proj_14.net205 ;
 wire \proj_14.net206 ;
 wire \proj_14.net207 ;
 wire \proj_14.net209 ;
 wire \proj_14.net210 ;
 wire \proj_14.net211 ;
 wire \proj_14.net212 ;
 wire \proj_14.net214 ;
 wire \proj_14.net215 ;
 wire \proj_14.net216 ;
 wire \proj_14.net217 ;
 wire \proj_14.net218 ;
 wire \proj_14.net219 ;
 wire \proj_14.net220 ;
 wire \proj_14.net221 ;
 wire \proj_14.net222 ;
 wire \proj_14.net223 ;
 wire \proj_14.net224 ;
 wire \proj_14.net226 ;
 wire \proj_14.net227 ;
 wire \proj_14.net228 ;
 wire \proj_14.net229 ;
 wire \proj_14.net23 ;
 wire \proj_14.net231 ;
 wire \proj_14.net232 ;
 wire \proj_14.net233 ;
 wire \proj_14.net234 ;
 wire \proj_14.net235 ;
 wire \proj_14.net236 ;
 wire \proj_14.net237 ;
 wire \proj_14.net238 ;
 wire \proj_14.net239 ;
 wire \proj_14.net240 ;
 wire \proj_14.net241 ;
 wire \proj_14.net242 ;
 wire \proj_14.net243 ;
 wire \proj_14.net244 ;
 wire \proj_14.net245 ;
 wire \proj_14.net246 ;
 wire \proj_14.net247 ;
 wire \proj_14.net248 ;
 wire \proj_14.net249 ;
 wire \proj_14.net25 ;
 wire \proj_14.net250 ;
 wire \proj_14.net251 ;
 wire \proj_14.net252 ;
 wire \proj_14.net253 ;
 wire \proj_14.net254 ;
 wire \proj_14.net255 ;
 wire \proj_14.net256 ;
 wire \proj_14.net257 ;
 wire \proj_14.net258 ;
 wire \proj_14.net259 ;
 wire \proj_14.net26 ;
 wire \proj_14.net260 ;
 wire \proj_14.net261 ;
 wire \proj_14.net262 ;
 wire \proj_14.net263 ;
 wire \proj_14.net264 ;
 wire \proj_14.net265 ;
 wire \proj_14.net266 ;
 wire \proj_14.net267 ;
 wire \proj_14.net268 ;
 wire \proj_14.net269 ;
 wire \proj_14.net27 ;
 wire \proj_14.net270 ;
 wire \proj_14.net271 ;
 wire \proj_14.net272 ;
 wire \proj_14.net273 ;
 wire \proj_14.net274 ;
 wire \proj_14.net275 ;
 wire \proj_14.net276 ;
 wire \proj_14.net277 ;
 wire \proj_14.net278 ;
 wire \proj_14.net279 ;
 wire \proj_14.net28 ;
 wire \proj_14.net280 ;
 wire \proj_14.net281 ;
 wire \proj_14.net282 ;
 wire \proj_14.net283 ;
 wire \proj_14.net284 ;
 wire \proj_14.net285 ;
 wire \proj_14.net286 ;
 wire \proj_14.net287 ;
 wire \proj_14.net288 ;
 wire \proj_14.net289 ;
 wire \proj_14.net29 ;
 wire \proj_14.net30 ;
 wire \proj_14.net31 ;
 wire \proj_14.net32 ;
 wire \proj_14.net33 ;
 wire \proj_14.net34 ;
 wire \proj_14.net36 ;
 wire \proj_14.net37 ;
 wire \proj_14.net38 ;
 wire \proj_14.net39 ;
 wire \proj_14.net40 ;
 wire \proj_14.net41 ;
 wire \proj_14.net42 ;
 wire \proj_14.net43 ;
 wire \proj_14.net44 ;
 wire \proj_14.net45 ;
 wire \proj_14.net46 ;
 wire \proj_14.net47 ;
 wire \proj_14.net48 ;
 wire \proj_14.net50 ;
 wire \proj_14.net51 ;
 wire \proj_14.net52 ;
 wire \proj_14.net53 ;
 wire \proj_14.net54 ;
 wire \proj_14.net55 ;
 wire \proj_14.net56 ;
 wire \proj_14.net57 ;
 wire \proj_14.net58 ;
 wire \proj_14.net59 ;
 wire \proj_14.net60 ;
 wire \proj_14.net61 ;
 wire \proj_14.net62 ;
 wire \proj_14.net63 ;
 wire \proj_14.net64 ;
 wire \proj_14.net65 ;
 wire \proj_14.net66 ;
 wire \proj_14.net67 ;
 wire \proj_14.net68 ;
 wire \proj_14.net69 ;
 wire \proj_14.net70 ;
 wire \proj_14.net71 ;
 wire \proj_14.net72 ;
 wire \proj_14.net73 ;
 wire \proj_14.net74 ;
 wire \proj_14.net75 ;
 wire \proj_14.net76 ;
 wire \proj_14.net77 ;
 wire \proj_14.net78 ;
 wire \proj_14.net79 ;
 wire \proj_14.net80 ;
 wire \proj_14.net81 ;
 wire \proj_14.net82 ;
 wire \proj_14.net83 ;
 wire \proj_14.net84 ;
 wire \proj_14.net85 ;
 wire \proj_14.net86 ;
 wire \proj_14.net87 ;
 wire \proj_14.net88 ;
 wire \proj_14.net89 ;
 wire \proj_14.net90 ;
 wire \proj_14.net91 ;
 wire \proj_14.net92 ;
 wire \proj_14.net93 ;
 wire \proj_14.net94 ;
 wire \proj_14.net95 ;
 wire \proj_14.net96 ;
 wire \proj_14.net97 ;
 wire \proj_14.net98 ;
 wire \proj_14.net99 ;
 wire \proj_15.net15 ;
 wire \proj_15.net16 ;
 wire \proj_15.net17 ;
 wire \proj_15.net18 ;
 wire \proj_15.net7 ;
 wire \proj_15.net8 ;
 wire \proj_15.net9 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__0.net9 ;
 wire \proj__1.net10 ;
 wire \proj__1.net16 ;
 wire \proj__1.net17 ;
 wire \proj__1.net18 ;
 wire \proj__1.net19 ;
 wire \proj__1.net20 ;
 wire \proj__1.net21 ;
 wire \proj__1.net22 ;
 wire \proj__1.net23 ;
 wire \proj__1.net24 ;
 wire \proj__1.net9 ;
 wire \proj__2.net10 ;
 wire \proj__2.net11 ;
 wire \proj__2.net12 ;
 wire \proj__2.net9 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net3 ;
 wire \proj__3.net4 ;
 wire \proj__3.net5 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net13 ;
 wire \proj__4.net14 ;
 wire \proj__4.net15 ;
 wire \proj__4.net16 ;
 wire \proj__4.net17 ;
 wire \proj__4.net18 ;
 wire \proj__5.net10 ;
 wire \proj__5.net11 ;
 wire \proj__5.net12 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net9 ;
 wire \proj__7.net14 ;
 wire \proj__7.net15 ;
 wire \proj__7.net5 ;
 wire \proj__7.net6 ;
 wire \proj__7.net7 ;
 wire \proj__7.net8 ;
 wire \proj__8.net7 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net13 ;
 wire \proj__9.net14 ;
 wire \proj__9.net15 ;
 wire \proj__9.net17 ;
 wire \proj__9.net5 ;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire \proj_10.nand1/b ;
 wire net241;
 wire \proj_13.flop1/notq ;
 wire net242;
 wire \proj_13.flop2/notq ;
 wire net243;
 wire \proj_13.flop3/notq ;
 wire \proj_14.flop1/_0_ ;
 wire \proj_14.flop1/_1_ ;
 wire net150;
 wire net151;
 wire \proj_14.flop10/_0_ ;
 wire \proj_14.flop10/_1_ ;
 wire net152;
 wire net153;
 wire \proj_14.flop11/_0_ ;
 wire \proj_14.flop11/_1_ ;
 wire net154;
 wire net155;
 wire \proj_14.flop12/_0_ ;
 wire \proj_14.flop12/_1_ ;
 wire net156;
 wire net157;
 wire \proj_14.flop13/_0_ ;
 wire \proj_14.flop13/_1_ ;
 wire net158;
 wire net159;
 wire \proj_14.flop14/_0_ ;
 wire \proj_14.flop14/_1_ ;
 wire net160;
 wire net161;
 wire \proj_14.flop15/_0_ ;
 wire \proj_14.flop15/_1_ ;
 wire net162;
 wire net163;
 wire \proj_14.flop16/_0_ ;
 wire \proj_14.flop16/_1_ ;
 wire net164;
 wire net165;
 wire \proj_14.flop17/_0_ ;
 wire \proj_14.flop17/_1_ ;
 wire net166;
 wire net167;
 wire \proj_14.flop18/_0_ ;
 wire \proj_14.flop18/_1_ ;
 wire net168;
 wire net169;
 wire \proj_14.flop19/_0_ ;
 wire \proj_14.flop19/_1_ ;
 wire net170;
 wire net171;
 wire \proj_14.flop2/_0_ ;
 wire \proj_14.flop2/_1_ ;
 wire net172;
 wire net173;
 wire \proj_14.flop20/_0_ ;
 wire \proj_14.flop20/_1_ ;
 wire net174;
 wire net175;
 wire \proj_14.flop21/_0_ ;
 wire \proj_14.flop21/_1_ ;
 wire net176;
 wire net177;
 wire \proj_14.flop22/_0_ ;
 wire \proj_14.flop22/_1_ ;
 wire net178;
 wire net179;
 wire \proj_14.flop23/_0_ ;
 wire \proj_14.flop23/_1_ ;
 wire net180;
 wire net181;
 wire \proj_14.flop24/_0_ ;
 wire \proj_14.flop24/_1_ ;
 wire net182;
 wire net183;
 wire \proj_14.flop25/_0_ ;
 wire \proj_14.flop25/_1_ ;
 wire net184;
 wire net185;
 wire \proj_14.flop25/notq ;
 wire \proj_14.flop26/_0_ ;
 wire \proj_14.flop26/_1_ ;
 wire net186;
 wire net187;
 wire \proj_14.flop26/notq ;
 wire \proj_14.flop27/_0_ ;
 wire \proj_14.flop27/_1_ ;
 wire net188;
 wire net189;
 wire \proj_14.flop27/q ;
 wire net244;
 wire \proj_14.flop28/notq ;
 wire \proj_14.flop29/_0_ ;
 wire \proj_14.flop29/_1_ ;
 wire net190;
 wire net191;
 wire \proj_14.flop3/_0_ ;
 wire \proj_14.flop3/_1_ ;
 wire net192;
 wire net193;
 wire \proj_14.flop30/_0_ ;
 wire \proj_14.flop30/_1_ ;
 wire net194;
 wire net195;
 wire \proj_14.flop31/_0_ ;
 wire \proj_14.flop31/_1_ ;
 wire net196;
 wire net197;
 wire \proj_14.flop31/notq ;
 wire \proj_14.flop32/_0_ ;
 wire \proj_14.flop32/_1_ ;
 wire net198;
 wire net199;
 wire \proj_14.flop32/notq ;
 wire \proj_14.flop33/_0_ ;
 wire \proj_14.flop33/_1_ ;
 wire net200;
 wire net201;
 wire \proj_14.flop33/notq ;
 wire \proj_14.flop34/_0_ ;
 wire \proj_14.flop34/_1_ ;
 wire net202;
 wire net203;
 wire \proj_14.flop34/notq ;
 wire \proj_14.flop35/_0_ ;
 wire \proj_14.flop35/_1_ ;
 wire net204;
 wire net205;
 wire \proj_14.flop35/notq ;
 wire \proj_14.flop36/_0_ ;
 wire \proj_14.flop36/_1_ ;
 wire net206;
 wire net207;
 wire \proj_14.flop36/notq ;
 wire \proj_14.flop37/_0_ ;
 wire \proj_14.flop37/_1_ ;
 wire net208;
 wire net209;
 wire \proj_14.flop37/notq ;
 wire \proj_14.flop4/_0_ ;
 wire \proj_14.flop4/_1_ ;
 wire net210;
 wire net211;
 wire net245;
 wire \proj_14.flop46/notq ;
 wire net246;
 wire \proj_14.flop47/notq ;
 wire net247;
 wire \proj_14.flop48/notq ;
 wire net248;
 wire \proj_14.flop49/notq ;
 wire \proj_14.flop5/_0_ ;
 wire \proj_14.flop5/_1_ ;
 wire net212;
 wire net213;
 wire net249;
 wire \proj_14.flop50/notq ;
 wire net250;
 wire \proj_14.flop51/notq ;
 wire net251;
 wire \proj_14.flop52/notq ;
 wire net252;
 wire \proj_14.flop53/notq ;
 wire net253;
 wire \proj_14.flop54/notq ;
 wire net254;
 wire \proj_14.flop55/notq ;
 wire net255;
 wire \proj_14.flop56/notq ;
 wire \proj_14.flop6/_0_ ;
 wire \proj_14.flop6/_1_ ;
 wire net214;
 wire net215;
 wire \proj_14.flop7/_0_ ;
 wire \proj_14.flop7/_1_ ;
 wire net216;
 wire net217;
 wire \proj_14.flop8/_0_ ;
 wire \proj_14.flop8/_1_ ;
 wire net218;
 wire net219;
 wire \proj_14.flop9/_0_ ;
 wire \proj_14.flop9/_1_ ;
 wire net220;
 wire net221;
 wire \proj__4.flop1/_0_ ;
 wire \proj__4.flop1/_1_ ;
 wire net222;
 wire net223;
 wire \proj__4.flop1/q ;
 wire \proj__4.flop1/s ;
 wire \proj__4.flop2/_0_ ;
 wire \proj__4.flop2/_1_ ;
 wire net224;
 wire net225;
 wire \proj__4.flop2/q ;
 wire \proj__4.flop2/s ;
 wire \proj__4.flop3/_0_ ;
 wire \proj__4.flop3/_1_ ;
 wire net226;
 wire net227;
 wire \proj__4.flop3/q ;
 wire \proj__4.flop3/s ;
 wire \proj__4.flop4/_0_ ;
 wire \proj__4.flop4/_1_ ;
 wire net228;
 wire net229;
 wire \proj__4.flop4/q ;
 wire \proj__4.flop4/s ;
 wire \proj__4.flop5/_0_ ;
 wire \proj__4.flop5/_1_ ;
 wire net230;
 wire net231;
 wire \proj__4.flop5/notq ;
 wire \proj__4.flop5/s ;
 wire \proj__4.flop6/_0_ ;
 wire \proj__4.flop6/_1_ ;
 wire net232;
 wire net233;
 wire \proj__4.flop6/notq ;
 wire \proj__4.flop6/s ;
 wire \proj__4.flop8/_0_ ;
 wire \proj__4.flop8/_1_ ;
 wire net234;
 wire net235;
 wire \proj__4.flop8/notq ;
 wire \proj__4.flop8/s ;
 wire \proj__4.flop9/_0_ ;
 wire \proj__4.flop9/_1_ ;
 wire net236;
 wire net237;
 wire \proj__4.flop9/notq ;
 wire \proj__4.flop9/s ;
 wire net256;
 wire net257;
 wire \proj__9.flop1/_0_ ;
 wire \proj__9.flop1/_1_ ;
 wire net238;
 wire net239;
 wire \proj__9.flop1/notq ;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;

 sg13g2_inv_1 _192_ (.Y(_056_),
    .A(\proj__0.net9 ));
 sg13g2_inv_1 _193_ (.Y(_057_),
    .A(\proj__0.net10 ));
 sg13g2_inv_1 _194_ (.Y(_058_),
    .A(\proj__0.net11 ));
 sg13g2_nor2b_2 _195_ (.A(net9),
    .B_N(net8),
    .Y(_059_));
 sg13g2_nor2b_2 _196_ (.A(net7),
    .B_N(net6),
    .Y(_060_));
 sg13g2_and2_1 _197_ (.A(_059_),
    .B(_060_),
    .X(_061_));
 sg13g2_and2_2 _198_ (.A(net8),
    .B(net9),
    .X(_062_));
 sg13g2_nor2b_1 _199_ (.A(net6),
    .B_N(net7),
    .Y(_063_));
 sg13g2_nand2b_1 _200_ (.Y(_064_),
    .B(net7),
    .A_N(net6));
 sg13g2_nor2_2 _201_ (.A(net7),
    .B(net6),
    .Y(_065_));
 sg13g2_or3_1 _202_ (.A(net7),
    .B(net6),
    .C(net8),
    .X(_066_));
 sg13g2_o21ai_1 _203_ (.B1(_066_),
    .Y(_067_),
    .A1(net9),
    .A2(_064_));
 sg13g2_a21o_1 _204_ (.A2(_062_),
    .A1(net6),
    .B1(_067_),
    .X(_068_));
 sg13g2_o21ai_1 _205_ (.B1(net5),
    .Y(_069_),
    .A1(_061_),
    .A2(_068_));
 sg13g2_nor2b_2 _206_ (.A(net8),
    .B_N(net9),
    .Y(_070_));
 sg13g2_and2_2 _207_ (.A(_063_),
    .B(_070_),
    .X(_071_));
 sg13g2_and2_1 _208_ (.A(net7),
    .B(net6),
    .X(_072_));
 sg13g2_and2_1 _209_ (.A(_059_),
    .B(_072_),
    .X(_073_));
 sg13g2_and2_2 _210_ (.A(_059_),
    .B(_065_),
    .X(_074_));
 sg13g2_nand2_1 _211_ (.Y(_075_),
    .A(\proj__4.net18 ),
    .B(_074_));
 sg13g2_a22oi_1 _212_ (.Y(_076_),
    .B1(_073_),
    .B2(\proj__7.net8 ),
    .A2(_071_),
    .A1(\proj_10.net13 ));
 sg13g2_nand3_1 _213_ (.B(_075_),
    .C(_076_),
    .A(_069_),
    .Y(uo_out[7]));
 sg13g2_nor2_2 _214_ (.A(net8),
    .B(net9),
    .Y(_077_));
 sg13g2_nor2_2 _215_ (.A(net9),
    .B(_066_),
    .Y(_078_));
 sg13g2_a21oi_1 _216_ (.A1(\proj_10.net9 ),
    .A2(_071_),
    .Y(_079_),
    .B1(_078_));
 sg13g2_nand2_1 _217_ (.Y(_080_),
    .A(\proj__4.net11 ),
    .B(_074_));
 sg13g2_nand3_1 _218_ (.B(_060_),
    .C(_077_),
    .A(\proj__1.net9 ),
    .Y(_081_));
 sg13g2_and2_1 _219_ (.A(_072_),
    .B(_077_),
    .X(_000_));
 sg13g2_a22oi_1 _220_ (.Y(_001_),
    .B1(_072_),
    .B2(_077_),
    .A2(net43),
    .A1(_059_));
 sg13g2_nor2b_1 _221_ (.A(_001_),
    .B_N(net52),
    .Y(_002_));
 sg13g2_and2_1 _222_ (.A(net43),
    .B(_077_),
    .X(_003_));
 sg13g2_and2_2 _223_ (.A(_062_),
    .B(net43),
    .X(_004_));
 sg13g2_nand3_1 _224_ (.B(_062_),
    .C(net43),
    .A(\proj_14.net11 ),
    .Y(_005_));
 sg13g2_and4_1 _225_ (.A(net7),
    .B(net6),
    .C(net8),
    .D(net9),
    .X(_006_));
 sg13g2_nand2_1 _226_ (.Y(_007_),
    .A(\proj_15.net7 ),
    .B(_006_));
 sg13g2_nand3_1 _227_ (.B(_060_),
    .C(_062_),
    .A(\proj_13.net7 ),
    .Y(_008_));
 sg13g2_and2_2 _228_ (.A(_062_),
    .B(_065_),
    .X(_009_));
 sg13g2_nand3_1 _229_ (.B(_062_),
    .C(_065_),
    .A(\proj_12.net9 ),
    .Y(_010_));
 sg13g2_nand3_1 _230_ (.B(_060_),
    .C(_070_),
    .A(\proj__9.net5 ),
    .Y(_011_));
 sg13g2_nand3_1 _231_ (.B(_065_),
    .C(_070_),
    .A(\proj__8.net7 ),
    .Y(_012_));
 sg13g2_nand3_1 _232_ (.B(_059_),
    .C(_060_),
    .A(\proj__5.net9 ),
    .Y(_013_));
 sg13g2_a22oi_1 _233_ (.Y(_014_),
    .B1(_003_),
    .B2(\proj__2.net9 ),
    .A2(_073_),
    .A1(\proj__7.net5 ));
 sg13g2_and3_1 _234_ (.X(_015_),
    .A(_079_),
    .B(_080_),
    .C(_014_));
 sg13g2_nand4_1 _235_ (.B(_005_),
    .C(_010_),
    .A(_081_),
    .Y(_016_),
    .D(_012_));
 sg13g2_nand4_1 _236_ (.B(_008_),
    .C(_011_),
    .A(_007_),
    .Y(_017_),
    .D(_013_));
 sg13g2_nor3_1 _237_ (.A(_002_),
    .B(_016_),
    .C(_017_),
    .Y(_018_));
 sg13g2_a22oi_1 _238_ (.Y(uo_out[0]),
    .B1(_015_),
    .B2(_018_),
    .A2(_078_),
    .A1(_056_));
 sg13g2_nand2_1 _239_ (.Y(_019_),
    .A(\proj__7.net6 ),
    .B(_073_));
 sg13g2_nand3_1 _240_ (.B(_060_),
    .C(_062_),
    .A(\proj_13.net8 ),
    .Y(_020_));
 sg13g2_nor2b_1 _241_ (.A(_001_),
    .B_N(net50),
    .Y(_021_));
 sg13g2_and2_1 _242_ (.A(\proj__2.net10 ),
    .B(_003_),
    .X(_022_));
 sg13g2_a221oi_1 _243_ (.B2(\proj__4.net12 ),
    .C1(_022_),
    .B1(_074_),
    .A1(net47),
    .Y(_023_),
    .A2(_071_));
 sg13g2_a21oi_1 _244_ (.A1(\proj_15.net8 ),
    .A2(_006_),
    .Y(_024_),
    .B1(_021_));
 sg13g2_a22oi_1 _245_ (.Y(_025_),
    .B1(_009_),
    .B2(\proj_12.net10 ),
    .A2(_004_),
    .A1(\proj_14.net12 ));
 sg13g2_and4_1 _246_ (.A(_012_),
    .B(_019_),
    .C(_020_),
    .D(_025_),
    .X(_026_));
 sg13g2_nand3_1 _247_ (.B(_024_),
    .C(_026_),
    .A(_023_),
    .Y(uo_out[1]));
 sg13g2_nand2_1 _248_ (.Y(_027_),
    .A(\proj_15.net9 ),
    .B(_006_));
 sg13g2_nand2_1 _249_ (.Y(_028_),
    .A(\proj__2.net11 ),
    .B(_003_));
 sg13g2_nand3_1 _250_ (.B(net43),
    .C(_070_),
    .A(net44),
    .Y(_029_));
 sg13g2_and2_1 _251_ (.A(_012_),
    .B(_029_),
    .X(_030_));
 sg13g2_nand3_1 _252_ (.B(_059_),
    .C(net43),
    .A(\proj__6.net9 ),
    .Y(_031_));
 sg13g2_a22oi_1 _253_ (.Y(_032_),
    .B1(_009_),
    .B2(\proj_12.net11 ),
    .A2(_074_),
    .A1(\proj__4.net13 ));
 sg13g2_and2_1 _254_ (.A(_028_),
    .B(_032_),
    .X(_033_));
 sg13g2_a21oi_1 _255_ (.A1(\proj_14.net13 ),
    .A2(_004_),
    .Y(_034_),
    .B1(_078_));
 sg13g2_and4_1 _256_ (.A(_027_),
    .B(_030_),
    .C(_031_),
    .D(_034_),
    .X(_035_));
 sg13g2_a22oi_1 _257_ (.Y(uo_out[2]),
    .B1(_033_),
    .B2(_035_),
    .A2(_078_),
    .A1(_057_));
 sg13g2_nand2_1 _258_ (.Y(_036_),
    .A(\proj__2.net12 ),
    .B(_003_));
 sg13g2_nand3_1 _259_ (.B(_059_),
    .C(net43),
    .A(\proj__6.net10 ),
    .Y(_037_));
 sg13g2_a22oi_1 _260_ (.Y(_038_),
    .B1(_009_),
    .B2(\proj_12.net12 ),
    .A2(_004_),
    .A1(\proj_14.net14 ));
 sg13g2_a21oi_1 _261_ (.A1(\proj__4.net14 ),
    .A2(_074_),
    .Y(_039_),
    .B1(_078_));
 sg13g2_and4_1 _262_ (.A(_036_),
    .B(_037_),
    .C(_038_),
    .D(_039_),
    .X(_040_));
 sg13g2_a22oi_1 _263_ (.Y(uo_out[3]),
    .B1(_030_),
    .B2(_040_),
    .A2(_078_),
    .A1(_058_));
 sg13g2_a22oi_1 _264_ (.Y(_041_),
    .B1(_072_),
    .B2(_059_),
    .A2(_062_),
    .A1(_060_));
 sg13g2_nand2b_1 _265_ (.Y(_042_),
    .B(_041_),
    .A_N(_067_));
 sg13g2_nand3_1 _266_ (.B(net43),
    .C(_070_),
    .A(\proj_10.net10 ),
    .Y(_043_));
 sg13g2_a22oi_1 _267_ (.Y(_044_),
    .B1(_074_),
    .B2(\proj__4.net15 ),
    .A2(_061_),
    .A1(\proj__5.net10 ));
 sg13g2_nand2_1 _268_ (.Y(_045_),
    .A(_081_),
    .B(_043_));
 sg13g2_a22oi_1 _269_ (.Y(_046_),
    .B1(_009_),
    .B2(\proj_12.net13 ),
    .A2(_000_),
    .A1(\proj__3.net3 ));
 sg13g2_a221oi_1 _270_ (.B2(net2),
    .C1(_045_),
    .B1(_042_),
    .A1(\proj_14.net15 ),
    .Y(_047_),
    .A2(_004_));
 sg13g2_nand3_1 _271_ (.B(_046_),
    .C(_047_),
    .A(_044_),
    .Y(uo_out[4]));
 sg13g2_nand2_1 _272_ (.Y(_048_),
    .A(\proj_14.net16 ),
    .B(_004_));
 sg13g2_a22oi_1 _273_ (.Y(_049_),
    .B1(_074_),
    .B2(\proj__4.net16 ),
    .A2(_071_),
    .A1(\proj_10.net11 ));
 sg13g2_a22oi_1 _274_ (.Y(_050_),
    .B1(_000_),
    .B2(\proj__3.net4 ),
    .A2(_061_),
    .A1(\proj__5.net11 ));
 sg13g2_nand4_1 _275_ (.B(_048_),
    .C(_049_),
    .A(_081_),
    .Y(_051_),
    .D(_050_));
 sg13g2_a21o_1 _276_ (.A2(_042_),
    .A1(net44),
    .B1(_051_),
    .X(uo_out[5]));
 sg13g2_nand2_1 _277_ (.Y(_052_),
    .A(net4),
    .B(_068_));
 sg13g2_a22oi_1 _278_ (.Y(_053_),
    .B1(_004_),
    .B2(\proj_14.net17 ),
    .A2(_000_),
    .A1(\proj__3.net5 ));
 sg13g2_a22oi_1 _279_ (.Y(_054_),
    .B1(_074_),
    .B2(\proj__4.net17 ),
    .A2(_071_),
    .A1(\proj_10.net12 ));
 sg13g2_a22oi_1 _280_ (.Y(_055_),
    .B1(_073_),
    .B2(\proj__7.net7 ),
    .A2(_061_),
    .A1(\proj__5.net12 ));
 sg13g2_nand4_1 _281_ (.B(_053_),
    .C(_054_),
    .A(_052_),
    .Y(uo_out[6]),
    .D(_055_));
 sg13g2_tiehi \proj_13.flop1/_1__226  (.L_HI(net240));
 sg13g2_tielo \proj_13.flop2/_1__11  (.L_LO(net11));
 sg13g2_tielo \proj_13.flop3/_1__12  (.L_LO(net12));
 sg13g2_tielo \proj_14.flop1/dffsr_13  (.L_LO(net13));
 sg13g2_tielo \proj_14.flop1/_4__14  (.L_LO(net14));
 sg13g2_tielo \proj_14.flop10/dffsr_15  (.L_LO(net15));
 sg13g2_tielo \proj_14.flop10/_4__16  (.L_LO(net16));
 sg13g2_tielo \proj_14.flop11/dffsr_17  (.L_LO(net17));
 sg13g2_tielo \proj_14.flop11/_4__18  (.L_LO(net18));
 sg13g2_tielo \proj_14.flop12/dffsr_19  (.L_LO(net19));
 sg13g2_tielo \proj_14.flop12/_4__20  (.L_LO(net20));
 sg13g2_tielo \proj_14.flop13/dffsr_21  (.L_LO(net21));
 sg13g2_tielo \proj_14.flop13/_4__22  (.L_LO(net22));
 sg13g2_tielo \proj_14.flop14/dffsr_23  (.L_LO(net23));
 sg13g2_tielo \proj_14.flop14/_4__24  (.L_LO(net24));
 sg13g2_tielo \proj_14.flop15/dffsr_25  (.L_LO(net25));
 sg13g2_tielo \proj_14.flop15/_4__26  (.L_LO(net26));
 sg13g2_tielo \proj_14.flop16/dffsr_27  (.L_LO(net27));
 sg13g2_tielo \proj_14.flop16/_4__28  (.L_LO(net28));
 sg13g2_tielo \proj_14.flop17/dffsr_29  (.L_LO(net29));
 sg13g2_tielo \proj_14.flop17/_4__30  (.L_LO(net30));
 sg13g2_tielo \proj_14.flop18/dffsr_31  (.L_LO(net31));
 sg13g2_tielo \proj_14.flop18/_4__32  (.L_LO(net32));
 sg13g2_tielo \proj_14.flop19/dffsr_33  (.L_LO(net33));
 sg13g2_tielo \proj_14.flop19/_4__34  (.L_LO(net34));
 sg13g2_tielo \proj_14.flop2/dffsr_35  (.L_LO(net35));
 sg13g2_tielo \proj_14.flop2/_4__36  (.L_LO(net36));
 sg13g2_tielo \proj_14.flop20/dffsr_37  (.L_LO(net37));
 sg13g2_tielo \proj_14.flop20/_4__38  (.L_LO(net38));
 sg13g2_tielo \proj_14.flop21/dffsr_39  (.L_LO(net39));
 sg13g2_tielo \proj_14.flop21/_4__40  (.L_LO(net40));
 sg13g2_tielo \proj_14.flop22/dffsr_41  (.L_LO(net41));
 sg13g2_tielo \proj_14.flop22/_4__42  (.L_LO(net42));
 sg13g2_tielo \proj_14.flop23/dffsr_43  (.L_LO(net57));
 sg13g2_tielo \proj_14.flop23/_4__44  (.L_LO(net58));
 sg13g2_tielo \proj_14.flop24/dffsr_45  (.L_LO(net59));
 sg13g2_tielo \proj_14.flop24/_4__46  (.L_LO(net60));
 sg13g2_tielo \proj_14.flop25/dffsr_47  (.L_LO(net61));
 sg13g2_tielo \proj_14.flop25/_4__48  (.L_LO(net62));
 sg13g2_tielo \proj_14.flop26/dffsr_49  (.L_LO(net63));
 sg13g2_tielo \proj_14.flop26/_4__50  (.L_LO(net64));
 sg13g2_tielo \proj_14.flop27/dffsr_51  (.L_LO(net65));
 sg13g2_tielo \proj_14.flop27/_4__52  (.L_LO(net66));
 sg13g2_tielo \proj_14.flop28/_1__53  (.L_LO(net67));
 sg13g2_tielo \proj_14.flop29/dffsr_54  (.L_LO(net68));
 sg13g2_tielo \proj_14.flop29/_4__55  (.L_LO(net69));
 sg13g2_tielo \proj_14.flop3/dffsr_56  (.L_LO(net70));
 sg13g2_tielo \proj_14.flop3/_4__57  (.L_LO(net71));
 sg13g2_tielo \proj_14.flop30/dffsr_58  (.L_LO(net72));
 sg13g2_tielo \proj_14.flop30/_4__59  (.L_LO(net73));
 sg13g2_tielo \proj_14.flop31/dffsr_60  (.L_LO(net74));
 sg13g2_tielo \proj_14.flop32/dffsr_61  (.L_LO(net75));
 sg13g2_tielo \proj_14.flop32/_4__62  (.L_LO(net76));
 sg13g2_tielo \proj_14.flop33/dffsr_63  (.L_LO(net77));
 sg13g2_tielo \proj_14.flop33/_4__64  (.L_LO(net78));
 sg13g2_tielo \proj_14.flop34/dffsr_65  (.L_LO(net79));
 sg13g2_tielo \proj_14.flop34/_4__66  (.L_LO(net80));
 sg13g2_tielo \proj_14.flop35/dffsr_67  (.L_LO(net81));
 sg13g2_tielo \proj_14.flop35/_5__68  (.L_LO(net82));
 sg13g2_tielo \proj_14.flop36/dffsr_69  (.L_LO(net83));
 sg13g2_tielo \proj_14.flop36/_4__70  (.L_LO(net84));
 sg13g2_tielo \proj_14.flop37/dffsr_71  (.L_LO(net85));
 sg13g2_tielo \proj_14.flop37/_5__72  (.L_LO(net86));
 sg13g2_tielo \proj_14.flop4/dffsr_73  (.L_LO(net87));
 sg13g2_tielo \proj_14.flop4/_5__74  (.L_LO(net88));
 sg13g2_tielo \proj_14.flop46/_1__75  (.L_LO(net89));
 sg13g2_tielo \proj_14.flop47/_1__76  (.L_LO(net90));
 sg13g2_tielo \proj_14.flop48/_1__77  (.L_LO(net91));
 sg13g2_tielo \proj_14.flop49/_1__78  (.L_LO(net92));
 sg13g2_tielo \proj_14.flop5/dffsr_79  (.L_LO(net93));
 sg13g2_tielo \proj_14.flop5/_4__80  (.L_LO(net94));
 sg13g2_tielo \proj_14.flop50/_1__81  (.L_LO(net95));
 sg13g2_tielo \proj_14.flop51/_1__82  (.L_LO(net96));
 sg13g2_tielo \proj_14.flop52/_1__83  (.L_LO(net97));
 sg13g2_tielo \proj_14.flop53/_1__84  (.L_LO(net98));
 sg13g2_tielo \proj_14.flop54/_1__85  (.L_LO(net99));
 sg13g2_tielo \proj_14.flop55/_1__86  (.L_LO(net100));
 sg13g2_tielo \proj_14.flop56/_1__87  (.L_LO(net101));
 sg13g2_tielo \proj_14.flop6/dffsr_88  (.L_LO(net102));
 sg13g2_tielo \proj_14.flop6/_5__89  (.L_LO(net103));
 sg13g2_tielo \proj_14.flop7/dffsr_90  (.L_LO(net104));
 sg13g2_tielo \proj_14.flop7/_4__91  (.L_LO(net105));
 sg13g2_tielo \proj_14.flop8/dffsr_92  (.L_LO(net106));
 sg13g2_tielo \proj_14.flop8/_4__93  (.L_LO(net107));
 sg13g2_tielo \proj_14.flop9/dffsr_94  (.L_LO(net108));
 sg13g2_tielo \proj_14.flop9/_5__95  (.L_LO(net109));
 sg13g2_tielo \proj_14.not1/_0__96  (.L_LO(net110));
 sg13g2_tielo \proj_14.not5/_0__97  (.L_LO(net111));
 sg13g2_tielo \proj__4.flop1/dffsr_98  (.L_LO(net112));
 sg13g2_tielo \proj__4.flop1/_5__99  (.L_LO(net113));
 sg13g2_tielo \proj__4.flop2/dffsr_100  (.L_LO(net114));
 sg13g2_tielo \proj__4.flop2/_5__101  (.L_LO(net115));
 sg13g2_tielo \proj__4.flop3/dffsr_102  (.L_LO(net116));
 sg13g2_tielo \proj__4.flop3/_5__103  (.L_LO(net117));
 sg13g2_tielo \proj__4.flop4/dffsr_104  (.L_LO(net118));
 sg13g2_tielo \proj__4.flop4/_5__105  (.L_LO(net119));
 sg13g2_tielo \proj__4.flop5/dffsr_106  (.L_LO(net120));
 sg13g2_tielo \proj__4.flop5/_5__107  (.L_LO(net121));
 sg13g2_tielo \proj__4.flop6/dffsr_108  (.L_LO(net122));
 sg13g2_tielo \proj__4.flop6/_5__109  (.L_LO(net123));
 sg13g2_tielo \proj__4.flop8/dffsr_110  (.L_LO(net124));
 sg13g2_tielo \proj__4.flop8/_5__111  (.L_LO(net125));
 sg13g2_tielo \proj__4.flop9/dffsr_112  (.L_LO(net126));
 sg13g2_tielo \proj__4.flop9/_5__113  (.L_LO(net127));
 sg13g2_tielo \proj__7.flop1/_1__114  (.L_LO(net128));
 sg13g2_tielo \proj__7.flop2/_1__115  (.L_LO(net129));
 sg13g2_tielo \proj__9.flop1/dffsr_116  (.L_LO(net130));
 sg13g2_tielo \proj__9.flop1/_4__117  (.L_LO(net131));
 sg13g2_tielo \proj__9.not3/_0__118  (.L_LO(net132));
 sg13g2_tielo tt_um_wokwi_group_3_119 (.L_LO(net133));
 sg13g2_tielo tt_um_wokwi_group_3_120 (.L_LO(net134));
 sg13g2_tielo tt_um_wokwi_group_3_121 (.L_LO(net135));
 sg13g2_tielo tt_um_wokwi_group_3_122 (.L_LO(net136));
 sg13g2_tielo tt_um_wokwi_group_3_123 (.L_LO(net137));
 sg13g2_tielo tt_um_wokwi_group_3_124 (.L_LO(net138));
 sg13g2_tielo tt_um_wokwi_group_3_125 (.L_LO(net139));
 sg13g2_tielo tt_um_wokwi_group_3_126 (.L_LO(net140));
 sg13g2_tielo tt_um_wokwi_group_3_127 (.L_LO(net141));
 sg13g2_tielo tt_um_wokwi_group_3_128 (.L_LO(net142));
 sg13g2_tielo tt_um_wokwi_group_3_129 (.L_LO(net143));
 sg13g2_tielo tt_um_wokwi_group_3_130 (.L_LO(net144));
 sg13g2_tielo tt_um_wokwi_group_3_131 (.L_LO(net145));
 sg13g2_tielo tt_um_wokwi_group_3_132 (.L_LO(net146));
 sg13g2_tielo tt_um_wokwi_group_3_133 (.L_LO(net147));
 sg13g2_tielo tt_um_wokwi_group_3_134 (.L_LO(net148));
 sg13g2_tielo \proj_14.flop1/dffsr_135  (.L_LO(net149));
 sg13g2_mux2_1 \proj_10.mux2/_0_  (.A0(net52),
    .A1(net49),
    .S(net48),
    .X(\proj_10.net9 ));
 sg13g2_nand2_1 \proj_10.nand1/_0_  (.Y(\proj_10.net10 ),
    .A(\proj_10.nand1/b ),
    .B(net45));
 sg13g2_inv_1 \proj_10.not1/_0_  (.Y(\proj_10.net12 ),
    .A(net4));
 sg13g2_inv_1 \proj_10.not2/_0_  (.Y(\proj_10.net13 ),
    .A(net5));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(net2),
    .A(net44),
    .X(\proj_10.net11 ));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net49),
    .B(net51),
    .X(\proj_12.net18 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(net45),
    .B(net47),
    .X(\proj_12.net20 ));
 sg13g2_and2_1 \proj_12.and4/_0_  (.A(\proj_12.net19 ),
    .B(\proj_12.net18 ),
    .X(\proj_12.net21 ));
 sg13g2_and2_1 \proj_12.and5/_0_  (.A(net44),
    .B(net2),
    .X(\proj_12.net24 ));
 sg13g2_and2_1 \proj_12.and6/_0_  (.A(\proj_12.net23 ),
    .B(\proj_12.net22 ),
    .X(\proj_12.net25 ));
 sg13g2_and2_1 \proj_12.and7/_0_  (.A(net5),
    .B(net4),
    .X(\proj_12.net28 ));
 sg13g2_and2_1 \proj_12.and8/_0_  (.A(\proj_12.net27 ),
    .B(\proj_12.net26 ),
    .X(\proj_12.net29 ));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net22 ),
    .B(\proj_12.net21 ),
    .A(\proj_12.net20 ));
 sg13g2_or2_1 \proj_12.or2/_0_  (.X(\proj_12.net26 ),
    .B(\proj_12.net25 ),
    .A(\proj_12.net24 ));
 sg13g2_or2_1 \proj_12.or3/_0_  (.X(\proj_12.net13 ),
    .B(\proj_12.net29 ),
    .A(\proj_12.net28 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net51),
    .A(net49),
    .X(\proj_12.net9 ));
 sg13g2_xor2_1 \proj_12.xor2/_0_  (.B(net47),
    .A(net45),
    .X(\proj_12.net19 ));
 sg13g2_xor2_1 \proj_12.xor3/_0_  (.B(\proj_12.net19 ),
    .A(\proj_12.net18 ),
    .X(\proj_12.net10 ));
 sg13g2_xor2_1 \proj_12.xor4/_0_  (.B(net2),
    .A(net44),
    .X(\proj_12.net23 ));
 sg13g2_xor2_1 \proj_12.xor5/_0_  (.B(\proj_12.net23 ),
    .A(\proj_12.net22 ),
    .X(\proj_12.net11 ));
 sg13g2_xor2_1 \proj_12.xor6/_0_  (.B(net4),
    .A(net5),
    .X(\proj_12.net27 ));
 sg13g2_xor2_1 \proj_12.xor7/_0_  (.B(\proj_12.net27 ),
    .A(\proj_12.net26 ),
    .X(\proj_12.net12 ));
 sg13g2_dfrbp_1 \proj_13.flop1/_1_  (.CLK(net10),
    .RESET_B(net240),
    .D(net53),
    .Q_N(\proj_13.flop1/notq ),
    .Q(\proj_13.net12 ));
 sg13g2_tiehi \proj_13.flop2/_1__227  (.L_HI(net241));
 sg13g2_dfrbp_1 \proj_13.flop2/_1_  (.CLK(net11),
    .RESET_B(net241),
    .D(\proj_13.net12 ),
    .Q_N(\proj_13.flop2/notq ),
    .Q(\proj_13.net13 ));
 sg13g2_tiehi \proj_13.flop3/_1__228  (.L_HI(net242));
 sg13g2_dfrbp_1 \proj_13.flop3/_1_  (.CLK(net12),
    .RESET_B(net242),
    .D(\proj_13.net13 ),
    .Q_N(\proj_13.flop3/notq ),
    .Q(\proj_13.net8 ));
 sg13g2_tiehi \proj_14.flop28/_1__229  (.L_HI(net243));
 sg13g2_inv_1 \proj_13.not5/_0_  (.Y(\proj_13.net7 ),
    .A(\proj_13.net13 ));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(\proj_14.net30 ),
    .B(\proj_14.net33 ),
    .X(\proj_14.net58 ));
 sg13g2_and2_1 \proj_14.and10/_0_  (.A(\proj_14.net32 ),
    .B(\proj_14.net30 ),
    .X(\proj_14.net64 ));
 sg13g2_and2_1 \proj_14.and11/_0_  (.A(\proj_14.net40 ),
    .B(\proj_14.net43 ),
    .X(\proj_14.net68 ));
 sg13g2_and2_1 \proj_14.and12/_0_  (.A(\proj_14.net68 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net69 ));
 sg13g2_and2_1 \proj_14.and13/_0_  (.A(\proj_14.net68 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net70 ));
 sg13g2_and2_1 \proj_14.and14/_0_  (.A(\proj_14.net39 ),
    .B(\proj_14.net43 ),
    .X(\proj_14.net71 ));
 sg13g2_and2_1 \proj_14.and15/_0_  (.A(\proj_14.net71 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net72 ));
 sg13g2_and2_1 \proj_14.and16/_0_  (.A(\proj_14.net71 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net73 ));
 sg13g2_and2_1 \proj_14.and17/_0_  (.A(\proj_14.net74 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net75 ));
 sg13g2_and2_1 \proj_14.and18/_0_  (.A(\proj_14.net74 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net76 ));
 sg13g2_and2_1 \proj_14.and19/_0_  (.A(\proj_14.net42 ),
    .B(\proj_14.net39 ),
    .X(\proj_14.net77 ));
 sg13g2_and2_1 \proj_14.and2/_0_  (.A(\proj_14.net58 ),
    .B(\proj_14.net27 ),
    .X(\proj_14.net59 ));
 sg13g2_and2_1 \proj_14.and20/_0_  (.A(\proj_14.net42 ),
    .B(\proj_14.net40 ),
    .X(\proj_14.net74 ));
 sg13g2_and2_1 \proj_14.and21/_0_  (.A(\proj_14.net54 ),
    .B(\proj_14.net57 ),
    .X(\proj_14.net78 ));
 sg13g2_and2_1 \proj_14.and22/_0_  (.A(\proj_14.net78 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net79 ));
 sg13g2_and2_1 \proj_14.and23/_0_  (.A(\proj_14.net78 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net80 ));
 sg13g2_and2_1 \proj_14.and24/_0_  (.A(\proj_14.net53 ),
    .B(\proj_14.net57 ),
    .X(\proj_14.net81 ));
 sg13g2_and2_1 \proj_14.and25/_0_  (.A(\proj_14.net81 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net82 ));
 sg13g2_and2_1 \proj_14.and26/_0_  (.A(\proj_14.net81 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net83 ));
 sg13g2_and2_1 \proj_14.and27/_0_  (.A(\proj_14.net84 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net85 ));
 sg13g2_and2_1 \proj_14.and28/_0_  (.A(\proj_14.net84 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net86 ));
 sg13g2_and2_1 \proj_14.and29/_0_  (.A(\proj_14.net56 ),
    .B(\proj_14.net53 ),
    .X(\proj_14.net87 ));
 sg13g2_and2_1 \proj_14.and3/_0_  (.A(\proj_14.net58 ),
    .B(\proj_14.net26 ),
    .X(\proj_14.net60 ));
 sg13g2_and2_1 \proj_14.and30/_0_  (.A(\proj_14.net56 ),
    .B(\proj_14.net54 ),
    .X(\proj_14.net84 ));
 sg13g2_and2_1 \proj_14.and31/_0_  (.A(\proj_14.net105 ),
    .B(\proj_14.net110 ),
    .X(\proj_14.net116 ));
 sg13g2_and2_1 \proj_14.and32/_0_  (.A(\proj_14.net116 ),
    .B(\proj_14.net114 ),
    .X(\proj_14.net121 ));
 sg13g2_and2_1 \proj_14.and33/_0_  (.A(\proj_14.net121 ),
    .B(\proj_14.net119 ),
    .X(\proj_14.net126 ));
 sg13g2_and2_1 \proj_14.and34/_0_  (.A(\proj_14.net126 ),
    .B(\proj_14.net124 ),
    .X(\proj_14.net131 ));
 sg13g2_and2_1 \proj_14.and35/_0_  (.A(\proj_14.net137 ),
    .B(\proj_14.net135 ),
    .X(\proj_14.net142 ));
 sg13g2_and2_1 \proj_14.and36/_0_  (.A(\proj_14.net142 ),
    .B(\proj_14.net140 ),
    .X(\proj_14.net147 ));
 sg13g2_and2_1 \proj_14.and37/_0_  (.A(\proj_14.net147 ),
    .B(\proj_14.net145 ),
    .X(\proj_14.net152 ));
 sg13g2_and2_1 \proj_14.and38/_0_  (.A(\proj_14.net152 ),
    .B(\proj_14.net150 ),
    .X(\proj_14.net157 ));
 sg13g2_and2_1 \proj_14.and39/_0_  (.A(\proj_14.net131 ),
    .B(\proj_14.net129 ),
    .X(\proj_14.net137 ));
 sg13g2_and2_1 \proj_14.and4/_0_  (.A(\proj_14.net29 ),
    .B(\proj_14.net33 ),
    .X(\proj_14.net61 ));
 sg13g2_and2_1 \proj_14.and40/_0_  (.A(\proj_14.net157 ),
    .B(\proj_14.net155 ),
    .X(\proj_14.net162 ));
 sg13g2_and2_1 \proj_14.and41/_0_  (.A(\proj_14.net162 ),
    .B(\proj_14.net160 ),
    .X(\proj_14.net167 ));
 sg13g2_and2_1 \proj_14.and42/_0_  (.A(\proj_14.net167 ),
    .B(\proj_14.net165 ),
    .X(\proj_14.net172 ));
 sg13g2_and2_1 \proj_14.and43/_0_  (.A(\proj_14.net172 ),
    .B(\proj_14.net170 ),
    .X(\proj_14.net177 ));
 sg13g2_and2_1 \proj_14.and44/_0_  (.A(\proj_14.net193 ),
    .B(\proj_14.net192 ),
    .X(\proj_14.net194 ));
 sg13g2_and2_1 \proj_14.and45/_0_  (.A(\proj_14.net196 ),
    .B(\proj_14.net195 ),
    .X(\proj_14.net197 ));
 sg13g2_and2_1 \proj_14.and46/_0_  (.A(\proj_14.net199 ),
    .B(\proj_14.net198 ),
    .X(\proj_14.net200 ));
 sg13g2_and2_1 \proj_14.and47/_0_  (.A(\proj_14.net202 ),
    .B(\proj_14.net201 ),
    .X(\proj_14.net203 ));
 sg13g2_and2_1 \proj_14.and48/_0_  (.A(\proj_14.net203 ),
    .B(\proj_14.net200 ),
    .X(\proj_14.net204 ));
 sg13g2_and2_1 \proj_14.and49/_0_  (.A(\proj_14.net197 ),
    .B(\proj_14.net205 ),
    .X(\proj_14.net206 ));
 sg13g2_and2_1 \proj_14.and5/_0_  (.A(\proj_14.net61 ),
    .B(\proj_14.net27 ),
    .X(\proj_14.net62 ));
 sg13g2_and2_1 \proj_14.and50/_0_  (.A(\proj_14.net204 ),
    .B(\proj_14.net206 ),
    .X(\proj_14.net178 ));
 sg13g2_and2_1 \proj_14.and51/_0_  (.A(\proj_14.net59 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net234 ));
 sg13g2_and2_1 \proj_14.and52/_0_  (.A(\proj_14.net60 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net235 ));
 sg13g2_and2_1 \proj_14.and53/_0_  (.A(\proj_14.net62 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net236 ));
 sg13g2_and2_1 \proj_14.and54/_0_  (.A(\proj_14.net63 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net237 ));
 sg13g2_and2_1 \proj_14.and55/_0_  (.A(\proj_14.net65 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net238 ));
 sg13g2_and2_1 \proj_14.and57/_0_  (.A(\proj_14.net67 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net239 ));
 sg13g2_and2_1 \proj_14.and58/_0_  (.A(\proj_14.net59 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net240 ));
 sg13g2_and2_1 \proj_14.and59/_0_  (.A(\proj_14.net60 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net241 ));
 sg13g2_and2_1 \proj_14.and6/_0_  (.A(\proj_14.net61 ),
    .B(\proj_14.net26 ),
    .X(\proj_14.net63 ));
 sg13g2_and2_1 \proj_14.and60/_0_  (.A(\proj_14.net62 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net242 ));
 sg13g2_and2_1 \proj_14.and61/_0_  (.A(\proj_14.net63 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net243 ));
 sg13g2_and2_1 \proj_14.and62/_0_  (.A(\proj_14.net65 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net244 ));
 sg13g2_and2_1 \proj_14.and63/_0_  (.A(\proj_14.net66 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net245 ));
 sg13g2_and2_1 \proj_14.and64/_0_  (.A(\proj_14.net182 ),
    .B(\proj_14.net181 ),
    .X(\proj_14.net183 ));
 sg13g2_and2_1 \proj_14.and65/_0_  (.A(\proj_14.net67 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net246 ));
 sg13g2_and2_1 \proj_14.and66/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net235 ),
    .X(\proj_14.net249 ));
 sg13g2_and2_1 \proj_14.and67/_0_  (.A(\proj_14.net235 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net248 ));
 sg13g2_and2_1 \proj_14.and68/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net238 ),
    .X(\proj_14.net252 ));
 sg13g2_and2_1 \proj_14.and69/_0_  (.A(\proj_14.net238 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net254 ));
 sg13g2_and2_1 \proj_14.and7/_0_  (.A(\proj_14.net64 ),
    .B(\proj_14.net27 ),
    .X(\proj_14.net65 ));
 sg13g2_and2_1 \proj_14.and70/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net239 ),
    .X(\proj_14.net258 ));
 sg13g2_and2_1 \proj_14.and71/_0_  (.A(\proj_14.net239 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net256 ));
 sg13g2_and2_1 \proj_14.and72/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net242 ),
    .X(\proj_14.net265 ));
 sg13g2_and2_1 \proj_14.and73/_0_  (.A(\proj_14.net242 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net261 ));
 sg13g2_and2_1 \proj_14.and74/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net245 ),
    .X(\proj_14.net267 ));
 sg13g2_and2_1 \proj_14.and75/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net246 ),
    .X(\proj_14.net259 ));
 sg13g2_and2_1 \proj_14.and76/_0_  (.A(\proj_14.net246 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net269 ));
 sg13g2_and2_1 \proj_14.and77/_0_  (.A(\proj_14.net194 ),
    .B(\proj_14.net135 ),
    .X(\proj_14.net205 ));
 sg13g2_and2_1 \proj_14.and8/_0_  (.A(\proj_14.net64 ),
    .B(\proj_14.net26 ),
    .X(\proj_14.net66 ));
 sg13g2_and2_1 \proj_14.and9/_0_  (.A(\proj_14.net32 ),
    .B(\proj_14.net29 ),
    .X(\proj_14.net67 ));
 sg13g2_inv_1 \proj_14.flop1/_4_  (.Y(\proj_14.flop1/_1_ ),
    .A(net14));
 sg13g2_inv_1 \proj_14.flop1/_5_  (.Y(\proj_14.flop1/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop1/dffsr_136  (.L_LO(net150));
 sg13g2_tielo \proj_14.flop10/dffsr_137  (.L_LO(net151));
 sg13g2_sdfbbp_1 \proj_14.flop1/dffsr  (.Q(\proj_14.net26 ),
    .Q_N(\proj_14.net27 ),
    .RESET_B(\proj_14.flop1/_0_ ),
    .SET_B(\proj_14.flop1/_1_ ),
    .D(\proj_14.net23 ),
    .SCE(net150),
    .SCD(net149),
    .CLK(net13));
 sg13g2_inv_1 \proj_14.flop10/_4_  (.Y(\proj_14.flop10/_1_ ),
    .A(net16));
 sg13g2_inv_1 \proj_14.flop10/_5_  (.Y(\proj_14.flop10/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop10/dffsr_138  (.L_LO(net152));
 sg13g2_tielo \proj_14.flop11/dffsr_139  (.L_LO(net153));
 sg13g2_sdfbbp_1 \proj_14.flop10/dffsr  (.Q(\proj_14.net105 ),
    .Q_N(\proj_14.net106 ),
    .RESET_B(\proj_14.flop10/_0_ ),
    .SET_B(\proj_14.flop10/_1_ ),
    .D(\proj_14.net102 ),
    .SCE(net152),
    .SCD(net151),
    .CLK(net15));
 sg13g2_inv_1 \proj_14.flop11/_4_  (.Y(\proj_14.flop11/_1_ ),
    .A(net18));
 sg13g2_inv_1 \proj_14.flop11/_5_  (.Y(\proj_14.flop11/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop11/dffsr_140  (.L_LO(net154));
 sg13g2_tielo \proj_14.flop12/dffsr_141  (.L_LO(net155));
 sg13g2_sdfbbp_1 \proj_14.flop11/dffsr  (.Q(\proj_14.net110 ),
    .Q_N(\proj_14.net111 ),
    .RESET_B(\proj_14.flop11/_0_ ),
    .SET_B(\proj_14.flop11/_1_ ),
    .D(\proj_14.net108 ),
    .SCE(net154),
    .SCD(net153),
    .CLK(net17));
 sg13g2_inv_1 \proj_14.flop12/_4_  (.Y(\proj_14.flop12/_1_ ),
    .A(net20));
 sg13g2_inv_1 \proj_14.flop12/_5_  (.Y(\proj_14.flop12/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop12/dffsr_142  (.L_LO(net156));
 sg13g2_tielo \proj_14.flop13/dffsr_143  (.L_LO(net157));
 sg13g2_sdfbbp_1 \proj_14.flop12/dffsr  (.Q(\proj_14.net114 ),
    .Q_N(\proj_14.net115 ),
    .RESET_B(\proj_14.flop12/_0_ ),
    .SET_B(\proj_14.flop12/_1_ ),
    .D(\proj_14.net112 ),
    .SCE(net156),
    .SCD(net155),
    .CLK(net19));
 sg13g2_inv_1 \proj_14.flop13/_4_  (.Y(\proj_14.flop13/_1_ ),
    .A(net22));
 sg13g2_inv_1 \proj_14.flop13/_5_  (.Y(\proj_14.flop13/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop13/dffsr_144  (.L_LO(net158));
 sg13g2_tielo \proj_14.flop14/dffsr_145  (.L_LO(net159));
 sg13g2_sdfbbp_1 \proj_14.flop13/dffsr  (.Q(\proj_14.net119 ),
    .Q_N(\proj_14.net120 ),
    .RESET_B(\proj_14.flop13/_0_ ),
    .SET_B(\proj_14.flop13/_1_ ),
    .D(\proj_14.net117 ),
    .SCE(net158),
    .SCD(net157),
    .CLK(net21));
 sg13g2_inv_1 \proj_14.flop14/_4_  (.Y(\proj_14.flop14/_1_ ),
    .A(net24));
 sg13g2_inv_1 \proj_14.flop14/_5_  (.Y(\proj_14.flop14/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop14/dffsr_146  (.L_LO(net160));
 sg13g2_tielo \proj_14.flop15/dffsr_147  (.L_LO(net161));
 sg13g2_sdfbbp_1 \proj_14.flop14/dffsr  (.Q(\proj_14.net124 ),
    .Q_N(\proj_14.net125 ),
    .RESET_B(\proj_14.flop14/_0_ ),
    .SET_B(\proj_14.flop14/_1_ ),
    .D(\proj_14.net122 ),
    .SCE(net160),
    .SCD(net159),
    .CLK(net23));
 sg13g2_inv_1 \proj_14.flop15/_4_  (.Y(\proj_14.flop15/_1_ ),
    .A(net26));
 sg13g2_inv_1 \proj_14.flop15/_5_  (.Y(\proj_14.flop15/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop15/dffsr_148  (.L_LO(net162));
 sg13g2_tielo \proj_14.flop16/dffsr_149  (.L_LO(net163));
 sg13g2_sdfbbp_1 \proj_14.flop15/dffsr  (.Q(\proj_14.net129 ),
    .Q_N(\proj_14.net130 ),
    .RESET_B(\proj_14.flop15/_0_ ),
    .SET_B(\proj_14.flop15/_1_ ),
    .D(\proj_14.net127 ),
    .SCE(net162),
    .SCD(net161),
    .CLK(net25));
 sg13g2_inv_1 \proj_14.flop16/_4_  (.Y(\proj_14.flop16/_1_ ),
    .A(net28));
 sg13g2_inv_1 \proj_14.flop16/_5_  (.Y(\proj_14.flop16/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop16/dffsr_150  (.L_LO(net164));
 sg13g2_tielo \proj_14.flop17/dffsr_151  (.L_LO(net165));
 sg13g2_sdfbbp_1 \proj_14.flop16/dffsr  (.Q(\proj_14.net135 ),
    .Q_N(\proj_14.net136 ),
    .RESET_B(\proj_14.flop16/_0_ ),
    .SET_B(\proj_14.flop16/_1_ ),
    .D(\proj_14.net133 ),
    .SCE(net164),
    .SCD(net163),
    .CLK(net27));
 sg13g2_inv_1 \proj_14.flop17/_4_  (.Y(\proj_14.flop17/_1_ ),
    .A(net30));
 sg13g2_inv_1 \proj_14.flop17/_5_  (.Y(\proj_14.flop17/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop17/dffsr_152  (.L_LO(net166));
 sg13g2_tielo \proj_14.flop18/dffsr_153  (.L_LO(net167));
 sg13g2_sdfbbp_1 \proj_14.flop17/dffsr  (.Q(\proj_14.net140 ),
    .Q_N(\proj_14.net141 ),
    .RESET_B(\proj_14.flop17/_0_ ),
    .SET_B(\proj_14.flop17/_1_ ),
    .D(\proj_14.net138 ),
    .SCE(net166),
    .SCD(net165),
    .CLK(net29));
 sg13g2_inv_1 \proj_14.flop18/_4_  (.Y(\proj_14.flop18/_1_ ),
    .A(net32));
 sg13g2_inv_1 \proj_14.flop18/_5_  (.Y(\proj_14.flop18/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop18/dffsr_154  (.L_LO(net168));
 sg13g2_tielo \proj_14.flop19/dffsr_155  (.L_LO(net169));
 sg13g2_sdfbbp_1 \proj_14.flop18/dffsr  (.Q(\proj_14.net145 ),
    .Q_N(\proj_14.net146 ),
    .RESET_B(\proj_14.flop18/_0_ ),
    .SET_B(\proj_14.flop18/_1_ ),
    .D(\proj_14.net143 ),
    .SCE(net168),
    .SCD(net167),
    .CLK(net31));
 sg13g2_inv_1 \proj_14.flop19/_4_  (.Y(\proj_14.flop19/_1_ ),
    .A(net34));
 sg13g2_inv_1 \proj_14.flop19/_5_  (.Y(\proj_14.flop19/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop19/dffsr_156  (.L_LO(net170));
 sg13g2_tielo \proj_14.flop2/dffsr_157  (.L_LO(net171));
 sg13g2_sdfbbp_1 \proj_14.flop19/dffsr  (.Q(\proj_14.net150 ),
    .Q_N(\proj_14.net151 ),
    .RESET_B(\proj_14.flop19/_0_ ),
    .SET_B(\proj_14.flop19/_1_ ),
    .D(\proj_14.net148 ),
    .SCE(net170),
    .SCD(net169),
    .CLK(net33));
 sg13g2_inv_1 \proj_14.flop2/_4_  (.Y(\proj_14.flop2/_1_ ),
    .A(net36));
 sg13g2_inv_1 \proj_14.flop2/_5_  (.Y(\proj_14.flop2/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop2/dffsr_158  (.L_LO(net172));
 sg13g2_tielo \proj_14.flop20/dffsr_159  (.L_LO(net173));
 sg13g2_sdfbbp_1 \proj_14.flop2/dffsr  (.Q(\proj_14.net29 ),
    .Q_N(\proj_14.net30 ),
    .RESET_B(\proj_14.flop2/_0_ ),
    .SET_B(\proj_14.flop2/_1_ ),
    .D(\proj_14.net28 ),
    .SCE(net172),
    .SCD(net171),
    .CLK(net35));
 sg13g2_inv_1 \proj_14.flop20/_4_  (.Y(\proj_14.flop20/_1_ ),
    .A(net38));
 sg13g2_inv_1 \proj_14.flop20/_5_  (.Y(\proj_14.flop20/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop20/dffsr_160  (.L_LO(net174));
 sg13g2_tielo \proj_14.flop21/dffsr_161  (.L_LO(net175));
 sg13g2_sdfbbp_1 \proj_14.flop20/dffsr  (.Q(\proj_14.net155 ),
    .Q_N(\proj_14.net156 ),
    .RESET_B(\proj_14.flop20/_0_ ),
    .SET_B(\proj_14.flop20/_1_ ),
    .D(\proj_14.net153 ),
    .SCE(net174),
    .SCD(net173),
    .CLK(net37));
 sg13g2_inv_1 \proj_14.flop21/_4_  (.Y(\proj_14.flop21/_1_ ),
    .A(net40));
 sg13g2_inv_1 \proj_14.flop21/_5_  (.Y(\proj_14.flop21/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop21/dffsr_162  (.L_LO(net176));
 sg13g2_tielo \proj_14.flop22/dffsr_163  (.L_LO(net177));
 sg13g2_sdfbbp_1 \proj_14.flop21/dffsr  (.Q(\proj_14.net160 ),
    .Q_N(\proj_14.net161 ),
    .RESET_B(\proj_14.flop21/_0_ ),
    .SET_B(\proj_14.flop21/_1_ ),
    .D(\proj_14.net158 ),
    .SCE(net176),
    .SCD(net175),
    .CLK(net39));
 sg13g2_inv_1 \proj_14.flop22/_4_  (.Y(\proj_14.flop22/_1_ ),
    .A(net42));
 sg13g2_inv_1 \proj_14.flop22/_5_  (.Y(\proj_14.flop22/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop22/dffsr_164  (.L_LO(net178));
 sg13g2_tielo \proj_14.flop23/dffsr_165  (.L_LO(net179));
 sg13g2_sdfbbp_1 \proj_14.flop22/dffsr  (.Q(\proj_14.net165 ),
    .Q_N(\proj_14.net166 ),
    .RESET_B(\proj_14.flop22/_0_ ),
    .SET_B(\proj_14.flop22/_1_ ),
    .D(\proj_14.net163 ),
    .SCE(net178),
    .SCD(net177),
    .CLK(net41));
 sg13g2_inv_1 \proj_14.flop23/_4_  (.Y(\proj_14.flop23/_1_ ),
    .A(net58));
 sg13g2_inv_1 \proj_14.flop23/_5_  (.Y(\proj_14.flop23/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop23/dffsr_166  (.L_LO(net180));
 sg13g2_tielo \proj_14.flop24/dffsr_167  (.L_LO(net181));
 sg13g2_sdfbbp_1 \proj_14.flop23/dffsr  (.Q(\proj_14.net170 ),
    .Q_N(\proj_14.net171 ),
    .RESET_B(\proj_14.flop23/_0_ ),
    .SET_B(\proj_14.flop23/_1_ ),
    .D(\proj_14.net168 ),
    .SCE(net180),
    .SCD(net179),
    .CLK(net57));
 sg13g2_inv_1 \proj_14.flop24/_4_  (.Y(\proj_14.flop24/_1_ ),
    .A(net60));
 sg13g2_inv_1 \proj_14.flop24/_5_  (.Y(\proj_14.flop24/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop24/dffsr_168  (.L_LO(net182));
 sg13g2_tielo \proj_14.flop25/dffsr_169  (.L_LO(net183));
 sg13g2_sdfbbp_1 \proj_14.flop24/dffsr  (.Q(\proj_14.net175 ),
    .Q_N(\proj_14.net176 ),
    .RESET_B(\proj_14.flop24/_0_ ),
    .SET_B(\proj_14.flop24/_1_ ),
    .D(\proj_14.net173 ),
    .SCE(net182),
    .SCD(net181),
    .CLK(net59));
 sg13g2_inv_1 \proj_14.flop25/_4_  (.Y(\proj_14.flop25/_1_ ),
    .A(net62));
 sg13g2_inv_1 \proj_14.flop25/_5_  (.Y(\proj_14.flop25/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop25/dffsr_170  (.L_LO(net184));
 sg13g2_tielo \proj_14.flop26/dffsr_171  (.L_LO(net185));
 sg13g2_sdfbbp_1 \proj_14.flop25/dffsr  (.Q(\proj_14.net180 ),
    .Q_N(\proj_14.flop25/notq ),
    .RESET_B(\proj_14.flop25/_0_ ),
    .SET_B(\proj_14.flop25/_1_ ),
    .D(\proj_14.net178 ),
    .SCE(net184),
    .SCD(net183),
    .CLK(net61));
 sg13g2_inv_1 \proj_14.flop26/_4_  (.Y(\proj_14.flop26/_1_ ),
    .A(net64));
 sg13g2_inv_1 \proj_14.flop26/_5_  (.Y(\proj_14.flop26/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop26/dffsr_172  (.L_LO(net186));
 sg13g2_tielo \proj_14.flop27/dffsr_173  (.L_LO(net187));
 sg13g2_sdfbbp_1 \proj_14.flop26/dffsr  (.Q(\proj_14.net181 ),
    .Q_N(\proj_14.flop26/notq ),
    .RESET_B(\proj_14.flop26/_0_ ),
    .SET_B(\proj_14.flop26/_1_ ),
    .D(\proj_14.net180 ),
    .SCE(net186),
    .SCD(net185),
    .CLK(net63));
 sg13g2_inv_1 \proj_14.flop27/_4_  (.Y(\proj_14.flop27/_1_ ),
    .A(net66));
 sg13g2_inv_1 \proj_14.flop27/_5_  (.Y(\proj_14.flop27/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop27/dffsr_174  (.L_LO(net188));
 sg13g2_tielo \proj_14.flop29/dffsr_175  (.L_LO(net189));
 sg13g2_sdfbbp_1 \proj_14.flop27/dffsr  (.Q(\proj_14.flop27/q ),
    .Q_N(\proj_14.net182 ),
    .RESET_B(\proj_14.flop27/_0_ ),
    .SET_B(\proj_14.flop27/_1_ ),
    .D(\proj_14.net181 ),
    .SCE(net188),
    .SCD(net187),
    .CLK(net65));
 sg13g2_dfrbp_1 \proj_14.flop28/_1_  (.CLK(net67),
    .RESET_B(net243),
    .D(\proj_14.net95 ),
    .Q_N(\proj_14.flop28/notq ),
    .Q(\proj_14.net11 ));
 sg13g2_tiehi \proj_14.flop46/_1__230  (.L_HI(net244));
 sg13g2_inv_1 \proj_14.flop29/_4_  (.Y(\proj_14.flop29/_1_ ),
    .A(net69));
 sg13g2_inv_1 \proj_14.flop29/_5_  (.Y(\proj_14.flop29/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop29/dffsr_176  (.L_LO(net190));
 sg13g2_tielo \proj_14.flop3/dffsr_177  (.L_LO(net191));
 sg13g2_sdfbbp_1 \proj_14.flop29/dffsr  (.Q(\proj_14.net209 ),
    .Q_N(\proj_14.net210 ),
    .RESET_B(\proj_14.flop29/_0_ ),
    .SET_B(\proj_14.flop29/_1_ ),
    .D(\proj_14.net207 ),
    .SCE(net190),
    .SCD(net189),
    .CLK(net68));
 sg13g2_inv_1 \proj_14.flop3/_4_  (.Y(\proj_14.flop3/_1_ ),
    .A(net71));
 sg13g2_inv_1 \proj_14.flop3/_5_  (.Y(\proj_14.flop3/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop3/dffsr_178  (.L_LO(net192));
 sg13g2_tielo \proj_14.flop30/dffsr_179  (.L_LO(net193));
 sg13g2_sdfbbp_1 \proj_14.flop3/dffsr  (.Q(\proj_14.net32 ),
    .Q_N(\proj_14.net33 ),
    .RESET_B(\proj_14.flop3/_0_ ),
    .SET_B(\proj_14.flop3/_1_ ),
    .D(\proj_14.net31 ),
    .SCE(net192),
    .SCD(net191),
    .CLK(net70));
 sg13g2_inv_1 \proj_14.flop30/_4_  (.Y(\proj_14.flop30/_1_ ),
    .A(net73));
 sg13g2_inv_1 \proj_14.flop30/_5_  (.Y(\proj_14.flop30/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop30/dffsr_180  (.L_LO(net194));
 sg13g2_tielo \proj_14.flop31/dffsr_181  (.L_LO(net195));
 sg13g2_sdfbbp_1 \proj_14.flop30/dffsr  (.Q(\proj_14.net214 ),
    .Q_N(\proj_14.net215 ),
    .RESET_B(\proj_14.flop30/_0_ ),
    .SET_B(\proj_14.flop30/_1_ ),
    .D(\proj_14.net212 ),
    .SCE(net194),
    .SCD(net193),
    .CLK(net72));
 sg13g2_inv_1 \proj_14.flop31/_4_  (.Y(\proj_14.flop31/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop31/_5_  (.Y(\proj_14.flop31/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop31/dffsr_182  (.L_LO(net196));
 sg13g2_tielo \proj_14.flop32/dffsr_183  (.L_LO(net197));
 sg13g2_sdfbbp_1 \proj_14.flop31/dffsr  (.Q(\proj_14.net217 ),
    .Q_N(\proj_14.flop31/notq ),
    .RESET_B(\proj_14.flop31/_0_ ),
    .SET_B(\proj_14.flop31/_1_ ),
    .D(\proj_14.net216 ),
    .SCE(net196),
    .SCD(net195),
    .CLK(net74));
 sg13g2_inv_1 \proj_14.flop32/_4_  (.Y(\proj_14.flop32/_1_ ),
    .A(net76));
 sg13g2_inv_1 \proj_14.flop32/_5_  (.Y(\proj_14.flop32/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop32/dffsr_184  (.L_LO(net198));
 sg13g2_tielo \proj_14.flop33/dffsr_185  (.L_LO(net199));
 sg13g2_sdfbbp_1 \proj_14.flop32/dffsr  (.Q(\proj_14.net219 ),
    .Q_N(\proj_14.flop32/notq ),
    .RESET_B(\proj_14.flop32/_0_ ),
    .SET_B(\proj_14.flop32/_1_ ),
    .D(\proj_14.net218 ),
    .SCE(net198),
    .SCD(net197),
    .CLK(net75));
 sg13g2_inv_1 \proj_14.flop33/_4_  (.Y(\proj_14.flop33/_1_ ),
    .A(net78));
 sg13g2_inv_1 \proj_14.flop33/_5_  (.Y(\proj_14.flop33/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop33/dffsr_186  (.L_LO(net200));
 sg13g2_tielo \proj_14.flop34/dffsr_187  (.L_LO(net201));
 sg13g2_sdfbbp_1 \proj_14.flop33/dffsr  (.Q(\proj_14.net221 ),
    .Q_N(\proj_14.flop33/notq ),
    .RESET_B(\proj_14.flop33/_0_ ),
    .SET_B(\proj_14.flop33/_1_ ),
    .D(\proj_14.net220 ),
    .SCE(net200),
    .SCD(net199),
    .CLK(net77));
 sg13g2_inv_1 \proj_14.flop34/_4_  (.Y(\proj_14.flop34/_1_ ),
    .A(net80));
 sg13g2_inv_1 \proj_14.flop34/_5_  (.Y(\proj_14.flop34/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop34/dffsr_188  (.L_LO(net202));
 sg13g2_tielo \proj_14.flop35/dffsr_189  (.L_LO(net203));
 sg13g2_sdfbbp_1 \proj_14.flop34/dffsr  (.Q(\proj_14.net223 ),
    .Q_N(\proj_14.flop34/notq ),
    .RESET_B(\proj_14.flop34/_0_ ),
    .SET_B(\proj_14.flop34/_1_ ),
    .D(\proj_14.net222 ),
    .SCE(net202),
    .SCD(net201),
    .CLK(net79));
 sg13g2_inv_1 \proj_14.flop35/_4_  (.Y(\proj_14.flop35/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop35/_5_  (.Y(\proj_14.flop35/_0_ ),
    .A(net82));
 sg13g2_tielo \proj_14.flop35/dffsr_190  (.L_LO(net204));
 sg13g2_tielo \proj_14.flop36/dffsr_191  (.L_LO(net205));
 sg13g2_sdfbbp_1 \proj_14.flop35/dffsr  (.Q(\proj_14.net226 ),
    .Q_N(\proj_14.flop35/notq ),
    .RESET_B(\proj_14.flop35/_0_ ),
    .SET_B(\proj_14.flop35/_1_ ),
    .D(\proj_14.net224 ),
    .SCE(net204),
    .SCD(net203),
    .CLK(net81));
 sg13g2_inv_1 \proj_14.flop36/_4_  (.Y(\proj_14.flop36/_1_ ),
    .A(net84));
 sg13g2_inv_1 \proj_14.flop36/_5_  (.Y(\proj_14.flop36/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop36/dffsr_192  (.L_LO(net206));
 sg13g2_tielo \proj_14.flop37/dffsr_193  (.L_LO(net207));
 sg13g2_sdfbbp_1 \proj_14.flop36/dffsr  (.Q(\proj_14.net228 ),
    .Q_N(\proj_14.flop36/notq ),
    .RESET_B(\proj_14.flop36/_0_ ),
    .SET_B(\proj_14.flop36/_1_ ),
    .D(\proj_14.net227 ),
    .SCE(net206),
    .SCD(net205),
    .CLK(net83));
 sg13g2_inv_1 \proj_14.flop37/_4_  (.Y(\proj_14.flop37/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop37/_5_  (.Y(\proj_14.flop37/_0_ ),
    .A(net86));
 sg13g2_tielo \proj_14.flop37/dffsr_194  (.L_LO(net208));
 sg13g2_tielo \proj_14.flop4/dffsr_195  (.L_LO(net209));
 sg13g2_sdfbbp_1 \proj_14.flop37/dffsr  (.Q(\proj_14.net231 ),
    .Q_N(\proj_14.flop37/notq ),
    .RESET_B(\proj_14.flop37/_0_ ),
    .SET_B(\proj_14.flop37/_1_ ),
    .D(\proj_14.net229 ),
    .SCE(net208),
    .SCD(net207),
    .CLK(net85));
 sg13g2_inv_1 \proj_14.flop4/_4_  (.Y(\proj_14.flop4/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop4/_5_  (.Y(\proj_14.flop4/_0_ ),
    .A(net88));
 sg13g2_tielo \proj_14.flop4/dffsr_196  (.L_LO(net210));
 sg13g2_tielo \proj_14.flop5/dffsr_197  (.L_LO(net211));
 sg13g2_sdfbbp_1 \proj_14.flop4/dffsr  (.Q(\proj_14.net36 ),
    .Q_N(\proj_14.net37 ),
    .RESET_B(\proj_14.flop4/_0_ ),
    .SET_B(\proj_14.flop4/_1_ ),
    .D(\proj_14.net34 ),
    .SCE(net210),
    .SCD(net209),
    .CLK(net87));
 sg13g2_dfrbp_1 \proj_14.flop46/_1_  (.CLK(net89),
    .RESET_B(net244),
    .D(\proj_14.net96 ),
    .Q_N(\proj_14.flop46/notq ),
    .Q(\proj_14.net12 ));
 sg13g2_tiehi \proj_14.flop47/_1__231  (.L_HI(net245));
 sg13g2_dfrbp_1 \proj_14.flop47/_1_  (.CLK(net90),
    .RESET_B(net245),
    .D(\proj_14.net97 ),
    .Q_N(\proj_14.flop47/notq ),
    .Q(\proj_14.net13 ));
 sg13g2_tiehi \proj_14.flop48/_1__232  (.L_HI(net246));
 sg13g2_dfrbp_1 \proj_14.flop48/_1_  (.CLK(net91),
    .RESET_B(net246),
    .D(\proj_14.net98 ),
    .Q_N(\proj_14.flop48/notq ),
    .Q(\proj_14.net14 ));
 sg13g2_tiehi \proj_14.flop49/_1__233  (.L_HI(net247));
 sg13g2_dfrbp_1 \proj_14.flop49/_1_  (.CLK(net92),
    .RESET_B(net247),
    .D(\proj_14.net99 ),
    .Q_N(\proj_14.flop49/notq ),
    .Q(\proj_14.net15 ));
 sg13g2_tiehi \proj_14.flop50/_1__234  (.L_HI(net248));
 sg13g2_inv_1 \proj_14.flop5/_4_  (.Y(\proj_14.flop5/_1_ ),
    .A(net94));
 sg13g2_inv_1 \proj_14.flop5/_5_  (.Y(\proj_14.flop5/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop5/dffsr_198  (.L_LO(net212));
 sg13g2_tielo \proj_14.flop6/dffsr_199  (.L_LO(net213));
 sg13g2_sdfbbp_1 \proj_14.flop5/dffsr  (.Q(\proj_14.net39 ),
    .Q_N(\proj_14.net40 ),
    .RESET_B(\proj_14.flop5/_0_ ),
    .SET_B(\proj_14.flop5/_1_ ),
    .D(\proj_14.net38 ),
    .SCE(net212),
    .SCD(net211),
    .CLK(net93));
 sg13g2_dfrbp_1 \proj_14.flop50/_1_  (.CLK(net95),
    .RESET_B(net248),
    .D(\proj_14.net100 ),
    .Q_N(\proj_14.flop50/notq ),
    .Q(\proj_14.net16 ));
 sg13g2_tiehi \proj_14.flop51/_1__235  (.L_HI(net249));
 sg13g2_dfrbp_1 \proj_14.flop51/_1_  (.CLK(net96),
    .RESET_B(net249),
    .D(\proj_14.net101 ),
    .Q_N(\proj_14.flop51/notq ),
    .Q(\proj_14.net17 ));
 sg13g2_tiehi \proj_14.flop52/_1__236  (.L_HI(net250));
 sg13g2_dfrbp_1 \proj_14.flop52/_1_  (.CLK(net97),
    .RESET_B(net250),
    .D(\proj_14.net183 ),
    .Q_N(\proj_14.flop52/notq ),
    .Q(\proj_14.net45 ));
 sg13g2_tiehi \proj_14.flop53/_1__237  (.L_HI(net251));
 sg13g2_dfrbp_1 \proj_14.flop53/_1_  (.CLK(net98),
    .RESET_B(net251),
    .D(\proj_14.net275 ),
    .Q_N(\proj_14.flop53/notq ),
    .Q(\proj_14.net44 ));
 sg13g2_tiehi \proj_14.flop54/_1__238  (.L_HI(net252));
 sg13g2_dfrbp_1 \proj_14.flop54/_1_  (.CLK(net99),
    .RESET_B(net252),
    .D(\proj_14.net277 ),
    .Q_N(\proj_14.flop54/notq ),
    .Q(\proj_14.net46 ));
 sg13g2_tiehi \proj_14.flop55/_1__239  (.L_HI(net253));
 sg13g2_dfrbp_1 \proj_14.flop55/_1_  (.CLK(net100),
    .RESET_B(net253),
    .D(\proj_14.net280 ),
    .Q_N(\proj_14.flop55/notq ),
    .Q(\proj_14.net47 ));
 sg13g2_tiehi \proj_14.flop56/_1__240  (.L_HI(net254));
 sg13g2_dfrbp_1 \proj_14.flop56/_1_  (.CLK(net101),
    .RESET_B(net254),
    .D(\proj_14.net281 ),
    .Q_N(\proj_14.flop56/notq ),
    .Q(\proj_14.net211 ));
 sg13g2_tiehi \proj__7.flop1/_1__241  (.L_HI(net255));
 sg13g2_inv_1 \proj_14.flop6/_4_  (.Y(\proj_14.flop6/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop6/_5_  (.Y(\proj_14.flop6/_0_ ),
    .A(net103));
 sg13g2_tielo \proj_14.flop6/dffsr_200  (.L_LO(net214));
 sg13g2_tielo \proj_14.flop7/dffsr_201  (.L_LO(net215));
 sg13g2_sdfbbp_1 \proj_14.flop6/dffsr  (.Q(\proj_14.net42 ),
    .Q_N(\proj_14.net43 ),
    .RESET_B(\proj_14.flop6/_0_ ),
    .SET_B(\proj_14.flop6/_1_ ),
    .D(\proj_14.net41 ),
    .SCE(net214),
    .SCD(net213),
    .CLK(net102));
 sg13g2_inv_1 \proj_14.flop7/_4_  (.Y(\proj_14.flop7/_1_ ),
    .A(net105));
 sg13g2_inv_1 \proj_14.flop7/_5_  (.Y(\proj_14.flop7/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop7/dffsr_202  (.L_LO(net216));
 sg13g2_tielo \proj_14.flop8/dffsr_203  (.L_LO(net217));
 sg13g2_sdfbbp_1 \proj_14.flop7/dffsr  (.Q(\proj_14.net50 ),
    .Q_N(\proj_14.net51 ),
    .RESET_B(\proj_14.flop7/_0_ ),
    .SET_B(\proj_14.flop7/_1_ ),
    .D(\proj_14.net48 ),
    .SCE(net216),
    .SCD(net215),
    .CLK(net104));
 sg13g2_inv_1 \proj_14.flop8/_4_  (.Y(\proj_14.flop8/_1_ ),
    .A(net107));
 sg13g2_inv_1 \proj_14.flop8/_5_  (.Y(\proj_14.flop8/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop8/dffsr_204  (.L_LO(net218));
 sg13g2_tielo \proj_14.flop9/dffsr_205  (.L_LO(net219));
 sg13g2_sdfbbp_1 \proj_14.flop8/dffsr  (.Q(\proj_14.net53 ),
    .Q_N(\proj_14.net54 ),
    .RESET_B(\proj_14.flop8/_0_ ),
    .SET_B(\proj_14.flop8/_1_ ),
    .D(\proj_14.net52 ),
    .SCE(net218),
    .SCD(net217),
    .CLK(net106));
 sg13g2_inv_1 \proj_14.flop9/_4_  (.Y(\proj_14.flop9/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop9/_5_  (.Y(\proj_14.flop9/_0_ ),
    .A(net109));
 sg13g2_tielo \proj_14.flop9/dffsr_206  (.L_LO(net220));
 sg13g2_tielo \proj__4.flop1/dffsr_207  (.L_LO(net221));
 sg13g2_sdfbbp_1 \proj_14.flop9/dffsr  (.Q(\proj_14.net56 ),
    .Q_N(\proj_14.net57 ),
    .RESET_B(\proj_14.flop9/_0_ ),
    .SET_B(\proj_14.flop9/_1_ ),
    .D(\proj_14.net55 ),
    .SCE(net220),
    .SCD(net219),
    .CLK(net108));
 sg13g2_mux2_1 \proj_14.mux1/_0_  (.A0(\proj_14.net23 ),
    .A1(\proj_14.net44 ),
    .S(net56),
    .X(\proj_14.net23 ));
 sg13g2_mux2_1 \proj_14.mux10/_0_  (.A0(\proj_14.net105 ),
    .A1(\proj_14.net106 ),
    .S(net239),
    .X(\proj_14.net102 ));
 sg13g2_mux2_1 \proj_14.mux11/_0_  (.A0(\proj_14.net110 ),
    .A1(\proj_14.net111 ),
    .S(\proj_14.net105 ),
    .X(\proj_14.net108 ));
 sg13g2_mux2_1 \proj_14.mux12/_0_  (.A0(\proj_14.net114 ),
    .A1(\proj_14.net115 ),
    .S(\proj_14.net116 ),
    .X(\proj_14.net112 ));
 sg13g2_mux2_1 \proj_14.mux13/_0_  (.A0(\proj_14.net119 ),
    .A1(\proj_14.net120 ),
    .S(\proj_14.net121 ),
    .X(\proj_14.net117 ));
 sg13g2_mux2_1 \proj_14.mux14/_0_  (.A0(\proj_14.net124 ),
    .A1(\proj_14.net125 ),
    .S(\proj_14.net126 ),
    .X(\proj_14.net122 ));
 sg13g2_mux2_1 \proj_14.mux15/_0_  (.A0(\proj_14.net129 ),
    .A1(\proj_14.net130 ),
    .S(\proj_14.net131 ),
    .X(\proj_14.net127 ));
 sg13g2_mux2_1 \proj_14.mux16/_0_  (.A0(\proj_14.net135 ),
    .A1(\proj_14.net136 ),
    .S(\proj_14.net137 ),
    .X(\proj_14.net133 ));
 sg13g2_mux2_1 \proj_14.mux17/_0_  (.A0(\proj_14.net140 ),
    .A1(\proj_14.net141 ),
    .S(\proj_14.net142 ),
    .X(\proj_14.net138 ));
 sg13g2_mux2_1 \proj_14.mux18/_0_  (.A0(\proj_14.net145 ),
    .A1(\proj_14.net146 ),
    .S(\proj_14.net147 ),
    .X(\proj_14.net143 ));
 sg13g2_mux2_1 \proj_14.mux19/_0_  (.A0(\proj_14.net150 ),
    .A1(\proj_14.net151 ),
    .S(\proj_14.net152 ),
    .X(\proj_14.net148 ));
 sg13g2_mux2_1 \proj_14.mux2/_0_  (.A0(\proj_14.net28 ),
    .A1(\proj_14.net46 ),
    .S(net56),
    .X(\proj_14.net28 ));
 sg13g2_mux2_1 \proj_14.mux20/_0_  (.A0(\proj_14.net155 ),
    .A1(\proj_14.net156 ),
    .S(\proj_14.net157 ),
    .X(\proj_14.net153 ));
 sg13g2_mux2_1 \proj_14.mux21/_0_  (.A0(\proj_14.net160 ),
    .A1(\proj_14.net161 ),
    .S(\proj_14.net162 ),
    .X(\proj_14.net158 ));
 sg13g2_mux2_1 \proj_14.mux22/_0_  (.A0(\proj_14.net165 ),
    .A1(\proj_14.net166 ),
    .S(\proj_14.net167 ),
    .X(\proj_14.net163 ));
 sg13g2_mux2_1 \proj_14.mux23/_0_  (.A0(\proj_14.net170 ),
    .A1(\proj_14.net171 ),
    .S(\proj_14.net172 ),
    .X(\proj_14.net168 ));
 sg13g2_mux2_1 \proj_14.mux24/_0_  (.A0(\proj_14.net175 ),
    .A1(\proj_14.net176 ),
    .S(\proj_14.net177 ),
    .X(\proj_14.net173 ));
 sg13g2_mux2_1 \proj_14.mux25/_0_  (.A0(\proj_14.net209 ),
    .A1(\proj_14.net211 ),
    .S(net56),
    .X(\proj_14.net207 ));
 sg13g2_mux2_1 \proj_14.mux26/_0_  (.A0(\proj_14.net214 ),
    .A1(\proj_14.net233 ),
    .S(net55),
    .X(\proj_14.net212 ));
 sg13g2_mux2_1 \proj_14.mux27/_0_  (.A0(\proj_14.net217 ),
    .A1(\proj_14.net214 ),
    .S(net54),
    .X(\proj_14.net216 ));
 sg13g2_mux2_1 \proj_14.mux28/_0_  (.A0(\proj_14.net219 ),
    .A1(\proj_14.net217 ),
    .S(net54),
    .X(\proj_14.net218 ));
 sg13g2_mux2_1 \proj_14.mux29/_0_  (.A0(\proj_14.net221 ),
    .A1(\proj_14.net219 ),
    .S(net54),
    .X(\proj_14.net220 ));
 sg13g2_mux2_1 \proj_14.mux3/_0_  (.A0(\proj_14.net31 ),
    .A1(\proj_14.net47 ),
    .S(net56),
    .X(\proj_14.net31 ));
 sg13g2_mux2_1 \proj_14.mux30/_0_  (.A0(\proj_14.net223 ),
    .A1(\proj_14.net221 ),
    .S(net54),
    .X(\proj_14.net222 ));
 sg13g2_mux2_1 \proj_14.mux31/_0_  (.A0(\proj_14.net226 ),
    .A1(\proj_14.net223 ),
    .S(net54),
    .X(\proj_14.net224 ));
 sg13g2_mux2_1 \proj_14.mux32/_0_  (.A0(\proj_14.net228 ),
    .A1(\proj_14.net226 ),
    .S(net54),
    .X(\proj_14.net227 ));
 sg13g2_mux2_1 \proj_14.mux33/_0_  (.A0(\proj_14.net231 ),
    .A1(\proj_14.net228 ),
    .S(net54),
    .X(\proj_14.net229 ));
 sg13g2_mux2_1 \proj_14.mux4/_0_  (.A0(\proj_14.net34 ),
    .A1(\proj_14.net26 ),
    .S(net56),
    .X(\proj_14.net34 ));
 sg13g2_mux2_1 \proj_14.mux5/_0_  (.A0(\proj_14.net38 ),
    .A1(\proj_14.net29 ),
    .S(net54),
    .X(\proj_14.net38 ));
 sg13g2_mux2_1 \proj_14.mux6/_0_  (.A0(\proj_14.net41 ),
    .A1(\proj_14.net32 ),
    .S(net55),
    .X(\proj_14.net41 ));
 sg13g2_mux2_1 \proj_14.mux7/_0_  (.A0(\proj_14.net48 ),
    .A1(\proj_14.net36 ),
    .S(net56),
    .X(\proj_14.net48 ));
 sg13g2_mux2_1 \proj_14.mux8/_0_  (.A0(\proj_14.net52 ),
    .A1(\proj_14.net39 ),
    .S(net55),
    .X(\proj_14.net52 ));
 sg13g2_mux2_1 \proj_14.mux9/_0_  (.A0(\proj_14.net55 ),
    .A1(\proj_14.net42 ),
    .S(net55),
    .X(\proj_14.net55 ));
 sg13g2_inv_1 \proj_14.not1/_0_  (.Y(\proj_14.net132 ),
    .A(net110));
 sg13g2_inv_1 \proj_14.not10/_0_  (.Y(\proj_14.net193 ),
    .A(\proj_14.net190 ));
 sg13g2_inv_1 \proj_14.not2/_0_  (.Y(\proj_14.net202 ),
    .A(\proj_14.net184 ));
 sg13g2_inv_1 \proj_14.not3/_0_  (.Y(\proj_14.net201 ),
    .A(\proj_14.net185 ));
 sg13g2_inv_1 \proj_14.not4/_0_  (.Y(\proj_14.net198 ),
    .A(\proj_14.net187 ));
 sg13g2_inv_1 \proj_14.not5/_0_  (.Y(\proj_14.net25 ),
    .A(net111));
 sg13g2_inv_1 \proj_14.not6/_0_  (.Y(\proj_14.net199 ),
    .A(\proj_14.net186 ));
 sg13g2_inv_1 \proj_14.not7/_0_  (.Y(\proj_14.net195 ),
    .A(\proj_14.net189 ));
 sg13g2_inv_1 \proj_14.not8/_0_  (.Y(\proj_14.net196 ),
    .A(\proj_14.net188 ));
 sg13g2_inv_1 \proj_14.not9/_0_  (.Y(\proj_14.net192 ),
    .A(\proj_14.net191 ));
 sg13g2_or2_1 \proj_14.or1/_0_  (.X(\proj_14.net104 ),
    .B(\proj_14.net132 ),
    .A(\proj_14.net183 ));
 sg13g2_or2_1 \proj_14.or10/_0_  (.X(\proj_14.net96 ),
    .B(\proj_14.net60 ),
    .A(\proj_14.net89 ));
 sg13g2_or2_1 \proj_14.or11/_0_  (.X(\proj_14.net97 ),
    .B(\proj_14.net62 ),
    .A(\proj_14.net90 ));
 sg13g2_or2_1 \proj_14.or12/_0_  (.X(\proj_14.net98 ),
    .B(\proj_14.net63 ),
    .A(\proj_14.net91 ));
 sg13g2_or2_1 \proj_14.or13/_0_  (.X(\proj_14.net99 ),
    .B(\proj_14.net65 ),
    .A(\proj_14.net92 ));
 sg13g2_or2_1 \proj_14.or14/_0_  (.X(\proj_14.net100 ),
    .B(\proj_14.net66 ),
    .A(\proj_14.net93 ));
 sg13g2_or2_1 \proj_14.or15/_0_  (.X(\proj_14.net101 ),
    .B(\proj_14.net67 ),
    .A(\proj_14.net94 ));
 sg13g2_or2_1 \proj_14.or16/_0_  (.X(\proj_14.net247 ),
    .B(\proj_14.net236 ),
    .A(\proj_14.net234 ));
 sg13g2_or2_1 \proj_14.or17/_0_  (.X(\proj_14.net250 ),
    .B(\proj_14.net248 ),
    .A(\proj_14.net249 ));
 sg13g2_or2_1 \proj_14.or18/_0_  (.X(\proj_14.net255 ),
    .B(\proj_14.net254 ),
    .A(\proj_14.net252 ));
 sg13g2_or2_1 \proj_14.or19/_0_  (.X(\proj_14.net251 ),
    .B(\proj_14.net237 ),
    .A(\proj_14.net248 ));
 sg13g2_or2_1 \proj_14.or2/_0_  (.X(\proj_14.net95 ),
    .B(\proj_14.net59 ),
    .A(\proj_14.net88 ));
 sg13g2_or2_1 \proj_14.or20/_0_  (.X(\proj_14.net253 ),
    .B(\proj_14.net252 ),
    .A(\proj_14.net236 ));
 sg13g2_or2_1 \proj_14.or21/_0_  (.X(\proj_14.net257 ),
    .B(\proj_14.net254 ),
    .A(\proj_14.net256 ));
 sg13g2_or2_1 \proj_14.or22/_0_  (.X(\proj_14.net272 ),
    .B(\proj_14.net253 ),
    .A(\proj_14.net250 ));
 sg13g2_or2_1 \proj_14.or23/_0_  (.X(\proj_14.net287 ),
    .B(\proj_14.net285 ),
    .A(\proj_14.net286 ));
 sg13g2_or2_1 \proj_14.or24/_0_  (.X(\proj_14.net260 ),
    .B(\proj_14.net259 ),
    .A(\proj_14.net240 ));
 sg13g2_or2_1 \proj_14.or25/_0_  (.X(\proj_14.net262 ),
    .B(\proj_14.net261 ),
    .A(\proj_14.net240 ));
 sg13g2_or2_1 \proj_14.or26/_0_  (.X(\proj_14.net263 ),
    .B(\proj_14.net243 ),
    .A(\proj_14.net261 ));
 sg13g2_or2_1 \proj_14.or27/_0_  (.X(\proj_14.net264 ),
    .B(\proj_14.net251 ),
    .A(\proj_14.net245 ));
 sg13g2_or2_1 \proj_14.or28/_0_  (.X(\proj_14.net266 ),
    .B(\proj_14.net244 ),
    .A(\proj_14.net265 ));
 sg13g2_or2_1 \proj_14.or29/_0_  (.X(\proj_14.net268 ),
    .B(\proj_14.net244 ),
    .A(\proj_14.net267 ));
 sg13g2_or2_1 \proj_14.or3/_0_  (.X(\proj_14.net88 ),
    .B(\proj_14.net69 ),
    .A(\proj_14.net79 ));
 sg13g2_or2_1 \proj_14.or30/_0_  (.X(\proj_14.net273 ),
    .B(\proj_14.net266 ),
    .A(\proj_14.net260 ));
 sg13g2_or2_1 \proj_14.or31/_0_  (.X(\proj_14.net270 ),
    .B(\proj_14.net269 ),
    .A(\proj_14.net268 ));
 sg13g2_or2_1 \proj_14.or32/_0_  (.X(\proj_14.net271 ),
    .B(\proj_14.net256 ),
    .A(\proj_14.net258 ));
 sg13g2_or2_1 \proj_14.or33/_0_  (.X(\proj_14.net274 ),
    .B(\proj_14.net257 ),
    .A(\proj_14.net247 ));
 sg13g2_or2_1 \proj_14.or34/_0_  (.X(\proj_14.net275 ),
    .B(\proj_14.net273 ),
    .A(\proj_14.net274 ));
 sg13g2_or2_1 \proj_14.or35/_0_  (.X(\proj_14.net276 ),
    .B(\proj_14.net263 ),
    .A(\proj_14.net272 ));
 sg13g2_or2_1 \proj_14.or36/_0_  (.X(\proj_14.net277 ),
    .B(\proj_14.net270 ),
    .A(\proj_14.net276 ));
 sg13g2_or2_1 \proj_14.or37/_0_  (.X(\proj_14.net278 ),
    .B(\proj_14.net271 ),
    .A(\proj_14.net262 ));
 sg13g2_or2_1 \proj_14.or38/_0_  (.X(\proj_14.net279 ),
    .B(\proj_14.net255 ),
    .A(\proj_14.net264 ));
 sg13g2_or2_1 \proj_14.or39/_0_  (.X(\proj_14.net280 ),
    .B(\proj_14.net278 ),
    .A(\proj_14.net279 ));
 sg13g2_or2_1 \proj_14.or4/_0_  (.X(\proj_14.net89 ),
    .B(\proj_14.net70 ),
    .A(\proj_14.net80 ));
 sg13g2_or2_1 \proj_14.or40/_0_  (.X(\proj_14.net283 ),
    .B(\proj_14.net240 ),
    .A(\proj_14.net241 ));
 sg13g2_or2_1 \proj_14.or41/_0_  (.X(\proj_14.net284 ),
    .B(\proj_14.net243 ),
    .A(\proj_14.net244 ));
 sg13g2_or2_1 \proj_14.or42/_0_  (.X(\proj_14.net285 ),
    .B(\proj_14.net283 ),
    .A(\proj_14.net284 ));
 sg13g2_or2_1 \proj_14.or43/_0_  (.X(\proj_14.net286 ),
    .B(\proj_14.net259 ),
    .A(\proj_14.net258 ));
 sg13g2_or2_1 \proj_14.or44/_0_  (.X(\proj_14.net288 ),
    .B(\proj_14.net265 ),
    .A(\proj_14.net252 ));
 sg13g2_or2_1 \proj_14.or45/_0_  (.X(\proj_14.net281 ),
    .B(\proj_14.net287 ),
    .A(\proj_14.net289 ));
 sg13g2_or2_1 \proj_14.or46/_0_  (.X(\proj_14.net289 ),
    .B(\proj_14.net245 ),
    .A(\proj_14.net288 ));
 sg13g2_or2_1 \proj_14.or5/_0_  (.X(\proj_14.net90 ),
    .B(\proj_14.net72 ),
    .A(\proj_14.net82 ));
 sg13g2_or2_1 \proj_14.or6/_0_  (.X(\proj_14.net91 ),
    .B(\proj_14.net73 ),
    .A(\proj_14.net83 ));
 sg13g2_or2_1 \proj_14.or7/_0_  (.X(\proj_14.net92 ),
    .B(\proj_14.net75 ),
    .A(\proj_14.net85 ));
 sg13g2_or2_1 \proj_14.or8/_0_  (.X(\proj_14.net93 ),
    .B(\proj_14.net76 ),
    .A(\proj_14.net86 ));
 sg13g2_or2_1 \proj_14.or9/_0_  (.X(\proj_14.net94 ),
    .B(\proj_14.net77 ),
    .A(\proj_14.net87 ));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(net5),
    .A(\proj_14.net175 ),
    .X(\proj_14.net184 ));
 sg13g2_xor2_1 \proj_14.xor10/_0_  (.B(\proj_14.net226 ),
    .A(\proj_14.net231 ),
    .X(\proj_14.net282 ));
 sg13g2_xor2_1 \proj_14.xor11/_0_  (.B(\proj_14.net221 ),
    .A(\proj_14.net232 ),
    .X(\proj_14.net233 ));
 sg13g2_xor2_1 \proj_14.xor2/_0_  (.B(net4),
    .A(\proj_14.net170 ),
    .X(\proj_14.net185 ));
 sg13g2_xor2_1 \proj_14.xor3/_0_  (.B(net3),
    .A(\proj_14.net165 ),
    .X(\proj_14.net186 ));
 sg13g2_xor2_1 \proj_14.xor4/_0_  (.B(net2),
    .A(\proj_14.net160 ),
    .X(\proj_14.net187 ));
 sg13g2_xor2_1 \proj_14.xor5/_0_  (.B(net46),
    .A(\proj_14.net155 ),
    .X(\proj_14.net188 ));
 sg13g2_xor2_1 \proj_14.xor6/_0_  (.B(net48),
    .A(\proj_14.net150 ),
    .X(\proj_14.net189 ));
 sg13g2_xor2_1 \proj_14.xor7/_0_  (.B(net50),
    .A(\proj_14.net145 ),
    .X(\proj_14.net190 ));
 sg13g2_xor2_1 \proj_14.xor8/_0_  (.B(net53),
    .A(\proj_14.net140 ),
    .X(\proj_14.net191 ));
 sg13g2_xor2_1 \proj_14.xor9/_0_  (.B(\proj_14.net223 ),
    .A(\proj_14.net282 ),
    .X(\proj_14.net232 ));
 sg13g2_and2_1 \proj_15.and1/_0_  (.A(net48),
    .B(net53),
    .X(\proj_15.net15 ));
 sg13g2_and2_1 \proj_15.and2/_0_  (.A(\proj_15.net15 ),
    .B(net1),
    .X(\proj_15.net18 ));
 sg13g2_and2_1 \proj_15.and3/_0_  (.A(net46),
    .B(\proj_15.net7 ),
    .X(\proj_15.net17 ));
 sg13g2_or2_1 \proj_15.or1/_0_  (.X(\proj_15.net9 ),
    .B(\proj_15.net17 ),
    .A(\proj_15.net18 ));
 sg13g2_xor2_1 \proj_15.xor1/_0_  (.B(net51),
    .A(net48),
    .X(\proj_15.net7 ));
 sg13g2_xor2_1 \proj_15.xor2/_0_  (.B(\proj_15.net15 ),
    .A(net1),
    .X(\proj_15.net16 ));
 sg13g2_xor2_1 \proj_15.xor3/_0_  (.B(\proj_15.net16 ),
    .A(net46),
    .X(\proj_15.net8 ));
 sg13g2_inv_1 \proj__0.not3/_0_  (.Y(\proj__0.net10 ),
    .A(net47));
 sg13g2_inv_1 \proj__0.not4/_0_  (.Y(\proj__0.net11 ),
    .A(net45));
 sg13g2_xor2_1 \proj__0.xor1/_0_  (.B(net51),
    .A(net49),
    .X(\proj__0.net9 ));
 sg13g2_and2_1 \proj__1.and1/_0_  (.A(\proj__1.net18 ),
    .B(net51),
    .X(\proj__1.net19 ));
 sg13g2_and2_1 \proj__1.and2/_0_  (.A(\proj__1.net16 ),
    .B(net48),
    .X(\proj__1.net20 ));
 sg13g2_and2_1 \proj__1.and3/_0_  (.A(\proj__1.net10 ),
    .B(net2),
    .X(\proj__1.net21 ));
 sg13g2_and2_1 \proj__1.and4/_0_  (.A(\proj__1.net17 ),
    .B(net4),
    .X(\proj__1.net22 ));
 sg13g2_and2_1 \proj__1.and5/_0_  (.A(\proj__1.net20 ),
    .B(\proj__1.net19 ),
    .X(\proj__1.net23 ));
 sg13g2_and2_1 \proj__1.and6/_0_  (.A(\proj__1.net22 ),
    .B(\proj__1.net21 ),
    .X(\proj__1.net24 ));
 sg13g2_and2_1 \proj__1.and7/_0_  (.A(\proj__1.net24 ),
    .B(\proj__1.net23 ),
    .X(\proj__1.net9 ));
 sg13g2_inv_1 \proj__1.not1/_0_  (.Y(\proj__1.net16 ),
    .A(net45));
 sg13g2_inv_1 \proj__1.not2/_0_  (.Y(\proj__1.net17 ),
    .A(net5));
 sg13g2_inv_1 \proj__1.not3/_0_  (.Y(\proj__1.net18 ),
    .A(net49));
 sg13g2_inv_1 \proj__1.not4/_0_  (.Y(\proj__1.net10 ),
    .A(net44));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net9 ),
    .A(net52));
 sg13g2_inv_1 \proj__2.not2/_0_  (.Y(\proj__2.net10 ),
    .A(net50));
 sg13g2_inv_1 \proj__2.not3/_0_  (.Y(\proj__2.net11 ),
    .A(net47));
 sg13g2_inv_1 \proj__2.not4/_0_  (.Y(\proj__2.net12 ),
    .A(net45));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net11 ),
    .B(net51),
    .X(\proj__3.net4 ));
 sg13g2_and2_1 \proj__3.and4/_0_  (.A(net49),
    .B(\proj__3.net12 ),
    .X(\proj__3.net3 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net11 ),
    .A(net49));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net12 ),
    .A(net51));
 sg13g2_inv_1 \proj__3.not6/_0_  (.Y(\proj__3.net5 ),
    .A(\proj__3.net13 ));
 sg13g2_or2_1 \proj__3.or4/_0_  (.X(\proj__3.net13 ),
    .B(\proj__3.net4 ),
    .A(\proj__3.net3 ));
 sg13g2_inv_1 \proj__4.flop1/_4_  (.Y(\proj__4.flop1/_1_ ),
    .A(\proj__4.flop1/s ));
 sg13g2_inv_1 \proj__4.flop1/_5_  (.Y(\proj__4.flop1/_0_ ),
    .A(net113));
 sg13g2_tielo \proj__4.flop1/dffsr_208  (.L_LO(net222));
 sg13g2_tielo \proj__4.flop2/dffsr_209  (.L_LO(net223));
 sg13g2_sdfbbp_1 \proj__4.flop1/dffsr  (.Q(\proj__4.flop1/q ),
    .Q_N(\proj__4.net11 ),
    .RESET_B(\proj__4.flop1/_0_ ),
    .SET_B(\proj__4.flop1/_1_ ),
    .D(net53),
    .SCE(net222),
    .SCD(net221),
    .CLK(net112));
 sg13g2_inv_1 \proj__4.flop2/_4_  (.Y(\proj__4.flop2/_1_ ),
    .A(\proj__4.flop2/s ));
 sg13g2_inv_1 \proj__4.flop2/_5_  (.Y(\proj__4.flop2/_0_ ),
    .A(net115));
 sg13g2_tielo \proj__4.flop2/dffsr_210  (.L_LO(net224));
 sg13g2_tielo \proj__4.flop3/dffsr_211  (.L_LO(net225));
 sg13g2_sdfbbp_1 \proj__4.flop2/dffsr  (.Q(\proj__4.flop2/q ),
    .Q_N(\proj__4.net12 ),
    .RESET_B(\proj__4.flop2/_0_ ),
    .SET_B(\proj__4.flop2/_1_ ),
    .D(net50),
    .SCE(net224),
    .SCD(net223),
    .CLK(net114));
 sg13g2_inv_1 \proj__4.flop3/_4_  (.Y(\proj__4.flop3/_1_ ),
    .A(\proj__4.flop3/s ));
 sg13g2_inv_1 \proj__4.flop3/_5_  (.Y(\proj__4.flop3/_0_ ),
    .A(net117));
 sg13g2_tielo \proj__4.flop3/dffsr_212  (.L_LO(net226));
 sg13g2_tielo \proj__4.flop4/dffsr_213  (.L_LO(net227));
 sg13g2_sdfbbp_1 \proj__4.flop3/dffsr  (.Q(\proj__4.flop3/q ),
    .Q_N(\proj__4.net13 ),
    .RESET_B(\proj__4.flop3/_0_ ),
    .SET_B(\proj__4.flop3/_1_ ),
    .D(net47),
    .SCE(net226),
    .SCD(net225),
    .CLK(net116));
 sg13g2_inv_1 \proj__4.flop4/_4_  (.Y(\proj__4.flop4/_1_ ),
    .A(\proj__4.flop4/s ));
 sg13g2_inv_1 \proj__4.flop4/_5_  (.Y(\proj__4.flop4/_0_ ),
    .A(net119));
 sg13g2_tielo \proj__4.flop4/dffsr_214  (.L_LO(net228));
 sg13g2_tielo \proj__4.flop5/dffsr_215  (.L_LO(net229));
 sg13g2_sdfbbp_1 \proj__4.flop4/dffsr  (.Q(\proj__4.flop4/q ),
    .Q_N(\proj__4.net14 ),
    .RESET_B(\proj__4.flop4/_0_ ),
    .SET_B(\proj__4.flop4/_1_ ),
    .D(net46),
    .SCE(net228),
    .SCD(net227),
    .CLK(net118));
 sg13g2_inv_1 \proj__4.flop5/_4_  (.Y(\proj__4.flop5/_1_ ),
    .A(\proj__4.flop5/s ));
 sg13g2_inv_1 \proj__4.flop5/_5_  (.Y(\proj__4.flop5/_0_ ),
    .A(net121));
 sg13g2_tielo \proj__4.flop5/dffsr_216  (.L_LO(net230));
 sg13g2_tielo \proj__4.flop6/dffsr_217  (.L_LO(net231));
 sg13g2_sdfbbp_1 \proj__4.flop5/dffsr  (.Q(\proj__4.net15 ),
    .Q_N(\proj__4.flop5/notq ),
    .RESET_B(\proj__4.flop5/_0_ ),
    .SET_B(\proj__4.flop5/_1_ ),
    .D(net2),
    .SCE(net230),
    .SCD(net229),
    .CLK(net120));
 sg13g2_inv_1 \proj__4.flop6/_4_  (.Y(\proj__4.flop6/_1_ ),
    .A(\proj__4.flop6/s ));
 sg13g2_inv_1 \proj__4.flop6/_5_  (.Y(\proj__4.flop6/_0_ ),
    .A(net123));
 sg13g2_tielo \proj__4.flop6/dffsr_218  (.L_LO(net232));
 sg13g2_tielo \proj__4.flop8/dffsr_219  (.L_LO(net233));
 sg13g2_sdfbbp_1 \proj__4.flop6/dffsr  (.Q(\proj__4.net16 ),
    .Q_N(\proj__4.flop6/notq ),
    .RESET_B(\proj__4.flop6/_0_ ),
    .SET_B(\proj__4.flop6/_1_ ),
    .D(net44),
    .SCE(net232),
    .SCD(net231),
    .CLK(net122));
 sg13g2_inv_1 \proj__4.flop8/_4_  (.Y(\proj__4.flop8/_1_ ),
    .A(\proj__4.flop8/s ));
 sg13g2_inv_1 \proj__4.flop8/_5_  (.Y(\proj__4.flop8/_0_ ),
    .A(net125));
 sg13g2_tielo \proj__4.flop8/dffsr_220  (.L_LO(net234));
 sg13g2_tielo \proj__4.flop9/dffsr_221  (.L_LO(net235));
 sg13g2_sdfbbp_1 \proj__4.flop8/dffsr  (.Q(\proj__4.net17 ),
    .Q_N(\proj__4.flop8/notq ),
    .RESET_B(\proj__4.flop8/_0_ ),
    .SET_B(\proj__4.flop8/_1_ ),
    .D(net4),
    .SCE(net234),
    .SCD(net233),
    .CLK(net124));
 sg13g2_inv_1 \proj__4.flop9/_4_  (.Y(\proj__4.flop9/_1_ ),
    .A(\proj__4.flop9/s ));
 sg13g2_inv_1 \proj__4.flop9/_5_  (.Y(\proj__4.flop9/_0_ ),
    .A(net127));
 sg13g2_tielo \proj__4.flop9/dffsr_222  (.L_LO(net236));
 sg13g2_tielo \proj__9.flop1/dffsr_223  (.L_LO(net237));
 sg13g2_sdfbbp_1 \proj__4.flop9/dffsr  (.Q(\proj__4.net18 ),
    .Q_N(\proj__4.flop9/notq ),
    .RESET_B(\proj__4.flop9/_0_ ),
    .SET_B(\proj__4.flop9/_1_ ),
    .D(net5),
    .SCE(net236),
    .SCD(net235),
    .CLK(net126));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net49),
    .B(net51),
    .X(\proj__5.net9 ));
 sg13g2_and2_1 \proj__5.and2/_0_  (.A(net45),
    .B(net47),
    .X(\proj__5.net12 ));
 sg13g2_inv_1 \proj__5.not1/_0_  (.Y(\proj__5.net10 ),
    .A(net4));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net11 ),
    .B(net2),
    .A(net44));
 sg13g2_inv_1 \proj__6.not3/_0_  (.Y(\proj__6.net9 ),
    .A(net47));
 sg13g2_inv_1 \proj__6.not4/_0_  (.Y(\proj__6.net10 ),
    .A(net45));
 sg13g2_dfrbp_1 \proj__7.flop1/_1_  (.CLK(net128),
    .RESET_B(net255),
    .D(net5),
    .Q_N(\proj__7.net6 ),
    .Q(\proj__7.net5 ));
 sg13g2_tiehi \proj__7.flop2/_1__242  (.L_HI(net256));
 sg13g2_dfrbp_1 \proj__7.flop2/_1_  (.CLK(net129),
    .RESET_B(net256),
    .D(\proj__7.net14 ),
    .Q_N(\proj__7.net14 ),
    .Q(\proj__7.net8 ));
 sg13g2_tiehi \proj__7.flop3/_1__243  (.L_HI(net257));
 sg13g2_dfrbp_1 \proj__7.flop3/_1_  (.CLK(\proj__7.net14 ),
    .RESET_B(net257),
    .D(\proj__7.net15 ),
    .Q_N(\proj__7.net15 ),
    .Q(\proj__7.net7 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(net50),
    .B(net52),
    .X(\proj__8.net7 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(\proj__9.net11 ),
    .B(net53),
    .X(\proj__9.net12 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(net50),
    .B(\proj__9.net13 ),
    .X(\proj__9.net14 ));
 sg13g2_inv_1 \proj__9.flop1/_4_  (.Y(\proj__9.flop1/_1_ ),
    .A(net131));
 sg13g2_inv_1 \proj__9.flop1/_5_  (.Y(\proj__9.flop1/_0_ ),
    .A(\proj__9.net17 ));
 sg13g2_tielo \proj__9.flop1/dffsr_224  (.L_LO(net238));
 sg13g2_tiehi \proj_14.mux10/_0__225  (.L_HI(net239));
 sg13g2_sdfbbp_1 \proj__9.flop1/dffsr  (.Q(\proj__9.net5 ),
    .Q_N(\proj__9.flop1/notq ),
    .RESET_B(\proj__9.flop1/_0_ ),
    .SET_B(\proj__9.flop1/_1_ ),
    .D(\proj__9.net15 ),
    .SCE(net238),
    .SCD(net237),
    .CLK(net130));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net11 ),
    .A(net50));
 sg13g2_inv_1 \proj__9.not2/_0_  (.Y(\proj__9.net13 ),
    .A(net53));
 sg13g2_inv_1 \proj__9.not3/_0_  (.Y(\proj__9.net17 ),
    .A(net132));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net15 ),
    .B(\proj__9.net12 ),
    .A(\proj__9.net14 ));
 sg13g2_buf_2 fanout43 (.A(_063_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(net3),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(ui_in[3]),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(ui_in[3]),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(ui_in[2]),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(net50),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(net1),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(net53),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net53),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(ui_in[0]),
    .X(net53));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(net55));
 sg13g2_buf_2 fanout55 (.A(net56),
    .X(net55));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(\proj_14.net45 ));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[4]));
 sg13g2_buf_2 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[6]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[7]));
 sg13g2_buf_2 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_tielo \proj_13.flop1/_1__10  (.L_LO(net10));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_2 FILLER_17_271 ();
 sg13g2_decap_4 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_fill_2 FILLER_17_291 ();
 sg13g2_fill_1 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_4 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_4 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_45 ();
 sg13g2_decap_4 FILLER_18_50 ();
 sg13g2_fill_2 FILLER_18_54 ();
 sg13g2_decap_4 FILLER_18_59 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_94 ();
 sg13g2_decap_8 FILLER_18_108 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_122 ();
 sg13g2_decap_8 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_decap_8 FILLER_18_185 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_213 ();
 sg13g2_decap_8 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_227 ();
 sg13g2_decap_8 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_decap_4 FILLER_18_255 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_fill_2 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_32 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_177 ();
 sg13g2_decap_4 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_230 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_4 FILLER_19_279 ();
 sg13g2_fill_2 FILLER_19_283 ();
 sg13g2_fill_1 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_327 ();
 sg13g2_decap_4 FILLER_19_333 ();
 sg13g2_fill_2 FILLER_19_337 ();
 sg13g2_fill_2 FILLER_19_345 ();
 sg13g2_decap_4 FILLER_19_374 ();
 sg13g2_fill_1 FILLER_19_378 ();
 sg13g2_decap_4 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_2 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_16 ();
 sg13g2_decap_4 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_25 ();
 sg13g2_decap_4 FILLER_20_31 ();
 sg13g2_fill_1 FILLER_20_35 ();
 sg13g2_decap_4 FILLER_20_39 ();
 sg13g2_fill_1 FILLER_20_43 ();
 sg13g2_decap_8 FILLER_20_54 ();
 sg13g2_decap_8 FILLER_20_61 ();
 sg13g2_decap_4 FILLER_20_68 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_2 FILLER_20_83 ();
 sg13g2_fill_1 FILLER_20_101 ();
 sg13g2_decap_4 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_114 ();
 sg13g2_fill_2 FILLER_20_121 ();
 sg13g2_fill_1 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_159 ();
 sg13g2_decap_8 FILLER_20_195 ();
 sg13g2_decap_8 FILLER_20_202 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_237 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_decap_8 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_4 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_314 ();
 sg13g2_decap_4 FILLER_20_358 ();
 sg13g2_fill_2 FILLER_20_362 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_2 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_fill_2 FILLER_21_72 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_167 ();
 sg13g2_decap_4 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_fill_2 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_fill_2 FILLER_21_221 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_fill_2 FILLER_21_228 ();
 sg13g2_decap_4 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_244 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_4 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_285 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_4 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_decap_4 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_fill_2 FILLER_21_378 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_388 ();
 sg13g2_fill_1 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_11 ();
 sg13g2_fill_2 FILLER_22_16 ();
 sg13g2_fill_1 FILLER_22_18 ();
 sg13g2_fill_2 FILLER_22_23 ();
 sg13g2_fill_1 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_33 ();
 sg13g2_fill_2 FILLER_22_40 ();
 sg13g2_fill_1 FILLER_22_52 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_decap_4 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_decap_4 FILLER_22_208 ();
 sg13g2_fill_2 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_4 FILLER_22_362 ();
 sg13g2_fill_2 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_372 ();
 sg13g2_decap_4 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_4 FILLER_22_387 ();
 sg13g2_fill_1 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_48 ();
 sg13g2_fill_2 FILLER_23_60 ();
 sg13g2_decap_8 FILLER_23_100 ();
 sg13g2_decap_4 FILLER_23_107 ();
 sg13g2_decap_8 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_decap_4 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_185 ();
 sg13g2_decap_4 FILLER_23_192 ();
 sg13g2_decap_4 FILLER_23_234 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_decap_4 FILLER_23_242 ();
 sg13g2_decap_4 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_decap_4 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_4 FILLER_23_305 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_decap_4 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_323 ();
 sg13g2_decap_4 FILLER_23_331 ();
 sg13g2_fill_2 FILLER_23_338 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_15 ();
 sg13g2_fill_1 FILLER_24_17 ();
 sg13g2_decap_4 FILLER_24_22 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_fill_2 FILLER_24_34 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_53 ();
 sg13g2_decap_4 FILLER_24_76 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_decap_8 FILLER_24_85 ();
 sg13g2_decap_4 FILLER_24_95 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_103 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_132 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_144 ();
 sg13g2_decap_4 FILLER_24_153 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_decap_4 FILLER_24_209 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_decap_4 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_decap_4 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_decap_4 FILLER_24_304 ();
 sg13g2_decap_4 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_4 FILLER_24_371 ();
 sg13g2_fill_2 FILLER_24_375 ();
 sg13g2_fill_1 FILLER_24_381 ();
 sg13g2_decap_4 FILLER_24_385 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_1 FILLER_25_54 ();
 sg13g2_fill_2 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_decap_4 FILLER_25_170 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_decap_8 FILLER_25_180 ();
 sg13g2_decap_8 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_fill_2 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_201 ();
 sg13g2_decap_4 FILLER_25_206 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_decap_4 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_decap_4 FILLER_25_263 ();
 sg13g2_decap_4 FILLER_25_270 ();
 sg13g2_fill_2 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_fill_2 FILLER_25_337 ();
 sg13g2_fill_1 FILLER_25_339 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_fill_2 FILLER_25_357 ();
 sg13g2_decap_4 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_fill_2 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_61 ();
 sg13g2_decap_4 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_72 ();
 sg13g2_fill_2 FILLER_26_81 ();
 sg13g2_decap_4 FILLER_26_87 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_104 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_157 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_decap_4 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_177 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_decap_4 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_257 ();
 sg13g2_fill_2 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_269 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_320 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_decap_4 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_fill_2 FILLER_26_385 ();
 sg13g2_fill_1 FILLER_26_387 ();
 sg13g2_fill_1 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_29 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_48 ();
 sg13g2_decap_8 FILLER_27_52 ();
 sg13g2_fill_2 FILLER_27_59 ();
 sg13g2_fill_2 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_292 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_4 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_decap_4 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_fill_1 FILLER_27_383 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_73 ();
 sg13g2_fill_2 FILLER_28_82 ();
 sg13g2_decap_4 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_92 ();
 sg13g2_decap_4 FILLER_28_96 ();
 sg13g2_fill_2 FILLER_28_100 ();
 sg13g2_decap_8 FILLER_28_106 ();
 sg13g2_fill_1 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_4 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_decap_4 FILLER_28_223 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_277 ();
 sg13g2_decap_4 FILLER_28_283 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_297 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_337 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_decap_4 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_358 ();
 sg13g2_decap_4 FILLER_28_365 ();
 sg13g2_fill_2 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_37 ();
 sg13g2_fill_2 FILLER_29_47 ();
 sg13g2_decap_8 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_72 ();
 sg13g2_decap_8 FILLER_29_79 ();
 sg13g2_decap_4 FILLER_29_86 ();
 sg13g2_fill_1 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_decap_4 FILLER_29_101 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_decap_4 FILLER_29_109 ();
 sg13g2_fill_2 FILLER_29_113 ();
 sg13g2_decap_8 FILLER_29_118 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_182 ();
 sg13g2_fill_1 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_315 ();
 sg13g2_decap_4 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_decap_4 FILLER_29_353 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_decap_4 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_88 ();
 sg13g2_decap_4 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_147 ();
 sg13g2_decap_4 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_fill_2 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_202 ();
 sg13g2_decap_4 FILLER_30_209 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_decap_4 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_decap_4 FILLER_30_231 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_fill_1 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_decap_4 FILLER_30_286 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_decap_4 FILLER_30_340 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_decap_4 FILLER_30_379 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_fill_2 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_31 ();
 sg13g2_fill_2 FILLER_31_36 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_46 ();
 sg13g2_decap_4 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_decap_4 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_87 ();
 sg13g2_fill_1 FILLER_31_89 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_decap_8 FILLER_31_106 ();
 sg13g2_decap_8 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_decap_4 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_170 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_208 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_decap_8 FILLER_31_247 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_decap_4 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_4 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_decap_4 FILLER_31_338 ();
 sg13g2_fill_2 FILLER_31_342 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_17 ();
 sg13g2_decap_4 FILLER_32_24 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_decap_8 FILLER_32_136 ();
 sg13g2_decap_8 FILLER_32_143 ();
 sg13g2_decap_4 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_decap_4 FILLER_32_224 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_fill_2 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_fill_2 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_fill_2 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_fill_2 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_fill_2 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_13 ();
 sg13g2_decap_4 FILLER_33_19 ();
 sg13g2_fill_1 FILLER_33_23 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_48 ();
 sg13g2_decap_4 FILLER_33_59 ();
 sg13g2_fill_2 FILLER_33_68 ();
 sg13g2_decap_8 FILLER_33_75 ();
 sg13g2_fill_1 FILLER_33_82 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_121 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_decap_8 FILLER_33_138 ();
 sg13g2_decap_4 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_decap_4 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_decap_4 FILLER_33_203 ();
 sg13g2_decap_4 FILLER_33_250 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_decap_4 FILLER_33_277 ();
 sg13g2_decap_4 FILLER_33_286 ();
 sg13g2_fill_2 FILLER_33_290 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_decap_4 FILLER_33_344 ();
 sg13g2_fill_2 FILLER_33_368 ();
 sg13g2_decap_4 FILLER_33_383 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_fill_2 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_30 ();
 sg13g2_fill_1 FILLER_34_37 ();
 sg13g2_decap_8 FILLER_34_48 ();
 sg13g2_fill_2 FILLER_34_55 ();
 sg13g2_fill_1 FILLER_34_57 ();
 sg13g2_fill_1 FILLER_34_68 ();
 sg13g2_fill_2 FILLER_34_74 ();
 sg13g2_fill_1 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_192 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_213 ();
 sg13g2_decap_4 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_222 ();
 sg13g2_fill_2 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_decap_4 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_decap_4 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_fill_1 FILLER_34_356 ();
 sg13g2_fill_2 FILLER_34_371 ();
 sg13g2_fill_1 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_55 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_decap_8 FILLER_35_124 ();
 sg13g2_decap_8 FILLER_35_131 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_159 ();
 sg13g2_decap_8 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_decap_4 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_fill_2 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_320 ();
 sg13g2_decap_8 FILLER_35_356 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_decap_4 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_4 FILLER_35_387 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_fill_2 FILLER_35_396 ();
 sg13g2_fill_1 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_25 ();
 sg13g2_fill_2 FILLER_36_31 ();
 sg13g2_decap_8 FILLER_36_37 ();
 sg13g2_decap_8 FILLER_36_44 ();
 sg13g2_decap_8 FILLER_36_51 ();
 sg13g2_decap_4 FILLER_36_58 ();
 sg13g2_fill_2 FILLER_36_62 ();
 sg13g2_decap_8 FILLER_36_69 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_4 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_decap_4 FILLER_36_106 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_145 ();
 sg13g2_decap_8 FILLER_36_152 ();
 sg13g2_decap_8 FILLER_36_159 ();
 sg13g2_decap_8 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_173 ();
 sg13g2_decap_8 FILLER_36_180 ();
 sg13g2_decap_8 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_219 ();
 sg13g2_decap_8 FILLER_36_225 ();
 sg13g2_decap_8 FILLER_36_232 ();
 sg13g2_decap_4 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_243 ();
 sg13g2_fill_2 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_254 ();
 sg13g2_decap_8 FILLER_36_265 ();
 sg13g2_decap_8 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_279 ();
 sg13g2_decap_8 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_decap_4 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_decap_4 FILLER_36_381 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_decap_4 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_393 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_4 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_128 ();
 sg13g2_decap_8 FILLER_37_134 ();
 sg13g2_decap_8 FILLER_37_141 ();
 sg13g2_decap_8 FILLER_37_148 ();
 sg13g2_decap_8 FILLER_37_155 ();
 sg13g2_decap_8 FILLER_37_162 ();
 sg13g2_decap_8 FILLER_37_169 ();
 sg13g2_decap_8 FILLER_37_176 ();
 sg13g2_decap_8 FILLER_37_183 ();
 sg13g2_decap_8 FILLER_37_190 ();
 sg13g2_decap_8 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_204 ();
 sg13g2_decap_8 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_decap_8 FILLER_37_225 ();
 sg13g2_decap_4 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_236 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_decap_4 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net133;
 assign uio_oe[1] = net134;
 assign uio_oe[2] = net135;
 assign uio_oe[3] = net136;
 assign uio_oe[4] = net137;
 assign uio_oe[5] = net138;
 assign uio_oe[6] = net139;
 assign uio_oe[7] = net140;
 assign uio_out[0] = net141;
 assign uio_out[1] = net142;
 assign uio_out[2] = net143;
 assign uio_out[3] = net144;
 assign uio_out[4] = net145;
 assign uio_out[5] = net146;
 assign uio_out[6] = net147;
 assign uio_out[7] = net148;
endmodule

module tt_um_pwm_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \PWM_Generador.DIV_FREQ.clk_out ;
 wire \PWM_Generador.DIV_FREQ.counter[0] ;
 wire \PWM_Generador.DIV_FREQ.counter[1] ;
 wire \PWM_Generador.DIV_FREQ.counter[2] ;
 wire \PWM_Generador.DIV_FREQ.counter[3] ;
 wire \PWM_Generador.DIV_FREQ.counter[4] ;
 wire \PWM_Generador.DIV_FREQ.counter[5] ;
 wire \PWM_Generador.DUTY_CYCLE[0] ;
 wire \PWM_Generador.DUTY_CYCLE[1] ;
 wire \PWM_Generador.DUTY_CYCLE[2] ;
 wire \PWM_Generador.DUTY_CYCLE[3] ;
 wire \PWM_Generador.PWM_DFF1.Q ;
 wire \PWM_Generador.PWM_DFF2.Q ;
 wire \PWM_Generador.PWM_DFF3.Q ;
 wire \PWM_Generador.PWM_DFF4.Q ;
 wire \PWM_Generador.counter_PWM[0] ;
 wire \PWM_Generador.counter_PWM[1] ;
 wire \PWM_Generador.counter_PWM[2] ;
 wire \PWM_Generador.counter_PWM[3] ;
 wire \PWM_Generador.counter_debounce[0] ;
 wire \PWM_Generador.counter_debounce[10] ;
 wire \PWM_Generador.counter_debounce[11] ;
 wire \PWM_Generador.counter_debounce[12] ;
 wire \PWM_Generador.counter_debounce[13] ;
 wire \PWM_Generador.counter_debounce[14] ;
 wire \PWM_Generador.counter_debounce[15] ;
 wire \PWM_Generador.counter_debounce[16] ;
 wire \PWM_Generador.counter_debounce[17] ;
 wire \PWM_Generador.counter_debounce[18] ;
 wire \PWM_Generador.counter_debounce[19] ;
 wire \PWM_Generador.counter_debounce[1] ;
 wire \PWM_Generador.counter_debounce[20] ;
 wire \PWM_Generador.counter_debounce[21] ;
 wire \PWM_Generador.counter_debounce[22] ;
 wire \PWM_Generador.counter_debounce[23] ;
 wire \PWM_Generador.counter_debounce[24] ;
 wire \PWM_Generador.counter_debounce[25] ;
 wire \PWM_Generador.counter_debounce[26] ;
 wire \PWM_Generador.counter_debounce[27] ;
 wire \PWM_Generador.counter_debounce[2] ;
 wire \PWM_Generador.counter_debounce[3] ;
 wire \PWM_Generador.counter_debounce[4] ;
 wire \PWM_Generador.counter_debounce[5] ;
 wire \PWM_Generador.counter_debounce[6] ;
 wire \PWM_Generador.counter_debounce[7] ;
 wire \PWM_Generador.counter_debounce[8] ;
 wire \PWM_Generador.counter_debounce[9] ;
 wire \PWM_Generador.pwm_out0 ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire net57;
 wire net56;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net66;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire net67;
 wire net68;
 wire net69;
 wire clknet_0_clk;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;

 sg13g2_inv_1 _226_ (.Y(_095_),
    .A(\PWM_Generador.counter_debounce[0] ));
 sg13g2_inv_1 _227_ (.Y(_096_),
    .A(net81));
 sg13g2_inv_1 _228_ (.Y(_097_),
    .A(_042_));
 sg13g2_inv_1 _229_ (.Y(_098_),
    .A(\PWM_Generador.PWM_DFF4.Q ));
 sg13g2_inv_1 _230_ (.Y(_099_),
    .A(\PWM_Generador.PWM_DFF3.Q ));
 sg13g2_inv_1 _231_ (.Y(_100_),
    .A(\PWM_Generador.counter_PWM[3] ));
 sg13g2_inv_1 _232_ (.Y(_101_),
    .A(\PWM_Generador.counter_PWM[2] ));
 sg13g2_inv_1 _233_ (.Y(_043_),
    .A(net54));
 sg13g2_nor4_1 _234_ (.A(\PWM_Generador.counter_debounce[12] ),
    .B(\PWM_Generador.counter_debounce[11] ),
    .C(\PWM_Generador.counter_debounce[10] ),
    .D(\PWM_Generador.counter_debounce[9] ),
    .Y(_102_));
 sg13g2_nor4_1 _235_ (.A(\PWM_Generador.counter_debounce[16] ),
    .B(\PWM_Generador.counter_debounce[15] ),
    .C(\PWM_Generador.counter_debounce[14] ),
    .D(\PWM_Generador.counter_debounce[13] ),
    .Y(_103_));
 sg13g2_or4_2 _236_ (.A(\PWM_Generador.counter_debounce[8] ),
    .B(\PWM_Generador.counter_debounce[7] ),
    .C(\PWM_Generador.counter_debounce[6] ),
    .D(\PWM_Generador.counter_debounce[5] ),
    .X(_104_));
 sg13g2_nor4_1 _237_ (.A(\PWM_Generador.counter_debounce[4] ),
    .B(\PWM_Generador.counter_debounce[3] ),
    .C(\PWM_Generador.counter_debounce[2] ),
    .D(\PWM_Generador.counter_debounce[1] ),
    .Y(_105_));
 sg13g2_nand3_1 _238_ (.B(_103_),
    .C(_105_),
    .A(_102_),
    .Y(_106_));
 sg13g2_nor2_1 _239_ (.A(_104_),
    .B(_106_),
    .Y(_107_));
 sg13g2_nor4_2 _240_ (.A(\PWM_Generador.counter_debounce[20] ),
    .B(\PWM_Generador.counter_debounce[19] ),
    .C(\PWM_Generador.counter_debounce[18] ),
    .Y(_108_),
    .D(\PWM_Generador.counter_debounce[17] ));
 sg13g2_nor4_1 _241_ (.A(\PWM_Generador.counter_debounce[24] ),
    .B(\PWM_Generador.counter_debounce[23] ),
    .C(\PWM_Generador.counter_debounce[22] ),
    .D(\PWM_Generador.counter_debounce[21] ),
    .Y(_109_));
 sg13g2_and2_1 _242_ (.A(_108_),
    .B(_109_),
    .X(_110_));
 sg13g2_nor3_1 _243_ (.A(\PWM_Generador.counter_debounce[26] ),
    .B(\PWM_Generador.counter_debounce[25] ),
    .C(\PWM_Generador.counter_debounce[27] ),
    .Y(_111_));
 sg13g2_nand4_1 _244_ (.B(_108_),
    .C(_109_),
    .A(\PWM_Generador.counter_debounce[0] ),
    .Y(_112_),
    .D(_111_));
 sg13g2_nor3_2 _245_ (.A(_104_),
    .B(_106_),
    .C(_112_),
    .Y(_113_));
 sg13g2_o21ai_1 _246_ (.B1(\PWM_Generador.DUTY_CYCLE[3] ),
    .Y(_114_),
    .A1(\PWM_Generador.DUTY_CYCLE[1] ),
    .A2(\PWM_Generador.DUTY_CYCLE[2] ));
 sg13g2_nand3b_1 _247_ (.B(\PWM_Generador.PWM_DFF1.Q ),
    .C(_114_),
    .Y(_115_),
    .A_N(\PWM_Generador.PWM_DFF2.Q ));
 sg13g2_nor4_2 _248_ (.A(_104_),
    .B(_106_),
    .C(_112_),
    .Y(_116_),
    .D(_115_));
 sg13g2_or4_1 _249_ (.A(_104_),
    .B(_106_),
    .C(_112_),
    .D(_115_),
    .X(_117_));
 sg13g2_or3_1 _250_ (.A(\PWM_Generador.DUTY_CYCLE[1] ),
    .B(\PWM_Generador.DUTY_CYCLE[0] ),
    .C(\PWM_Generador.DUTY_CYCLE[2] ),
    .X(_118_));
 sg13g2_nor2b_1 _251_ (.A(_116_),
    .B_N(\PWM_Generador.DUTY_CYCLE[1] ),
    .Y(_119_));
 sg13g2_xnor2_1 _252_ (.Y(_120_),
    .A(\PWM_Generador.DUTY_CYCLE[1] ),
    .B(_116_));
 sg13g2_and2_1 _253_ (.A(\PWM_Generador.DUTY_CYCLE[0] ),
    .B(_120_),
    .X(_121_));
 sg13g2_xnor2_1 _254_ (.Y(_122_),
    .A(\PWM_Generador.DUTY_CYCLE[2] ),
    .B(_116_));
 sg13g2_o21ai_1 _255_ (.B1(_122_),
    .Y(_123_),
    .A1(_119_),
    .A2(_121_));
 sg13g2_nand2_1 _256_ (.Y(_124_),
    .A(\PWM_Generador.PWM_DFF3.Q ),
    .B(_113_));
 sg13g2_nor2_1 _257_ (.A(\PWM_Generador.DUTY_CYCLE[3] ),
    .B(_118_),
    .Y(_125_));
 sg13g2_nor3_1 _258_ (.A(\PWM_Generador.PWM_DFF4.Q ),
    .B(_124_),
    .C(_125_),
    .Y(_126_));
 sg13g2_o21ai_1 _259_ (.B1(_117_),
    .Y(_127_),
    .A1(\PWM_Generador.DUTY_CYCLE[2] ),
    .A2(_126_));
 sg13g2_a22oi_1 _260_ (.Y(_128_),
    .B1(_123_),
    .B2(_127_),
    .A2(_118_),
    .A1(_117_));
 sg13g2_xor2_1 _261_ (.B(_128_),
    .A(\PWM_Generador.DUTY_CYCLE[3] ),
    .X(_094_));
 sg13g2_nor2_2 _262_ (.A(_116_),
    .B(_126_),
    .Y(_129_));
 sg13g2_nand2_1 _263_ (.Y(_130_),
    .A(_221_),
    .B(_129_));
 sg13g2_or3_1 _264_ (.A(_119_),
    .B(_121_),
    .C(_122_),
    .X(_131_));
 sg13g2_and2_1 _265_ (.A(_123_),
    .B(_131_),
    .X(_132_));
 sg13g2_o21ai_1 _266_ (.B1(_130_),
    .Y(_093_),
    .A1(_129_),
    .A2(_132_));
 sg13g2_nand2_1 _267_ (.Y(_133_),
    .A(\PWM_Generador.DUTY_CYCLE[1] ),
    .B(_129_));
 sg13g2_xnor2_1 _268_ (.Y(_134_),
    .A(\PWM_Generador.DUTY_CYCLE[0] ),
    .B(_120_));
 sg13g2_o21ai_1 _269_ (.B1(_133_),
    .Y(_092_),
    .A1(_129_),
    .A2(_134_));
 sg13g2_mux2_1 _270_ (.A0(\PWM_Generador.DUTY_CYCLE[0] ),
    .A1(_220_),
    .S(_129_),
    .X(_091_));
 sg13g2_nor3_2 _271_ (.A(net5),
    .B(net3),
    .C(net4),
    .Y(_135_));
 sg13g2_nor2b_1 _272_ (.A(net6),
    .B_N(_135_),
    .Y(_136_));
 sg13g2_nand2b_1 _273_ (.Y(_137_),
    .B(_136_),
    .A_N(net7));
 sg13g2_nor2_1 _274_ (.A(net8),
    .B(_137_),
    .Y(_138_));
 sg13g2_xnor2_1 _275_ (.Y(_139_),
    .A(net6),
    .B(_135_));
 sg13g2_xnor2_1 _276_ (.Y(_140_),
    .A(\PWM_Generador.DIV_FREQ.counter[2] ),
    .B(_139_));
 sg13g2_or2_1 _277_ (.X(_141_),
    .B(net71),
    .A(net83));
 sg13g2_nand2_1 _278_ (.Y(_142_),
    .A(net3),
    .B(net4));
 sg13g2_xor2_1 _279_ (.B(net4),
    .A(net3),
    .X(_143_));
 sg13g2_nand2_1 _280_ (.Y(_144_),
    .A(net83),
    .B(net71));
 sg13g2_o21ai_1 _281_ (.B1(net5),
    .Y(_145_),
    .A1(net3),
    .A2(net4));
 sg13g2_a21oi_1 _282_ (.A1(\PWM_Generador.DIV_FREQ.counter[1] ),
    .A2(_142_),
    .Y(_146_),
    .B1(_145_));
 sg13g2_o21ai_1 _283_ (.B1(_144_),
    .Y(_147_),
    .A1(_135_),
    .A2(_146_));
 sg13g2_o21ai_1 _284_ (.B1(_147_),
    .Y(_148_),
    .A1(_141_),
    .A2(_143_));
 sg13g2_xnor2_1 _285_ (.Y(_149_),
    .A(net7),
    .B(_136_));
 sg13g2_a22oi_1 _286_ (.Y(_150_),
    .B1(_149_),
    .B2(_096_),
    .A2(_139_),
    .A1(_097_));
 sg13g2_o21ai_1 _287_ (.B1(_150_),
    .Y(_151_),
    .A1(_140_),
    .A2(_148_));
 sg13g2_nand2_1 _288_ (.Y(_152_),
    .A(net8),
    .B(_137_));
 sg13g2_nand2b_1 _289_ (.Y(_153_),
    .B(_040_),
    .A_N(_149_));
 sg13g2_xor2_1 _290_ (.B(_152_),
    .A(\PWM_Generador.DIV_FREQ.counter[4] ),
    .X(_154_));
 sg13g2_nand3_1 _291_ (.B(_153_),
    .C(_154_),
    .A(_151_),
    .Y(_155_));
 sg13g2_a21oi_1 _292_ (.A1(net8),
    .A2(_137_),
    .Y(_156_),
    .B1(net76));
 sg13g2_nor2b_1 _293_ (.A(_156_),
    .B_N(net73),
    .Y(_157_));
 sg13g2_a21oi_2 _294_ (.B1(_138_),
    .Y(_158_),
    .A2(_157_),
    .A1(_155_));
 sg13g2_mux2_1 _295_ (.A0(net47),
    .A1(net70),
    .S(_158_),
    .X(_090_));
 sg13g2_nor2_1 _296_ (.A(net71),
    .B(_158_),
    .Y(_032_));
 sg13g2_nand2_1 _297_ (.Y(_159_),
    .A(_141_),
    .B(_144_));
 sg13g2_nor2_1 _298_ (.A(_158_),
    .B(_159_),
    .Y(_033_));
 sg13g2_and2_1 _299_ (.A(net79),
    .B(_144_),
    .X(_160_));
 sg13g2_nor2_1 _300_ (.A(net79),
    .B(_144_),
    .Y(_161_));
 sg13g2_nor3_1 _301_ (.A(_158_),
    .B(net80),
    .C(_161_),
    .Y(_034_));
 sg13g2_xnor2_1 _302_ (.Y(_162_),
    .A(_096_),
    .B(_161_));
 sg13g2_nor2_1 _303_ (.A(_158_),
    .B(net82),
    .Y(_035_));
 sg13g2_nand4_1 _304_ (.B(\PWM_Generador.DIV_FREQ.counter[2] ),
    .C(\PWM_Generador.DIV_FREQ.counter[1] ),
    .A(\PWM_Generador.DIV_FREQ.counter[3] ),
    .Y(_163_),
    .D(net71));
 sg13g2_nor2_1 _305_ (.A(net76),
    .B(_163_),
    .Y(_164_));
 sg13g2_and2_1 _306_ (.A(net76),
    .B(_163_),
    .X(_165_));
 sg13g2_nor3_1 _307_ (.A(_158_),
    .B(_164_),
    .C(net77),
    .Y(_036_));
 sg13g2_xor2_1 _308_ (.B(_164_),
    .A(net73),
    .X(_166_));
 sg13g2_nor2_1 _309_ (.A(_158_),
    .B(net74),
    .Y(_037_));
 sg13g2_and4_1 _310_ (.A(_095_),
    .B(_107_),
    .C(_110_),
    .D(_111_),
    .X(_004_));
 sg13g2_nor2_1 _311_ (.A(\PWM_Generador.counter_PWM[0] ),
    .B(\PWM_Generador.counter_PWM[1] ),
    .Y(_167_));
 sg13g2_a21oi_1 _312_ (.A1(_101_),
    .A2(_167_),
    .Y(_168_),
    .B1(_100_));
 sg13g2_nor2_1 _313_ (.A(\PWM_Generador.counter_PWM[0] ),
    .B(_168_),
    .Y(_000_));
 sg13g2_and2_1 _314_ (.A(\PWM_Generador.counter_PWM[0] ),
    .B(\PWM_Generador.counter_PWM[1] ),
    .X(_169_));
 sg13g2_nor3_1 _315_ (.A(\PWM_Generador.counter_PWM[3] ),
    .B(_167_),
    .C(_169_),
    .Y(_001_));
 sg13g2_a21oi_1 _316_ (.A1(\PWM_Generador.counter_PWM[2] ),
    .A2(_169_),
    .Y(_170_),
    .B1(\PWM_Generador.counter_PWM[3] ));
 sg13g2_o21ai_1 _317_ (.B1(_170_),
    .Y(_171_),
    .A1(\PWM_Generador.counter_PWM[2] ),
    .A2(_169_));
 sg13g2_inv_1 _318_ (.Y(_002_),
    .A(_171_));
 sg13g2_nor2_1 _319_ (.A(_168_),
    .B(_170_),
    .Y(_003_));
 sg13g2_nand2_1 _320_ (.Y(_172_),
    .A(\PWM_Generador.DUTY_CYCLE[3] ),
    .B(_100_));
 sg13g2_nand2b_1 _321_ (.Y(_173_),
    .B(\PWM_Generador.counter_PWM[1] ),
    .A_N(\PWM_Generador.DUTY_CYCLE[1] ));
 sg13g2_nor2b_1 _322_ (.A(\PWM_Generador.counter_PWM[0] ),
    .B_N(\PWM_Generador.DUTY_CYCLE[0] ),
    .Y(_174_));
 sg13g2_nor2b_1 _323_ (.A(\PWM_Generador.counter_PWM[1] ),
    .B_N(\PWM_Generador.DUTY_CYCLE[1] ),
    .Y(_175_));
 sg13g2_a221oi_1 _324_ (.B2(_174_),
    .C1(_175_),
    .B1(_173_),
    .A1(\PWM_Generador.DUTY_CYCLE[2] ),
    .Y(_176_),
    .A2(_101_));
 sg13g2_nand2b_1 _325_ (.Y(_177_),
    .B(\PWM_Generador.counter_PWM[3] ),
    .A_N(\PWM_Generador.DUTY_CYCLE[3] ));
 sg13g2_o21ai_1 _326_ (.B1(_177_),
    .Y(_178_),
    .A1(\PWM_Generador.DUTY_CYCLE[2] ),
    .A2(_101_));
 sg13g2_o21ai_1 _327_ (.B1(_172_),
    .Y(\PWM_Generador.pwm_out0 ),
    .A1(_176_),
    .A2(_178_));
 sg13g2_o21ai_1 _328_ (.B1(_124_),
    .Y(_086_),
    .A1(_098_),
    .A2(_113_));
 sg13g2_nand2_1 _329_ (.Y(_179_),
    .A(net2),
    .B(_113_));
 sg13g2_o21ai_1 _330_ (.B1(_179_),
    .Y(_087_),
    .A1(_099_),
    .A2(_113_));
 sg13g2_mux2_1 _331_ (.A0(\PWM_Generador.PWM_DFF2.Q ),
    .A1(\PWM_Generador.PWM_DFF1.Q ),
    .S(_113_),
    .X(_088_));
 sg13g2_mux2_1 _332_ (.A0(\PWM_Generador.PWM_DFF1.Q ),
    .A1(net1),
    .S(_113_),
    .X(_089_));
 sg13g2_inv_1 _333_ (.Y(_044_),
    .A(net55));
 sg13g2_inv_1 _334_ (.Y(_045_),
    .A(net50));
 sg13g2_inv_1 _335_ (.Y(_046_),
    .A(net55));
 sg13g2_inv_1 _336_ (.Y(_047_),
    .A(net51));
 sg13g2_inv_1 _337_ (.Y(_048_),
    .A(net54));
 sg13g2_inv_1 _338_ (.Y(_049_),
    .A(net54));
 sg13g2_inv_1 _339_ (.Y(_050_),
    .A(net54));
 sg13g2_inv_1 _340_ (.Y(_051_),
    .A(net54));
 sg13g2_inv_1 _341_ (.Y(_052_),
    .A(net51));
 sg13g2_inv_1 _342_ (.Y(_053_),
    .A(net54));
 sg13g2_inv_1 _343_ (.Y(_054_),
    .A(net51));
 sg13g2_inv_1 _344_ (.Y(_055_),
    .A(net51));
 sg13g2_inv_1 _345_ (.Y(_056_),
    .A(net51));
 sg13g2_inv_1 _346_ (.Y(_057_),
    .A(net51));
 sg13g2_inv_1 _347_ (.Y(_058_),
    .A(net52));
 sg13g2_inv_1 _348_ (.Y(_059_),
    .A(net49));
 sg13g2_inv_1 _349_ (.Y(_060_),
    .A(net49));
 sg13g2_inv_1 _350_ (.Y(_061_),
    .A(net49));
 sg13g2_inv_1 _351_ (.Y(_062_),
    .A(net49));
 sg13g2_inv_1 _352_ (.Y(_063_),
    .A(net50));
 sg13g2_inv_1 _353_ (.Y(_064_),
    .A(net53));
 sg13g2_inv_1 _354_ (.Y(_065_),
    .A(net53));
 sg13g2_inv_1 _355_ (.Y(_066_),
    .A(net53));
 sg13g2_inv_1 _356_ (.Y(_067_),
    .A(net50));
 sg13g2_inv_1 _357_ (.Y(_068_),
    .A(net50));
 sg13g2_inv_1 _358_ (.Y(_069_),
    .A(net50));
 sg13g2_inv_1 _359_ (.Y(_070_),
    .A(net50));
 sg13g2_inv_1 _360_ (.Y(_071_),
    .A(net49));
 sg13g2_inv_1 _361_ (.Y(_072_),
    .A(net49));
 sg13g2_inv_1 _362_ (.Y(_073_),
    .A(net49));
 sg13g2_inv_1 _363_ (.Y(_074_),
    .A(net49));
 sg13g2_inv_1 _364_ (.Y(_075_),
    .A(net52));
 sg13g2_inv_1 _365_ (.Y(_076_),
    .A(net53));
 sg13g2_inv_1 _366_ (.Y(_077_),
    .A(net52));
 sg13g2_inv_1 _367_ (.Y(_078_),
    .A(net53));
 sg13g2_inv_1 _368_ (.Y(_079_),
    .A(net52));
 sg13g2_inv_1 _369_ (.Y(_080_),
    .A(net52));
 sg13g2_inv_1 _370_ (.Y(_081_),
    .A(net52));
 sg13g2_inv_1 _371_ (.Y(_082_),
    .A(net52));
 sg13g2_inv_1 _372_ (.Y(_083_),
    .A(net53));
 sg13g2_inv_1 _373_ (.Y(_084_),
    .A(net52));
 sg13g2_inv_1 _374_ (.Y(_085_),
    .A(net54));
 sg13g2_dfrbp_1 _375_ (.CLK(net47),
    .RESET_B(net66),
    .D(_086_),
    .Q_N(_219_),
    .Q(\PWM_Generador.PWM_DFF4.Q ));
 sg13g2_dfrbp_1 _376_ (.CLK(net47),
    .RESET_B(net69),
    .D(_087_),
    .Q_N(_218_),
    .Q(\PWM_Generador.PWM_DFF3.Q ));
 sg13g2_dfrbp_1 _377_ (.CLK(net47),
    .RESET_B(net68),
    .D(_088_),
    .Q_N(_217_),
    .Q(\PWM_Generador.PWM_DFF2.Q ));
 sg13g2_dfrbp_1 _378_ (.CLK(net47),
    .RESET_B(net67),
    .D(_089_),
    .Q_N(_216_),
    .Q(\PWM_Generador.PWM_DFF1.Q ));
 sg13g2_dfrbp_1 _379_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(_043_),
    .D(_090_),
    .Q_N(_038_),
    .Q(\PWM_Generador.DIV_FREQ.clk_out ));
 sg13g2_dfrbp_1 _380_ (.CLK(net48),
    .RESET_B(_044_),
    .D(_091_),
    .Q_N(\PWM_Generador.DUTY_CYCLE[0] ),
    .Q(_220_));
 sg13g2_dfrbp_1 _381_ (.CLK(net48),
    .RESET_B(_045_),
    .D(_092_),
    .Q_N(_215_),
    .Q(\PWM_Generador.DUTY_CYCLE[1] ));
 sg13g2_dfrbp_1 _382_ (.CLK(net44),
    .RESET_B(_046_),
    .D(_093_),
    .Q_N(\PWM_Generador.DUTY_CYCLE[2] ),
    .Q(_221_));
 sg13g2_dfrbp_1 _383_ (.CLK(net44),
    .RESET_B(_047_),
    .D(_094_),
    .Q_N(_214_),
    .Q(\PWM_Generador.DUTY_CYCLE[3] ));
 sg13g2_dfrbp_1 _384_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(_048_),
    .D(net72),
    .Q_N(_213_),
    .Q(\PWM_Generador.DIV_FREQ.counter[0] ));
 sg13g2_dfrbp_1 _385_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(_049_),
    .D(_033_),
    .Q_N(_212_),
    .Q(\PWM_Generador.DIV_FREQ.counter[1] ));
 sg13g2_dfrbp_1 _386_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(_050_),
    .D(_034_),
    .Q_N(_042_),
    .Q(\PWM_Generador.DIV_FREQ.counter[2] ));
 sg13g2_dfrbp_1 _387_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(_051_),
    .D(_035_),
    .Q_N(_040_),
    .Q(\PWM_Generador.DIV_FREQ.counter[3] ));
 sg13g2_dfrbp_1 _388_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(_052_),
    .D(net78),
    .Q_N(_041_),
    .Q(\PWM_Generador.DIV_FREQ.counter[4] ));
 sg13g2_dfrbp_1 _389_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(_053_),
    .D(net75),
    .Q_N(_039_),
    .Q(\PWM_Generador.DIV_FREQ.counter[5] ));
 sg13g2_dfrbp_1 _390_ (.CLK(net44),
    .RESET_B(_054_),
    .D(_000_),
    .Q_N(_211_),
    .Q(\PWM_Generador.counter_PWM[0] ));
 sg13g2_dfrbp_1 _391_ (.CLK(net44),
    .RESET_B(_055_),
    .D(_001_),
    .Q_N(_210_),
    .Q(\PWM_Generador.counter_PWM[1] ));
 sg13g2_dfrbp_1 _392_ (.CLK(net44),
    .RESET_B(_056_),
    .D(_002_),
    .Q_N(_209_),
    .Q(\PWM_Generador.counter_PWM[2] ));
 sg13g2_dfrbp_1 _393_ (.CLK(net44),
    .RESET_B(_057_),
    .D(_003_),
    .Q_N(_208_),
    .Q(\PWM_Generador.counter_PWM[3] ));
 sg13g2_dfrbp_1 _394_ (.CLK(net46),
    .RESET_B(_058_),
    .D(_004_),
    .Q_N(_207_),
    .Q(\PWM_Generador.counter_debounce[0] ));
 sg13g2_dfrbp_1 _395_ (.CLK(net42),
    .RESET_B(_059_),
    .D(net65),
    .Q_N(_206_),
    .Q(\PWM_Generador.counter_debounce[1] ));
 sg13g2_dfrbp_1 _396_ (.CLK(net42),
    .RESET_B(_060_),
    .D(net64),
    .Q_N(_205_),
    .Q(\PWM_Generador.counter_debounce[2] ));
 sg13g2_dfrbp_1 _397_ (.CLK(net42),
    .RESET_B(_061_),
    .D(net63),
    .Q_N(_204_),
    .Q(\PWM_Generador.counter_debounce[3] ));
 sg13g2_dfrbp_1 _398_ (.CLK(net42),
    .RESET_B(_062_),
    .D(net62),
    .Q_N(_203_),
    .Q(\PWM_Generador.counter_debounce[4] ));
 sg13g2_dfrbp_1 _399_ (.CLK(net43),
    .RESET_B(_063_),
    .D(net61),
    .Q_N(_202_),
    .Q(\PWM_Generador.counter_debounce[5] ));
 sg13g2_dfrbp_1 _400_ (.CLK(net45),
    .RESET_B(_064_),
    .D(net60),
    .Q_N(_201_),
    .Q(\PWM_Generador.counter_debounce[6] ));
 sg13g2_dfrbp_1 _401_ (.CLK(net45),
    .RESET_B(_065_),
    .D(net59),
    .Q_N(_200_),
    .Q(\PWM_Generador.counter_debounce[7] ));
 sg13g2_dfrbp_1 _402_ (.CLK(net45),
    .RESET_B(_066_),
    .D(net58),
    .Q_N(_199_),
    .Q(\PWM_Generador.counter_debounce[8] ));
 sg13g2_dfrbp_1 _403_ (.CLK(net43),
    .RESET_B(_067_),
    .D(net57),
    .Q_N(_198_),
    .Q(\PWM_Generador.counter_debounce[9] ));
 sg13g2_dfrbp_1 _404_ (.CLK(net43),
    .RESET_B(_068_),
    .D(net56),
    .Q_N(_197_),
    .Q(\PWM_Generador.counter_debounce[10] ));
 sg13g2_dfrbp_1 _405_ (.CLK(net43),
    .RESET_B(_069_),
    .D(net41),
    .Q_N(_196_),
    .Q(\PWM_Generador.counter_debounce[11] ));
 sg13g2_dfrbp_1 _406_ (.CLK(net43),
    .RESET_B(_070_),
    .D(net40),
    .Q_N(_195_),
    .Q(\PWM_Generador.counter_debounce[12] ));
 sg13g2_dfrbp_1 _407_ (.CLK(net42),
    .RESET_B(_071_),
    .D(net39),
    .Q_N(_194_),
    .Q(\PWM_Generador.counter_debounce[13] ));
 sg13g2_dfrbp_1 _408_ (.CLK(net42),
    .RESET_B(_072_),
    .D(net38),
    .Q_N(_193_),
    .Q(\PWM_Generador.counter_debounce[14] ));
 sg13g2_dfrbp_1 _409_ (.CLK(net42),
    .RESET_B(_073_),
    .D(net37),
    .Q_N(_192_),
    .Q(\PWM_Generador.counter_debounce[15] ));
 sg13g2_dfrbp_1 _410_ (.CLK(net42),
    .RESET_B(_074_),
    .D(net36),
    .Q_N(_191_),
    .Q(\PWM_Generador.counter_debounce[16] ));
 sg13g2_dfrbp_1 _411_ (.CLK(net46),
    .RESET_B(_075_),
    .D(net35),
    .Q_N(_190_),
    .Q(\PWM_Generador.counter_debounce[17] ));
 sg13g2_dfrbp_1 _412_ (.CLK(net45),
    .RESET_B(_076_),
    .D(net34),
    .Q_N(_189_),
    .Q(\PWM_Generador.counter_debounce[18] ));
 sg13g2_dfrbp_1 _413_ (.CLK(net45),
    .RESET_B(_077_),
    .D(net33),
    .Q_N(_188_),
    .Q(\PWM_Generador.counter_debounce[19] ));
 sg13g2_dfrbp_1 _414_ (.CLK(net45),
    .RESET_B(_078_),
    .D(net32),
    .Q_N(_187_),
    .Q(\PWM_Generador.counter_debounce[20] ));
 sg13g2_dfrbp_1 _415_ (.CLK(net46),
    .RESET_B(_079_),
    .D(net31),
    .Q_N(_186_),
    .Q(\PWM_Generador.counter_debounce[21] ));
 sg13g2_dfrbp_1 _416_ (.CLK(net46),
    .RESET_B(_080_),
    .D(net30),
    .Q_N(_185_),
    .Q(\PWM_Generador.counter_debounce[22] ));
 sg13g2_dfrbp_1 _417_ (.CLK(net45),
    .RESET_B(_081_),
    .D(net29),
    .Q_N(_184_),
    .Q(\PWM_Generador.counter_debounce[23] ));
 sg13g2_dfrbp_1 _418_ (.CLK(net45),
    .RESET_B(_082_),
    .D(net28),
    .Q_N(_183_),
    .Q(\PWM_Generador.counter_debounce[24] ));
 sg13g2_dfrbp_1 _419_ (.CLK(net48),
    .RESET_B(_083_),
    .D(net27),
    .Q_N(_182_),
    .Q(\PWM_Generador.counter_debounce[25] ));
 sg13g2_dfrbp_1 _420_ (.CLK(net47),
    .RESET_B(_084_),
    .D(net26),
    .Q_N(_181_),
    .Q(\PWM_Generador.counter_debounce[26] ));
 sg13g2_dfrbp_1 _421_ (.CLK(net48),
    .RESET_B(_085_),
    .D(net25),
    .Q_N(_180_),
    .Q(\PWM_Generador.counter_debounce[27] ));
 sg13g2_tiehi _378__53 (.L_HI(net67));
 sg13g2_tiehi _377__54 (.L_HI(net68));
 sg13g2_tiehi _376__55 (.L_HI(net69));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_pwm_top_10 (.L_LO(net10));
 sg13g2_tielo tt_um_pwm_top_11 (.L_LO(net11));
 sg13g2_tielo tt_um_pwm_top_12 (.L_LO(net12));
 sg13g2_tielo tt_um_pwm_top_13 (.L_LO(net13));
 sg13g2_tielo tt_um_pwm_top_14 (.L_LO(net14));
 sg13g2_tielo tt_um_pwm_top_15 (.L_LO(net15));
 sg13g2_tielo tt_um_pwm_top_16 (.L_LO(net16));
 sg13g2_tielo tt_um_pwm_top_17 (.L_LO(net17));
 sg13g2_tielo tt_um_pwm_top_18 (.L_LO(net18));
 sg13g2_tielo tt_um_pwm_top_19 (.L_LO(net19));
 sg13g2_tielo tt_um_pwm_top_20 (.L_LO(net20));
 sg13g2_tielo tt_um_pwm_top_21 (.L_LO(net21));
 sg13g2_tielo tt_um_pwm_top_22 (.L_LO(net22));
 sg13g2_tielo tt_um_pwm_top_23 (.L_LO(net23));
 sg13g2_tielo tt_um_pwm_top_24 (.L_LO(net24));
 sg13g2_tielo _421__25 (.L_LO(net25));
 sg13g2_tielo _420__26 (.L_LO(net26));
 sg13g2_tielo _419__27 (.L_LO(net27));
 sg13g2_tielo _418__28 (.L_LO(net28));
 sg13g2_tielo _417__29 (.L_LO(net29));
 sg13g2_tielo _416__30 (.L_LO(net30));
 sg13g2_tielo _415__31 (.L_LO(net31));
 sg13g2_tielo _414__32 (.L_LO(net32));
 sg13g2_tielo _413__33 (.L_LO(net33));
 sg13g2_tielo _412__34 (.L_LO(net34));
 sg13g2_tielo _411__35 (.L_LO(net35));
 sg13g2_tielo _410__36 (.L_LO(net36));
 sg13g2_tielo _409__37 (.L_LO(net37));
 sg13g2_tielo _408__38 (.L_LO(net38));
 sg13g2_tielo _407__39 (.L_LO(net39));
 sg13g2_tielo _406__40 (.L_LO(net40));
 sg13g2_tielo _405__41 (.L_LO(net41));
 sg13g2_tielo _404__42 (.L_LO(net56));
 sg13g2_tielo _403__43 (.L_LO(net57));
 sg13g2_tielo _402__44 (.L_LO(net58));
 sg13g2_tielo _401__45 (.L_LO(net59));
 sg13g2_tielo _400__46 (.L_LO(net60));
 sg13g2_tielo _399__47 (.L_LO(net61));
 sg13g2_tielo _398__48 (.L_LO(net62));
 sg13g2_tielo _397__49 (.L_LO(net63));
 sg13g2_tielo _396__50 (.L_LO(net64));
 sg13g2_tielo _395__51 (.L_LO(net65));
 sg13g2_tiehi _375__52 (.L_HI(net66));
 sg13g2_buf_1 _469_ (.A(\PWM_Generador.pwm_out0 ),
    .X(uo_out[0]));
 sg13g2_buf_1 _470_ (.A(\PWM_Generador.pwm_out0 ),
    .X(uo_out[1]));
 sg13g2_buf_1 _471_ (.A(\PWM_Generador.pwm_out0 ),
    .X(uo_out[2]));
 sg13g2_buf_1 _472_ (.A(\PWM_Generador.pwm_out0 ),
    .X(uo_out[3]));
 sg13g2_buf_1 _473_ (.A(\PWM_Generador.pwm_out0 ),
    .X(uo_out[4]));
 sg13g2_buf_1 _474_ (.A(\PWM_Generador.pwm_out0 ),
    .X(uo_out[5]));
 sg13g2_buf_1 _475_ (.A(\PWM_Generador.pwm_out0 ),
    .X(uo_out[6]));
 sg13g2_buf_1 _476_ (.A(\PWM_Generador.pwm_out0 ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout42 (.A(net44),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(net44),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(net48),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(net47),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(\PWM_Generador.DIV_FREQ.clk_out ),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(net51),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(net51),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(net55),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(net53),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(net54),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(rst_n),
    .X(net55));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_pwm_top_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_038_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold2 (.A(\PWM_Generador.DIV_FREQ.counter[0] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold3 (.A(_032_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold4 (.A(_039_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold5 (.A(_166_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold6 (.A(_037_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold7 (.A(_041_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold8 (.A(_165_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold9 (.A(_036_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold10 (.A(_042_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold11 (.A(_160_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold12 (.A(_040_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold13 (.A(_162_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold14 (.A(\PWM_Generador.DIV_FREQ.counter[1] ),
    .X(net83));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_fill_2 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_4 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_275 ();
 sg13g2_decap_8 FILLER_21_282 ();
 sg13g2_decap_8 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_296 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_307 ();
 sg13g2_fill_2 FILLER_21_314 ();
 sg13g2_fill_1 FILLER_21_316 ();
 sg13g2_fill_2 FILLER_21_321 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_4 FILLER_21_334 ();
 sg13g2_decap_4 FILLER_21_364 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_4 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_4 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_fill_2 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_4 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_4 FILLER_24_210 ();
 sg13g2_fill_2 FILLER_24_214 ();
 sg13g2_decap_4 FILLER_24_294 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_367 ();
 sg13g2_decap_4 FILLER_24_374 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_decap_8 FILLER_25_230 ();
 sg13g2_decap_4 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_246 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_259 ();
 sg13g2_decap_4 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_298 ();
 sg13g2_decap_4 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_fill_2 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_decap_4 FILLER_26_174 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_decap_4 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_241 ();
 sg13g2_decap_8 FILLER_26_248 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_decap_4 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_331 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_decap_4 FILLER_26_348 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_decap_4 FILLER_27_247 ();
 sg13g2_decap_4 FILLER_27_277 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_decap_4 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_4 FILLER_28_154 ();
 sg13g2_fill_1 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_fill_2 FILLER_28_229 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_fill_2 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_decap_4 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_decap_4 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_4 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_fill_2 FILLER_29_163 ();
 sg13g2_fill_1 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_fill_2 FILLER_29_186 ();
 sg13g2_fill_1 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_215 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_decap_4 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_decap_4 FILLER_29_277 ();
 sg13g2_fill_2 FILLER_29_304 ();
 sg13g2_decap_4 FILLER_29_332 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_decap_4 FILLER_30_185 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_decap_4 FILLER_30_194 ();
 sg13g2_fill_1 FILLER_30_198 ();
 sg13g2_decap_4 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_decap_4 FILLER_30_220 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_236 ();
 sg13g2_decap_4 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_262 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_decap_4 FILLER_30_285 ();
 sg13g2_decap_4 FILLER_30_297 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_314 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_4 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_158 ();
 sg13g2_decap_4 FILLER_31_216 ();
 sg13g2_decap_4 FILLER_31_230 ();
 sg13g2_fill_1 FILLER_31_234 ();
 sg13g2_decap_4 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_372 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_398 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_4 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_195 ();
 sg13g2_decap_8 FILLER_32_202 ();
 sg13g2_decap_8 FILLER_32_209 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_4 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_293 ();
 sg13g2_decap_4 FILLER_32_303 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_4 FILLER_33_224 ();
 sg13g2_fill_2 FILLER_33_228 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_4 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_decap_4 FILLER_34_280 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_288 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_303 ();
 sg13g2_decap_8 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_231 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_decap_4 FILLER_35_371 ();
 sg13g2_fill_1 FILLER_35_375 ();
 sg13g2_fill_2 FILLER_35_383 ();
 sg13g2_fill_2 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_4 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_4 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_332 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

module tt_um_roy1707018 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire \ascon_inst.en ;
 wire \buffer_out[0] ;
 wire \buffer_out[1] ;
 wire \buffer_out[2] ;
 wire \buffer_out[3] ;
 wire \buffer_out[4] ;
 wire \buffer_out[5] ;
 wire \buffer_out[6] ;
 wire \buffer_out[7] ;
 wire \ro_buffer_counter_inst.ro1_A.cq4 ;
 wire \ro_buffer_counter_inst.ro1_A.en ;
 wire \ro_buffer_counter_inst.ro1_A.q ;
 wire \ro_buffer_counter_inst.ro1_A.q0 ;
 wire \ro_buffer_counter_inst.ro1_A.q1 ;
 wire \ro_buffer_counter_inst.ro1_A.q2 ;
 wire \ro_buffer_counter_inst.ro1_A.q3 ;
 wire \ro_buffer_counter_inst.ro1_A.q4 ;
 wire \ro_buffer_counter_inst.ro1_B.cq4 ;
 wire \ro_buffer_counter_inst.ro1_B.q ;
 wire \ro_buffer_counter_inst.ro1_B.q0 ;
 wire \ro_buffer_counter_inst.ro1_B.q1 ;
 wire \ro_buffer_counter_inst.ro1_B.q2 ;
 wire \ro_buffer_counter_inst.ro1_B.q3 ;
 wire \ro_buffer_counter_inst.ro1_B.q4 ;
 wire \ro_buffer_counter_inst.ro1_C.cq4 ;
 wire \ro_buffer_counter_inst.ro1_C.q ;
 wire \ro_buffer_counter_inst.ro1_C.q0 ;
 wire \ro_buffer_counter_inst.ro1_C.q1 ;
 wire \ro_buffer_counter_inst.ro1_C.q2 ;
 wire \ro_buffer_counter_inst.ro1_C.q3 ;
 wire \ro_buffer_counter_inst.ro1_C.q4 ;
 wire \ro_buffer_counter_inst.ro1_D.cq4 ;
 wire \ro_buffer_counter_inst.ro1_D.q ;
 wire \ro_buffer_counter_inst.ro1_D.q0 ;
 wire \ro_buffer_counter_inst.ro1_D.q1 ;
 wire \ro_buffer_counter_inst.ro1_D.q2 ;
 wire \ro_buffer_counter_inst.ro1_D.q3 ;
 wire \ro_buffer_counter_inst.ro1_D.q4 ;
 wire \ro_buffer_counter_inst.ro1_E.cq4 ;
 wire \ro_buffer_counter_inst.ro1_E.q ;
 wire \ro_buffer_counter_inst.ro1_E.q0 ;
 wire \ro_buffer_counter_inst.ro1_E.q1 ;
 wire \ro_buffer_counter_inst.ro1_E.q2 ;
 wire \ro_buffer_counter_inst.ro1_E.q3 ;
 wire \ro_buffer_counter_inst.ro1_E.q4 ;
 wire \ro_buffer_counter_inst.ro1_F.cq4 ;
 wire \ro_buffer_counter_inst.ro1_F.q ;
 wire \ro_buffer_counter_inst.ro1_F.q0 ;
 wire \ro_buffer_counter_inst.ro1_F.q1 ;
 wire \ro_buffer_counter_inst.ro1_F.q2 ;
 wire \ro_buffer_counter_inst.ro1_F.q3 ;
 wire \ro_buffer_counter_inst.ro1_F.q4 ;
 wire \ro_buffer_counter_inst.ro1_G.cq4 ;
 wire \ro_buffer_counter_inst.ro1_G.q ;
 wire \ro_buffer_counter_inst.ro1_G.q0 ;
 wire \ro_buffer_counter_inst.ro1_G.q1 ;
 wire \ro_buffer_counter_inst.ro1_G.q2 ;
 wire \ro_buffer_counter_inst.ro1_G.q3 ;
 wire \ro_buffer_counter_inst.ro1_G.q4 ;
 wire \ro_buffer_counter_inst.ro1_H.cq4 ;
 wire \ro_buffer_counter_inst.ro1_H.q ;
 wire \ro_buffer_counter_inst.ro1_H.q0 ;
 wire \ro_buffer_counter_inst.ro1_H.q1 ;
 wire \ro_buffer_counter_inst.ro1_H.q2 ;
 wire \ro_buffer_counter_inst.ro1_H.q3 ;
 wire \ro_buffer_counter_inst.ro1_H.q4 ;
 wire \ro_buffer_counter_inst.ro2_A.cq4 ;
 wire \ro_buffer_counter_inst.ro2_A.en ;
 wire \ro_buffer_counter_inst.ro2_A.q ;
 wire \ro_buffer_counter_inst.ro2_A.q0 ;
 wire \ro_buffer_counter_inst.ro2_A.q1 ;
 wire \ro_buffer_counter_inst.ro2_A.q2 ;
 wire \ro_buffer_counter_inst.ro2_A.q3 ;
 wire \ro_buffer_counter_inst.ro2_A.q4 ;
 wire \ro_buffer_counter_inst.ro2_B.cq4 ;
 wire \ro_buffer_counter_inst.ro2_B.q ;
 wire \ro_buffer_counter_inst.ro2_B.q0 ;
 wire \ro_buffer_counter_inst.ro2_B.q1 ;
 wire \ro_buffer_counter_inst.ro2_B.q2 ;
 wire \ro_buffer_counter_inst.ro2_B.q3 ;
 wire \ro_buffer_counter_inst.ro2_B.q4 ;
 wire \ro_buffer_counter_inst.ro2_C.cq4 ;
 wire \ro_buffer_counter_inst.ro2_C.q ;
 wire \ro_buffer_counter_inst.ro2_C.q0 ;
 wire \ro_buffer_counter_inst.ro2_C.q1 ;
 wire \ro_buffer_counter_inst.ro2_C.q2 ;
 wire \ro_buffer_counter_inst.ro2_C.q3 ;
 wire \ro_buffer_counter_inst.ro2_C.q4 ;
 wire \ro_buffer_counter_inst.ro2_D.cq4 ;
 wire \ro_buffer_counter_inst.ro2_D.q ;
 wire \ro_buffer_counter_inst.ro2_D.q0 ;
 wire \ro_buffer_counter_inst.ro2_D.q1 ;
 wire \ro_buffer_counter_inst.ro2_D.q2 ;
 wire \ro_buffer_counter_inst.ro2_D.q3 ;
 wire \ro_buffer_counter_inst.ro2_D.q4 ;
 wire \ro_buffer_counter_inst.ro2_E.cq4 ;
 wire \ro_buffer_counter_inst.ro2_E.q ;
 wire \ro_buffer_counter_inst.ro2_E.q0 ;
 wire \ro_buffer_counter_inst.ro2_E.q1 ;
 wire \ro_buffer_counter_inst.ro2_E.q2 ;
 wire \ro_buffer_counter_inst.ro2_E.q3 ;
 wire \ro_buffer_counter_inst.ro2_E.q4 ;
 wire \ro_buffer_counter_inst.ro2_F.cq4 ;
 wire \ro_buffer_counter_inst.ro2_F.q ;
 wire \ro_buffer_counter_inst.ro2_F.q0 ;
 wire \ro_buffer_counter_inst.ro2_F.q1 ;
 wire \ro_buffer_counter_inst.ro2_F.q2 ;
 wire \ro_buffer_counter_inst.ro2_F.q3 ;
 wire \ro_buffer_counter_inst.ro2_F.q4 ;
 wire \ro_buffer_counter_inst.ro2_G.cq4 ;
 wire \ro_buffer_counter_inst.ro2_G.q ;
 wire \ro_buffer_counter_inst.ro2_G.q0 ;
 wire \ro_buffer_counter_inst.ro2_G.q1 ;
 wire \ro_buffer_counter_inst.ro2_G.q2 ;
 wire \ro_buffer_counter_inst.ro2_G.q3 ;
 wire \ro_buffer_counter_inst.ro2_G.q4 ;
 wire \ro_buffer_counter_inst.ro2_H.cq4 ;
 wire \ro_buffer_counter_inst.ro2_H.q ;
 wire \ro_buffer_counter_inst.ro2_H.q0 ;
 wire \ro_buffer_counter_inst.ro2_H.q1 ;
 wire \ro_buffer_counter_inst.ro2_H.q2 ;
 wire \ro_buffer_counter_inst.ro2_H.q3 ;
 wire \ro_buffer_counter_inst.ro2_H.q4 ;
 wire \ro_buffer_counter_inst.ro_1_reg_A ;
 wire \ro_buffer_counter_inst.ro_1_reg_B ;
 wire \ro_buffer_counter_inst.ro_1_reg_C ;
 wire \ro_buffer_counter_inst.ro_1_reg_D ;
 wire \ro_buffer_counter_inst.ro_1_reg_E ;
 wire \ro_buffer_counter_inst.ro_1_reg_F ;
 wire \ro_buffer_counter_inst.ro_1_reg_G ;
 wire \ro_buffer_counter_inst.ro_1_reg_H ;
 wire \ro_buffer_counter_inst.ro_2_reg_A ;
 wire \ro_buffer_counter_inst.ro_2_reg_B ;
 wire \ro_buffer_counter_inst.ro_2_reg_C ;
 wire \ro_buffer_counter_inst.ro_2_reg_D ;
 wire \ro_buffer_counter_inst.ro_2_reg_E ;
 wire \ro_buffer_counter_inst.ro_2_reg_F ;
 wire \ro_buffer_counter_inst.ro_2_reg_G ;
 wire \ro_buffer_counter_inst.ro_2_reg_H ;
 wire \ro_buffer_counter_inst.shift_register[0] ;
 wire \ro_buffer_counter_inst.shift_register[10] ;
 wire \ro_buffer_counter_inst.shift_register[11] ;
 wire \ro_buffer_counter_inst.shift_register[12] ;
 wire \ro_buffer_counter_inst.shift_register[13] ;
 wire \ro_buffer_counter_inst.shift_register[14] ;
 wire \ro_buffer_counter_inst.shift_register[15] ;
 wire \ro_buffer_counter_inst.shift_register[16] ;
 wire \ro_buffer_counter_inst.shift_register[17] ;
 wire \ro_buffer_counter_inst.shift_register[18] ;
 wire \ro_buffer_counter_inst.shift_register[19] ;
 wire \ro_buffer_counter_inst.shift_register[1] ;
 wire \ro_buffer_counter_inst.shift_register[20] ;
 wire \ro_buffer_counter_inst.shift_register[21] ;
 wire \ro_buffer_counter_inst.shift_register[22] ;
 wire \ro_buffer_counter_inst.shift_register[23] ;
 wire \ro_buffer_counter_inst.shift_register[24] ;
 wire \ro_buffer_counter_inst.shift_register[25] ;
 wire \ro_buffer_counter_inst.shift_register[26] ;
 wire \ro_buffer_counter_inst.shift_register[27] ;
 wire \ro_buffer_counter_inst.shift_register[28] ;
 wire \ro_buffer_counter_inst.shift_register[29] ;
 wire \ro_buffer_counter_inst.shift_register[2] ;
 wire \ro_buffer_counter_inst.shift_register[30] ;
 wire \ro_buffer_counter_inst.shift_register[31] ;
 wire \ro_buffer_counter_inst.shift_register[32] ;
 wire \ro_buffer_counter_inst.shift_register[33] ;
 wire \ro_buffer_counter_inst.shift_register[34] ;
 wire \ro_buffer_counter_inst.shift_register[35] ;
 wire \ro_buffer_counter_inst.shift_register[36] ;
 wire \ro_buffer_counter_inst.shift_register[37] ;
 wire \ro_buffer_counter_inst.shift_register[38] ;
 wire \ro_buffer_counter_inst.shift_register[39] ;
 wire \ro_buffer_counter_inst.shift_register[3] ;
 wire \ro_buffer_counter_inst.shift_register[40] ;
 wire \ro_buffer_counter_inst.shift_register[41] ;
 wire \ro_buffer_counter_inst.shift_register[42] ;
 wire \ro_buffer_counter_inst.shift_register[43] ;
 wire \ro_buffer_counter_inst.shift_register[44] ;
 wire \ro_buffer_counter_inst.shift_register[45] ;
 wire \ro_buffer_counter_inst.shift_register[46] ;
 wire \ro_buffer_counter_inst.shift_register[47] ;
 wire \ro_buffer_counter_inst.shift_register[48] ;
 wire \ro_buffer_counter_inst.shift_register[49] ;
 wire \ro_buffer_counter_inst.shift_register[4] ;
 wire \ro_buffer_counter_inst.shift_register[50] ;
 wire \ro_buffer_counter_inst.shift_register[51] ;
 wire \ro_buffer_counter_inst.shift_register[52] ;
 wire \ro_buffer_counter_inst.shift_register[53] ;
 wire \ro_buffer_counter_inst.shift_register[54] ;
 wire \ro_buffer_counter_inst.shift_register[55] ;
 wire \ro_buffer_counter_inst.shift_register[56] ;
 wire \ro_buffer_counter_inst.shift_register[57] ;
 wire \ro_buffer_counter_inst.shift_register[58] ;
 wire \ro_buffer_counter_inst.shift_register[59] ;
 wire \ro_buffer_counter_inst.shift_register[5] ;
 wire \ro_buffer_counter_inst.shift_register[60] ;
 wire \ro_buffer_counter_inst.shift_register[61] ;
 wire \ro_buffer_counter_inst.shift_register[62] ;
 wire \ro_buffer_counter_inst.shift_register[63] ;
 wire \ro_buffer_counter_inst.shift_register[6] ;
 wire \ro_buffer_counter_inst.shift_register[7] ;
 wire \ro_buffer_counter_inst.shift_register[8] ;
 wire \ro_buffer_counter_inst.shift_register[9] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_0_clk;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;

 sg13g2_nor2_2 _283_ (.A(net123),
    .B(_090_),
    .Y(_091_));
 sg13g2_a22oi_1 _284_ (.Y(_092_),
    .B1(_089_),
    .B2(\ro_buffer_counter_inst.shift_register[8] ),
    .A2(_086_),
    .A1(\ro_buffer_counter_inst.shift_register[0] ));
 sg13g2_a22oi_1 _285_ (.Y(_093_),
    .B1(_091_),
    .B2(\ro_buffer_counter_inst.shift_register[24] ),
    .A2(_085_),
    .A1(\ro_buffer_counter_inst.shift_register[16] ));
 sg13g2_nand3_1 _286_ (.B(_092_),
    .C(_093_),
    .A(_083_),
    .Y(_094_));
 sg13g2_and2_1 _287_ (.A(net123),
    .B(_087_),
    .X(_095_));
 sg13g2_nand2b_1 _288_ (.Y(_096_),
    .B(net107),
    .A_N(\ro_buffer_counter_inst.shift_register[32] ));
 sg13g2_and2_2 _289_ (.A(net123),
    .B(_084_),
    .X(_097_));
 sg13g2_nand2_2 _290_ (.Y(_098_),
    .A(net124),
    .B(_084_));
 sg13g2_a221oi_1 _291_ (.B2(_094_),
    .C1(_097_),
    .B1(_096_),
    .A1(net45),
    .Y(_099_),
    .A2(net109));
 sg13g2_and3_1 _292_ (.X(_100_),
    .A(net3),
    .B(net4),
    .C(net124));
 sg13g2_nand3_1 _293_ (.B(net4),
    .C(net124),
    .A(net3),
    .Y(_101_));
 sg13g2_o21ai_1 _294_ (.B1(_101_),
    .Y(_102_),
    .A1(\ro_buffer_counter_inst.shift_register[48] ),
    .A2(_098_));
 sg13g2_nand2_1 _295_ (.Y(_103_),
    .A(net46),
    .B(net122));
 sg13g2_o21ai_1 _296_ (.B1(_103_),
    .Y(_000_),
    .A1(_099_),
    .A2(_102_));
 sg13g2_a22oi_1 _297_ (.Y(_104_),
    .B1(_089_),
    .B2(\ro_buffer_counter_inst.shift_register[9] ),
    .A2(_086_),
    .A1(net103));
 sg13g2_a221oi_1 _298_ (.B2(net144),
    .C1(net108),
    .B1(_091_),
    .A1(net83),
    .Y(_105_),
    .A2(_085_));
 sg13g2_a22oi_1 _299_ (.Y(_106_),
    .B1(_104_),
    .B2(_105_),
    .A2(net108),
    .A1(_072_));
 sg13g2_a21oi_1 _300_ (.A1(net54),
    .A2(_095_),
    .Y(_107_),
    .B1(net148));
 sg13g2_a21oi_1 _301_ (.A1(net80),
    .A2(_097_),
    .Y(_108_),
    .B1(_100_));
 sg13g2_a22oi_1 _302_ (.Y(_001_),
    .B1(_107_),
    .B2(_108_),
    .A2(net122),
    .A1(_073_));
 sg13g2_a22oi_1 _303_ (.Y(_109_),
    .B1(_091_),
    .B2(\ro_buffer_counter_inst.shift_register[26] ),
    .A2(_085_),
    .A1(\ro_buffer_counter_inst.shift_register[18] ));
 sg13g2_a22oi_1 _304_ (.Y(_110_),
    .B1(_089_),
    .B2(\ro_buffer_counter_inst.shift_register[10] ),
    .A2(_086_),
    .A1(\ro_buffer_counter_inst.shift_register[2] ));
 sg13g2_nand3_1 _305_ (.B(_109_),
    .C(_110_),
    .A(_083_),
    .Y(_111_));
 sg13g2_nand2b_1 _306_ (.Y(_112_),
    .B(net108),
    .A_N(\ro_buffer_counter_inst.shift_register[34] ));
 sg13g2_a221oi_1 _307_ (.B2(_112_),
    .C1(_097_),
    .B1(_111_),
    .A1(\ro_buffer_counter_inst.shift_register[42] ),
    .Y(_113_),
    .A2(net109));
 sg13g2_o21ai_1 _308_ (.B1(_101_),
    .Y(_114_),
    .A1(net37),
    .A2(_098_));
 sg13g2_nand2_1 _309_ (.Y(_115_),
    .A(net27),
    .B(net122));
 sg13g2_o21ai_1 _310_ (.B1(_115_),
    .Y(_002_),
    .A1(_113_),
    .A2(_114_));
 sg13g2_a22oi_1 _311_ (.Y(_116_),
    .B1(_089_),
    .B2(\ro_buffer_counter_inst.shift_register[11] ),
    .A2(_086_),
    .A1(\ro_buffer_counter_inst.shift_register[3] ));
 sg13g2_a221oi_1 _312_ (.B2(\ro_buffer_counter_inst.shift_register[27] ),
    .C1(net107),
    .B1(_091_),
    .A1(\ro_buffer_counter_inst.shift_register[19] ),
    .Y(_117_),
    .A2(_085_));
 sg13g2_a22oi_1 _313_ (.Y(_118_),
    .B1(_116_),
    .B2(_117_),
    .A2(net108),
    .A1(_074_));
 sg13g2_a221oi_1 _314_ (.B2(\ro_buffer_counter_inst.shift_register[43] ),
    .C1(_118_),
    .B1(net109),
    .A1(net123),
    .Y(_119_),
    .A2(_084_));
 sg13g2_o21ai_1 _315_ (.B1(_101_),
    .Y(_120_),
    .A1(\ro_buffer_counter_inst.shift_register[51] ),
    .A2(_098_));
 sg13g2_nand2_1 _316_ (.Y(_121_),
    .A(net39),
    .B(net122));
 sg13g2_o21ai_1 _317_ (.B1(_121_),
    .Y(_003_),
    .A1(_119_),
    .A2(_120_));
 sg13g2_a22oi_1 _318_ (.Y(_122_),
    .B1(_089_),
    .B2(\ro_buffer_counter_inst.shift_register[12] ),
    .A2(_086_),
    .A1(\ro_buffer_counter_inst.shift_register[4] ));
 sg13g2_a221oi_1 _319_ (.B2(\ro_buffer_counter_inst.shift_register[28] ),
    .C1(net107),
    .B1(_091_),
    .A1(\ro_buffer_counter_inst.shift_register[20] ),
    .Y(_123_),
    .A2(_085_));
 sg13g2_a22oi_1 _320_ (.Y(_124_),
    .B1(_122_),
    .B2(_123_),
    .A2(net107),
    .A1(_075_));
 sg13g2_a221oi_1 _321_ (.B2(\ro_buffer_counter_inst.shift_register[44] ),
    .C1(_124_),
    .B1(net109),
    .A1(net123),
    .Y(_125_),
    .A2(_084_));
 sg13g2_o21ai_1 _322_ (.B1(_101_),
    .Y(_126_),
    .A1(\ro_buffer_counter_inst.shift_register[52] ),
    .A2(_098_));
 sg13g2_nand2_1 _323_ (.Y(_127_),
    .A(net41),
    .B(net122));
 sg13g2_o21ai_1 _324_ (.B1(_127_),
    .Y(_004_),
    .A1(_125_),
    .A2(_126_));
 sg13g2_a22oi_1 _325_ (.Y(_128_),
    .B1(_091_),
    .B2(\ro_buffer_counter_inst.shift_register[29] ),
    .A2(_085_),
    .A1(\ro_buffer_counter_inst.shift_register[21] ));
 sg13g2_a22oi_1 _326_ (.Y(_129_),
    .B1(_089_),
    .B2(\ro_buffer_counter_inst.shift_register[13] ),
    .A2(_086_),
    .A1(\ro_buffer_counter_inst.shift_register[5] ));
 sg13g2_nand3_1 _327_ (.B(_128_),
    .C(_129_),
    .A(_083_),
    .Y(_130_));
 sg13g2_a21oi_1 _328_ (.A1(_076_),
    .A2(net107),
    .Y(_131_),
    .B1(net109));
 sg13g2_a22oi_1 _329_ (.Y(_132_),
    .B1(_130_),
    .B2(_131_),
    .A2(net109),
    .A1(net92));
 sg13g2_a21oi_1 _330_ (.A1(net93),
    .A2(_097_),
    .Y(_133_),
    .B1(net122));
 sg13g2_a22oi_1 _331_ (.Y(_005_),
    .B1(_132_),
    .B2(_133_),
    .A2(net122),
    .A1(_077_));
 sg13g2_nor2_1 _332_ (.A(net31),
    .B(_101_),
    .Y(_134_));
 sg13g2_a22oi_1 _333_ (.Y(_135_),
    .B1(_089_),
    .B2(\ro_buffer_counter_inst.shift_register[14] ),
    .A2(_086_),
    .A1(\ro_buffer_counter_inst.shift_register[6] ));
 sg13g2_a221oi_1 _334_ (.B2(\ro_buffer_counter_inst.shift_register[30] ),
    .C1(net107),
    .B1(_091_),
    .A1(\ro_buffer_counter_inst.shift_register[22] ),
    .Y(_136_),
    .A2(_085_));
 sg13g2_a22oi_1 _335_ (.Y(_137_),
    .B1(_135_),
    .B2(_136_),
    .A2(net107),
    .A1(_078_));
 sg13g2_a221oi_1 _336_ (.B2(\ro_buffer_counter_inst.shift_register[54] ),
    .C1(_137_),
    .B1(_097_),
    .A1(net48),
    .Y(_138_),
    .A2(net109));
 sg13g2_a21oi_1 _337_ (.A1(_101_),
    .A2(net49),
    .Y(_006_),
    .B1(_134_));
 sg13g2_a22oi_1 _338_ (.Y(_139_),
    .B1(_089_),
    .B2(\ro_buffer_counter_inst.shift_register[15] ),
    .A2(_086_),
    .A1(\ro_buffer_counter_inst.shift_register[7] ));
 sg13g2_a22oi_1 _339_ (.Y(_140_),
    .B1(_091_),
    .B2(\ro_buffer_counter_inst.shift_register[31] ),
    .A2(_085_),
    .A1(\ro_buffer_counter_inst.shift_register[23] ));
 sg13g2_nand3_1 _340_ (.B(_139_),
    .C(_140_),
    .A(_083_),
    .Y(_141_));
 sg13g2_nand2b_1 _341_ (.Y(_142_),
    .B(net107),
    .A_N(\ro_buffer_counter_inst.shift_register[39] ));
 sg13g2_a221oi_1 _342_ (.B2(_142_),
    .C1(_097_),
    .B1(_141_),
    .A1(\ro_buffer_counter_inst.shift_register[47] ),
    .Y(_143_),
    .A2(net109));
 sg13g2_o21ai_1 _343_ (.B1(_101_),
    .Y(_144_),
    .A1(\ro_buffer_counter_inst.shift_register[55] ),
    .A2(_098_));
 sg13g2_nand2_1 _344_ (.Y(_145_),
    .A(net33),
    .B(net122));
 sg13g2_o21ai_1 _345_ (.B1(_145_),
    .Y(_007_),
    .A1(_143_),
    .A2(_144_));
 sg13g2_and2_1 _346_ (.A(\ro_buffer_counter_inst.ro2_H.q ),
    .B(net153),
    .X(\ro_buffer_counter_inst.ro2_H.cq4 ));
 sg13g2_and2_1 _347_ (.A(net153),
    .B(\ro_buffer_counter_inst.ro2_G.q ),
    .X(\ro_buffer_counter_inst.ro2_G.cq4 ));
 sg13g2_and2_1 _348_ (.A(net153),
    .B(\ro_buffer_counter_inst.ro2_F.q ),
    .X(\ro_buffer_counter_inst.ro2_F.cq4 ));
 sg13g2_and2_1 _349_ (.A(net153),
    .B(\ro_buffer_counter_inst.ro2_E.q ),
    .X(\ro_buffer_counter_inst.ro2_E.cq4 ));
 sg13g2_and2_1 _350_ (.A(net153),
    .B(\ro_buffer_counter_inst.ro2_D.q ),
    .X(\ro_buffer_counter_inst.ro2_D.cq4 ));
 sg13g2_and2_1 _351_ (.A(net153),
    .B(\ro_buffer_counter_inst.ro2_C.q ),
    .X(\ro_buffer_counter_inst.ro2_C.cq4 ));
 sg13g2_and2_1 _352_ (.A(net153),
    .B(\ro_buffer_counter_inst.ro2_B.q ),
    .X(\ro_buffer_counter_inst.ro2_B.cq4 ));
 sg13g2_and2_1 _353_ (.A(net153),
    .B(\ro_buffer_counter_inst.ro2_A.q ),
    .X(\ro_buffer_counter_inst.ro2_A.cq4 ));
 sg13g2_and2_1 _354_ (.A(\ro_buffer_counter_inst.ro1_H.q ),
    .B(net154),
    .X(\ro_buffer_counter_inst.ro1_H.cq4 ));
 sg13g2_and2_1 _355_ (.A(net154),
    .B(\ro_buffer_counter_inst.ro1_G.q ),
    .X(\ro_buffer_counter_inst.ro1_G.cq4 ));
 sg13g2_and2_1 _356_ (.A(net154),
    .B(\ro_buffer_counter_inst.ro1_F.q ),
    .X(\ro_buffer_counter_inst.ro1_F.cq4 ));
 sg13g2_and2_1 _357_ (.A(net154),
    .B(\ro_buffer_counter_inst.ro1_E.q ),
    .X(\ro_buffer_counter_inst.ro1_E.cq4 ));
 sg13g2_and2_1 _358_ (.A(net154),
    .B(\ro_buffer_counter_inst.ro1_D.q ),
    .X(\ro_buffer_counter_inst.ro1_D.cq4 ));
 sg13g2_and2_1 _359_ (.A(net154),
    .B(\ro_buffer_counter_inst.ro1_C.q ),
    .X(\ro_buffer_counter_inst.ro1_C.cq4 ));
 sg13g2_and2_1 _360_ (.A(net154),
    .B(\ro_buffer_counter_inst.ro1_B.q ),
    .X(\ro_buffer_counter_inst.ro1_B.cq4 ));
 sg13g2_and2_1 _361_ (.A(net154),
    .B(\ro_buffer_counter_inst.ro1_A.q ),
    .X(\ro_buffer_counter_inst.ro1_A.cq4 ));
 sg13g2_nor2_1 _362_ (.A(_084_),
    .B(_087_),
    .Y(_146_));
 sg13g2_xnor2_1 _363_ (.Y(_147_),
    .A(net3),
    .B(net7));
 sg13g2_nand2_1 _364_ (.Y(_148_),
    .A(net6),
    .B(_147_));
 sg13g2_xnor2_1 _365_ (.Y(_149_),
    .A(_146_),
    .B(_148_));
 sg13g2_nor2_1 _366_ (.A(_080_),
    .B(_149_),
    .Y(_150_));
 sg13g2_xor2_1 _367_ (.B(_150_),
    .A(\buffer_out[0] ),
    .X(uo_out[0]));
 sg13g2_o21ai_1 _368_ (.B1(_088_),
    .Y(_151_),
    .A1(net7),
    .A2(_084_));
 sg13g2_nand2b_1 _369_ (.Y(_152_),
    .B(net124),
    .A_N(net6));
 sg13g2_xnor2_1 _370_ (.Y(_153_),
    .A(net124),
    .B(net6));
 sg13g2_xor2_1 _371_ (.B(_153_),
    .A(_087_),
    .X(_154_));
 sg13g2_o21ai_1 _372_ (.B1(\ascon_inst.en ),
    .Y(_155_),
    .A1(_151_),
    .A2(_153_));
 sg13g2_a21oi_1 _373_ (.A1(_151_),
    .A2(_154_),
    .Y(_156_),
    .B1(_155_));
 sg13g2_xor2_1 _374_ (.B(_156_),
    .A(\buffer_out[1] ),
    .X(uo_out[1]));
 sg13g2_nand2_1 _375_ (.Y(_157_),
    .A(\ascon_inst.en ),
    .B(_154_));
 sg13g2_xnor2_1 _376_ (.Y(uo_out[2]),
    .A(\buffer_out[2] ),
    .B(_157_));
 sg13g2_mux2_1 _377_ (.A0(_079_),
    .A1(net124),
    .S(net4),
    .X(_158_));
 sg13g2_xnor2_1 _378_ (.Y(_159_),
    .A(_147_),
    .B(_152_));
 sg13g2_nand2_1 _379_ (.Y(_160_),
    .A(_158_),
    .B(_159_));
 sg13g2_o21ai_1 _380_ (.B1(_160_),
    .Y(_161_),
    .A1(_147_),
    .A2(_158_));
 sg13g2_nor2_1 _381_ (.A(_080_),
    .B(_161_),
    .Y(_162_));
 sg13g2_xor2_1 _382_ (.B(_162_),
    .A(\buffer_out[3] ),
    .X(uo_out[3]));
 sg13g2_o21ai_1 _383_ (.B1(\ascon_inst.en ),
    .Y(_163_),
    .A1(_149_),
    .A2(_159_));
 sg13g2_a21oi_1 _384_ (.A1(_149_),
    .A2(_159_),
    .Y(_164_),
    .B1(_163_));
 sg13g2_xor2_1 _385_ (.B(_164_),
    .A(\buffer_out[4] ),
    .X(uo_out[4]));
 sg13g2_nor2_2 _386_ (.A(net2),
    .B(net1),
    .Y(_165_));
 sg13g2_xnor2_1 _387_ (.Y(_166_),
    .A(\ro_buffer_counter_inst.ro_2_reg_A ),
    .B(\ro_buffer_counter_inst.ro_2_reg_D ));
 sg13g2_xnor2_1 _388_ (.Y(_167_),
    .A(\ro_buffer_counter_inst.ro_2_reg_F ),
    .B(\ro_buffer_counter_inst.ro_1_reg_H ));
 sg13g2_xnor2_1 _389_ (.Y(_168_),
    .A(_166_),
    .B(_167_));
 sg13g2_xnor2_1 _390_ (.Y(_169_),
    .A(\ro_buffer_counter_inst.ro_2_reg_C ),
    .B(_168_));
 sg13g2_xnor2_1 _391_ (.Y(_170_),
    .A(\ro_buffer_counter_inst.ro_1_reg_A ),
    .B(\ro_buffer_counter_inst.ro_2_reg_E ));
 sg13g2_xor2_1 _392_ (.B(\ro_buffer_counter_inst.ro_1_reg_G ),
    .A(\ro_buffer_counter_inst.ro_1_reg_C ),
    .X(_171_));
 sg13g2_xnor2_1 _393_ (.Y(_172_),
    .A(\ro_buffer_counter_inst.ro_2_reg_H ),
    .B(_171_));
 sg13g2_xnor2_1 _394_ (.Y(_173_),
    .A(_170_),
    .B(_172_));
 sg13g2_xor2_1 _395_ (.B(\ro_buffer_counter_inst.ro_2_reg_G ),
    .A(\ro_buffer_counter_inst.ro_1_reg_F ),
    .X(_174_));
 sg13g2_xor2_1 _396_ (.B(\ro_buffer_counter_inst.ro_2_reg_B ),
    .A(\ro_buffer_counter_inst.ro_1_reg_B ),
    .X(_175_));
 sg13g2_xnor2_1 _397_ (.Y(_176_),
    .A(_174_),
    .B(_175_));
 sg13g2_xnor2_1 _398_ (.Y(_177_),
    .A(\ro_buffer_counter_inst.ro_1_reg_D ),
    .B(\ro_buffer_counter_inst.ro_1_reg_E ));
 sg13g2_xnor2_1 _399_ (.Y(_178_),
    .A(_176_),
    .B(_177_));
 sg13g2_xnor2_1 _400_ (.Y(_179_),
    .A(_173_),
    .B(_178_));
 sg13g2_xnor2_1 _401_ (.Y(_180_),
    .A(_169_),
    .B(_179_));
 sg13g2_mux2_1 _402_ (.A0(_180_),
    .A1(net56),
    .S(net120),
    .X(_008_));
 sg13g2_mux2_1 _403_ (.A0(net56),
    .A1(\ro_buffer_counter_inst.shift_register[1] ),
    .S(net120),
    .X(_009_));
 sg13g2_mux2_1 _404_ (.A0(net103),
    .A1(net84),
    .S(net120),
    .X(_010_));
 sg13g2_mux2_1 _405_ (.A0(net84),
    .A1(net68),
    .S(net121),
    .X(_011_));
 sg13g2_mux2_1 _406_ (.A0(net68),
    .A1(net58),
    .S(net119),
    .X(_012_));
 sg13g2_mux2_1 _407_ (.A0(net58),
    .A1(net50),
    .S(net119),
    .X(_013_));
 sg13g2_mux2_1 _408_ (.A0(net50),
    .A1(\ro_buffer_counter_inst.shift_register[6] ),
    .S(net118),
    .X(_014_));
 sg13g2_mux2_1 _409_ (.A0(net59),
    .A1(\ro_buffer_counter_inst.shift_register[7] ),
    .S(net121),
    .X(_015_));
 sg13g2_mux2_1 _410_ (.A0(net72),
    .A1(\ro_buffer_counter_inst.shift_register[8] ),
    .S(net120),
    .X(_016_));
 sg13g2_mux2_1 _411_ (.A0(net90),
    .A1(\ro_buffer_counter_inst.shift_register[9] ),
    .S(net120),
    .X(_017_));
 sg13g2_mux2_1 _412_ (.A0(net150),
    .A1(net62),
    .S(net120),
    .X(_018_));
 sg13g2_mux2_1 _413_ (.A0(net62),
    .A1(\ro_buffer_counter_inst.shift_register[11] ),
    .S(net121),
    .X(_019_));
 sg13g2_mux2_1 _414_ (.A0(net106),
    .A1(net79),
    .S(net121),
    .X(_020_));
 sg13g2_mux2_1 _415_ (.A0(net79),
    .A1(net66),
    .S(net118),
    .X(_021_));
 sg13g2_mux2_1 _416_ (.A0(net66),
    .A1(\ro_buffer_counter_inst.shift_register[14] ),
    .S(net118),
    .X(_022_));
 sg13g2_mux2_1 _417_ (.A0(net98),
    .A1(\ro_buffer_counter_inst.shift_register[15] ),
    .S(net118),
    .X(_023_));
 sg13g2_mux2_1 _418_ (.A0(net145),
    .A1(net95),
    .S(net118),
    .X(_024_));
 sg13g2_mux2_1 _419_ (.A0(net95),
    .A1(net83),
    .S(net118),
    .X(_025_));
 sg13g2_mux2_1 _420_ (.A0(net83),
    .A1(net76),
    .S(net118),
    .X(_026_));
 sg13g2_mux2_1 _421_ (.A0(net76),
    .A1(\ro_buffer_counter_inst.shift_register[19] ),
    .S(net118),
    .X(_027_));
 sg13g2_mux2_1 _422_ (.A0(net104),
    .A1(\ro_buffer_counter_inst.shift_register[20] ),
    .S(net111),
    .X(_028_));
 sg13g2_mux2_1 _423_ (.A0(net149),
    .A1(net89),
    .S(net111),
    .X(_029_));
 sg13g2_mux2_1 _424_ (.A0(net89),
    .A1(net85),
    .S(net110),
    .X(_030_));
 sg13g2_mux2_1 _425_ (.A0(net85),
    .A1(net81),
    .S(net110),
    .X(_031_));
 sg13g2_mux2_1 _426_ (.A0(net81),
    .A1(\ro_buffer_counter_inst.shift_register[24] ),
    .S(net111),
    .X(_032_));
 sg13g2_mux2_1 _427_ (.A0(net151),
    .A1(net144),
    .S(net111),
    .X(_033_));
 sg13g2_mux2_1 _428_ (.A0(net144),
    .A1(net142),
    .S(net111),
    .X(_034_));
 sg13g2_mux2_1 _429_ (.A0(net142),
    .A1(net88),
    .S(net111),
    .X(_035_));
 sg13g2_mux2_1 _430_ (.A0(net88),
    .A1(net86),
    .S(net111),
    .X(_036_));
 sg13g2_mux2_1 _431_ (.A0(net86),
    .A1(net70),
    .S(net111),
    .X(_037_));
 sg13g2_mux2_1 _432_ (.A0(net70),
    .A1(\ro_buffer_counter_inst.shift_register[30] ),
    .S(net110),
    .X(_038_));
 sg13g2_mux2_1 _433_ (.A0(net74),
    .A1(\ro_buffer_counter_inst.shift_register[31] ),
    .S(net110),
    .X(_039_));
 sg13g2_mux2_1 _434_ (.A0(net100),
    .A1(net64),
    .S(net110),
    .X(_040_));
 sg13g2_nor2_1 _435_ (.A(net64),
    .B(net112),
    .Y(_181_));
 sg13g2_a21oi_1 _436_ (.A1(_072_),
    .A2(net112),
    .Y(_041_),
    .B1(_181_));
 sg13g2_nand2_1 _437_ (.Y(_182_),
    .A(net29),
    .B(net112));
 sg13g2_o21ai_1 _438_ (.B1(_182_),
    .Y(_042_),
    .A1(_072_),
    .A2(net112));
 sg13g2_nor2_1 _439_ (.A(net29),
    .B(net119),
    .Y(_183_));
 sg13g2_a21oi_1 _440_ (.A1(_074_),
    .A2(net119),
    .Y(_043_),
    .B1(_183_));
 sg13g2_nor2_1 _441_ (.A(net43),
    .B(net119),
    .Y(_184_));
 sg13g2_a21oi_1 _442_ (.A1(_075_),
    .A2(net112),
    .Y(_044_),
    .B1(_184_));
 sg13g2_nor2_1 _443_ (.A(net53),
    .B(net112),
    .Y(_185_));
 sg13g2_a21oi_1 _444_ (.A1(_076_),
    .A2(net113),
    .Y(_045_),
    .B1(_185_));
 sg13g2_nor2_1 _445_ (.A(net35),
    .B(net110),
    .Y(_186_));
 sg13g2_a21oi_1 _446_ (.A1(_078_),
    .A2(net110),
    .Y(_046_),
    .B1(_186_));
 sg13g2_nand2_1 _447_ (.Y(_187_),
    .A(net25),
    .B(net113));
 sg13g2_o21ai_1 _448_ (.B1(_187_),
    .Y(_047_),
    .A1(_078_),
    .A2(net110));
 sg13g2_mux2_1 _449_ (.A0(net25),
    .A1(net45),
    .S(net113),
    .X(_048_));
 sg13g2_mux2_1 _450_ (.A0(net45),
    .A1(net54),
    .S(net116),
    .X(_049_));
 sg13g2_mux2_1 _451_ (.A0(net54),
    .A1(\ro_buffer_counter_inst.shift_register[42] ),
    .S(net116),
    .X(_050_));
 sg13g2_mux2_1 _452_ (.A0(net96),
    .A1(\ro_buffer_counter_inst.shift_register[43] ),
    .S(net121),
    .X(_051_));
 sg13g2_mux2_1 _453_ (.A0(net152),
    .A1(net101),
    .S(net121),
    .X(_052_));
 sg13g2_mux2_1 _454_ (.A0(net101),
    .A1(net92),
    .S(net115),
    .X(_053_));
 sg13g2_mux2_1 _455_ (.A0(net92),
    .A1(net48),
    .S(net115),
    .X(_054_));
 sg13g2_mux2_1 _456_ (.A0(net48),
    .A1(net52),
    .S(net115),
    .X(_055_));
 sg13g2_mux2_1 _457_ (.A0(net52),
    .A1(net61),
    .S(net115),
    .X(_056_));
 sg13g2_mux2_1 _458_ (.A0(net61),
    .A1(net80),
    .S(net115),
    .X(_057_));
 sg13g2_mux2_1 _459_ (.A0(net80),
    .A1(net37),
    .S(net117),
    .X(_058_));
 sg13g2_mux2_1 _460_ (.A0(net37),
    .A1(net146),
    .S(net114),
    .X(_059_));
 sg13g2_mux2_1 _461_ (.A0(net146),
    .A1(net143),
    .S(net114),
    .X(_060_));
 sg13g2_mux2_1 _462_ (.A0(net143),
    .A1(net93),
    .S(net114),
    .X(_061_));
 sg13g2_mux2_1 _463_ (.A0(net93),
    .A1(\ro_buffer_counter_inst.shift_register[54] ),
    .S(net115),
    .X(_062_));
 sg13g2_mux2_1 _464_ (.A0(net102),
    .A1(net69),
    .S(net115),
    .X(_063_));
 sg13g2_mux2_1 _465_ (.A0(net69),
    .A1(net46),
    .S(net114),
    .X(_064_));
 sg13g2_nor2_1 _466_ (.A(net46),
    .B(net116),
    .Y(_188_));
 sg13g2_a21oi_1 _467_ (.A1(_073_),
    .A2(net116),
    .Y(_065_),
    .B1(_188_));
 sg13g2_nand2_1 _468_ (.Y(_189_),
    .A(net27),
    .B(net116));
 sg13g2_o21ai_1 _469_ (.B1(_189_),
    .Y(_066_),
    .A1(_073_),
    .A2(net116));
 sg13g2_mux2_1 _470_ (.A0(net27),
    .A1(net39),
    .S(net116),
    .X(_067_));
 sg13g2_mux2_1 _471_ (.A0(net39),
    .A1(net41),
    .S(net116),
    .X(_068_));
 sg13g2_nor2_1 _472_ (.A(net41),
    .B(net117),
    .Y(_190_));
 sg13g2_a21oi_1 _473_ (.A1(_077_),
    .A2(net114),
    .Y(_069_),
    .B1(_190_));
 sg13g2_nand2_1 _474_ (.Y(_191_),
    .A(net31),
    .B(net114));
 sg13g2_o21ai_1 _475_ (.B1(_191_),
    .Y(_070_),
    .A1(_077_),
    .A2(net114));
 sg13g2_mux2_1 _476_ (.A0(net31),
    .A1(net33),
    .S(net114),
    .X(_071_));
 sg13g2_inv_1 _477_ (.Y(_072_),
    .A(net147));
 sg13g2_inv_1 _478_ (.Y(_073_),
    .A(net87));
 sg13g2_inv_1 _479_ (.Y(_074_),
    .A(net43));
 sg13g2_inv_1 _480_ (.Y(_075_),
    .A(\ro_buffer_counter_inst.shift_register[36] ));
 sg13g2_inv_1 _481_ (.Y(_076_),
    .A(net35));
 sg13g2_inv_1 _482_ (.Y(_077_),
    .A(net78));
 sg13g2_inv_1 _483_ (.Y(_078_),
    .A(\ro_buffer_counter_inst.shift_register[38] ));
 sg13g2_inv_1 _484_ (.Y(_079_),
    .A(net6));
 sg13g2_inv_1 _485_ (.Y(_080_),
    .A(\ascon_inst.en ));
 sg13g2_nor2_1 _486_ (.A(net3),
    .B(net4),
    .Y(_081_));
 sg13g2_and2_1 _487_ (.A(net123),
    .B(_081_),
    .X(_082_));
 sg13g2_nand2_2 _488_ (.Y(_083_),
    .A(net123),
    .B(_081_));
 sg13g2_nor2b_2 _489_ (.A(net3),
    .B_N(net4),
    .Y(_084_));
 sg13g2_nor2b_2 _490_ (.A(net123),
    .B_N(_084_),
    .Y(_085_));
 sg13g2_nor3_2 _491_ (.A(net3),
    .B(net4),
    .C(net5),
    .Y(_086_));
 sg13g2_nor2b_2 _492_ (.A(net4),
    .B_N(net3),
    .Y(_087_));
 sg13g2_inv_1 _493_ (.Y(_088_),
    .A(_087_));
 sg13g2_nor2b_2 _494_ (.A(net124),
    .B_N(_087_),
    .Y(_089_));
 sg13g2_nand2_1 _495_ (.Y(_090_),
    .A(net3),
    .B(net4));
 sg13g2_dfrbp_1 _496_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net137),
    .D(_008_),
    .Q_N(_255_),
    .Q(\ro_buffer_counter_inst.shift_register[0] ));
 sg13g2_dfrbp_1 _497_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net136),
    .D(net57),
    .Q_N(_254_),
    .Q(\ro_buffer_counter_inst.shift_register[1] ));
 sg13g2_dfrbp_1 _498_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net135),
    .D(_010_),
    .Q_N(_253_),
    .Q(\ro_buffer_counter_inst.shift_register[2] ));
 sg13g2_dfrbp_1 _499_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net135),
    .D(_011_),
    .Q_N(_252_),
    .Q(\ro_buffer_counter_inst.shift_register[3] ));
 sg13g2_dfrbp_1 _500_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net134),
    .D(_012_),
    .Q_N(_251_),
    .Q(\ro_buffer_counter_inst.shift_register[4] ));
 sg13g2_dfrbp_1 _501_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net135),
    .D(_013_),
    .Q_N(_250_),
    .Q(\ro_buffer_counter_inst.shift_register[5] ));
 sg13g2_dfrbp_1 _502_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net134),
    .D(net51),
    .Q_N(_249_),
    .Q(\ro_buffer_counter_inst.shift_register[6] ));
 sg13g2_dfrbp_1 _503_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net134),
    .D(net60),
    .Q_N(_248_),
    .Q(\ro_buffer_counter_inst.shift_register[7] ));
 sg13g2_dfrbp_1 _504_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net136),
    .D(net73),
    .Q_N(_247_),
    .Q(\ro_buffer_counter_inst.shift_register[8] ));
 sg13g2_dfrbp_1 _505_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net137),
    .D(net91),
    .Q_N(_246_),
    .Q(\ro_buffer_counter_inst.shift_register[9] ));
 sg13g2_dfrbp_1 _506_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net136),
    .D(_018_),
    .Q_N(_245_),
    .Q(\ro_buffer_counter_inst.shift_register[10] ));
 sg13g2_dfrbp_1 _507_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net140),
    .D(net63),
    .Q_N(_244_),
    .Q(\ro_buffer_counter_inst.shift_register[11] ));
 sg13g2_dfrbp_1 _508_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net140),
    .D(_020_),
    .Q_N(_243_),
    .Q(\ro_buffer_counter_inst.shift_register[12] ));
 sg13g2_dfrbp_1 _509_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net135),
    .D(_021_),
    .Q_N(_242_),
    .Q(\ro_buffer_counter_inst.shift_register[13] ));
 sg13g2_dfrbp_1 _510_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net134),
    .D(net67),
    .Q_N(_241_),
    .Q(\ro_buffer_counter_inst.shift_register[14] ));
 sg13g2_dfrbp_1 _511_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net134),
    .D(net99),
    .Q_N(_240_),
    .Q(\ro_buffer_counter_inst.shift_register[15] ));
 sg13g2_dfrbp_1 _512_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net134),
    .D(_024_),
    .Q_N(_239_),
    .Q(\ro_buffer_counter_inst.shift_register[16] ));
 sg13g2_dfrbp_1 _513_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net127),
    .D(_025_),
    .Q_N(_238_),
    .Q(\ro_buffer_counter_inst.shift_register[17] ));
 sg13g2_dfrbp_1 _514_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net134),
    .D(_026_),
    .Q_N(_237_),
    .Q(\ro_buffer_counter_inst.shift_register[18] ));
 sg13g2_dfrbp_1 _515_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net134),
    .D(net77),
    .Q_N(_236_),
    .Q(\ro_buffer_counter_inst.shift_register[19] ));
 sg13g2_dfrbp_1 _516_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net127),
    .D(net105),
    .Q_N(_235_),
    .Q(\ro_buffer_counter_inst.shift_register[20] ));
 sg13g2_dfrbp_1 _517_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net127),
    .D(_029_),
    .Q_N(_234_),
    .Q(\ro_buffer_counter_inst.shift_register[21] ));
 sg13g2_dfrbp_1 _518_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net125),
    .D(_030_),
    .Q_N(_233_),
    .Q(\ro_buffer_counter_inst.shift_register[22] ));
 sg13g2_dfrbp_1 _519_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net125),
    .D(_031_),
    .Q_N(_232_),
    .Q(\ro_buffer_counter_inst.shift_register[23] ));
 sg13g2_dfrbp_1 _520_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net127),
    .D(net82),
    .Q_N(_231_),
    .Q(\ro_buffer_counter_inst.shift_register[24] ));
 sg13g2_dfrbp_1 _521_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net127),
    .D(_033_),
    .Q_N(_230_),
    .Q(\ro_buffer_counter_inst.shift_register[25] ));
 sg13g2_dfrbp_1 _522_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net127),
    .D(_034_),
    .Q_N(_229_),
    .Q(\ro_buffer_counter_inst.shift_register[26] ));
 sg13g2_dfrbp_1 _523_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net127),
    .D(_035_),
    .Q_N(_228_),
    .Q(\ro_buffer_counter_inst.shift_register[27] ));
 sg13g2_dfrbp_1 _524_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net127),
    .D(_036_),
    .Q_N(_227_),
    .Q(\ro_buffer_counter_inst.shift_register[28] ));
 sg13g2_dfrbp_1 _525_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net125),
    .D(_037_),
    .Q_N(_226_),
    .Q(\ro_buffer_counter_inst.shift_register[29] ));
 sg13g2_dfrbp_1 _526_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net125),
    .D(net71),
    .Q_N(_225_),
    .Q(\ro_buffer_counter_inst.shift_register[30] ));
 sg13g2_dfrbp_1 _527_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net125),
    .D(net75),
    .Q_N(_224_),
    .Q(\ro_buffer_counter_inst.shift_register[31] ));
 sg13g2_dfrbp_1 _528_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(_040_),
    .Q_N(_223_),
    .Q(\ro_buffer_counter_inst.shift_register[32] ));
 sg13g2_dfrbp_1 _529_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(net65),
    .Q_N(_222_),
    .Q(\ro_buffer_counter_inst.shift_register[33] ));
 sg13g2_dfrbp_1 _530_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net128),
    .D(net30),
    .Q_N(_221_),
    .Q(\ro_buffer_counter_inst.shift_register[34] ));
 sg13g2_dfrbp_1 _531_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net128),
    .D(_043_),
    .Q_N(_220_),
    .Q(\ro_buffer_counter_inst.shift_register[35] ));
 sg13g2_dfrbp_1 _532_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net128),
    .D(net44),
    .Q_N(_219_),
    .Q(\ro_buffer_counter_inst.shift_register[36] ));
 sg13g2_dfrbp_1 _533_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(_045_),
    .Q_N(_218_),
    .Q(\ro_buffer_counter_inst.shift_register[37] ));
 sg13g2_dfrbp_1 _534_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net125),
    .D(net36),
    .Q_N(_217_),
    .Q(\ro_buffer_counter_inst.shift_register[38] ));
 sg13g2_dfrbp_1 _535_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(net26),
    .Q_N(_216_),
    .Q(\ro_buffer_counter_inst.shift_register[39] ));
 sg13g2_dfrbp_1 _536_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(_048_),
    .Q_N(_215_),
    .Q(\ro_buffer_counter_inst.shift_register[40] ));
 sg13g2_dfrbp_1 _537_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net128),
    .D(_049_),
    .Q_N(_214_),
    .Q(\ro_buffer_counter_inst.shift_register[41] ));
 sg13g2_dfrbp_1 _538_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net132),
    .D(net55),
    .Q_N(_213_),
    .Q(\ro_buffer_counter_inst.shift_register[42] ));
 sg13g2_dfrbp_1 _539_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net132),
    .D(net97),
    .Q_N(_212_),
    .Q(\ro_buffer_counter_inst.shift_register[43] ));
 sg13g2_dfrbp_1 _540_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net140),
    .D(_052_),
    .Q_N(_211_),
    .Q(\ro_buffer_counter_inst.shift_register[44] ));
 sg13g2_dfrbp_1 _541_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net125),
    .D(_053_),
    .Q_N(_210_),
    .Q(\ro_buffer_counter_inst.shift_register[45] ));
 sg13g2_dfrbp_1 _542_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net126),
    .D(_054_),
    .Q_N(_209_),
    .Q(\ro_buffer_counter_inst.shift_register[46] ));
 sg13g2_dfrbp_1 _543_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net125),
    .D(_055_),
    .Q_N(_208_),
    .Q(\ro_buffer_counter_inst.shift_register[47] ));
 sg13g2_dfrbp_1 _544_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net131),
    .D(_056_),
    .Q_N(_207_),
    .Q(\ro_buffer_counter_inst.shift_register[48] ));
 sg13g2_dfrbp_1 _545_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net131),
    .D(_057_),
    .Q_N(_206_),
    .Q(\ro_buffer_counter_inst.shift_register[49] ));
 sg13g2_dfrbp_1 _546_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net132),
    .D(_058_),
    .Q_N(_205_),
    .Q(\ro_buffer_counter_inst.shift_register[50] ));
 sg13g2_dfrbp_1 _547_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net130),
    .D(_059_),
    .Q_N(_204_),
    .Q(\ro_buffer_counter_inst.shift_register[51] ));
 sg13g2_dfrbp_1 _548_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net130),
    .D(_060_),
    .Q_N(_203_),
    .Q(\ro_buffer_counter_inst.shift_register[52] ));
 sg13g2_dfrbp_1 _549_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net131),
    .D(_061_),
    .Q_N(_202_),
    .Q(\ro_buffer_counter_inst.shift_register[53] ));
 sg13g2_dfrbp_1 _550_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net131),
    .D(net94),
    .Q_N(_201_),
    .Q(\ro_buffer_counter_inst.shift_register[54] ));
 sg13g2_dfrbp_1 _551_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net131),
    .D(_063_),
    .Q_N(_200_),
    .Q(\ro_buffer_counter_inst.shift_register[55] ));
 sg13g2_dfrbp_1 _552_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net131),
    .D(_064_),
    .Q_N(_199_),
    .Q(\ro_buffer_counter_inst.shift_register[56] ));
 sg13g2_dfrbp_1 _553_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net132),
    .D(_065_),
    .Q_N(_198_),
    .Q(\ro_buffer_counter_inst.shift_register[57] ));
 sg13g2_dfrbp_1 _554_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net132),
    .D(net28),
    .Q_N(_197_),
    .Q(\ro_buffer_counter_inst.shift_register[58] ));
 sg13g2_dfrbp_1 _555_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net133),
    .D(_067_),
    .Q_N(_196_),
    .Q(\ro_buffer_counter_inst.shift_register[59] ));
 sg13g2_dfrbp_1 _556_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net130),
    .D(_068_),
    .Q_N(_195_),
    .Q(\ro_buffer_counter_inst.shift_register[60] ));
 sg13g2_dfrbp_1 _557_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net130),
    .D(_069_),
    .Q_N(_194_),
    .Q(\ro_buffer_counter_inst.shift_register[61] ));
 sg13g2_dfrbp_1 _558_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net130),
    .D(net32),
    .Q_N(_193_),
    .Q(\ro_buffer_counter_inst.shift_register[62] ));
 sg13g2_dfrbp_1 _559_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net130),
    .D(_071_),
    .Q_N(_256_),
    .Q(\ro_buffer_counter_inst.shift_register[63] ));
 sg13g2_dfrbp_1 _560_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net139),
    .D(net2),
    .Q_N(_257_),
    .Q(\ro_buffer_counter_inst.ro2_A.en ));
 sg13g2_dfrbp_1 _561_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net139),
    .D(net1),
    .Q_N(_258_),
    .Q(\ro_buffer_counter_inst.ro1_A.en ));
 sg13g2_dfrbp_1 _562_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net138),
    .D(\ro_buffer_counter_inst.ro2_G.cq4 ),
    .Q_N(_259_),
    .Q(\ro_buffer_counter_inst.ro_2_reg_G ));
 sg13g2_dfrbp_1 _563_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net139),
    .D(\ro_buffer_counter_inst.ro1_D.cq4 ),
    .Q_N(_260_),
    .Q(\ro_buffer_counter_inst.ro_1_reg_D ));
 sg13g2_dfrbp_1 _564_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net136),
    .D(\ro_buffer_counter_inst.ro2_F.cq4 ),
    .Q_N(_261_),
    .Q(\ro_buffer_counter_inst.ro_2_reg_F ));
 sg13g2_dfrbp_1 _565_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net138),
    .D(\ro_buffer_counter_inst.ro1_A.cq4 ),
    .Q_N(_262_),
    .Q(\ro_buffer_counter_inst.ro_1_reg_A ));
 sg13g2_dfrbp_1 _566_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net138),
    .D(\ro_buffer_counter_inst.ro2_E.cq4 ),
    .Q_N(_263_),
    .Q(\ro_buffer_counter_inst.ro_2_reg_E ));
 sg13g2_dfrbp_1 _567_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net139),
    .D(\ro_buffer_counter_inst.ro1_E.cq4 ),
    .Q_N(_264_),
    .Q(\ro_buffer_counter_inst.ro_1_reg_E ));
 sg13g2_dfrbp_1 _568_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net136),
    .D(\ro_buffer_counter_inst.ro2_D.cq4 ),
    .Q_N(_265_),
    .Q(\ro_buffer_counter_inst.ro_2_reg_D ));
 sg13g2_dfrbp_1 _569_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net138),
    .D(\ro_buffer_counter_inst.ro1_C.cq4 ),
    .Q_N(_266_),
    .Q(\ro_buffer_counter_inst.ro_1_reg_C ));
 sg13g2_dfrbp_1 _570_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net136),
    .D(\ro_buffer_counter_inst.ro2_C.cq4 ),
    .Q_N(_267_),
    .Q(\ro_buffer_counter_inst.ro_2_reg_C ));
 sg13g2_dfrbp_1 _571_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net138),
    .D(\ro_buffer_counter_inst.ro1_F.cq4 ),
    .Q_N(_268_),
    .Q(\ro_buffer_counter_inst.ro_1_reg_F ));
 sg13g2_dfrbp_1 _572_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net139),
    .D(\ro_buffer_counter_inst.ro2_B.cq4 ),
    .Q_N(_269_),
    .Q(\ro_buffer_counter_inst.ro_2_reg_B ));
 sg13g2_dfrbp_1 _573_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net138),
    .D(\ro_buffer_counter_inst.ro2_H.cq4 ),
    .Q_N(_270_),
    .Q(\ro_buffer_counter_inst.ro_2_reg_H ));
 sg13g2_dfrbp_1 _574_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net136),
    .D(\ro_buffer_counter_inst.ro2_A.cq4 ),
    .Q_N(_271_),
    .Q(\ro_buffer_counter_inst.ro_2_reg_A ));
 sg13g2_dfrbp_1 _575_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net138),
    .D(\ro_buffer_counter_inst.ro1_G.cq4 ),
    .Q_N(_272_),
    .Q(\ro_buffer_counter_inst.ro_1_reg_G ));
 sg13g2_dfrbp_1 _576_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net138),
    .D(\ro_buffer_counter_inst.ro1_B.cq4 ),
    .Q_N(_273_),
    .Q(\ro_buffer_counter_inst.ro_1_reg_B ));
 sg13g2_dfrbp_1 _577_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net133),
    .D(net47),
    .Q_N(_274_),
    .Q(\buffer_out[0] ));
 sg13g2_dfrbp_1 _578_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net133),
    .D(_001_),
    .Q_N(_275_),
    .Q(\buffer_out[1] ));
 sg13g2_dfrbp_1 _579_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net132),
    .D(net38),
    .Q_N(_276_),
    .Q(\buffer_out[2] ));
 sg13g2_dfrbp_1 _580_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net132),
    .D(net40),
    .Q_N(_277_),
    .Q(\buffer_out[3] ));
 sg13g2_dfrbp_1 _581_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net132),
    .D(net42),
    .Q_N(_278_),
    .Q(\buffer_out[4] ));
 sg13g2_dfrbp_1 _582_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net131),
    .D(_005_),
    .Q_N(_279_),
    .Q(\buffer_out[5] ));
 sg13g2_dfrbp_1 _583_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net130),
    .D(_006_),
    .Q_N(_280_),
    .Q(\buffer_out[6] ));
 sg13g2_dfrbp_1 _584_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net130),
    .D(net34),
    .Q_N(_281_),
    .Q(\buffer_out[7] ));
 sg13g2_dfrbp_1 _585_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net136),
    .D(\ro_buffer_counter_inst.ro1_H.cq4 ),
    .Q_N(_282_),
    .Q(\ro_buffer_counter_inst.ro_1_reg_H ));
 sg13g2_dfrbp_1 _586_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net140),
    .D(net8),
    .Q_N(_192_),
    .Q(\ascon_inst.en ));
 sg13g2_tielo tt_um_roy1707018_10 (.L_LO(net10));
 sg13g2_tielo tt_um_roy1707018_11 (.L_LO(net11));
 sg13g2_tielo tt_um_roy1707018_12 (.L_LO(net12));
 sg13g2_tielo tt_um_roy1707018_13 (.L_LO(net13));
 sg13g2_tielo tt_um_roy1707018_14 (.L_LO(net14));
 sg13g2_tielo tt_um_roy1707018_15 (.L_LO(net15));
 sg13g2_tielo tt_um_roy1707018_16 (.L_LO(net16));
 sg13g2_tielo tt_um_roy1707018_17 (.L_LO(net17));
 sg13g2_tielo tt_um_roy1707018_18 (.L_LO(net18));
 sg13g2_tielo tt_um_roy1707018_19 (.L_LO(net19));
 sg13g2_tielo tt_um_roy1707018_20 (.L_LO(net20));
 sg13g2_tielo tt_um_roy1707018_21 (.L_LO(net21));
 sg13g2_tielo tt_um_roy1707018_22 (.L_LO(net22));
 sg13g2_tielo tt_um_roy1707018_23 (.L_LO(net23));
 sg13g2_tielo tt_um_roy1707018_24 (.L_LO(net24));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _603_ (.A(\ro_buffer_counter_inst.ro1_A.q ),
    .X(\ro_buffer_counter_inst.ro1_A.q4 ));
 sg13g2_buf_1 _604_ (.A(\ro_buffer_counter_inst.ro1_B.q ),
    .X(\ro_buffer_counter_inst.ro1_B.q4 ));
 sg13g2_buf_1 _605_ (.A(\ro_buffer_counter_inst.ro1_C.q ),
    .X(\ro_buffer_counter_inst.ro1_C.q4 ));
 sg13g2_buf_1 _606_ (.A(\ro_buffer_counter_inst.ro1_D.q ),
    .X(\ro_buffer_counter_inst.ro1_D.q4 ));
 sg13g2_buf_1 _607_ (.A(\ro_buffer_counter_inst.ro1_E.q ),
    .X(\ro_buffer_counter_inst.ro1_E.q4 ));
 sg13g2_buf_1 _608_ (.A(\ro_buffer_counter_inst.ro1_F.q ),
    .X(\ro_buffer_counter_inst.ro1_F.q4 ));
 sg13g2_buf_1 _609_ (.A(\ro_buffer_counter_inst.ro1_G.q ),
    .X(\ro_buffer_counter_inst.ro1_G.q4 ));
 sg13g2_buf_1 _610_ (.A(\ro_buffer_counter_inst.ro1_H.q ),
    .X(\ro_buffer_counter_inst.ro1_H.q4 ));
 sg13g2_buf_1 _611_ (.A(\ro_buffer_counter_inst.ro2_A.q ),
    .X(\ro_buffer_counter_inst.ro2_A.q4 ));
 sg13g2_buf_1 _612_ (.A(\ro_buffer_counter_inst.ro2_B.q ),
    .X(\ro_buffer_counter_inst.ro2_B.q4 ));
 sg13g2_buf_1 _613_ (.A(\ro_buffer_counter_inst.ro2_C.q ),
    .X(\ro_buffer_counter_inst.ro2_C.q4 ));
 sg13g2_buf_1 _614_ (.A(\ro_buffer_counter_inst.ro2_D.q ),
    .X(\ro_buffer_counter_inst.ro2_D.q4 ));
 sg13g2_buf_1 _615_ (.A(\ro_buffer_counter_inst.ro2_E.q ),
    .X(\ro_buffer_counter_inst.ro2_E.q4 ));
 sg13g2_buf_1 _616_ (.A(\ro_buffer_counter_inst.ro2_F.q ),
    .X(\ro_buffer_counter_inst.ro2_F.q4 ));
 sg13g2_buf_1 _617_ (.A(\ro_buffer_counter_inst.ro2_G.q ),
    .X(\ro_buffer_counter_inst.ro2_G.q4 ));
 sg13g2_buf_1 _618_ (.A(\ro_buffer_counter_inst.ro2_H.q ),
    .X(\ro_buffer_counter_inst.ro2_H.q4 ));
 sg13g2_buf_1 _619_ (.A(\buffer_out[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _620_ (.A(\buffer_out[6] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _621_ (.A(\buffer_out[7] ),
    .X(uo_out[7]));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_A.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro1_A.q0 ),
    .A(\ro_buffer_counter_inst.ro1_A.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_A.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro1_A.q1 ),
    .A(\ro_buffer_counter_inst.ro1_A.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_A.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro1_A.q2 ),
    .A(\ro_buffer_counter_inst.ro1_A.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_A.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro1_A.q3 ),
    .A(\ro_buffer_counter_inst.ro1_A.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_A.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro1_A.q ),
    .A(\ro_buffer_counter_inst.ro1_A.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_B.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro1_B.q0 ),
    .A(\ro_buffer_counter_inst.ro1_B.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_B.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro1_B.q1 ),
    .A(\ro_buffer_counter_inst.ro1_B.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_B.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro1_B.q2 ),
    .A(\ro_buffer_counter_inst.ro1_B.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_B.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro1_B.q3 ),
    .A(\ro_buffer_counter_inst.ro1_B.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_B.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro1_B.q ),
    .A(\ro_buffer_counter_inst.ro1_B.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_C.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro1_C.q0 ),
    .A(\ro_buffer_counter_inst.ro1_C.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_C.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro1_C.q1 ),
    .A(\ro_buffer_counter_inst.ro1_C.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_C.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro1_C.q2 ),
    .A(\ro_buffer_counter_inst.ro1_C.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_C.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro1_C.q3 ),
    .A(\ro_buffer_counter_inst.ro1_C.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_C.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro1_C.q ),
    .A(\ro_buffer_counter_inst.ro1_C.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_D.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro1_D.q0 ),
    .A(\ro_buffer_counter_inst.ro1_D.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_D.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro1_D.q1 ),
    .A(\ro_buffer_counter_inst.ro1_D.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_D.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro1_D.q2 ),
    .A(\ro_buffer_counter_inst.ro1_D.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_D.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro1_D.q3 ),
    .A(\ro_buffer_counter_inst.ro1_D.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_D.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro1_D.q ),
    .A(\ro_buffer_counter_inst.ro1_D.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_E.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro1_E.q0 ),
    .A(\ro_buffer_counter_inst.ro1_E.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_E.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro1_E.q1 ),
    .A(\ro_buffer_counter_inst.ro1_E.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_E.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro1_E.q2 ),
    .A(\ro_buffer_counter_inst.ro1_E.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_E.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro1_E.q3 ),
    .A(\ro_buffer_counter_inst.ro1_E.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_E.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro1_E.q ),
    .A(\ro_buffer_counter_inst.ro1_E.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_F.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro1_F.q0 ),
    .A(\ro_buffer_counter_inst.ro1_F.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_F.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro1_F.q1 ),
    .A(\ro_buffer_counter_inst.ro1_F.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_F.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro1_F.q2 ),
    .A(\ro_buffer_counter_inst.ro1_F.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_F.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro1_F.q3 ),
    .A(\ro_buffer_counter_inst.ro1_F.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_F.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro1_F.q ),
    .A(\ro_buffer_counter_inst.ro1_F.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_G.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro1_G.q0 ),
    .A(\ro_buffer_counter_inst.ro1_G.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_G.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro1_G.q1 ),
    .A(\ro_buffer_counter_inst.ro1_G.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_G.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro1_G.q2 ),
    .A(\ro_buffer_counter_inst.ro1_G.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_G.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro1_G.q3 ),
    .A(\ro_buffer_counter_inst.ro1_G.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_G.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro1_G.q ),
    .A(\ro_buffer_counter_inst.ro1_G.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_H.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro1_H.q0 ),
    .A(\ro_buffer_counter_inst.ro1_H.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_H.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro1_H.q1 ),
    .A(\ro_buffer_counter_inst.ro1_H.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_H.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro1_H.q2 ),
    .A(\ro_buffer_counter_inst.ro1_H.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_H.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro1_H.q3 ),
    .A(\ro_buffer_counter_inst.ro1_H.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro1_H.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro1_H.q ),
    .A(\ro_buffer_counter_inst.ro1_H.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_A.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro2_A.q0 ),
    .A(\ro_buffer_counter_inst.ro2_A.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_A.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro2_A.q1 ),
    .A(\ro_buffer_counter_inst.ro2_A.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_A.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro2_A.q2 ),
    .A(\ro_buffer_counter_inst.ro2_A.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_A.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro2_A.q3 ),
    .A(\ro_buffer_counter_inst.ro2_A.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_A.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro2_A.q ),
    .A(\ro_buffer_counter_inst.ro2_A.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_B.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro2_B.q0 ),
    .A(\ro_buffer_counter_inst.ro2_B.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_B.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro2_B.q1 ),
    .A(\ro_buffer_counter_inst.ro2_B.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_B.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro2_B.q2 ),
    .A(\ro_buffer_counter_inst.ro2_B.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_B.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro2_B.q3 ),
    .A(\ro_buffer_counter_inst.ro2_B.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_B.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro2_B.q ),
    .A(\ro_buffer_counter_inst.ro2_B.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_C.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro2_C.q0 ),
    .A(\ro_buffer_counter_inst.ro2_C.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_C.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro2_C.q1 ),
    .A(\ro_buffer_counter_inst.ro2_C.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_C.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro2_C.q2 ),
    .A(\ro_buffer_counter_inst.ro2_C.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_C.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro2_C.q3 ),
    .A(\ro_buffer_counter_inst.ro2_C.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_C.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro2_C.q ),
    .A(\ro_buffer_counter_inst.ro2_C.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_D.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro2_D.q0 ),
    .A(\ro_buffer_counter_inst.ro2_D.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_D.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro2_D.q1 ),
    .A(\ro_buffer_counter_inst.ro2_D.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_D.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro2_D.q2 ),
    .A(\ro_buffer_counter_inst.ro2_D.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_D.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro2_D.q3 ),
    .A(\ro_buffer_counter_inst.ro2_D.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_D.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro2_D.q ),
    .A(\ro_buffer_counter_inst.ro2_D.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_E.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro2_E.q0 ),
    .A(\ro_buffer_counter_inst.ro2_E.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_E.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro2_E.q1 ),
    .A(\ro_buffer_counter_inst.ro2_E.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_E.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro2_E.q2 ),
    .A(\ro_buffer_counter_inst.ro2_E.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_E.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro2_E.q3 ),
    .A(\ro_buffer_counter_inst.ro2_E.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_E.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro2_E.q ),
    .A(\ro_buffer_counter_inst.ro2_E.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_F.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro2_F.q0 ),
    .A(\ro_buffer_counter_inst.ro2_F.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_F.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro2_F.q1 ),
    .A(\ro_buffer_counter_inst.ro2_F.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_F.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro2_F.q2 ),
    .A(\ro_buffer_counter_inst.ro2_F.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_F.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro2_F.q3 ),
    .A(\ro_buffer_counter_inst.ro2_F.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_F.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro2_F.q ),
    .A(\ro_buffer_counter_inst.ro2_F.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_G.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro2_G.q0 ),
    .A(\ro_buffer_counter_inst.ro2_G.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_G.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro2_G.q1 ),
    .A(\ro_buffer_counter_inst.ro2_G.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_G.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro2_G.q2 ),
    .A(\ro_buffer_counter_inst.ro2_G.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_G.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro2_G.q3 ),
    .A(\ro_buffer_counter_inst.ro2_G.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_G.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro2_G.q ),
    .A(\ro_buffer_counter_inst.ro2_G.q3 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_H.cinv1/_0_  (.Y(\ro_buffer_counter_inst.ro2_H.q0 ),
    .A(\ro_buffer_counter_inst.ro2_H.cq4 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_H.cinv2/_0_  (.Y(\ro_buffer_counter_inst.ro2_H.q1 ),
    .A(\ro_buffer_counter_inst.ro2_H.q0 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_H.cinv3/_0_  (.Y(\ro_buffer_counter_inst.ro2_H.q2 ),
    .A(\ro_buffer_counter_inst.ro2_H.q1 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_H.cinv4/_0_  (.Y(\ro_buffer_counter_inst.ro2_H.q3 ),
    .A(\ro_buffer_counter_inst.ro2_H.q2 ));
 sg13g2_inv_1 \ro_buffer_counter_inst.ro2_H.cinv5/_0_  (.Y(\ro_buffer_counter_inst.ro2_H.q ),
    .A(\ro_buffer_counter_inst.ro2_H.q3 ));
 sg13g2_buf_2 fanout107 (.A(_082_),
    .X(net107));
 sg13g2_buf_1 fanout108 (.A(_082_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_095_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(net113),
    .X(net110));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(net113));
 sg13g2_buf_2 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_165_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(net115),
    .X(net114));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(net117));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(net117));
 sg13g2_buf_1 fanout117 (.A(_165_),
    .X(net117));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(net120));
 sg13g2_buf_2 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(net121));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(_165_));
 sg13g2_buf_2 fanout122 (.A(_100_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(net124),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(net5),
    .X(net124));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(net129));
 sg13g2_buf_2 fanout126 (.A(net129),
    .X(net126));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(net129));
 sg13g2_buf_2 fanout128 (.A(net129),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(net141),
    .X(net129));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(net131));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(net133));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(net133));
 sg13g2_buf_2 fanout133 (.A(net141),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net137));
 sg13g2_buf_2 fanout135 (.A(net137),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net137));
 sg13g2_buf_2 fanout137 (.A(net141),
    .X(net137));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net140));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(rst_n),
    .X(net141));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[3]));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_roy1707018_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ro_buffer_counter_inst.shift_register[39] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold2 (.A(_047_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ro_buffer_counter_inst.shift_register[58] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold4 (.A(_066_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ro_buffer_counter_inst.shift_register[34] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold6 (.A(_042_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold7 (.A(\ro_buffer_counter_inst.shift_register[62] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold8 (.A(_070_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ro_buffer_counter_inst.shift_register[63] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold10 (.A(_007_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold11 (.A(\ro_buffer_counter_inst.shift_register[37] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold12 (.A(_046_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ro_buffer_counter_inst.shift_register[50] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold14 (.A(_002_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold15 (.A(\ro_buffer_counter_inst.shift_register[59] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold16 (.A(_003_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ro_buffer_counter_inst.shift_register[60] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold18 (.A(_004_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ro_buffer_counter_inst.shift_register[35] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold20 (.A(_044_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold21 (.A(\ro_buffer_counter_inst.shift_register[40] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ro_buffer_counter_inst.shift_register[56] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold23 (.A(_000_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ro_buffer_counter_inst.shift_register[46] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold25 (.A(_138_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ro_buffer_counter_inst.shift_register[5] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold27 (.A(_014_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold28 (.A(\ro_buffer_counter_inst.shift_register[47] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ro_buffer_counter_inst.shift_register[36] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ro_buffer_counter_inst.shift_register[41] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold31 (.A(_050_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ro_buffer_counter_inst.shift_register[0] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold33 (.A(_009_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ro_buffer_counter_inst.shift_register[4] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold35 (.A(\ro_buffer_counter_inst.shift_register[6] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold36 (.A(_015_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold37 (.A(\ro_buffer_counter_inst.shift_register[48] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold38 (.A(\ro_buffer_counter_inst.shift_register[10] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold39 (.A(_019_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold40 (.A(\ro_buffer_counter_inst.shift_register[32] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold41 (.A(_041_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold42 (.A(\ro_buffer_counter_inst.shift_register[13] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold43 (.A(_022_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold44 (.A(\ro_buffer_counter_inst.shift_register[3] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold45 (.A(\ro_buffer_counter_inst.shift_register[55] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold46 (.A(\ro_buffer_counter_inst.shift_register[29] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold47 (.A(_038_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ro_buffer_counter_inst.shift_register[7] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold49 (.A(_016_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ro_buffer_counter_inst.shift_register[30] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold51 (.A(_039_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ro_buffer_counter_inst.shift_register[18] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold53 (.A(_027_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ro_buffer_counter_inst.shift_register[61] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold55 (.A(\ro_buffer_counter_inst.shift_register[12] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold56 (.A(\ro_buffer_counter_inst.shift_register[49] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ro_buffer_counter_inst.shift_register[23] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold58 (.A(_032_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold59 (.A(\ro_buffer_counter_inst.shift_register[17] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold60 (.A(\ro_buffer_counter_inst.shift_register[2] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold61 (.A(\ro_buffer_counter_inst.shift_register[22] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ro_buffer_counter_inst.shift_register[28] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold63 (.A(\ro_buffer_counter_inst.shift_register[57] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ro_buffer_counter_inst.shift_register[27] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold65 (.A(\ro_buffer_counter_inst.shift_register[21] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold66 (.A(\ro_buffer_counter_inst.shift_register[8] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold67 (.A(_017_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold68 (.A(\ro_buffer_counter_inst.shift_register[45] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ro_buffer_counter_inst.shift_register[53] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold70 (.A(_062_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ro_buffer_counter_inst.shift_register[16] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold72 (.A(\ro_buffer_counter_inst.shift_register[42] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold73 (.A(_051_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold74 (.A(\ro_buffer_counter_inst.shift_register[14] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold75 (.A(_023_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold76 (.A(\ro_buffer_counter_inst.shift_register[31] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ro_buffer_counter_inst.shift_register[44] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ro_buffer_counter_inst.shift_register[54] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ro_buffer_counter_inst.shift_register[1] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold80 (.A(\ro_buffer_counter_inst.shift_register[19] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold81 (.A(_028_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ro_buffer_counter_inst.shift_register[11] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold83 (.A(\ro_buffer_counter_inst.shift_register[26] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold84 (.A(\ro_buffer_counter_inst.shift_register[52] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold85 (.A(\ro_buffer_counter_inst.shift_register[25] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold86 (.A(\ro_buffer_counter_inst.shift_register[15] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold87 (.A(\ro_buffer_counter_inst.shift_register[51] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold88 (.A(\ro_buffer_counter_inst.shift_register[33] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold89 (.A(_106_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold90 (.A(\ro_buffer_counter_inst.shift_register[20] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ro_buffer_counter_inst.shift_register[9] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold92 (.A(\ro_buffer_counter_inst.shift_register[24] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold93 (.A(\ro_buffer_counter_inst.shift_register[43] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold94 (.A(\ro_buffer_counter_inst.ro2_A.en ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold95 (.A(\ro_buffer_counter_inst.ro1_A.en ),
    .X(net154));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_decap_8 FILLER_18_166 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_decap_8 FILLER_18_180 ();
 sg13g2_decap_4 FILLER_18_187 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_4 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_130 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_decap_4 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_decap_4 FILLER_19_246 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_decap_4 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_4 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_114 ();
 sg13g2_fill_2 FILLER_20_145 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_4 FILLER_21_77 ();
 sg13g2_fill_1 FILLER_21_81 ();
 sg13g2_fill_2 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_110 ();
 sg13g2_decap_4 FILLER_21_137 ();
 sg13g2_fill_2 FILLER_21_141 ();
 sg13g2_decap_4 FILLER_21_169 ();
 sg13g2_fill_1 FILLER_21_173 ();
 sg13g2_decap_4 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_decap_8 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_decap_4 FILLER_21_278 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_112 ();
 sg13g2_decap_4 FILLER_22_142 ();
 sg13g2_fill_2 FILLER_22_146 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_190 ();
 sg13g2_decap_8 FILLER_22_237 ();
 sg13g2_decap_4 FILLER_22_280 ();
 sg13g2_fill_2 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_96 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_136 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_decap_4 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_217 ();
 sg13g2_fill_2 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_229 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_4 FILLER_24_70 ();
 sg13g2_fill_1 FILLER_24_129 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_decap_4 FILLER_24_227 ();
 sg13g2_decap_4 FILLER_24_251 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_65 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_135 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_decap_4 FILLER_25_316 ();
 sg13g2_fill_2 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_110 ();
 sg13g2_fill_2 FILLER_26_138 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_67 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_142 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_229 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_2 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_2 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_235 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_fill_2 FILLER_28_341 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_fill_2 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_210 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_309 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_fill_2 FILLER_29_391 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_89 ();
 sg13g2_fill_1 FILLER_30_96 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_decap_4 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_decap_8 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_decap_4 FILLER_31_264 ();
 sg13g2_fill_1 FILLER_31_268 ();
 sg13g2_decap_4 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_345 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_decap_4 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_369 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_4 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_157 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_fill_2 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_294 ();
 sg13g2_decap_4 FILLER_32_308 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_345 ();
 sg13g2_decap_4 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_60 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_320 ();
 sg13g2_decap_4 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_decap_8 FILLER_33_369 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_383 ();
 sg13g2_decap_4 FILLER_33_390 ();
 sg13g2_fill_2 FILLER_33_394 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_4 FILLER_34_340 ();
 sg13g2_decap_4 FILLER_34_347 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_2 FILLER_34_394 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_fill_2 FILLER_35_56 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_fill_2 FILLER_35_107 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_decap_4 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_207 ();
 sg13g2_fill_1 FILLER_35_248 ();
 sg13g2_decap_8 FILLER_35_275 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_decap_4 FILLER_35_296 ();
 sg13g2_decap_4 FILLER_35_335 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_67 ();
 sg13g2_fill_2 FILLER_36_82 ();
 sg13g2_fill_1 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_decap_8 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_decap_4 FILLER_36_300 ();
 sg13g2_decap_8 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_fill_2 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_140 ();
 sg13g2_fill_1 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_fill_2 FILLER_37_180 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_decap_4 FILLER_37_252 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_2 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_395 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_fill_1 FILLER_38_186 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_decap_8 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

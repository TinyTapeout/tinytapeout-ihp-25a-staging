module tt_um_dlmiles_poc_fskmodem_hdlctrx (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire clknet_leaf_0_clk;
 wire \latched[0] ;
 wire \latched[12] ;
 wire \latched[14] ;
 wire \latched[15] ;
 wire \latched[1] ;
 wire \latched[3] ;
 wire \latched[5] ;
 wire \latched[6] ;
 wire \latched[7] ;
 wire \modem.analog_rxDac8[7] ;
 wire \modem.cfgAddrDirection ;
 wire \modem.cfgRxClockDirection ;
 wire \modem.cfgUpDownSource ;
 wire \modem.control._zz_ ;
 wire \modem.control._zz__1 ;
 wire \modem.control._zz__1_regNext ;
 wire \modem.control._zz__2 ;
 wire \modem.control._zz__2_regNext ;
 wire \modem.control._zz__3 ;
 wire \modem.control._zz__3_regNext ;
 wire \modem.control._zz__regNext ;
 wire \modem.control._zz_txClockInternalFallStb ;
 wire \modem.control._zz_txClockInternalFallStb_regNext ;
 wire \modem.control.io_rxClock ;
 wire \modem.control.io_txClockStb ;
 wire \modem.control.io_upDownOut ;
 wire \modem.control.phase[0] ;
 wire \modem.control.rst_n ;
 wire \modem.control.rxAddr[0] ;
 wire \modem.control.rxAddr[10] ;
 wire \modem.control.rxAddr[11] ;
 wire \modem.control.rxAddr[1] ;
 wire \modem.control.rxAddr[4] ;
 wire \modem.control.rxAddr[5] ;
 wire \modem.control.rxAddr[6] ;
 wire \modem.control.rxAddr[7] ;
 wire \modem.control.rxAddr[8] ;
 wire \modem.control.rxAddr[9] ;
 wire \modem.control.rxRcrDacTmp[3] ;
 wire \modem.control.scrambler_1.io_dataIn ;
 wire \modem.control.scrambler_1.io_vecOut[0] ;
 wire \modem.control.scrambler_1.io_vecOut[10] ;
 wire \modem.control.scrambler_1.io_vecOut[11] ;
 wire \modem.control.scrambler_1.io_vecOut[12] ;
 wire \modem.control.scrambler_1.io_vecOut[13] ;
 wire \modem.control.scrambler_1.io_vecOut[14] ;
 wire \modem.control.scrambler_1.io_vecOut[15] ;
 wire \modem.control.scrambler_1.io_vecOut[16] ;
 wire \modem.control.scrambler_1.io_vecOut[1] ;
 wire \modem.control.scrambler_1.io_vecOut[2] ;
 wire \modem.control.scrambler_1.io_vecOut[3] ;
 wire \modem.control.scrambler_1.io_vecOut[4] ;
 wire \modem.control.scrambler_1.io_vecOut[5] ;
 wire \modem.control.scrambler_1.io_vecOut[6] ;
 wire \modem.control.scrambler_1.io_vecOut[7] ;
 wire \modem.control.scrambler_1.io_vecOut[8] ;
 wire \modem.control.scrambler_1.io_vecOut[9] ;
 wire \modem.control.tablePhase[3] ;
 wire \modem.control.zeroCrossDet_0 ;
 wire \modem.control.zeroCrossDet_1 ;
 wire \modem.control.zeroCrossDet_2 ;
 wire \modem.control.zeroCrossDet_3 ;
 wire \modem.control.zeroCrossDet_4 ;
 wire \modem.control.zeroCrossDet_5 ;
 wire \modem.control.zeroCrossDet_6 ;
 wire \modem.control.zeroCrossDet_7 ;
 wire \modem.dcd ;
 wire \modem.dcdHistory_1 ;
 wire \modem.dcdHistory_2 ;
 wire \modem.dcdHistory_3 ;
 wire \modem.dcdHistory_4 ;
 wire \modem.dcdHistory_5 ;
 wire \modem.dcdHistory_6 ;
 wire \modem.dcdHistory_7 ;
 wire \modem.uart.descram.io_dataIn ;
 wire \modem.uart.io_isSending ;
 wire \modem.uart.io_uartCtsOut ;
 wire \modem.uart.io_uartTxOut ;
 wire \modem.uart.rxFifo.count[0] ;
 wire \modem.uart.rxFifo.count[1] ;
 wire \modem.uart.rxFifo.count[2] ;
 wire \modem.uart.rxFifo.count[3] ;
 wire \modem.uart.rxFifo.fifo_0[0] ;
 wire \modem.uart.rxFifo.fifo_0[1] ;
 wire \modem.uart.rxFifo.fifo_0[2] ;
 wire \modem.uart.rxFifo.fifo_0[3] ;
 wire \modem.uart.rxFifo.fifo_0[4] ;
 wire \modem.uart.rxFifo.fifo_0[5] ;
 wire \modem.uart.rxFifo.fifo_0[6] ;
 wire \modem.uart.rxFifo.fifo_0[7] ;
 wire \modem.uart.rxFifo.fifo_1[0] ;
 wire \modem.uart.rxFifo.fifo_1[1] ;
 wire \modem.uart.rxFifo.fifo_1[2] ;
 wire \modem.uart.rxFifo.fifo_1[3] ;
 wire \modem.uart.rxFifo.fifo_1[4] ;
 wire \modem.uart.rxFifo.fifo_1[5] ;
 wire \modem.uart.rxFifo.fifo_1[6] ;
 wire \modem.uart.rxFifo.fifo_1[7] ;
 wire \modem.uart.rxFifo.fifo_2[0] ;
 wire \modem.uart.rxFifo.fifo_2[1] ;
 wire \modem.uart.rxFifo.fifo_2[2] ;
 wire \modem.uart.rxFifo.fifo_2[3] ;
 wire \modem.uart.rxFifo.fifo_2[4] ;
 wire \modem.uart.rxFifo.fifo_2[5] ;
 wire \modem.uart.rxFifo.fifo_2[6] ;
 wire \modem.uart.rxFifo.fifo_2[7] ;
 wire \modem.uart.rxFifo.fifo_3[0] ;
 wire \modem.uart.rxFifo.fifo_3[1] ;
 wire \modem.uart.rxFifo.fifo_3[2] ;
 wire \modem.uart.rxFifo.fifo_3[3] ;
 wire \modem.uart.rxFifo.fifo_3[4] ;
 wire \modem.uart.rxFifo.fifo_3[5] ;
 wire \modem.uart.rxFifo.fifo_3[6] ;
 wire \modem.uart.rxFifo.fifo_3[7] ;
 wire \modem.uart.rxFifo.fifo_4[0] ;
 wire \modem.uart.rxFifo.fifo_4[1] ;
 wire \modem.uart.rxFifo.fifo_4[2] ;
 wire \modem.uart.rxFifo.fifo_4[3] ;
 wire \modem.uart.rxFifo.fifo_4[4] ;
 wire \modem.uart.rxFifo.fifo_4[5] ;
 wire \modem.uart.rxFifo.fifo_4[6] ;
 wire \modem.uart.rxFifo.fifo_4[7] ;
 wire \modem.uart.rxFifo.fifo_5[0] ;
 wire \modem.uart.rxFifo.fifo_5[1] ;
 wire \modem.uart.rxFifo.fifo_5[2] ;
 wire \modem.uart.rxFifo.fifo_5[3] ;
 wire \modem.uart.rxFifo.fifo_5[4] ;
 wire \modem.uart.rxFifo.fifo_5[5] ;
 wire \modem.uart.rxFifo.fifo_5[6] ;
 wire \modem.uart.rxFifo.fifo_5[7] ;
 wire \modem.uart.rxFifo.fifo_6[0] ;
 wire \modem.uart.rxFifo.fifo_6[1] ;
 wire \modem.uart.rxFifo.fifo_6[2] ;
 wire \modem.uart.rxFifo.fifo_6[3] ;
 wire \modem.uart.rxFifo.fifo_6[4] ;
 wire \modem.uart.rxFifo.fifo_6[5] ;
 wire \modem.uart.rxFifo.fifo_6[6] ;
 wire \modem.uart.rxFifo.fifo_6[7] ;
 wire \modem.uart.rxFifo.fifo_7[0] ;
 wire \modem.uart.rxFifo.fifo_7[1] ;
 wire \modem.uart.rxFifo.fifo_7[2] ;
 wire \modem.uart.rxFifo.fifo_7[3] ;
 wire \modem.uart.rxFifo.fifo_7[4] ;
 wire \modem.uart.rxFifo.fifo_7[5] ;
 wire \modem.uart.rxFifo.fifo_7[6] ;
 wire \modem.uart.rxFifo.fifo_7[7] ;
 wire \modem.uart.rxFifo.io_dataInEn ;
 wire \modem.uart.rxFifo.io_dataIn[0] ;
 wire \modem.uart.rxFifo.io_dataIn[1] ;
 wire \modem.uart.rxFifo.io_dataIn[2] ;
 wire \modem.uart.rxFifo.io_dataIn[3] ;
 wire \modem.uart.rxFifo.io_dataIn[4] ;
 wire \modem.uart.rxFifo.io_dataIn[5] ;
 wire \modem.uart.rxFifo.io_dataIn[6] ;
 wire \modem.uart.rxFifo.io_dataIn[7] ;
 wire \modem.uart.rxFifo.nextIn[0] ;
 wire \modem.uart.rxFifo.nextIn[1] ;
 wire \modem.uart.rxFifo.nextIn[2] ;
 wire \modem.uart.rxFifo.nextOut[0] ;
 wire \modem.uart.rxFifo.nextOut[1] ;
 wire \modem.uart.rxFifo.nextOut[2] ;
 wire \modem.uart.rxHdlc.canInhibit ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_bit[0] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_bit[1] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_bit[2] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_rxByte[0] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_rxByte[1] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_rxByte[2] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_rxByte[3] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_rxByte[4] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_rxByte[5] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_rxByte[6] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_stateReg[0] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_stateReg[1] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_stateReg[2] ;
 wire \modem.uart.rxHdlc.fsmHdlcRx_stateReg[3] ;
 wire \modem.uart.rxHdlc.io_payload[0] ;
 wire \modem.uart.rxHdlc.io_payload[1] ;
 wire \modem.uart.rxHdlc.io_payload[2] ;
 wire \modem.uart.rxHdlc.io_payload[3] ;
 wire \modem.uart.rxHdlc.io_payload[4] ;
 wire \modem.uart.rxHdlc.io_payload[5] ;
 wire \modem.uart.rxHdlc.io_payload[6] ;
 wire \modem.uart.rxHdlc.io_payload[7] ;
 wire \modem.uart.rxHdlc.io_valid ;
 wire \modem.uart.rxHdlc.oneBitCount[0] ;
 wire \modem.uart.rxHdlc.oneBitCount[1] ;
 wire \modem.uart.rxHdlc.oneBitCount[2] ;
 wire \modem.uart.rxHdlc.regNextRxDataIn ;
 wire \modem.uart.rxUart._zz_sampleValue_29 ;
 wire \modem.uart.rxUart.bitId[0] ;
 wire \modem.uart.rxUart.bitId[1] ;
 wire \modem.uart.rxUart.bitId[2] ;
 wire \modem.uart.rxUart.fsmUartRx_stateReg[1] ;
 wire \modem.uart.rxUart.fsmUartRx_stateReg[2] ;
 wire \modem.uart.rxUart.fsmUartRx_stateReg[3] ;
 wire \modem.uart.rxUart.fsmUartRx_stateReg[4] ;
 wire \modem.uart.rxUart.fsmUartRx_stateReg[5] ;
 wire \modem.uart.rxUart.io_uartRxIn_buffercc.buffers_0 ;
 wire \modem.uart.rxUart.io_uartRxIn_buffercc.buffers_1 ;
 wire \modem.uart.rxUart.sampleTimer_counter[0] ;
 wire \modem.uart.rxUart.sampleTimer_counter[1] ;
 wire \modem.uart.rxUart.sampleTimer_counter[2] ;
 wire \modem.uart.rxUart.samples_2 ;
 wire \modem.uart.rxUart.samples_3 ;
 wire \modem.uart.rxUart.samples_4 ;
 wire \modem.uart.rxUart.samples_5 ;
 wire \modem.uart.rxUart.samples_6 ;
 wire \modem.uart.tx.bitId[0] ;
 wire \modem.uart.tx.bitId[1] ;
 wire \modem.uart.tx.bitId[2] ;
 wire \modem.uart.tx.fsmUartTx_stateReg[1] ;
 wire \modem.uart.tx.fsmUartTx_stateReg[2] ;
 wire \modem.uart.tx.fsmUartTx_stateReg[3] ;
 wire \modem.uart.tx.fsmUartTx_stateReg[4] ;
 wire \modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[1] ;
 wire \modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[2] ;
 wire \modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[3] ;
 wire \modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[4] ;
 wire \modem.uart.txCommandDecoder.io_valid ;
 wire \modem.uart.txCommandDecoder.io_wantTx ;
 wire \modem.uart.txFifo.count[0] ;
 wire \modem.uart.txFifo.count[1] ;
 wire \modem.uart.txFifo.count[2] ;
 wire \modem.uart.txFifo.fifo_0[0] ;
 wire \modem.uart.txFifo.fifo_0[1] ;
 wire \modem.uart.txFifo.fifo_0[2] ;
 wire \modem.uart.txFifo.fifo_0[3] ;
 wire \modem.uart.txFifo.fifo_0[4] ;
 wire \modem.uart.txFifo.fifo_0[5] ;
 wire \modem.uart.txFifo.fifo_0[6] ;
 wire \modem.uart.txFifo.fifo_0[7] ;
 wire \modem.uart.txFifo.fifo_1[0] ;
 wire \modem.uart.txFifo.fifo_1[1] ;
 wire \modem.uart.txFifo.fifo_1[2] ;
 wire \modem.uart.txFifo.fifo_1[3] ;
 wire \modem.uart.txFifo.fifo_1[4] ;
 wire \modem.uart.txFifo.fifo_1[5] ;
 wire \modem.uart.txFifo.fifo_1[6] ;
 wire \modem.uart.txFifo.fifo_1[7] ;
 wire \modem.uart.txFifo.fifo_2[0] ;
 wire \modem.uart.txFifo.fifo_2[1] ;
 wire \modem.uart.txFifo.fifo_2[2] ;
 wire \modem.uart.txFifo.fifo_2[3] ;
 wire \modem.uart.txFifo.fifo_2[4] ;
 wire \modem.uart.txFifo.fifo_2[5] ;
 wire \modem.uart.txFifo.fifo_2[6] ;
 wire \modem.uart.txFifo.fifo_2[7] ;
 wire \modem.uart.txFifo.fifo_3[0] ;
 wire \modem.uart.txFifo.fifo_3[1] ;
 wire \modem.uart.txFifo.fifo_3[2] ;
 wire \modem.uart.txFifo.fifo_3[3] ;
 wire \modem.uart.txFifo.fifo_3[4] ;
 wire \modem.uart.txFifo.fifo_3[5] ;
 wire \modem.uart.txFifo.fifo_3[6] ;
 wire \modem.uart.txFifo.fifo_3[7] ;
 wire \modem.uart.txFifo.nextIn[0] ;
 wire \modem.uart.txFifo.nextIn[1] ;
 wire \modem.uart.txFifo.nextOut[0] ;
 wire \modem.uart.txFifo.nextOut[1] ;
 wire \modem.uart.txHdlc.bit8[0] ;
 wire \modem.uart.txHdlc.bit8[1] ;
 wire \modem.uart.txHdlc.bit8[2] ;
 wire \modem.uart.txHdlc.bitstuffCnt[0] ;
 wire \modem.uart.txHdlc.bitstuffCnt[1] ;
 wire \modem.uart.txHdlc.bitstuffCnt[2] ;
 wire \modem.uart.txHdlc.isAbort ;
 wire \modem.uart.txHdlc.isCRC ;
 wire \modem.uart.txHdlc.txCrc.crcNext_1 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_10 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_11 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_13 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_14 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_15 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_2 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_3 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_4 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_6 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_7 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_8 ;
 wire \modem.uart.txHdlc.txCrc.crcNext_9 ;
 wire \modem.uart.txHdlc.txCrc.crc[11] ;
 wire \modem.uart.txHdlc.txCrc.crc[15] ;
 wire \modem.uart.txHdlc.txCrc.crc[4] ;
 wire \modem.uart.txHdlc.wantFrameEnd ;
 wire \modem.uart.txHdlc.when_ModemTop_l593 ;
 wire \modem.uart.txPacketUpper.fsmKissDecoder_stateReg[1] ;
 wire \modem.uart.txPacketUpper.fsmKissDecoder_stateReg[2] ;
 wire \modem.uart.txPacketUpper.fsmKissDecoder_stateReg[3] ;
 wire \modem.uart.txPacketUpper.fsmKissDecoder_stateReg[4] ;
 wire \modem.uart.txPacketUpper.fsmKissDecoder_stateReg[5] ;
 wire \modem.uart.txPacketUpper.fsmKissDecoder_stateReg[6] ;
 wire \modem.uart.txPacketUpper.io_ready ;
 wire \modem.uart.uart_txCommandDecoder_io_wantTx_regNext ;
 wire \modem.uart.uart_txPacketUpper_io_ready_regNext ;
 wire net13;
 wire net14;
 wire net15;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;

 sg13g2_inv_1 _1790_ (.Y(_0943_),
    .A(net493));
 sg13g2_inv_1 _1791_ (.Y(_0944_),
    .A(net417));
 sg13g2_inv_1 _1792_ (.Y(_0945_),
    .A(net841));
 sg13g2_inv_1 _1793_ (.Y(_0946_),
    .A(\modem.dcdHistory_4 ));
 sg13g2_inv_1 _1794_ (.Y(_0947_),
    .A(net817));
 sg13g2_inv_1 _1795_ (.Y(_0948_),
    .A(net776));
 sg13g2_inv_1 _1796_ (.Y(_0949_),
    .A(net866));
 sg13g2_inv_1 _1797_ (.Y(_0950_),
    .A(net482));
 sg13g2_inv_1 _1798_ (.Y(_0951_),
    .A(net531));
 sg13g2_inv_1 _1799_ (.Y(_0952_),
    .A(net521));
 sg13g2_inv_1 _1800_ (.Y(_0953_),
    .A(net659));
 sg13g2_inv_1 _1801_ (.Y(_0954_),
    .A(net681));
 sg13g2_inv_1 _1802_ (.Y(_0955_),
    .A(net324));
 sg13g2_inv_1 _1803_ (.Y(_0956_),
    .A(net520));
 sg13g2_inv_1 _1804_ (.Y(_0957_),
    .A(net489));
 sg13g2_inv_1 _1805_ (.Y(_0958_),
    .A(net655));
 sg13g2_inv_1 _1806_ (.Y(_0959_),
    .A(net674));
 sg13g2_inv_1 _1807_ (.Y(_0960_),
    .A(net555));
 sg13g2_inv_1 _1808_ (.Y(_0961_),
    .A(net670));
 sg13g2_inv_1 _1809_ (.Y(_0962_),
    .A(net690));
 sg13g2_inv_1 _1810_ (.Y(_0963_),
    .A(net700));
 sg13g2_inv_1 _1811_ (.Y(_0964_),
    .A(net760));
 sg13g2_inv_1 _1812_ (.Y(_0965_),
    .A(net703));
 sg13g2_inv_1 _1813_ (.Y(_0966_),
    .A(\modem.control._zz_txClockInternalFallStb ));
 sg13g2_inv_1 _1814_ (.Y(_0967_),
    .A(\modem.control.rxAddr[1] ));
 sg13g2_inv_1 _1815_ (.Y(_0968_),
    .A(net307));
 sg13g2_inv_1 _1816_ (.Y(_0969_),
    .A(\modem.control.rxAddr[5] ));
 sg13g2_inv_1 _1817_ (.Y(_0970_),
    .A(net622));
 sg13g2_inv_1 _1818_ (.Y(_0971_),
    .A(net431));
 sg13g2_inv_1 _1819_ (.Y(_0972_),
    .A(net340));
 sg13g2_inv_2 _1820_ (.Y(_0973_),
    .A(net835));
 sg13g2_inv_2 _1821_ (.Y(_0974_),
    .A(\modem.uart.rxHdlc.io_payload[6] ));
 sg13g2_inv_2 _1822_ (.Y(_0975_),
    .A(\modem.uart.rxHdlc.io_payload[5] ));
 sg13g2_inv_2 _1823_ (.Y(_0976_),
    .A(\modem.uart.rxHdlc.io_payload[4] ));
 sg13g2_inv_2 _1824_ (.Y(_0977_),
    .A(\modem.uart.rxHdlc.io_payload[3] ));
 sg13g2_inv_2 _1825_ (.Y(_0978_),
    .A(\modem.uart.rxHdlc.io_payload[2] ));
 sg13g2_inv_2 _1826_ (.Y(_0979_),
    .A(\modem.uart.rxHdlc.io_payload[1] ));
 sg13g2_inv_2 _1827_ (.Y(_0980_),
    .A(\modem.uart.rxHdlc.io_payload[0] ));
 sg13g2_inv_1 _1828_ (.Y(_0981_),
    .A(net305));
 sg13g2_inv_1 _1829_ (.Y(_0982_),
    .A(\modem.uart.txFifo.nextIn[0] ));
 sg13g2_inv_1 _1830_ (.Y(_0983_),
    .A(net794));
 sg13g2_inv_1 _1831_ (.Y(_0984_),
    .A(net691));
 sg13g2_inv_2 _1832_ (.Y(_0985_),
    .A(net429));
 sg13g2_inv_4 _1833_ (.A(net715),
    .Y(_0986_));
 sg13g2_inv_4 _1834_ (.A(net728),
    .Y(_0987_));
 sg13g2_inv_4 _1835_ (.A(net757),
    .Y(_0988_));
 sg13g2_inv_4 _1836_ (.A(net769),
    .Y(_0989_));
 sg13g2_inv_1 _1837_ (.Y(_0990_),
    .A(net606));
 sg13g2_inv_4 _1838_ (.A(net720),
    .Y(_0991_));
 sg13g2_inv_4 _1839_ (.A(\modem.uart.rxFifo.io_dataIn[1] ),
    .Y(_0992_));
 sg13g2_inv_1 _1840_ (.Y(_0993_),
    .A(net542));
 sg13g2_inv_1 _1841_ (.Y(_0994_),
    .A(net319));
 sg13g2_inv_1 _1842_ (.Y(_0995_),
    .A(net418));
 sg13g2_inv_1 _1843_ (.Y(_0996_),
    .A(net313));
 sg13g2_inv_1 _1844_ (.Y(_0997_),
    .A(net684));
 sg13g2_inv_1 _1845_ (.Y(_0998_),
    .A(\modem.uart.rxUart.samples_4 ));
 sg13g2_inv_1 _1846_ (.Y(_0999_),
    .A(net897));
 sg13g2_inv_1 _1847_ (.Y(_1000_),
    .A(net742));
 sg13g2_inv_1 _1848_ (.Y(_1001_),
    .A(net445));
 sg13g2_inv_1 _1849_ (.Y(_1002_),
    .A(\modem.uart.tx.fsmUartTx_stateReg[2] ));
 sg13g2_inv_1 _1850_ (.Y(_1003_),
    .A(net676));
 sg13g2_inv_1 _1851_ (.Y(_1004_),
    .A(net799));
 sg13g2_inv_1 _1852_ (.Y(_1005_),
    .A(\modem.uart.rxUart.bitId[0] ));
 sg13g2_inv_2 _1853_ (.Y(_1006_),
    .A(\modem.uart.tx.bitId[0] ));
 sg13g2_inv_1 _1854_ (.Y(_1007_),
    .A(\modem.uart.rxHdlc.oneBitCount[0] ));
 sg13g2_inv_1 _1855_ (.Y(_1008_),
    .A(_0054_));
 sg13g2_inv_2 _1856_ (.Y(_1009_),
    .A(net424));
 sg13g2_inv_2 _1857_ (.Y(_1010_),
    .A(net422));
 sg13g2_inv_1 _1858_ (.Y(_1011_),
    .A(\modem.uart.txHdlc.wantFrameEnd ));
 sg13g2_inv_1 _1859_ (.Y(_1012_),
    .A(\modem.uart.io_isSending ));
 sg13g2_inv_1 _1860_ (.Y(_1013_),
    .A(net412));
 sg13g2_inv_1 _1861_ (.Y(_1014_),
    .A(_0035_));
 sg13g2_inv_1 _1862_ (.Y(_1015_),
    .A(_0034_));
 sg13g2_inv_1 _1863_ (.Y(_1016_),
    .A(_0033_));
 sg13g2_inv_1 _1864_ (.Y(_1017_),
    .A(net3));
 sg13g2_inv_1 _1865_ (.Y(_1018_),
    .A(\modem.uart.txFifo.fifo_3[0] ));
 sg13g2_inv_1 _1866_ (.Y(_1019_),
    .A(net870));
 sg13g2_inv_1 _1867_ (.Y(\modem.cfgAddrDirection ),
    .A(\latched[7] ));
 sg13g2_inv_1 _1868_ (.Y(\modem.cfgUpDownSource ),
    .A(\latched[6] ));
 sg13g2_inv_1 _1869_ (.Y(\modem.cfgRxClockDirection ),
    .A(\latched[5] ));
 sg13g2_inv_1 _1870_ (.Y(_1020_),
    .A(net852));
 sg13g2_inv_1 _1871_ (.Y(_1021_),
    .A(\modem.uart.rxUart.bitId[2] ));
 sg13g2_inv_1 _1872_ (.Y(_1022_),
    .A(net302));
 sg13g2_inv_1 _1873_ (.Y(_1023_),
    .A(net434));
 sg13g2_inv_1 _1874_ (.Y(_1024_),
    .A(_0075_));
 sg13g2_inv_1 _1875_ (.Y(_1025_),
    .A(_0058_));
 sg13g2_inv_1 _1876_ (.Y(_1026_),
    .A(net630));
 sg13g2_and2_1 _1877_ (.A(\latched[6] ),
    .B(\modem.analog_rxDac8[7] ),
    .X(_1027_));
 sg13g2_a21oi_1 _1878_ (.A1(\modem.cfgUpDownSource ),
    .A2(net8),
    .Y(_1028_),
    .B1(_1027_));
 sg13g2_inv_1 _1879_ (.Y(\modem.control.io_upDownOut ),
    .A(net369));
 sg13g2_nor2b_1 _1880_ (.A(\modem.control._zz__1_regNext ),
    .B_N(\latched[1] ),
    .Y(_1029_));
 sg13g2_nor3_1 _1881_ (.A(_1022_),
    .B(\modem.control._zz__regNext ),
    .C(\latched[1] ),
    .Y(_1030_));
 sg13g2_a21oi_2 _1882_ (.B1(_1030_),
    .Y(_1031_),
    .A2(_1029_),
    .A1(\modem.control._zz__1 ));
 sg13g2_a21o_2 _1883_ (.A2(_1029_),
    .A1(\modem.control._zz__1 ),
    .B1(_1030_),
    .X(_1032_));
 sg13g2_nor2_2 _1884_ (.A(net885),
    .B(net368),
    .Y(_1033_));
 sg13g2_nand2b_2 _1885_ (.Y(_1034_),
    .B(net366),
    .A_N(\modem.uart.txHdlc.isAbort ));
 sg13g2_nor3_2 _1886_ (.A(net430),
    .B(_0057_),
    .C(_1034_),
    .Y(_1035_));
 sg13g2_and2_2 _1887_ (.A(net425),
    .B(net423),
    .X(_1036_));
 sg13g2_nand2_1 _1888_ (.Y(_1037_),
    .A(net427),
    .B(net424));
 sg13g2_nor3_2 _1889_ (.A(_1010_),
    .B(\modem.uart.txHdlc.when_ModemTop_l593 ),
    .C(_1037_),
    .Y(_1038_));
 sg13g2_nand2_1 _1890_ (.Y(_1039_),
    .A(net816),
    .B(_1038_));
 sg13g2_nand3_1 _1891_ (.B(_1035_),
    .C(_1038_),
    .A(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[4] ),
    .Y(_1040_));
 sg13g2_nor2_1 _1892_ (.A(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[2] ),
    .B(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[3] ),
    .Y(_1041_));
 sg13g2_nand3_1 _1893_ (.B(_1040_),
    .C(_1041_),
    .A(\modem.uart.txCommandDecoder.io_valid ),
    .Y(_1042_));
 sg13g2_nor2_2 _1894_ (.A(net405),
    .B(_1042_),
    .Y(_1043_));
 sg13g2_nor4_2 _1895_ (.A(\modem.uart.rxFifo.count[3] ),
    .B(\modem.uart.rxFifo.count[2] ),
    .C(\modem.uart.rxFifo.count[1] ),
    .Y(_1044_),
    .D(\modem.uart.rxFifo.count[0] ));
 sg13g2_nor2_2 _1896_ (.A(net439),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_nor2b_1 _1897_ (.A(\modem.uart.rxFifo.nextOut[0] ),
    .B_N(\modem.uart.rxFifo.nextOut[1] ),
    .Y(_1046_));
 sg13g2_and2_1 _1898_ (.A(net433),
    .B(net399),
    .X(_1047_));
 sg13g2_nor2_2 _1899_ (.A(\modem.uart.rxFifo.nextOut[1] ),
    .B(\modem.uart.rxFifo.nextOut[0] ),
    .Y(_1048_));
 sg13g2_and2_2 _1900_ (.A(net436),
    .B(_1048_),
    .X(_1049_));
 sg13g2_nor3_2 _1901_ (.A(net435),
    .B(\modem.uart.rxFifo.nextOut[1] ),
    .C(\modem.uart.rxFifo.nextOut[0] ),
    .Y(_1050_));
 sg13g2_and2_1 _1902_ (.A(\modem.uart.rxFifo.fifo_0[5] ),
    .B(_1050_),
    .X(_1051_));
 sg13g2_a221oi_1 _1903_ (.B2(\modem.uart.rxFifo.fifo_4[5] ),
    .C1(_1051_),
    .B1(_1049_),
    .A1(\modem.uart.rxFifo.fifo_2[5] ),
    .Y(_1052_),
    .A2(_1047_));
 sg13g2_nor2b_1 _1904_ (.A(\modem.uart.rxFifo.nextOut[1] ),
    .B_N(\modem.uart.rxFifo.nextOut[0] ),
    .Y(_1053_));
 sg13g2_and2_2 _1905_ (.A(net402),
    .B(net397),
    .X(_1054_));
 sg13g2_nand3_1 _1906_ (.B(\modem.uart.rxFifo.fifo_5[5] ),
    .C(net397),
    .A(net402),
    .Y(_1055_));
 sg13g2_and2_1 _1907_ (.A(\modem.uart.rxFifo.nextOut[1] ),
    .B(\modem.uart.rxFifo.nextOut[0] ),
    .X(_1056_));
 sg13g2_and2_1 _1908_ (.A(net436),
    .B(net396),
    .X(_1057_));
 sg13g2_o21ai_1 _1909_ (.B1(net396),
    .Y(_1058_),
    .A1(net436),
    .A2(\modem.uart.rxFifo.fifo_3[5] ));
 sg13g2_nand3_1 _1910_ (.B(\modem.uart.rxFifo.fifo_1[5] ),
    .C(net397),
    .A(net433),
    .Y(_1059_));
 sg13g2_nand3_1 _1911_ (.B(\modem.uart.rxFifo.fifo_6[5] ),
    .C(net399),
    .A(net402),
    .Y(_1060_));
 sg13g2_and4_1 _1912_ (.A(_1055_),
    .B(_1058_),
    .C(_1059_),
    .D(_1060_),
    .X(_1061_));
 sg13g2_and2_1 _1913_ (.A(_0041_),
    .B(net388),
    .X(_1062_));
 sg13g2_a21o_1 _1914_ (.A2(_1061_),
    .A1(_1052_),
    .B1(_1062_),
    .X(_1063_));
 sg13g2_nand2_1 _1915_ (.Y(_1064_),
    .A(\modem.uart.rxFifo.fifo_0[7] ),
    .B(_1050_));
 sg13g2_and3_1 _1916_ (.X(_1065_),
    .A(net433),
    .B(\modem.uart.rxFifo.fifo_1[7] ),
    .C(net397));
 sg13g2_o21ai_1 _1917_ (.B1(_1056_),
    .Y(_1066_),
    .A1(net436),
    .A2(\modem.uart.rxFifo.fifo_3[7] ));
 sg13g2_nand3_1 _1918_ (.B(\modem.uart.rxFifo.fifo_5[7] ),
    .C(net398),
    .A(net402),
    .Y(_1067_));
 sg13g2_nand3_1 _1919_ (.B(\modem.uart.rxFifo.fifo_6[7] ),
    .C(net400),
    .A(net402),
    .Y(_1068_));
 sg13g2_a221oi_1 _1920_ (.B2(\modem.uart.rxFifo.fifo_4[7] ),
    .C1(_1065_),
    .B1(_1049_),
    .A1(\modem.uart.rxFifo.fifo_2[7] ),
    .Y(_1069_),
    .A2(_1047_));
 sg13g2_and4_1 _1921_ (.A(_1064_),
    .B(_1066_),
    .C(_1067_),
    .D(_1068_),
    .X(_1070_));
 sg13g2_a22oi_1 _1922_ (.Y(_1071_),
    .B1(_1069_),
    .B2(_1070_),
    .A2(net388),
    .A1(_0039_));
 sg13g2_and2_1 _1923_ (.A(_1063_),
    .B(_1071_),
    .X(_1072_));
 sg13g2_and3_1 _1924_ (.X(_1073_),
    .A(net433),
    .B(\modem.uart.rxFifo.fifo_1[6] ),
    .C(net397));
 sg13g2_a221oi_1 _1925_ (.B2(\modem.uart.rxFifo.fifo_5[6] ),
    .C1(_1073_),
    .B1(_1054_),
    .A1(\modem.uart.rxFifo.fifo_2[6] ),
    .Y(_1074_),
    .A2(_1047_));
 sg13g2_nand3_1 _1926_ (.B(\modem.uart.rxFifo.fifo_4[6] ),
    .C(_1048_),
    .A(net435),
    .Y(_1075_));
 sg13g2_o21ai_1 _1927_ (.B1(_1056_),
    .Y(_1076_),
    .A1(net435),
    .A2(\modem.uart.rxFifo.fifo_3[6] ));
 sg13g2_nand2_1 _1928_ (.Y(_1077_),
    .A(\modem.uart.rxFifo.fifo_0[6] ),
    .B(_1050_));
 sg13g2_nand3_1 _1929_ (.B(\modem.uart.rxFifo.fifo_6[6] ),
    .C(net400),
    .A(net403),
    .Y(_1078_));
 sg13g2_and4_1 _1930_ (.A(_1075_),
    .B(_1076_),
    .C(_1077_),
    .D(_1078_),
    .X(_1079_));
 sg13g2_a22oi_1 _1931_ (.Y(_1080_),
    .B1(_1074_),
    .B2(_1079_),
    .A2(net388),
    .A1(_0040_));
 sg13g2_nand3_1 _1932_ (.B(\modem.uart.rxFifo.fifo_6[4] ),
    .C(net399),
    .A(net402),
    .Y(_1081_));
 sg13g2_and3_1 _1933_ (.X(_1082_),
    .A(net433),
    .B(\modem.uart.rxFifo.fifo_1[4] ),
    .C(net397));
 sg13g2_o21ai_1 _1934_ (.B1(net396),
    .Y(_1083_),
    .A1(net436),
    .A2(\modem.uart.rxFifo.fifo_3[4] ));
 sg13g2_nand3_1 _1935_ (.B(\modem.uart.rxFifo.fifo_2[4] ),
    .C(net399),
    .A(net433),
    .Y(_1084_));
 sg13g2_nand2_1 _1936_ (.Y(_1085_),
    .A(\modem.uart.rxFifo.fifo_0[4] ),
    .B(_1050_));
 sg13g2_a221oi_1 _1937_ (.B2(\modem.uart.rxFifo.fifo_5[4] ),
    .C1(_1082_),
    .B1(_1054_),
    .A1(\modem.uart.rxFifo.fifo_4[4] ),
    .Y(_1086_),
    .A2(_1049_));
 sg13g2_and4_1 _1938_ (.A(_1081_),
    .B(_1083_),
    .C(_1084_),
    .D(_1085_),
    .X(_1087_));
 sg13g2_a22oi_1 _1939_ (.Y(_1088_),
    .B1(_1086_),
    .B2(_1087_),
    .A2(net388),
    .A1(_0042_));
 sg13g2_and4_1 _1940_ (.A(_1063_),
    .B(_1071_),
    .C(_1080_),
    .D(_1088_),
    .X(_1089_));
 sg13g2_nand4_1 _1941_ (.B(_1071_),
    .C(_1080_),
    .A(_1063_),
    .Y(_1090_),
    .D(_1088_));
 sg13g2_and3_1 _1942_ (.X(_1091_),
    .A(net434),
    .B(\modem.uart.rxFifo.fifo_1[2] ),
    .C(net398));
 sg13g2_a221oi_1 _1943_ (.B2(\modem.uart.rxFifo.fifo_5[2] ),
    .C1(_1091_),
    .B1(_1054_),
    .A1(\modem.uart.rxFifo.fifo_0[2] ),
    .Y(_1092_),
    .A2(_1050_));
 sg13g2_nand3_1 _1944_ (.B(\modem.uart.rxFifo.fifo_4[2] ),
    .C(_1048_),
    .A(net435),
    .Y(_1093_));
 sg13g2_o21ai_1 _1945_ (.B1(net396),
    .Y(_1094_),
    .A1(net435),
    .A2(\modem.uart.rxFifo.fifo_3[2] ));
 sg13g2_nand3_1 _1946_ (.B(\modem.uart.rxFifo.fifo_2[2] ),
    .C(net400),
    .A(net434),
    .Y(_1095_));
 sg13g2_nand3_1 _1947_ (.B(\modem.uart.rxFifo.fifo_6[2] ),
    .C(net400),
    .A(net403),
    .Y(_1096_));
 sg13g2_and4_1 _1948_ (.A(_1093_),
    .B(_1094_),
    .C(_1095_),
    .D(_1096_),
    .X(_1097_));
 sg13g2_a22oi_1 _1949_ (.Y(_1098_),
    .B1(_1092_),
    .B2(_1097_),
    .A2(net388),
    .A1(_0044_));
 sg13g2_and2_1 _1950_ (.A(\modem.uart.rxFifo.fifo_0[0] ),
    .B(_1050_),
    .X(_1099_));
 sg13g2_a221oi_1 _1951_ (.B2(\modem.uart.rxFifo.fifo_5[0] ),
    .C1(_1099_),
    .B1(_1054_),
    .A1(\modem.uart.rxFifo.fifo_4[0] ),
    .Y(_1100_),
    .A2(_1049_));
 sg13g2_nand3_1 _1952_ (.B(\modem.uart.rxFifo.fifo_1[0] ),
    .C(net398),
    .A(net434),
    .Y(_1101_));
 sg13g2_o21ai_1 _1953_ (.B1(net396),
    .Y(_1102_),
    .A1(net435),
    .A2(\modem.uart.rxFifo.fifo_3[0] ));
 sg13g2_nand3_1 _1954_ (.B(\modem.uart.rxFifo.fifo_2[0] ),
    .C(net399),
    .A(net434),
    .Y(_1103_));
 sg13g2_nand3_1 _1955_ (.B(\modem.uart.rxFifo.fifo_6[0] ),
    .C(net399),
    .A(net402),
    .Y(_1104_));
 sg13g2_and4_1 _1956_ (.A(_1101_),
    .B(_1102_),
    .C(_1103_),
    .D(_1104_),
    .X(_1105_));
 sg13g2_and2_1 _1957_ (.A(_0046_),
    .B(_1057_),
    .X(_1106_));
 sg13g2_a21o_2 _1958_ (.A2(_1105_),
    .A1(_1100_),
    .B1(_1106_),
    .X(_1107_));
 sg13g2_nand2_1 _1959_ (.Y(_1108_),
    .A(\modem.uart.rxFifo.fifo_0[3] ),
    .B(_1050_));
 sg13g2_and3_1 _1960_ (.X(_1109_),
    .A(net433),
    .B(\modem.uart.rxFifo.fifo_1[3] ),
    .C(net397));
 sg13g2_o21ai_1 _1961_ (.B1(_1056_),
    .Y(_1110_),
    .A1(net435),
    .A2(\modem.uart.rxFifo.fifo_3[3] ));
 sg13g2_nand3_1 _1962_ (.B(\modem.uart.rxFifo.fifo_5[3] ),
    .C(net398),
    .A(net403),
    .Y(_1111_));
 sg13g2_nand3_1 _1963_ (.B(\modem.uart.rxFifo.fifo_6[3] ),
    .C(net400),
    .A(net403),
    .Y(_1112_));
 sg13g2_a221oi_1 _1964_ (.B2(\modem.uart.rxFifo.fifo_4[3] ),
    .C1(_1109_),
    .B1(_1049_),
    .A1(\modem.uart.rxFifo.fifo_2[3] ),
    .Y(_1113_),
    .A2(_1047_));
 sg13g2_and4_1 _1965_ (.A(_1108_),
    .B(_1110_),
    .C(_1111_),
    .D(_1112_),
    .X(_1114_));
 sg13g2_a22oi_1 _1966_ (.Y(_1115_),
    .B1(_1113_),
    .B2(_1114_),
    .A2(net388),
    .A1(_0043_));
 sg13g2_and2_1 _1967_ (.A(\modem.uart.rxFifo.fifo_0[1] ),
    .B(_1050_),
    .X(_1116_));
 sg13g2_a221oi_1 _1968_ (.B2(\modem.uart.rxFifo.fifo_5[1] ),
    .C1(_1116_),
    .B1(_1054_),
    .A1(\modem.uart.rxFifo.fifo_4[1] ),
    .Y(_1117_),
    .A2(_1049_));
 sg13g2_nand3_1 _1969_ (.B(\modem.uart.rxFifo.fifo_1[1] ),
    .C(net397),
    .A(net434),
    .Y(_1118_));
 sg13g2_o21ai_1 _1970_ (.B1(net396),
    .Y(_1119_),
    .A1(net436),
    .A2(\modem.uart.rxFifo.fifo_3[1] ));
 sg13g2_nand3_1 _1971_ (.B(\modem.uart.rxFifo.fifo_2[1] ),
    .C(net399),
    .A(net433),
    .Y(_1120_));
 sg13g2_nand3_1 _1972_ (.B(\modem.uart.rxFifo.fifo_6[1] ),
    .C(net399),
    .A(net402),
    .Y(_1121_));
 sg13g2_and4_1 _1973_ (.A(_1118_),
    .B(_1119_),
    .C(_1120_),
    .D(_1121_),
    .X(_1122_));
 sg13g2_and2_1 _1974_ (.A(_0045_),
    .B(net388),
    .X(_1123_));
 sg13g2_a21o_1 _1975_ (.A2(_1122_),
    .A1(_1117_),
    .B1(_1123_),
    .X(_1124_));
 sg13g2_nor3_1 _1976_ (.A(_1098_),
    .B(_1107_),
    .C(_1124_),
    .Y(_1125_));
 sg13g2_nand3_1 _1977_ (.B(_1115_),
    .C(_1125_),
    .A(_1089_),
    .Y(_1126_));
 sg13g2_and2_1 _1978_ (.A(_1107_),
    .B(_1124_),
    .X(_1127_));
 sg13g2_nor2_1 _1979_ (.A(_1098_),
    .B(_1115_),
    .Y(_1128_));
 sg13g2_and2_1 _1980_ (.A(_1127_),
    .B(_1128_),
    .X(_1129_));
 sg13g2_nor2b_1 _1981_ (.A(_1088_),
    .B_N(_1080_),
    .Y(_1130_));
 sg13g2_nand3_1 _1982_ (.B(_1129_),
    .C(_1130_),
    .A(_1072_),
    .Y(_1131_));
 sg13g2_nand2_1 _1983_ (.Y(_1132_),
    .A(_1126_),
    .B(_1131_));
 sg13g2_nand3_1 _1984_ (.B(_1126_),
    .C(_1131_),
    .A(net897),
    .Y(_1133_));
 sg13g2_nor3_1 _1985_ (.A(net439),
    .B(net401),
    .C(_1133_),
    .Y(_1134_));
 sg13g2_a21o_1 _1986_ (.A2(_1043_),
    .A1(net610),
    .B1(_1134_),
    .X(_0021_));
 sg13g2_and2_1 _1987_ (.A(_1098_),
    .B(_1115_),
    .X(_1135_));
 sg13g2_nand3_1 _1988_ (.B(_1127_),
    .C(_1135_),
    .A(_1089_),
    .Y(_1136_));
 sg13g2_nor2_1 _1989_ (.A(_1000_),
    .B(net401),
    .Y(_1137_));
 sg13g2_nand2_1 _1990_ (.Y(_1138_),
    .A(net742),
    .B(_1045_));
 sg13g2_nand2_1 _1991_ (.Y(_1139_),
    .A(net723),
    .B(_1043_));
 sg13g2_o21ai_1 _1992_ (.B1(net724),
    .Y(_0020_),
    .A1(_1136_),
    .A2(_1138_));
 sg13g2_nor2_1 _1993_ (.A(net401),
    .B(_1131_),
    .Y(_1140_));
 sg13g2_nand3b_1 _1994_ (.B(net705),
    .C(net442),
    .Y(_1141_),
    .A_N(_1140_));
 sg13g2_nand3_1 _1995_ (.B(_1115_),
    .C(_1124_),
    .A(_1098_),
    .Y(_1142_));
 sg13g2_or2_2 _1996_ (.X(_1143_),
    .B(_1142_),
    .A(_1090_));
 sg13g2_nand2_2 _1997_ (.Y(_1144_),
    .A(_1137_),
    .B(_1143_));
 sg13g2_nand2_2 _1998_ (.Y(_1145_),
    .A(net445),
    .B(net772));
 sg13g2_o21ai_1 _1999_ (.B1(_1145_),
    .Y(_1146_),
    .A1(net439),
    .A2(_1144_));
 sg13g2_nand2b_1 _2000_ (.Y(_0019_),
    .B(_1141_),
    .A_N(_1146_));
 sg13g2_nor2b_1 _2001_ (.A(_0082_),
    .B_N(\modem.uart.rxUart.samples_6 ),
    .Y(_1147_));
 sg13g2_nand2_1 _2002_ (.Y(_1148_),
    .A(\modem.uart.rxUart.io_uartRxIn_buffercc.buffers_1 ),
    .B(\modem.uart.rxUart._zz_sampleValue_29 ));
 sg13g2_nor2_1 _2003_ (.A(_0069_),
    .B(_1148_),
    .Y(_1149_));
 sg13g2_a22oi_1 _2004_ (.Y(_1150_),
    .B1(_1149_),
    .B2(\modem.uart.rxUart.samples_2 ),
    .A2(_1147_),
    .A1(\modem.uart.rxUart.samples_4 ));
 sg13g2_nor3_1 _2005_ (.A(\modem.uart.rxUart.io_uartRxIn_buffercc.buffers_1 ),
    .B(\modem.uart.rxUart._zz_sampleValue_29 ),
    .C(\modem.uart.rxUart.samples_2 ),
    .Y(_1151_));
 sg13g2_nor2b_1 _2006_ (.A(\modem.uart.rxUart.samples_3 ),
    .B_N(_1151_),
    .Y(_1152_));
 sg13g2_o21ai_1 _2007_ (.B1(\modem.uart.rxUart.samples_2 ),
    .Y(_1153_),
    .A1(\modem.uart.rxUart.io_uartRxIn_buffercc.buffers_1 ),
    .A2(\modem.uart.rxUart._zz_sampleValue_29 ));
 sg13g2_o21ai_1 _2008_ (.B1(_1153_),
    .Y(_1154_),
    .A1(_0069_),
    .A2(_1148_));
 sg13g2_nor2_1 _2009_ (.A(\modem.uart.rxUart.samples_5 ),
    .B(\modem.uart.rxUart.samples_6 ),
    .Y(_1155_));
 sg13g2_a22oi_1 _2010_ (.Y(_1156_),
    .B1(_1155_),
    .B2(_0998_),
    .A2(_1148_),
    .A1(_0069_));
 sg13g2_nand2b_1 _2011_ (.Y(_1157_),
    .B(\modem.uart.rxUart.samples_3 ),
    .A_N(_1151_));
 sg13g2_nand3_1 _2012_ (.B(_1153_),
    .C(_1157_),
    .A(_1148_),
    .Y(_1158_));
 sg13g2_nor2_1 _2013_ (.A(_0068_),
    .B(_1155_),
    .Y(_1159_));
 sg13g2_or2_1 _2014_ (.X(_1160_),
    .B(_1159_),
    .A(_1147_));
 sg13g2_a22oi_1 _2015_ (.Y(_1161_),
    .B1(_1158_),
    .B2(_1160_),
    .A2(_1156_),
    .A1(_1154_));
 sg13g2_o21ai_1 _2016_ (.B1(_1161_),
    .Y(_1162_),
    .A1(_1150_),
    .A2(_1152_));
 sg13g2_inv_2 _2017_ (.Y(_1163_),
    .A(_1162_));
 sg13g2_nor3_1 _2018_ (.A(_1013_),
    .B(\modem.control._zz__2_regNext ),
    .C(\latched[0] ),
    .Y(_1164_));
 sg13g2_nand2b_2 _2019_ (.Y(_1165_),
    .B(net626),
    .A_N(\modem.control._zz__3_regNext ));
 sg13g2_inv_2 _2020_ (.Y(\modem.control.io_txClockStb ),
    .A(_1165_));
 sg13g2_a21oi_2 _2021_ (.B1(_1164_),
    .Y(_1166_),
    .A2(\modem.control.io_txClockStb ),
    .A1(\latched[0] ));
 sg13g2_inv_1 _2022_ (.Y(_1167_),
    .A(net364));
 sg13g2_nor2_1 _2023_ (.A(_1162_),
    .B(net364),
    .Y(_1168_));
 sg13g2_nand2_1 _2024_ (.Y(_1169_),
    .A(\modem.uart.rxUart.fsmUartRx_stateReg[2] ),
    .B(_1168_));
 sg13g2_inv_1 _2025_ (.Y(_1170_),
    .A(_1169_));
 sg13g2_nor3_1 _2026_ (.A(\modem.uart.rxUart.sampleTimer_counter[0] ),
    .B(net751),
    .C(net365),
    .Y(_1171_));
 sg13g2_inv_1 _2027_ (.Y(_1172_),
    .A(_1171_));
 sg13g2_nor2_1 _2028_ (.A(\modem.uart.rxUart.sampleTimer_counter[2] ),
    .B(_1172_),
    .Y(_1173_));
 sg13g2_inv_1 _2029_ (.Y(_1174_),
    .A(_1173_));
 sg13g2_nor2_1 _2030_ (.A(net440),
    .B(_1173_),
    .Y(_1175_));
 sg13g2_a22oi_1 _2031_ (.Y(_1176_),
    .B1(_1175_),
    .B2(net653),
    .A2(_1170_),
    .A1(net443));
 sg13g2_inv_1 _2032_ (.Y(_0007_),
    .A(net654));
 sg13g2_nor2_2 _2033_ (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[5] ),
    .B(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[3] ),
    .Y(_1177_));
 sg13g2_and2_1 _2034_ (.A(_0075_),
    .B(_1177_),
    .X(_1178_));
 sg13g2_or2_1 _2035_ (.X(_1179_),
    .B(_1178_),
    .A(_0076_));
 sg13g2_nor2_2 _2036_ (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[1] ),
    .B(_1178_),
    .Y(_1180_));
 sg13g2_inv_1 _2037_ (.Y(_1181_),
    .A(_1180_));
 sg13g2_nor2_1 _2038_ (.A(net401),
    .B(_1178_),
    .Y(_1182_));
 sg13g2_nand4_1 _2039_ (.B(_1127_),
    .C(_1135_),
    .A(_1089_),
    .Y(_1183_),
    .D(_1182_));
 sg13g2_nand3_1 _2040_ (.B(_1181_),
    .C(_1183_),
    .A(_1088_),
    .Y(_1184_));
 sg13g2_and2_1 _2041_ (.A(_1179_),
    .B(_1184_),
    .X(_1185_));
 sg13g2_nor4_1 _2042_ (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[5] ),
    .B(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[3] ),
    .C(_1080_),
    .D(_1180_),
    .Y(_1186_));
 sg13g2_nand4_1 _2043_ (.B(_1129_),
    .C(_1185_),
    .A(_1072_),
    .Y(_1187_),
    .D(_1186_));
 sg13g2_nand2_1 _2044_ (.Y(_1188_),
    .A(net444),
    .B(net860));
 sg13g2_nand3_1 _2045_ (.B(net860),
    .C(\modem.uart.txCommandDecoder.io_valid ),
    .A(net444),
    .Y(_1189_));
 sg13g2_nor3_2 _2046_ (.A(_0999_),
    .B(net401),
    .C(_1131_),
    .Y(_1190_));
 sg13g2_nor2_1 _2047_ (.A(net439),
    .B(_1190_),
    .Y(_1191_));
 sg13g2_nand2_1 _2048_ (.Y(_1192_),
    .A(net518),
    .B(_1191_));
 sg13g2_o21ai_1 _2049_ (.B1(_1192_),
    .Y(_0013_),
    .A1(_1187_),
    .A2(_1189_));
 sg13g2_a21oi_1 _2050_ (.A1(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[4] ),
    .A2(_1190_),
    .Y(_1193_),
    .B1(net784));
 sg13g2_nand2_2 _2051_ (.Y(_1194_),
    .A(\modem.uart.txCommandDecoder.io_valid ),
    .B(_1039_));
 sg13g2_nor3_1 _2052_ (.A(net439),
    .B(net785),
    .C(_1194_),
    .Y(_0012_));
 sg13g2_nor2_2 _2053_ (.A(net408),
    .B(_1031_),
    .Y(_1195_));
 sg13g2_nand2_2 _2054_ (.Y(_1196_),
    .A(net438),
    .B(net437));
 sg13g2_nor2_2 _2055_ (.A(_0070_),
    .B(_1196_),
    .Y(_1197_));
 sg13g2_nand2b_1 _2056_ (.Y(_1198_),
    .B(\modem.uart.tx.fsmUartTx_stateReg[4] ),
    .A_N(net440));
 sg13g2_a21oi_1 _2057_ (.A1(net367),
    .A2(_1197_),
    .Y(_1199_),
    .B1(_1198_));
 sg13g2_a21o_1 _2058_ (.A2(_1195_),
    .A1(net693),
    .B1(_1199_),
    .X(_0011_));
 sg13g2_a21oi_1 _2059_ (.A1(net604),
    .A2(net367),
    .Y(_1200_),
    .B1(net710));
 sg13g2_nor2_1 _2060_ (.A(\modem.uart.txFifo.count[1] ),
    .B(\modem.uart.txFifo.count[0] ),
    .Y(_1201_));
 sg13g2_nor3_1 _2061_ (.A(net624),
    .B(\modem.uart.txFifo.count[1] ),
    .C(\modem.uart.txFifo.count[0] ),
    .Y(_1202_));
 sg13g2_nand2_1 _2062_ (.Y(_1203_),
    .A(net444),
    .B(_1202_));
 sg13g2_o21ai_1 _2063_ (.B1(_1145_),
    .Y(_0010_),
    .A1(_1200_),
    .A2(_1203_));
 sg13g2_nor2_2 _2064_ (.A(net440),
    .B(net367),
    .Y(_1204_));
 sg13g2_nor3_1 _2065_ (.A(net440),
    .B(_1200_),
    .C(_1202_),
    .Y(_1205_));
 sg13g2_a21o_1 _2066_ (.A2(_1204_),
    .A1(net693),
    .B1(_1205_),
    .X(_0009_));
 sg13g2_a21o_1 _2067_ (.A2(\modem.uart.rxFifo.count[1] ),
    .A1(\modem.uart.rxFifo.count[2] ),
    .B1(\modem.uart.rxFifo.count[3] ),
    .X(\modem.uart.io_uartCtsOut ));
 sg13g2_and3_2 _2068_ (.X(_1206_),
    .A(\modem.uart.tx.fsmUartTx_stateReg[4] ),
    .B(net367),
    .C(_1197_));
 sg13g2_a22oi_1 _2069_ (.Y(_1207_),
    .B1(_1206_),
    .B2(net452),
    .A2(_1204_),
    .A1(net604));
 sg13g2_inv_1 _2070_ (.Y(_0008_),
    .A(net605));
 sg13g2_xnor2_1 _2071_ (.Y(_1208_),
    .A(net431),
    .B(net630));
 sg13g2_nand2b_1 _2072_ (.Y(_1209_),
    .B(\modem.uart.rxHdlc.canInhibit ),
    .A_N(_0085_));
 sg13g2_nor4_2 _2073_ (.A(_1007_),
    .B(\modem.uart.rxHdlc.oneBitCount[1] ),
    .C(_1208_),
    .Y(_1210_),
    .D(_1209_));
 sg13g2_nand2_1 _2074_ (.Y(_1211_),
    .A(net685),
    .B(\modem.uart.rxHdlc.fsmHdlcRx_bit[1] ));
 sg13g2_nor2_2 _2075_ (.A(net854),
    .B(_1211_),
    .Y(_1212_));
 sg13g2_or2_1 _2076_ (.X(_1213_),
    .B(_1212_),
    .A(_1210_));
 sg13g2_nand2_1 _2077_ (.Y(_1214_),
    .A(\modem.uart.rxHdlc.oneBitCount[0] ),
    .B(\modem.uart.rxHdlc.oneBitCount[1] ));
 sg13g2_nor2_1 _2078_ (.A(net876),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_or2_1 _2079_ (.X(_1216_),
    .B(_1214_),
    .A(_0085_));
 sg13g2_nand2_1 _2080_ (.Y(_1217_),
    .A(net431),
    .B(net367));
 sg13g2_nand2_1 _2081_ (.Y(_1218_),
    .A(net432),
    .B(_1195_));
 sg13g2_nand3_1 _2082_ (.B(_1195_),
    .C(_1216_),
    .A(net431),
    .Y(_1219_));
 sg13g2_o21ai_1 _2083_ (.B1(_1195_),
    .Y(_1220_),
    .A1(_0971_),
    .A2(_1216_));
 sg13g2_a21oi_1 _2084_ (.A1(_1195_),
    .A2(_1210_),
    .Y(_1221_),
    .B1(_1204_));
 sg13g2_o21ai_1 _2085_ (.B1(_1221_),
    .Y(_1222_),
    .A1(_1213_),
    .A2(_1220_));
 sg13g2_nand2_1 _2086_ (.Y(_1223_),
    .A(net676),
    .B(_1212_));
 sg13g2_inv_1 _2087_ (.Y(_1224_),
    .A(_1223_));
 sg13g2_nand3_1 _2088_ (.B(net697),
    .C(\modem.uart.rxHdlc.oneBitCount[1] ),
    .A(_1007_),
    .Y(_1225_));
 sg13g2_inv_1 _2089_ (.Y(_1226_),
    .A(_1225_));
 sg13g2_nor3_2 _2090_ (.A(_1210_),
    .B(_1223_),
    .C(_1226_),
    .Y(_1227_));
 sg13g2_nor2_2 _2091_ (.A(net431),
    .B(_1225_),
    .Y(_1228_));
 sg13g2_nand3_1 _2092_ (.B(_1032_),
    .C(_1228_),
    .A(net799),
    .Y(_1229_));
 sg13g2_nand3_1 _2093_ (.B(_0067_),
    .C(_1195_),
    .A(_0971_),
    .Y(_1230_));
 sg13g2_o21ai_1 _2094_ (.B1(_1230_),
    .Y(_1231_),
    .A1(\modem.uart.rxHdlc.io_valid ),
    .A2(_1219_));
 sg13g2_a22oi_1 _2095_ (.Y(_1232_),
    .B1(_1227_),
    .B2(_1231_),
    .A2(_1222_),
    .A1(net676));
 sg13g2_o21ai_1 _2096_ (.B1(_1232_),
    .Y(_0000_),
    .A1(net406),
    .A2(net800));
 sg13g2_nor2_1 _2097_ (.A(net658),
    .B(_1173_),
    .Y(_1233_));
 sg13g2_nand2_2 _2098_ (.Y(_1234_),
    .A(\modem.uart.rxUart.bitId[0] ),
    .B(\modem.uart.rxUart.bitId[1] ));
 sg13g2_nor2_1 _2099_ (.A(net812),
    .B(_1234_),
    .Y(_1235_));
 sg13g2_a21oi_1 _2100_ (.A1(net807),
    .A2(_1235_),
    .Y(_1236_),
    .B1(_1174_));
 sg13g2_nor3_1 _2101_ (.A(net440),
    .B(_1233_),
    .C(_1236_),
    .Y(_0006_));
 sg13g2_nor2_1 _2102_ (.A(net408),
    .B(_1174_),
    .Y(_1237_));
 sg13g2_nand3_1 _2103_ (.B(net678),
    .C(net364),
    .A(net443),
    .Y(_1238_));
 sg13g2_a22oi_1 _2104_ (.Y(_1239_),
    .B1(_1237_),
    .B2(net658),
    .A2(net678),
    .A1(net443));
 sg13g2_o21ai_1 _2105_ (.B1(_1145_),
    .Y(_1240_),
    .A1(_1162_),
    .A2(_1239_));
 sg13g2_nand2b_1 _2106_ (.Y(_0005_),
    .B(net679),
    .A_N(_1240_));
 sg13g2_nand2_1 _2107_ (.Y(_1241_),
    .A(net505),
    .B(_1163_));
 sg13g2_nand2_1 _2108_ (.Y(_1242_),
    .A(\modem.uart.rxUart.fsmUartRx_stateReg[5] ),
    .B(_1237_));
 sg13g2_a21oi_1 _2109_ (.A1(net419),
    .A2(net505),
    .Y(_1243_),
    .B1(_1242_));
 sg13g2_and2_1 _2110_ (.A(_1241_),
    .B(_1243_),
    .X(_1244_));
 sg13g2_a21oi_1 _2111_ (.A1(net678),
    .A2(_1167_),
    .Y(_1245_),
    .B1(net892));
 sg13g2_nor3_1 _2112_ (.A(net440),
    .B(_1168_),
    .C(_1245_),
    .Y(_1246_));
 sg13g2_and3_1 _2113_ (.X(_0243_),
    .A(net658),
    .B(_1162_),
    .C(_1237_));
 sg13g2_or3_1 _2114_ (.A(_1244_),
    .B(_1246_),
    .C(_0243_),
    .X(_0004_));
 sg13g2_nor3_1 _2115_ (.A(net408),
    .B(_1174_),
    .C(_1235_),
    .Y(_1247_));
 sg13g2_o21ai_1 _2116_ (.B1(\modem.uart.rxUart.fsmUartRx_stateReg[1] ),
    .Y(_1248_),
    .A1(_1175_),
    .A2(_1247_));
 sg13g2_o21ai_1 _2117_ (.B1(_1248_),
    .Y(_0003_),
    .A1(_1241_),
    .A2(_1242_));
 sg13g2_a21oi_1 _2118_ (.A1(_1224_),
    .A2(_1226_),
    .Y(_1249_),
    .B1(net701));
 sg13g2_a21oi_1 _2119_ (.A1(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[1] ),
    .A2(_1032_),
    .Y(_1250_),
    .B1(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[2] ));
 sg13g2_o21ai_1 _2120_ (.B1(_1215_),
    .Y(_1251_),
    .A1(net432),
    .A2(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[2] ));
 sg13g2_nor2_1 _2121_ (.A(_1250_),
    .B(_1251_),
    .Y(_1252_));
 sg13g2_a22oi_1 _2122_ (.Y(_1253_),
    .B1(_1252_),
    .B2(_1195_),
    .A2(_1204_),
    .A1(net701));
 sg13g2_o21ai_1 _2123_ (.B1(_1253_),
    .Y(_0002_),
    .A1(_1218_),
    .A2(_1249_));
 sg13g2_nand2_1 _2124_ (.Y(_1254_),
    .A(\modem.dcdHistory_7 ),
    .B(\modem.dcdHistory_6 ));
 sg13g2_or2_1 _2125_ (.X(_1255_),
    .B(\modem.dcdHistory_6 ),
    .A(\modem.dcdHistory_7 ));
 sg13g2_xnor2_1 _2126_ (.Y(_1256_),
    .A(_0027_),
    .B(net360));
 sg13g2_nor2_1 _2127_ (.A(\modem.dcdHistory_1 ),
    .B(net360),
    .Y(_1257_));
 sg13g2_a22oi_1 _2128_ (.Y(_1258_),
    .B1(_1257_),
    .B2(\modem.dcdHistory_2 ),
    .A2(_1256_),
    .A1(_0028_));
 sg13g2_and2_1 _2129_ (.A(_0028_),
    .B(_1257_),
    .X(_1259_));
 sg13g2_nand2_1 _2130_ (.Y(_1260_),
    .A(_0028_),
    .B(_1257_));
 sg13g2_nor3_1 _2131_ (.A(_0947_),
    .B(\modem.dcdHistory_2 ),
    .C(net369),
    .Y(_1261_));
 sg13g2_a21o_1 _2132_ (.A2(_1256_),
    .A1(\modem.dcdHistory_2 ),
    .B1(_1261_),
    .X(_1262_));
 sg13g2_o21ai_1 _2133_ (.B1(_1258_),
    .Y(_1263_),
    .A1(_1259_),
    .A2(_1262_));
 sg13g2_nand2_1 _2134_ (.Y(_1264_),
    .A(\modem.dcdHistory_4 ),
    .B(\modem.dcdHistory_3 ));
 sg13g2_a21oi_1 _2135_ (.A1(\modem.dcdHistory_4 ),
    .A2(\modem.dcdHistory_3 ),
    .Y(_1265_),
    .B1(_0026_));
 sg13g2_nand3_1 _2136_ (.B(_0949_),
    .C(_0026_),
    .A(_0946_),
    .Y(_1266_));
 sg13g2_o21ai_1 _2137_ (.B1(\modem.dcdHistory_5 ),
    .Y(_1267_),
    .A1(\modem.dcdHistory_4 ),
    .A2(\modem.dcdHistory_3 ));
 sg13g2_nand3_1 _2138_ (.B(_1266_),
    .C(_1267_),
    .A(_1264_),
    .Y(_1268_));
 sg13g2_o21ai_1 _2139_ (.B1(_1268_),
    .Y(_1269_),
    .A1(_0945_),
    .A2(_1265_));
 sg13g2_and2_1 _2140_ (.A(_1263_),
    .B(_1269_),
    .X(_1270_));
 sg13g2_a21oi_1 _2141_ (.A1(_1258_),
    .A2(_1260_),
    .Y(_1271_),
    .B1(_1262_));
 sg13g2_a21o_1 _2142_ (.A2(_1264_),
    .A1(_0026_),
    .B1(\modem.dcdHistory_5 ),
    .X(_1272_));
 sg13g2_and2_1 _2143_ (.A(_1267_),
    .B(_1272_),
    .X(_1273_));
 sg13g2_and3_1 _2144_ (.X(_1274_),
    .A(_1254_),
    .B(_1271_),
    .C(_1273_));
 sg13g2_nor2_1 _2145_ (.A(_1271_),
    .B(_1273_),
    .Y(_1275_));
 sg13g2_a21oi_1 _2146_ (.A1(_1271_),
    .A2(_1273_),
    .Y(_1276_),
    .B1(_1254_));
 sg13g2_nor2_1 _2147_ (.A(_1275_),
    .B(_1276_),
    .Y(_1277_));
 sg13g2_nor2_1 _2148_ (.A(_1263_),
    .B(_1269_),
    .Y(_1278_));
 sg13g2_a22oi_1 _2149_ (.Y(_1279_),
    .B1(_1277_),
    .B2(_1278_),
    .A2(_1274_),
    .A1(_1270_));
 sg13g2_a21oi_1 _2150_ (.A1(_1254_),
    .A2(_1255_),
    .Y(_1280_),
    .B1(_1279_));
 sg13g2_nand2_1 _2151_ (.Y(_1281_),
    .A(_1255_),
    .B(_1275_));
 sg13g2_a21oi_1 _2152_ (.A1(_1254_),
    .A2(_1278_),
    .Y(_1282_),
    .B1(_1281_));
 sg13g2_nor2_1 _2153_ (.A(_1270_),
    .B(_1274_),
    .Y(_1283_));
 sg13g2_a21oi_1 _2154_ (.A1(_1270_),
    .A2(_1277_),
    .Y(_1284_),
    .B1(_1283_));
 sg13g2_nor3_1 _2155_ (.A(_1280_),
    .B(_1282_),
    .C(_1284_),
    .Y(\modem.dcd ));
 sg13g2_xor2_1 _2156_ (.B(net364),
    .A(net858),
    .X(_1285_));
 sg13g2_nor2_1 _2157_ (.A(_1170_),
    .B(_1285_),
    .Y(_0023_));
 sg13g2_o21ai_1 _2158_ (.B1(net751),
    .Y(_1286_),
    .A1(\modem.uart.rxUart.sampleTimer_counter[0] ),
    .A2(net364));
 sg13g2_nand3_1 _2159_ (.B(_1172_),
    .C(net752),
    .A(_1169_),
    .Y(_0024_));
 sg13g2_xor2_1 _2160_ (.B(_1171_),
    .A(net500),
    .X(_0326_));
 sg13g2_nor2_1 _2161_ (.A(_1170_),
    .B(net501),
    .Y(_0025_));
 sg13g2_or2_1 _2162_ (.X(_0327_),
    .B(_1210_),
    .A(net368));
 sg13g2_o21ai_1 _2163_ (.B1(_0327_),
    .Y(_0328_),
    .A1(net565),
    .A2(net366));
 sg13g2_o21ai_1 _2164_ (.B1(_0328_),
    .Y(_0329_),
    .A1(\modem.uart.rxHdlc.canInhibit ),
    .A2(_1217_));
 sg13g2_inv_1 _2165_ (.Y(_0022_),
    .A(net566));
 sg13g2_nor2_2 _2166_ (.A(net413),
    .B(net411),
    .Y(_0330_));
 sg13g2_and2_1 _2167_ (.A(net414),
    .B(net411),
    .X(_0331_));
 sg13g2_nand2b_2 _2168_ (.Y(_0332_),
    .B(net412),
    .A_N(net414));
 sg13g2_nor2b_2 _2169_ (.A(net411),
    .B_N(net414),
    .Y(_0333_));
 sg13g2_nand2_1 _2170_ (.Y(_0334_),
    .A(net414),
    .B(_1013_));
 sg13g2_mux4_1 _2171_ (.S0(net411),
    .A0(\modem.control.scrambler_1.io_vecOut[4] ),
    .A1(_1014_),
    .A2(net417),
    .A3(\modem.control.rxAddr[0] ),
    .S1(net413),
    .X(uio_out[2]));
 sg13g2_o21ai_1 _2172_ (.B1(net411),
    .Y(_0335_),
    .A1(net413),
    .A2(_1015_));
 sg13g2_a22oi_1 _2173_ (.Y(_0336_),
    .B1(_0333_),
    .B2(\modem.control._zz_txClockInternalFallStb ),
    .A2(_0330_),
    .A1(\modem.control.scrambler_1.io_vecOut[5] ));
 sg13g2_a22oi_1 _2174_ (.Y(uio_out[3]),
    .B1(_0335_),
    .B2(_0336_),
    .A2(_0331_),
    .A1(_0967_));
 sg13g2_nand2_1 _2175_ (.Y(_0337_),
    .A(\modem.control.scrambler_1.io_vecOut[6] ),
    .B(_0330_));
 sg13g2_nand2_1 _2176_ (.Y(_0338_),
    .A(_0965_),
    .B(_1013_));
 sg13g2_nor2_1 _2177_ (.A(_0033_),
    .B(_0332_),
    .Y(_0339_));
 sg13g2_a21oi_1 _2178_ (.A1(net413),
    .A2(_0338_),
    .Y(_0340_),
    .B1(_0339_));
 sg13g2_a22oi_1 _2179_ (.Y(uio_out[4]),
    .B1(_0337_),
    .B2(_0340_),
    .A2(_0331_),
    .A1(_0944_));
 sg13g2_o21ai_1 _2180_ (.B1(net413),
    .Y(_0341_),
    .A1(\modem.control.scrambler_1.io_vecOut[1] ),
    .A2(net411));
 sg13g2_nor2_1 _2181_ (.A(_0032_),
    .B(_0332_),
    .Y(_0342_));
 sg13g2_a21oi_1 _2182_ (.A1(\modem.control.scrambler_1.io_vecOut[7] ),
    .A2(_0330_),
    .Y(_0343_),
    .B1(_0342_));
 sg13g2_a22oi_1 _2183_ (.Y(uio_out[5]),
    .B1(_0341_),
    .B2(_0343_),
    .A2(_0331_),
    .A1(_0966_));
 sg13g2_nand2_1 _2184_ (.Y(_0344_),
    .A(net411),
    .B(_0031_));
 sg13g2_a21oi_1 _2185_ (.A1(_0338_),
    .A2(_0344_),
    .Y(_0345_),
    .B1(net413));
 sg13g2_a221oi_1 _2186_ (.B2(_0963_),
    .C1(_0345_),
    .B1(_0333_),
    .A1(_0970_),
    .Y(uio_out[6]),
    .A2(_0331_));
 sg13g2_o21ai_1 _2187_ (.B1(net411),
    .Y(_0346_),
    .A1(\modem.control.rxAddr[11] ),
    .A2(net413));
 sg13g2_a22oi_1 _2188_ (.Y(_0347_),
    .B1(_0330_),
    .B2(\modem.control.scrambler_1.io_vecOut[1] ),
    .A2(net413),
    .A1(\modem.control.scrambler_1.io_vecOut[3] ));
 sg13g2_a22oi_1 _2189_ (.Y(uio_out[7]),
    .B1(_0346_),
    .B2(_0347_),
    .A2(_0331_),
    .A1(_0969_));
 sg13g2_nor2b_2 _2190_ (.A(\modem.uart.txFifo.nextOut[0] ),
    .B_N(net420),
    .Y(_0348_));
 sg13g2_nor2b_2 _2191_ (.A(net420),
    .B_N(\modem.uart.txFifo.nextOut[0] ),
    .Y(_0349_));
 sg13g2_nor2_2 _2192_ (.A(net420),
    .B(\modem.uart.txFifo.nextOut[0] ),
    .Y(_0350_));
 sg13g2_nand2_1 _2193_ (.Y(_0351_),
    .A(_1006_),
    .B(\modem.uart.tx.bitId[1] ));
 sg13g2_a22oi_1 _2194_ (.Y(_0352_),
    .B1(_0350_),
    .B2(\modem.uart.txFifo.fifo_0[0] ),
    .A2(_0349_),
    .A1(\modem.uart.txFifo.fifo_1[0] ));
 sg13g2_a21oi_1 _2195_ (.A1(\modem.uart.txFifo.fifo_2[0] ),
    .A2(_0348_),
    .Y(_0353_),
    .B1(net438));
 sg13g2_a22oi_1 _2196_ (.Y(_0354_),
    .B1(_0349_),
    .B2(\modem.uart.txFifo.fifo_1[1] ),
    .A2(_0348_),
    .A1(\modem.uart.txFifo.fifo_2[1] ));
 sg13g2_a21oi_1 _2197_ (.A1(\modem.uart.txFifo.fifo_0[1] ),
    .A2(_0350_),
    .Y(_0355_),
    .B1(_1006_));
 sg13g2_a221oi_1 _2198_ (.B2(_0355_),
    .C1(net437),
    .B1(_0354_),
    .A1(_0352_),
    .Y(_0356_),
    .A2(_0353_));
 sg13g2_a22oi_1 _2199_ (.Y(_0357_),
    .B1(_0349_),
    .B2(\modem.uart.txFifo.fifo_1[3] ),
    .A2(_0348_),
    .A1(\modem.uart.txFifo.fifo_2[3] ));
 sg13g2_a21oi_1 _2200_ (.A1(\modem.uart.txFifo.fifo_0[3] ),
    .A2(_0350_),
    .Y(_0358_),
    .B1(_1006_));
 sg13g2_a22oi_1 _2201_ (.Y(_0359_),
    .B1(_0350_),
    .B2(\modem.uart.txFifo.fifo_0[2] ),
    .A2(_0349_),
    .A1(\modem.uart.txFifo.fifo_1[2] ));
 sg13g2_a21oi_1 _2202_ (.A1(\modem.uart.txFifo.fifo_2[2] ),
    .A2(_0348_),
    .Y(_0360_),
    .B1(net438));
 sg13g2_a22oi_1 _2203_ (.Y(_0361_),
    .B1(_0359_),
    .B2(_0360_),
    .A2(_0358_),
    .A1(_0357_));
 sg13g2_a21oi_1 _2204_ (.A1(net437),
    .A2(_0361_),
    .Y(_0362_),
    .B1(_0356_));
 sg13g2_nand2_1 _2205_ (.Y(_0363_),
    .A(net420),
    .B(\modem.uart.txFifo.nextOut[0] ));
 sg13g2_a22oi_1 _2206_ (.Y(_0364_),
    .B1(_0350_),
    .B2(\modem.uart.txFifo.fifo_0[5] ),
    .A2(_0349_),
    .A1(\modem.uart.txFifo.fifo_1[5] ));
 sg13g2_a21oi_1 _2207_ (.A1(\modem.uart.txFifo.fifo_2[5] ),
    .A2(_0348_),
    .Y(_0365_),
    .B1(_1006_));
 sg13g2_a22oi_1 _2208_ (.Y(_0366_),
    .B1(\modem.uart.txFifo.fifo_1[4] ),
    .B2(_0349_),
    .A2(\modem.uart.txFifo.fifo_2[4] ),
    .A1(net420));
 sg13g2_a21oi_1 _2209_ (.A1(\modem.uart.txFifo.fifo_0[4] ),
    .A2(_0350_),
    .Y(_0367_),
    .B1(net438));
 sg13g2_a221oi_1 _2210_ (.B2(_0367_),
    .C1(net437),
    .B1(_0366_),
    .A1(_0364_),
    .Y(_0368_),
    .A2(_0365_));
 sg13g2_a21oi_1 _2211_ (.A1(\modem.uart.txFifo.fifo_2[6] ),
    .A2(_0348_),
    .Y(_0369_),
    .B1(net438));
 sg13g2_a22oi_1 _2212_ (.Y(_0370_),
    .B1(_0350_),
    .B2(\modem.uart.txFifo.fifo_0[6] ),
    .A2(_0349_),
    .A1(\modem.uart.txFifo.fifo_1[6] ));
 sg13g2_nand2_1 _2213_ (.Y(_0371_),
    .A(\modem.uart.txFifo.fifo_1[7] ),
    .B(_0349_));
 sg13g2_a22oi_1 _2214_ (.Y(_0372_),
    .B1(_0350_),
    .B2(\modem.uart.txFifo.fifo_0[7] ),
    .A2(\modem.uart.txFifo.fifo_2[7] ),
    .A1(net420));
 sg13g2_nand3_1 _2215_ (.B(_0371_),
    .C(_0372_),
    .A(net438),
    .Y(_0373_));
 sg13g2_nand2_1 _2216_ (.Y(_0374_),
    .A(net437),
    .B(_0373_));
 sg13g2_a21oi_1 _2217_ (.A1(_0369_),
    .A2(_0370_),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_nor3_1 _2218_ (.A(_1019_),
    .B(_0368_),
    .C(_0375_),
    .Y(_0376_));
 sg13g2_a221oi_1 _2219_ (.B2(_0362_),
    .C1(_0376_),
    .B1(_1019_),
    .A1(\modem.uart.txFifo.nextOut[1] ),
    .Y(_0377_),
    .A2(\modem.uart.txFifo.nextOut[0] ));
 sg13g2_a21oi_1 _2220_ (.A1(net438),
    .A2(\modem.uart.txFifo.fifo_3[1] ),
    .Y(_0378_),
    .B1(net437));
 sg13g2_o21ai_1 _2221_ (.B1(_0378_),
    .Y(_0379_),
    .A1(\modem.uart.tx.bitId[0] ),
    .A2(_1018_));
 sg13g2_nor2_1 _2222_ (.A(\modem.uart.txFifo.fifo_3[3] ),
    .B(_1196_),
    .Y(_0380_));
 sg13g2_o21ai_1 _2223_ (.B1(_1019_),
    .Y(_0381_),
    .A1(\modem.uart.txFifo.fifo_3[2] ),
    .A2(_0351_));
 sg13g2_nor2_1 _2224_ (.A(_0380_),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_nand2_1 _2225_ (.Y(_0383_),
    .A(\modem.uart.tx.bitId[0] ),
    .B(\modem.uart.txFifo.fifo_3[5] ));
 sg13g2_a21oi_1 _2226_ (.A1(_1006_),
    .A2(\modem.uart.txFifo.fifo_3[4] ),
    .Y(_0384_),
    .B1(net437));
 sg13g2_or2_1 _2227_ (.X(_0385_),
    .B(_1196_),
    .A(\modem.uart.txFifo.fifo_3[7] ));
 sg13g2_o21ai_1 _2228_ (.B1(\modem.uart.tx.bitId[2] ),
    .Y(_0386_),
    .A1(\modem.uart.txFifo.fifo_3[6] ),
    .A2(_0351_));
 sg13g2_a21oi_1 _2229_ (.A1(_0383_),
    .A2(_0384_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_a22oi_1 _2230_ (.Y(_0388_),
    .B1(_0385_),
    .B2(_0387_),
    .A2(_0382_),
    .A1(_0379_));
 sg13g2_o21ai_1 _2231_ (.B1(\modem.uart.tx.fsmUartTx_stateReg[4] ),
    .Y(_0389_),
    .A1(_0363_),
    .A2(_0388_));
 sg13g2_or2_1 _2232_ (.X(_0390_),
    .B(_0078_),
    .A(\modem.uart.tx.fsmUartTx_stateReg[4] ));
 sg13g2_o21ai_1 _2233_ (.B1(_0390_),
    .Y(_0391_),
    .A1(_0377_),
    .A2(_0389_));
 sg13g2_inv_1 _2234_ (.Y(\modem.uart.io_uartTxOut ),
    .A(_0391_));
 sg13g2_nor3_1 _2235_ (.A(_1107_),
    .B(_1138_),
    .C(_1143_),
    .Y(_0392_));
 sg13g2_a21o_1 _2236_ (.A2(_1043_),
    .A1(net755),
    .B1(_0392_),
    .X(_0018_));
 sg13g2_nand2b_1 _2237_ (.Y(_0393_),
    .B(_1177_),
    .A_N(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[6] ));
 sg13g2_and2_1 _2238_ (.A(_1042_),
    .B(_0393_),
    .X(_0394_));
 sg13g2_a21oi_1 _2239_ (.A1(net880),
    .A2(net401),
    .Y(_0395_),
    .B1(_0394_));
 sg13g2_o21ai_1 _2240_ (.B1(_1045_),
    .Y(_0396_),
    .A1(net880),
    .A2(net705));
 sg13g2_or2_1 _2241_ (.X(_0397_),
    .B(_0396_),
    .A(_1131_));
 sg13g2_o21ai_1 _2242_ (.B1(_0397_),
    .Y(_0017_),
    .A1(net405),
    .A2(_0395_));
 sg13g2_nand2_1 _2243_ (.Y(_0398_),
    .A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[2] ),
    .B(_1045_));
 sg13g2_nand3_1 _2244_ (.B(net442),
    .C(net401),
    .A(net742),
    .Y(_0399_));
 sg13g2_o21ai_1 _2245_ (.B1(_0399_),
    .Y(_0016_),
    .A1(_1126_),
    .A2(_0398_));
 sg13g2_nor2b_1 _2246_ (.A(_1189_),
    .B_N(_1187_),
    .Y(_0400_));
 sg13g2_a21o_1 _2247_ (.A2(_1191_),
    .A1(net884),
    .B1(_0400_),
    .X(_0015_));
 sg13g2_nand2_1 _2248_ (.Y(_0401_),
    .A(net444),
    .B(_1194_));
 sg13g2_and2_1 _2249_ (.A(net444),
    .B(net518),
    .X(_0402_));
 sg13g2_o21ai_1 _2250_ (.B1(_1145_),
    .Y(_0403_),
    .A1(\modem.uart.txCommandDecoder.io_valid ),
    .A2(_1188_));
 sg13g2_a21oi_1 _2251_ (.A1(_1190_),
    .A2(_0402_),
    .Y(_0404_),
    .B1(net861));
 sg13g2_o21ai_1 _2252_ (.B1(_0404_),
    .Y(_0014_),
    .A1(net785),
    .A2(_0401_));
 sg13g2_nor2_1 _2253_ (.A(_0067_),
    .B(_1218_),
    .Y(_0405_));
 sg13g2_nor2_1 _2254_ (.A(_1004_),
    .B(_1228_),
    .Y(_0406_));
 sg13g2_a22oi_1 _2255_ (.Y(_0407_),
    .B1(_0406_),
    .B2(_1195_),
    .A2(_0405_),
    .A1(_1227_));
 sg13g2_a221oi_1 _2256_ (.B2(_1224_),
    .C1(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[3] ),
    .B1(_1228_),
    .A1(\modem.uart.rxHdlc.io_valid ),
    .Y(_0408_),
    .A2(_1227_));
 sg13g2_nor4_1 _2257_ (.A(net432),
    .B(net408),
    .C(_1031_),
    .D(_0408_),
    .Y(_0409_));
 sg13g2_a221oi_1 _2258_ (.B2(net799),
    .C1(_0409_),
    .B1(_1204_),
    .A1(net445),
    .Y(_0410_),
    .A2(net772));
 sg13g2_o21ai_1 _2259_ (.B1(_0410_),
    .Y(_0001_),
    .A1(_1215_),
    .A2(_0407_));
 sg13g2_nand3b_1 _2260_ (.B(_1132_),
    .C(net880),
    .Y(_0411_),
    .A_N(_1044_));
 sg13g2_a21oi_1 _2261_ (.A1(net705),
    .A2(_1140_),
    .Y(_0412_),
    .B1(_0394_));
 sg13g2_nand2_1 _2262_ (.Y(\modem.uart.txPacketUpper.io_ready ),
    .A(_0411_),
    .B(_0412_));
 sg13g2_xor2_1 _2263_ (.B(\modem.control.scrambler_1.io_dataIn ),
    .A(\modem.control.scrambler_1.io_vecOut[11] ),
    .X(_0413_));
 sg13g2_o21ai_1 _2264_ (.B1(net446),
    .Y(_0414_),
    .A1(net332),
    .A2(_0413_));
 sg13g2_a21oi_1 _2265_ (.A1(net332),
    .A2(_0413_),
    .Y(_0086_),
    .B1(_0414_));
 sg13g2_a21oi_1 _2266_ (.A1(net367),
    .A2(_1228_),
    .Y(_0415_),
    .B1(_1004_));
 sg13g2_nor3_2 _2267_ (.A(_1210_),
    .B(_1250_),
    .C(_0415_),
    .Y(_0416_));
 sg13g2_nor3_1 _2268_ (.A(_0997_),
    .B(net778),
    .C(_1212_),
    .Y(_0417_));
 sg13g2_mux2_1 _2269_ (.A0(net685),
    .A1(_0417_),
    .S(_0416_),
    .X(_0087_));
 sg13g2_xnor2_1 _2270_ (.Y(_0418_),
    .A(\modem.uart.rxHdlc.fsmHdlcRx_bit[0] ),
    .B(\modem.uart.rxHdlc.fsmHdlcRx_bit[1] ));
 sg13g2_nor2_1 _2271_ (.A(net778),
    .B(_0418_),
    .Y(_0419_));
 sg13g2_mux2_1 _2272_ (.A0(net849),
    .A1(_0419_),
    .S(_0416_),
    .X(_0088_));
 sg13g2_nor2b_1 _2273_ (.A(_1211_),
    .B_N(_0416_),
    .Y(_0420_));
 sg13g2_o21ai_1 _2274_ (.B1(_0416_),
    .Y(_0421_),
    .A1(net778),
    .A2(_1212_));
 sg13g2_o21ai_1 _2275_ (.B1(net779),
    .Y(_0422_),
    .A1(net689),
    .A2(_0420_));
 sg13g2_a21oi_1 _2276_ (.A1(net689),
    .A2(_0420_),
    .Y(_0089_),
    .B1(net780));
 sg13g2_nand2_1 _2277_ (.Y(_0423_),
    .A(net495),
    .B(net365));
 sg13g2_o21ai_1 _2278_ (.B1(_0423_),
    .Y(_0090_),
    .A1(_0998_),
    .A2(net365));
 sg13g2_mux2_1 _2279_ (.A0(net495),
    .A1(net688),
    .S(net365),
    .X(_0091_));
 sg13g2_a221oi_1 _2280_ (.B2(\modem.uart.tx.fsmUartTx_stateReg[4] ),
    .C1(net368),
    .B1(_1197_),
    .A1(_1002_),
    .Y(_0424_),
    .A2(_0079_));
 sg13g2_nand3_1 _2281_ (.B(net310),
    .C(_0424_),
    .A(\modem.uart.tx.fsmUartTx_stateReg[4] ),
    .Y(_0425_));
 sg13g2_o21ai_1 _2282_ (.B1(net311),
    .Y(_0092_),
    .A1(_1006_),
    .A2(_0424_));
 sg13g2_nand2_1 _2283_ (.Y(_0426_),
    .A(\modem.uart.tx.fsmUartTx_stateReg[4] ),
    .B(_1196_));
 sg13g2_and2_1 _2284_ (.A(_0424_),
    .B(_0426_),
    .X(_0427_));
 sg13g2_a21oi_1 _2285_ (.A1(net438),
    .A2(_0424_),
    .Y(_0428_),
    .B1(net437));
 sg13g2_nor2_1 _2286_ (.A(_0427_),
    .B(net891),
    .Y(_0093_));
 sg13g2_nor2_1 _2287_ (.A(net870),
    .B(_1196_),
    .Y(_0429_));
 sg13g2_nand3_1 _2288_ (.B(_0424_),
    .C(_0429_),
    .A(\modem.uart.tx.fsmUartTx_stateReg[4] ),
    .Y(_0430_));
 sg13g2_o21ai_1 _2289_ (.B1(net871),
    .Y(_0094_),
    .A1(_1019_),
    .A2(_0427_));
 sg13g2_nor2_2 _2290_ (.A(net864),
    .B(_1174_),
    .Y(_0431_));
 sg13g2_nor3_2 _2291_ (.A(\modem.uart.rxUart.bitId[0] ),
    .B(\modem.uart.rxUart.bitId[1] ),
    .C(\modem.uart.rxUart.bitId[2] ),
    .Y(_0432_));
 sg13g2_nand2_1 _2292_ (.Y(_0433_),
    .A(_0431_),
    .B(_0432_));
 sg13g2_nor2_1 _2293_ (.A(_1162_),
    .B(_0433_),
    .Y(_0434_));
 sg13g2_a21oi_1 _2294_ (.A1(_0993_),
    .A2(_0433_),
    .Y(_0095_),
    .B1(_0434_));
 sg13g2_a21oi_1 _2295_ (.A1(_1005_),
    .A2(_1020_),
    .Y(_0435_),
    .B1(_1021_));
 sg13g2_nor2_1 _2296_ (.A(_0432_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_nand2_2 _2297_ (.Y(_0437_),
    .A(_0431_),
    .B(_0436_));
 sg13g2_nand2_1 _2298_ (.Y(_0438_),
    .A(\modem.uart.rxUart.bitId[0] ),
    .B(_1020_));
 sg13g2_nand2_1 _2299_ (.Y(_0439_),
    .A(_1005_),
    .B(\modem.uart.rxUart.bitId[1] ));
 sg13g2_nand2_1 _2300_ (.Y(_0440_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_nand3b_1 _2301_ (.B(_1162_),
    .C(_0440_),
    .Y(_0441_),
    .A_N(net497));
 sg13g2_o21ai_1 _2302_ (.B1(net843),
    .Y(_0442_),
    .A1(_0437_),
    .A2(_0438_));
 sg13g2_o21ai_1 _2303_ (.B1(net844),
    .Y(_0096_),
    .A1(_0437_),
    .A2(_0441_));
 sg13g2_nor2_1 _2304_ (.A(_0437_),
    .B(_0439_),
    .Y(_0443_));
 sg13g2_nor2_1 _2305_ (.A(net720),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_a21oi_1 _2306_ (.A1(_1163_),
    .A2(_0443_),
    .Y(_0097_),
    .B1(net721));
 sg13g2_or4_1 _2307_ (.A(net497),
    .B(_1163_),
    .C(_0432_),
    .D(_0440_),
    .X(_0445_));
 sg13g2_nor2_1 _2308_ (.A(\modem.uart.rxUart.bitId[2] ),
    .B(_1234_),
    .Y(_0446_));
 sg13g2_a21o_1 _2309_ (.A2(_0446_),
    .A1(_0431_),
    .B1(net410),
    .X(_0447_));
 sg13g2_o21ai_1 _2310_ (.B1(_0447_),
    .Y(_0098_),
    .A1(_0437_),
    .A2(_0445_));
 sg13g2_nor2_1 _2311_ (.A(_1021_),
    .B(_0437_),
    .Y(_0448_));
 sg13g2_nor2_1 _2312_ (.A(net769),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_a21oi_1 _2313_ (.A1(_1163_),
    .A2(_0448_),
    .Y(_0099_),
    .B1(net770));
 sg13g2_nand2b_2 _2314_ (.Y(_0450_),
    .B(_0431_),
    .A_N(_0436_));
 sg13g2_o21ai_1 _2315_ (.B1(net757),
    .Y(_0451_),
    .A1(_0438_),
    .A2(_0450_));
 sg13g2_o21ai_1 _2316_ (.B1(net758),
    .Y(_0100_),
    .A1(_0441_),
    .A2(_0450_));
 sg13g2_nor2_1 _2317_ (.A(_0439_),
    .B(_0450_),
    .Y(_0452_));
 sg13g2_nor2_1 _2318_ (.A(net728),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_a21oi_1 _2319_ (.A1(_1163_),
    .A2(_0452_),
    .Y(_0101_),
    .B1(net729));
 sg13g2_o21ai_1 _2320_ (.B1(net715),
    .Y(_0454_),
    .A1(_1234_),
    .A2(_0450_));
 sg13g2_o21ai_1 _2321_ (.B1(net716),
    .Y(_0102_),
    .A1(_0445_),
    .A2(_0450_));
 sg13g2_mux2_1 _2322_ (.A0(net761),
    .A1(\modem.uart.rxUart._zz_sampleValue_29 ),
    .S(net364),
    .X(_0103_));
 sg13g2_mux2_1 _2323_ (.A0(net836),
    .A1(net823),
    .S(net364),
    .X(_0104_));
 sg13g2_mux2_1 _2324_ (.A0(net823),
    .A1(net736),
    .S(net364),
    .X(_0105_));
 sg13g2_nor2_1 _2325_ (.A(net736),
    .B(net365),
    .Y(_0455_));
 sg13g2_a21oi_1 _2326_ (.A1(_0998_),
    .A2(net365),
    .Y(_0106_),
    .B1(_0455_));
 sg13g2_nor3_1 _2327_ (.A(_1223_),
    .B(_1228_),
    .C(_0327_),
    .Y(_0456_));
 sg13g2_nand2_2 _2328_ (.Y(_0457_),
    .A(net624),
    .B(_1201_));
 sg13g2_and2_1 _2329_ (.A(\modem.uart.rxHdlc.io_valid ),
    .B(_0457_),
    .X(_0458_));
 sg13g2_nand2_2 _2330_ (.Y(_0459_),
    .A(\modem.uart.rxHdlc.io_valid ),
    .B(_0457_));
 sg13g2_o21ai_1 _2331_ (.B1(_0459_),
    .Y(_0460_),
    .A1(\modem.uart.rxHdlc.io_valid ),
    .A2(_1225_));
 sg13g2_nor2_1 _2332_ (.A(net881),
    .B(_0457_),
    .Y(_0461_));
 sg13g2_o21ai_1 _2333_ (.B1(net445),
    .Y(_0462_),
    .A1(_0456_),
    .A2(_0461_));
 sg13g2_a21oi_1 _2334_ (.A1(_0456_),
    .A2(_0460_),
    .Y(_0107_),
    .B1(_0462_));
 sg13g2_o21ai_1 _2335_ (.B1(net443),
    .Y(_0463_),
    .A1(net418),
    .A2(\modem.uart.rxFifo.nextIn[0] ));
 sg13g2_a21oi_1 _2336_ (.A1(net418),
    .A2(_0996_),
    .Y(_0108_),
    .B1(_0463_));
 sg13g2_a21oi_1 _2337_ (.A1(net418),
    .A2(\modem.uart.rxFifo.nextIn[0] ),
    .Y(_0464_),
    .B1(net862));
 sg13g2_nand3_1 _2338_ (.B(net862),
    .C(\modem.uart.rxFifo.nextIn[0] ),
    .A(net418),
    .Y(_0465_));
 sg13g2_inv_1 _2339_ (.Y(_0466_),
    .A(_0465_));
 sg13g2_nor3_1 _2340_ (.A(net406),
    .B(net863),
    .C(_0466_),
    .Y(_0109_));
 sg13g2_xor2_1 _2341_ (.B(_0465_),
    .A(net872),
    .X(_0467_));
 sg13g2_nor2_1 _2342_ (.A(net406),
    .B(_0467_),
    .Y(_0110_));
 sg13g2_a21oi_1 _2343_ (.A1(_0411_),
    .A2(_0412_),
    .Y(_0468_),
    .B1(\modem.uart.uart_txPacketUpper_io_ready_regNext ));
 sg13g2_o21ai_1 _2344_ (.B1(net442),
    .Y(_0469_),
    .A1(\modem.uart.rxFifo.nextOut[0] ),
    .A2(net346));
 sg13g2_a21oi_1 _2345_ (.A1(_0994_),
    .A2(net346),
    .Y(_0111_),
    .B1(_0469_));
 sg13g2_a21oi_1 _2346_ (.A1(\modem.uart.rxFifo.nextOut[0] ),
    .A2(net346),
    .Y(_0470_),
    .B1(net833));
 sg13g2_a21oi_1 _2347_ (.A1(net396),
    .A2(net346),
    .Y(_0471_),
    .B1(net405));
 sg13g2_nor2b_1 _2348_ (.A(net834),
    .B_N(_0471_),
    .Y(_0112_));
 sg13g2_a21oi_1 _2349_ (.A1(net396),
    .A2(net346),
    .Y(_0472_),
    .B1(net435));
 sg13g2_a21oi_1 _2350_ (.A1(net388),
    .A2(net346),
    .Y(_0473_),
    .B1(net405));
 sg13g2_nor2b_1 _2351_ (.A(_0472_),
    .B_N(_0473_),
    .Y(_0113_));
 sg13g2_nand2_2 _2352_ (.Y(_0474_),
    .A(net418),
    .B(net441));
 sg13g2_nand2b_1 _2353_ (.Y(_0475_),
    .B(\modem.uart.rxFifo.nextIn[1] ),
    .A_N(\modem.uart.rxFifo.nextIn[0] ));
 sg13g2_nor3_2 _2354_ (.A(_0065_),
    .B(_0474_),
    .C(_0475_),
    .Y(_0476_));
 sg13g2_nor2_1 _2355_ (.A(net589),
    .B(net387),
    .Y(_0477_));
 sg13g2_a21oi_1 _2356_ (.A1(net409),
    .A2(net387),
    .Y(_0114_),
    .B1(_0477_));
 sg13g2_nor2_1 _2357_ (.A(net540),
    .B(net386),
    .Y(_0478_));
 sg13g2_a21oi_1 _2358_ (.A1(_0992_),
    .A2(net386),
    .Y(_0115_),
    .B1(_0478_));
 sg13g2_nor2_1 _2359_ (.A(net585),
    .B(net387),
    .Y(_0479_));
 sg13g2_a21oi_1 _2360_ (.A1(_0991_),
    .A2(net387),
    .Y(_0116_),
    .B1(_0479_));
 sg13g2_nor2_1 _2361_ (.A(net597),
    .B(net387),
    .Y(_0480_));
 sg13g2_a21oi_1 _2362_ (.A1(net410),
    .A2(net387),
    .Y(_0117_),
    .B1(_0480_));
 sg13g2_nor2_1 _2363_ (.A(net601),
    .B(net386),
    .Y(_0481_));
 sg13g2_a21oi_1 _2364_ (.A1(_0989_),
    .A2(net386),
    .Y(_0118_),
    .B1(_0481_));
 sg13g2_nor2_1 _2365_ (.A(net523),
    .B(net386),
    .Y(_0482_));
 sg13g2_a21oi_1 _2366_ (.A1(_0988_),
    .A2(net386),
    .Y(_0119_),
    .B1(_0482_));
 sg13g2_nor2_1 _2367_ (.A(net577),
    .B(net387),
    .Y(_0483_));
 sg13g2_a21oi_1 _2368_ (.A1(_0987_),
    .A2(net387),
    .Y(_0120_),
    .B1(_0483_));
 sg13g2_nor2_1 _2369_ (.A(net534),
    .B(net386),
    .Y(_0484_));
 sg13g2_a21oi_1 _2370_ (.A1(_0986_),
    .A2(net386),
    .Y(_0121_),
    .B1(_0484_));
 sg13g2_nand2b_1 _2371_ (.Y(_0485_),
    .B(\modem.uart.rxFifo.nextIn[0] ),
    .A_N(\modem.uart.rxFifo.nextIn[1] ));
 sg13g2_nor3_2 _2372_ (.A(_0065_),
    .B(_0474_),
    .C(_0485_),
    .Y(_0486_));
 sg13g2_nor2_1 _2373_ (.A(net632),
    .B(net385),
    .Y(_0487_));
 sg13g2_a21oi_1 _2374_ (.A1(net409),
    .A2(net385),
    .Y(_0122_),
    .B1(_0487_));
 sg13g2_nor2_1 _2375_ (.A(net567),
    .B(net384),
    .Y(_0488_));
 sg13g2_a21oi_1 _2376_ (.A1(_0992_),
    .A2(net384),
    .Y(_0123_),
    .B1(_0488_));
 sg13g2_nor2_1 _2377_ (.A(net672),
    .B(net385),
    .Y(_0489_));
 sg13g2_a21oi_1 _2378_ (.A1(_0991_),
    .A2(net385),
    .Y(_0124_),
    .B1(_0489_));
 sg13g2_nor2_1 _2379_ (.A(net631),
    .B(net385),
    .Y(_0490_));
 sg13g2_a21oi_1 _2380_ (.A1(net410),
    .A2(net385),
    .Y(_0125_),
    .B1(_0490_));
 sg13g2_nor2_1 _2381_ (.A(net571),
    .B(net384),
    .Y(_0491_));
 sg13g2_a21oi_1 _2382_ (.A1(_0989_),
    .A2(net384),
    .Y(_0126_),
    .B1(_0491_));
 sg13g2_nor2_1 _2383_ (.A(net536),
    .B(net385),
    .Y(_0492_));
 sg13g2_a21oi_1 _2384_ (.A1(_0988_),
    .A2(net384),
    .Y(_0127_),
    .B1(_0492_));
 sg13g2_nor2_1 _2385_ (.A(net573),
    .B(net384),
    .Y(_0493_));
 sg13g2_a21oi_1 _2386_ (.A1(_0987_),
    .A2(net384),
    .Y(_0128_),
    .B1(_0493_));
 sg13g2_nor2_1 _2387_ (.A(net667),
    .B(_0486_),
    .Y(_0494_));
 sg13g2_a21oi_1 _2388_ (.A1(_0986_),
    .A2(net384),
    .Y(_0129_),
    .B1(net668));
 sg13g2_nor4_2 _2389_ (.A(\modem.uart.rxFifo.nextIn[1] ),
    .B(\modem.uart.rxFifo.nextIn[0] ),
    .C(_0065_),
    .Y(_0495_),
    .D(_0474_));
 sg13g2_nor2_1 _2390_ (.A(net687),
    .B(net383),
    .Y(_0496_));
 sg13g2_a21oi_1 _2391_ (.A1(net409),
    .A2(net383),
    .Y(_0130_),
    .B1(_0496_));
 sg13g2_nor2_1 _2392_ (.A(net579),
    .B(net382),
    .Y(_0497_));
 sg13g2_a21oi_1 _2393_ (.A1(_0992_),
    .A2(net383),
    .Y(_0131_),
    .B1(_0497_));
 sg13g2_nor2_1 _2394_ (.A(net593),
    .B(net383),
    .Y(_0498_));
 sg13g2_a21oi_1 _2395_ (.A1(_0991_),
    .A2(_0495_),
    .Y(_0132_),
    .B1(_0498_));
 sg13g2_nor2_1 _2396_ (.A(net649),
    .B(net383),
    .Y(_0499_));
 sg13g2_a21oi_1 _2397_ (.A1(net410),
    .A2(net382),
    .Y(_0133_),
    .B1(_0499_));
 sg13g2_nor2_1 _2398_ (.A(net637),
    .B(net382),
    .Y(_0500_));
 sg13g2_a21oi_1 _2399_ (.A1(_0989_),
    .A2(net382),
    .Y(_0134_),
    .B1(_0500_));
 sg13g2_nor2_1 _2400_ (.A(net557),
    .B(net382),
    .Y(_0501_));
 sg13g2_a21oi_1 _2401_ (.A1(_0988_),
    .A2(net382),
    .Y(_0135_),
    .B1(_0501_));
 sg13g2_nor2_1 _2402_ (.A(net544),
    .B(net383),
    .Y(_0502_));
 sg13g2_a21oi_1 _2403_ (.A1(_0987_),
    .A2(net383),
    .Y(_0136_),
    .B1(_0502_));
 sg13g2_nor2_1 _2404_ (.A(net656),
    .B(net382),
    .Y(_0503_));
 sg13g2_a21oi_1 _2405_ (.A1(_0986_),
    .A2(net382),
    .Y(_0137_),
    .B1(_0503_));
 sg13g2_nand3_1 _2406_ (.B(\modem.uart.rxFifo.nextIn[0] ),
    .C(_0065_),
    .A(\modem.uart.rxFifo.nextIn[1] ),
    .Y(_0504_));
 sg13g2_nor2_1 _2407_ (.A(_0474_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_nor2_1 _2408_ (.A(net677),
    .B(net380),
    .Y(_0506_));
 sg13g2_a21oi_1 _2409_ (.A1(net409),
    .A2(net380),
    .Y(_0138_),
    .B1(_0506_));
 sg13g2_nor2_1 _2410_ (.A(net740),
    .B(net381),
    .Y(_0507_));
 sg13g2_a21oi_1 _2411_ (.A1(_0992_),
    .A2(net381),
    .Y(_0139_),
    .B1(_0507_));
 sg13g2_nor2_1 _2412_ (.A(net628),
    .B(net380),
    .Y(_0508_));
 sg13g2_a21oi_1 _2413_ (.A1(_0991_),
    .A2(net380),
    .Y(_0140_),
    .B1(_0508_));
 sg13g2_nor2_1 _2414_ (.A(\modem.uart.rxFifo.fifo_3[3] ),
    .B(_0505_),
    .Y(_0509_));
 sg13g2_a21oi_1 _2415_ (.A1(_0990_),
    .A2(net380),
    .Y(_0141_),
    .B1(_0509_));
 sg13g2_nor2_1 _2416_ (.A(net608),
    .B(net381),
    .Y(_0510_));
 sg13g2_a21oi_1 _2417_ (.A1(_0989_),
    .A2(net381),
    .Y(_0142_),
    .B1(_0510_));
 sg13g2_nor2_1 _2418_ (.A(net651),
    .B(net381),
    .Y(_0511_));
 sg13g2_a21oi_1 _2419_ (.A1(_0988_),
    .A2(net381),
    .Y(_0143_),
    .B1(_0511_));
 sg13g2_nor2_1 _2420_ (.A(net644),
    .B(net380),
    .Y(_0512_));
 sg13g2_a21oi_1 _2421_ (.A1(_0987_),
    .A2(net380),
    .Y(_0144_),
    .B1(_0512_));
 sg13g2_nor2_1 _2422_ (.A(net695),
    .B(net380),
    .Y(_0513_));
 sg13g2_a21oi_1 _2423_ (.A1(_0986_),
    .A2(net381),
    .Y(_0145_),
    .B1(_0513_));
 sg13g2_nor3_1 _2424_ (.A(\modem.uart.rxFifo.nextIn[2] ),
    .B(_0474_),
    .C(_0475_),
    .Y(_0514_));
 sg13g2_nor2_1 _2425_ (.A(net590),
    .B(net379),
    .Y(_0515_));
 sg13g2_a21oi_1 _2426_ (.A1(net409),
    .A2(net379),
    .Y(_0146_),
    .B1(_0515_));
 sg13g2_nor2_1 _2427_ (.A(net549),
    .B(net377),
    .Y(_0516_));
 sg13g2_a21oi_1 _2428_ (.A1(_0992_),
    .A2(net377),
    .Y(_0147_),
    .B1(_0516_));
 sg13g2_nor2_1 _2429_ (.A(net527),
    .B(net379),
    .Y(_0517_));
 sg13g2_a21oi_1 _2430_ (.A1(_0991_),
    .A2(net379),
    .Y(_0148_),
    .B1(_0517_));
 sg13g2_nor2_1 _2431_ (.A(net666),
    .B(net377),
    .Y(_0518_));
 sg13g2_a21oi_1 _2432_ (.A1(net410),
    .A2(net377),
    .Y(_0149_),
    .B1(_0518_));
 sg13g2_nor2_1 _2433_ (.A(net538),
    .B(net377),
    .Y(_0519_));
 sg13g2_a21oi_1 _2434_ (.A1(_0989_),
    .A2(net377),
    .Y(_0150_),
    .B1(_0519_));
 sg13g2_nor2_1 _2435_ (.A(net575),
    .B(net378),
    .Y(_0520_));
 sg13g2_a21oi_1 _2436_ (.A1(_0988_),
    .A2(net378),
    .Y(_0151_),
    .B1(_0520_));
 sg13g2_nor2_1 _2437_ (.A(net616),
    .B(net378),
    .Y(_0521_));
 sg13g2_a21oi_1 _2438_ (.A1(_0987_),
    .A2(net378),
    .Y(_0152_),
    .B1(_0521_));
 sg13g2_nor2_1 _2439_ (.A(net591),
    .B(net377),
    .Y(_0522_));
 sg13g2_a21oi_1 _2440_ (.A1(_0986_),
    .A2(net377),
    .Y(_0153_),
    .B1(_0522_));
 sg13g2_nor3_1 _2441_ (.A(\modem.uart.rxFifo.nextIn[2] ),
    .B(_0474_),
    .C(_0485_),
    .Y(_0523_));
 sg13g2_nor2_1 _2442_ (.A(net603),
    .B(net376),
    .Y(_0524_));
 sg13g2_a21oi_1 _2443_ (.A1(net409),
    .A2(net376),
    .Y(_0154_),
    .B1(_0524_));
 sg13g2_nor2_1 _2444_ (.A(net682),
    .B(net375),
    .Y(_0525_));
 sg13g2_a21oi_1 _2445_ (.A1(_0992_),
    .A2(net375),
    .Y(_0155_),
    .B1(_0525_));
 sg13g2_nor2_1 _2446_ (.A(net529),
    .B(net376),
    .Y(_0526_));
 sg13g2_a21oi_1 _2447_ (.A1(_0991_),
    .A2(net376),
    .Y(_0156_),
    .B1(_0526_));
 sg13g2_nor2_1 _2448_ (.A(net559),
    .B(net374),
    .Y(_0527_));
 sg13g2_a21oi_1 _2449_ (.A1(net410),
    .A2(net374),
    .Y(_0157_),
    .B1(_0527_));
 sg13g2_nor2_1 _2450_ (.A(net641),
    .B(net375),
    .Y(_0528_));
 sg13g2_a21oi_1 _2451_ (.A1(_0989_),
    .A2(net374),
    .Y(_0158_),
    .B1(_0528_));
 sg13g2_nor2_1 _2452_ (.A(net551),
    .B(net374),
    .Y(_0529_));
 sg13g2_a21oi_1 _2453_ (.A1(_0988_),
    .A2(net374),
    .Y(_0159_),
    .B1(_0529_));
 sg13g2_nor2_1 _2454_ (.A(net614),
    .B(net374),
    .Y(_0530_));
 sg13g2_a21oi_1 _2455_ (.A1(_0987_),
    .A2(net374),
    .Y(_0160_),
    .B1(_0530_));
 sg13g2_nor2_1 _2456_ (.A(net612),
    .B(net374),
    .Y(_0531_));
 sg13g2_a21oi_1 _2457_ (.A1(_0986_),
    .A2(net375),
    .Y(_0161_),
    .B1(_0531_));
 sg13g2_mux2_1 _2458_ (.A0(net660),
    .A1(net635),
    .S(\modem.control.io_txClockStb ),
    .X(_0162_));
 sg13g2_nor4_1 _2459_ (.A(\modem.uart.rxFifo.nextIn[2] ),
    .B(_0995_),
    .C(\modem.uart.rxFifo.nextIn[1] ),
    .D(\modem.uart.rxFifo.nextIn[0] ),
    .Y(_0532_));
 sg13g2_o21ai_1 _2460_ (.B1(net442),
    .Y(_0533_),
    .A1(net806),
    .A2(net373));
 sg13g2_a21oi_1 _2461_ (.A1(net409),
    .A2(net373),
    .Y(_0163_),
    .B1(_0533_));
 sg13g2_o21ai_1 _2462_ (.B1(net441),
    .Y(_0534_),
    .A1(net810),
    .A2(net373));
 sg13g2_a21oi_1 _2463_ (.A1(_0992_),
    .A2(net373),
    .Y(_0164_),
    .B1(_0534_));
 sg13g2_o21ai_1 _2464_ (.B1(net441),
    .Y(_0535_),
    .A1(net840),
    .A2(net372));
 sg13g2_a21oi_1 _2465_ (.A1(_0991_),
    .A2(net372),
    .Y(_0165_),
    .B1(_0535_));
 sg13g2_o21ai_1 _2466_ (.B1(net441),
    .Y(_0536_),
    .A1(net798),
    .A2(net372));
 sg13g2_a21oi_1 _2467_ (.A1(net410),
    .A2(net372),
    .Y(_0166_),
    .B1(_0536_));
 sg13g2_o21ai_1 _2468_ (.B1(net441),
    .Y(_0537_),
    .A1(net829),
    .A2(net372));
 sg13g2_a21oi_1 _2469_ (.A1(_0989_),
    .A2(net372),
    .Y(_0167_),
    .B1(_0537_));
 sg13g2_o21ai_1 _2470_ (.B1(net442),
    .Y(_0538_),
    .A1(net814),
    .A2(net373));
 sg13g2_a21oi_1 _2471_ (.A1(_0988_),
    .A2(net373),
    .Y(_0168_),
    .B1(_0538_));
 sg13g2_o21ai_1 _2472_ (.B1(net441),
    .Y(_0539_),
    .A1(net846),
    .A2(net372));
 sg13g2_a21oi_1 _2473_ (.A1(_0987_),
    .A2(net372),
    .Y(_0169_),
    .B1(_0539_));
 sg13g2_o21ai_1 _2474_ (.B1(net441),
    .Y(_0540_),
    .A1(net803),
    .A2(net373));
 sg13g2_a21oi_1 _2475_ (.A1(_0986_),
    .A2(net373),
    .Y(_0170_),
    .B1(_0540_));
 sg13g2_xnor2_1 _2476_ (.Y(_0541_),
    .A(_0995_),
    .B(_0468_));
 sg13g2_nor2_1 _2477_ (.A(\modem.uart.rxFifo.count[0] ),
    .B(_0541_),
    .Y(_0542_));
 sg13g2_nor2b_1 _2478_ (.A(net487),
    .B_N(_0541_),
    .Y(_0543_));
 sg13g2_nor3_1 _2479_ (.A(net406),
    .B(_0542_),
    .C(_0543_),
    .Y(_0171_));
 sg13g2_nor2b_1 _2480_ (.A(net418),
    .B_N(\modem.uart.rxFifo.count[1] ),
    .Y(_0544_));
 sg13g2_nand2b_1 _2481_ (.Y(_0545_),
    .B(net418),
    .A_N(\modem.uart.rxFifo.count[1] ));
 sg13g2_nor2b_1 _2482_ (.A(_0544_),
    .B_N(_0545_),
    .Y(_0546_));
 sg13g2_xnor2_1 _2483_ (.Y(_0547_),
    .A(net487),
    .B(_0546_));
 sg13g2_mux2_1 _2484_ (.A0(net893),
    .A1(_0547_),
    .S(_0541_),
    .X(_0548_));
 sg13g2_and2_1 _2485_ (.A(net443),
    .B(_0548_),
    .X(_0172_));
 sg13g2_o21ai_1 _2486_ (.B1(_0545_),
    .Y(_0549_),
    .A1(\modem.uart.rxFifo.count[0] ),
    .A2(_0544_));
 sg13g2_xor2_1 _2487_ (.B(net419),
    .A(\modem.uart.rxFifo.count[2] ),
    .X(_0550_));
 sg13g2_xnor2_1 _2488_ (.Y(_0551_),
    .A(_0549_),
    .B(_0550_));
 sg13g2_nand2_1 _2489_ (.Y(_0552_),
    .A(_0541_),
    .B(_0551_));
 sg13g2_o21ai_1 _2490_ (.B1(_0552_),
    .Y(_0553_),
    .A1(net883),
    .A2(_0541_));
 sg13g2_nor2_1 _2491_ (.A(net406),
    .B(_0553_),
    .Y(_0173_));
 sg13g2_nor4_1 _2492_ (.A(_0995_),
    .B(net346),
    .C(_0549_),
    .D(_0550_),
    .Y(_0554_));
 sg13g2_nor4_1 _2493_ (.A(\modem.uart.rxFifo.count[2] ),
    .B(\modem.uart.rxFifo.count[1] ),
    .C(\modem.uart.rxFifo.count[0] ),
    .D(net419),
    .Y(_0555_));
 sg13g2_a21o_1 _2494_ (.A2(_0555_),
    .A1(net346),
    .B1(_0554_),
    .X(_0556_));
 sg13g2_o21ai_1 _2495_ (.B1(net443),
    .Y(_0557_),
    .A1(net662),
    .A2(_0556_));
 sg13g2_a21oi_1 _2496_ (.A1(net662),
    .A2(_0556_),
    .Y(_0174_),
    .B1(_0557_));
 sg13g2_nor2_1 _2497_ (.A(net430),
    .B(_1012_),
    .Y(_0558_));
 sg13g2_nand2_1 _2498_ (.Y(_0559_),
    .A(_0985_),
    .B(\modem.uart.io_isSending ));
 sg13g2_a21oi_1 _2499_ (.A1(_1179_),
    .A2(_1184_),
    .Y(_0560_),
    .B1(net426));
 sg13g2_nor2b_1 _2500_ (.A(_1180_),
    .B_N(net426),
    .Y(_0561_));
 sg13g2_nand2_1 _2501_ (.Y(_0562_),
    .A(net426),
    .B(_1181_));
 sg13g2_o21ai_1 _2502_ (.B1(_1009_),
    .Y(_0563_),
    .A1(_1063_),
    .A2(_0562_));
 sg13g2_nand3b_1 _2503_ (.B(_1080_),
    .C(_1181_),
    .Y(_0564_),
    .A_N(net426));
 sg13g2_nand3_1 _2504_ (.B(_1177_),
    .C(_0564_),
    .A(net424),
    .Y(_0565_));
 sg13g2_a21o_1 _2505_ (.A2(_0561_),
    .A1(_1071_),
    .B1(_0565_),
    .X(_0566_));
 sg13g2_and2_1 _2506_ (.A(net422),
    .B(_0566_),
    .X(_0567_));
 sg13g2_o21ai_1 _2507_ (.B1(_0567_),
    .Y(_0568_),
    .A1(_0560_),
    .A2(_0563_));
 sg13g2_o21ai_1 _2508_ (.B1(_1179_),
    .Y(_0569_),
    .A1(_1107_),
    .A2(_1180_));
 sg13g2_nor2_1 _2509_ (.A(net426),
    .B(_0569_),
    .Y(_0570_));
 sg13g2_nand2b_1 _2510_ (.Y(_0571_),
    .B(_1137_),
    .A_N(_1178_));
 sg13g2_nor4_1 _2511_ (.A(_1090_),
    .B(_1107_),
    .C(_1142_),
    .D(_0571_),
    .Y(_0572_));
 sg13g2_and2_1 _2512_ (.A(net426),
    .B(_1179_),
    .X(_0573_));
 sg13g2_o21ai_1 _2513_ (.B1(_0573_),
    .Y(_0574_),
    .A1(_1124_),
    .A2(_1180_));
 sg13g2_nor2_1 _2514_ (.A(_0572_),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_o21ai_1 _2515_ (.B1(_1009_),
    .Y(_0576_),
    .A1(_0570_),
    .A2(_0575_));
 sg13g2_nand3_1 _2516_ (.B(_1181_),
    .C(_1183_),
    .A(_1115_),
    .Y(_0577_));
 sg13g2_nand3_1 _2517_ (.B(_0573_),
    .C(_0577_),
    .A(net424),
    .Y(_0578_));
 sg13g2_nor2_2 _2518_ (.A(net426),
    .B(_1009_),
    .Y(_0579_));
 sg13g2_nor2b_1 _2519_ (.A(_1143_),
    .B_N(_1182_),
    .Y(_0580_));
 sg13g2_o21ai_1 _2520_ (.B1(_1098_),
    .Y(_0581_),
    .A1(_1024_),
    .A2(_1177_));
 sg13g2_o21ai_1 _2521_ (.B1(_0579_),
    .Y(_0582_),
    .A1(_0580_),
    .A2(_0581_));
 sg13g2_nand4_1 _2522_ (.B(_0576_),
    .C(_0578_),
    .A(_1010_),
    .Y(_0583_),
    .D(_0582_));
 sg13g2_and2_2 _2523_ (.A(_0568_),
    .B(_0583_),
    .X(_0584_));
 sg13g2_nand2b_1 _2524_ (.Y(_0585_),
    .B(\modem.uart.txHdlc.bitstuffCnt[0] ),
    .A_N(_0053_));
 sg13g2_nor2_2 _2525_ (.A(\modem.uart.txHdlc.bitstuffCnt[1] ),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_inv_1 _2526_ (.Y(_0587_),
    .A(_0586_));
 sg13g2_and2_1 _2527_ (.A(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[4] ),
    .B(\modem.uart.txCommandDecoder.io_valid ),
    .X(_0588_));
 sg13g2_nand2_2 _2528_ (.Y(_0589_),
    .A(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[4] ),
    .B(\modem.uart.txCommandDecoder.io_valid ));
 sg13g2_nor4_1 _2529_ (.A(_0559_),
    .B(_0584_),
    .C(_0586_),
    .D(_0589_),
    .Y(_0590_));
 sg13g2_nand2b_1 _2530_ (.Y(_0591_),
    .B(net428),
    .A_N(\modem.uart.txHdlc.txCrc.crcNext_2 ));
 sg13g2_o21ai_1 _2531_ (.B1(_0591_),
    .Y(_0592_),
    .A1(\modem.uart.txHdlc.txCrc.crcNext_1 ),
    .A2(net425));
 sg13g2_a22oi_1 _2532_ (.Y(_0593_),
    .B1(_0579_),
    .B2(\modem.uart.txHdlc.txCrc.crcNext_3 ),
    .A2(_1036_),
    .A1(\modem.uart.txHdlc.txCrc.crcNext_4 ));
 sg13g2_o21ai_1 _2533_ (.B1(_0593_),
    .Y(_0594_),
    .A1(net423),
    .A2(_0592_));
 sg13g2_nor2b_1 _2534_ (.A(net425),
    .B_N(\modem.uart.txHdlc.txCrc.crc[4] ),
    .Y(_0595_));
 sg13g2_a21oi_1 _2535_ (.A1(\modem.uart.txHdlc.txCrc.crcNext_6 ),
    .A2(net425),
    .Y(_0596_),
    .B1(_0595_));
 sg13g2_a221oi_1 _2536_ (.B2(\modem.uart.txHdlc.txCrc.crcNext_7 ),
    .C1(_1010_),
    .B1(_0579_),
    .A1(\modem.uart.txHdlc.txCrc.crcNext_8 ),
    .Y(_0597_),
    .A2(_1036_));
 sg13g2_o21ai_1 _2537_ (.B1(_0597_),
    .Y(_0598_),
    .A1(net423),
    .A2(_0596_));
 sg13g2_o21ai_1 _2538_ (.B1(_0598_),
    .Y(_0599_),
    .A1(net422),
    .A2(_0594_));
 sg13g2_nor2b_1 _2539_ (.A(\modem.uart.txHdlc.bit8[2] ),
    .B_N(net421),
    .Y(_0600_));
 sg13g2_nor2b_1 _2540_ (.A(net425),
    .B_N(\modem.uart.txHdlc.txCrc.crcNext_9 ),
    .Y(_0601_));
 sg13g2_a21oi_1 _2541_ (.A1(\modem.uart.txHdlc.txCrc.crcNext_10 ),
    .A2(net425),
    .Y(_0602_),
    .B1(_0601_));
 sg13g2_a22oi_1 _2542_ (.Y(_0603_),
    .B1(_0579_),
    .B2(\modem.uart.txHdlc.txCrc.crcNext_11 ),
    .A2(_1036_),
    .A1(\modem.uart.txHdlc.txCrc.crc[11] ));
 sg13g2_o21ai_1 _2543_ (.B1(_0603_),
    .Y(_0604_),
    .A1(net423),
    .A2(_0602_));
 sg13g2_nor2b_1 _2544_ (.A(net425),
    .B_N(\modem.uart.txHdlc.txCrc.crcNext_13 ),
    .Y(_0605_));
 sg13g2_a21oi_1 _2545_ (.A1(\modem.uart.txHdlc.txCrc.crcNext_14 ),
    .A2(net425),
    .Y(_0606_),
    .B1(_0605_));
 sg13g2_a22oi_1 _2546_ (.Y(_0607_),
    .B1(_0579_),
    .B2(\modem.uart.txHdlc.txCrc.crcNext_15 ),
    .A2(_1036_),
    .A1(\modem.uart.txHdlc.txCrc.crc[15] ));
 sg13g2_o21ai_1 _2547_ (.B1(_0607_),
    .Y(_0608_),
    .A1(net423),
    .A2(_0606_));
 sg13g2_nand3_1 _2548_ (.B(net421),
    .C(_0608_),
    .A(net422),
    .Y(_0609_));
 sg13g2_o21ai_1 _2549_ (.B1(_0609_),
    .Y(_0610_),
    .A1(net421),
    .A2(_0599_));
 sg13g2_a21oi_2 _2550_ (.B1(_0610_),
    .Y(_0611_),
    .A2(_0604_),
    .A1(_0600_));
 sg13g2_nand2_1 _2551_ (.Y(_0612_),
    .A(net429),
    .B(_0611_));
 sg13g2_nand2_1 _2552_ (.Y(_0613_),
    .A(_0558_),
    .B(_0589_));
 sg13g2_nand3_1 _2553_ (.B(_0558_),
    .C(_0589_),
    .A(net878),
    .Y(_0614_));
 sg13g2_nor2_2 _2554_ (.A(net430),
    .B(\modem.uart.io_isSending ),
    .Y(_0615_));
 sg13g2_and2_1 _2555_ (.A(_0054_),
    .B(_0615_),
    .X(_0616_));
 sg13g2_o21ai_1 _2556_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_1009_),
    .A2(_1010_));
 sg13g2_nand2_1 _2557_ (.Y(_0618_),
    .A(\modem.uart.txHdlc.wantFrameEnd ),
    .B(_0611_));
 sg13g2_o21ai_1 _2558_ (.B1(_0618_),
    .Y(_0619_),
    .A1(net431),
    .A2(\modem.uart.txHdlc.wantFrameEnd ));
 sg13g2_nor2_1 _2559_ (.A(_0613_),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_o21ai_1 _2560_ (.B1(_0617_),
    .Y(_0621_),
    .A1(_0586_),
    .A2(_0612_));
 sg13g2_nor3_1 _2561_ (.A(_0590_),
    .B(_0620_),
    .C(_0621_),
    .Y(_0622_));
 sg13g2_or2_1 _2562_ (.X(_0623_),
    .B(_0622_),
    .A(\modem.uart.txHdlc.isAbort ));
 sg13g2_o21ai_1 _2563_ (.B1(\modem.uart.txHdlc.when_ModemTop_l593 ),
    .Y(_0624_),
    .A1(net424),
    .A2(net422));
 sg13g2_nor4_1 _2564_ (.A(net427),
    .B(net423),
    .C(net422),
    .D(net421),
    .Y(_0625_));
 sg13g2_nand2_1 _2565_ (.Y(_0626_),
    .A(\modem.uart.txHdlc.isAbort ),
    .B(_0624_));
 sg13g2_nor2_2 _2566_ (.A(_0625_),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_nor3_1 _2567_ (.A(net868),
    .B(net368),
    .C(_0627_),
    .Y(_0628_));
 sg13g2_a221oi_1 _2568_ (.B2(_0628_),
    .C1(net405),
    .B1(_0623_),
    .A1(_0971_),
    .Y(_0175_),
    .A2(net368));
 sg13g2_mux2_1 _2569_ (.A0(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[4] ),
    .A1(_1194_),
    .S(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[1] ),
    .X(_0629_));
 sg13g2_or3_1 _2570_ (.A(net303),
    .B(\modem.uart.txCommandDecoder.io_valid ),
    .C(_1190_),
    .X(_0630_));
 sg13g2_nand2_1 _2571_ (.Y(_0631_),
    .A(_1190_),
    .B(_1194_));
 sg13g2_nand3_1 _2572_ (.B(_0630_),
    .C(_0631_),
    .A(net316),
    .Y(_0632_));
 sg13g2_o21ai_1 _2573_ (.B1(net444),
    .Y(_0633_),
    .A1(net303),
    .A2(_0629_));
 sg13g2_a21oi_1 _2574_ (.A1(_0629_),
    .A2(_0632_),
    .Y(_0176_),
    .B1(_0633_));
 sg13g2_a21oi_2 _2575_ (.B1(_0587_),
    .Y(_0634_),
    .A2(_0583_),
    .A1(_0568_));
 sg13g2_nand2_1 _2576_ (.Y(_0635_),
    .A(_0060_),
    .B(_0589_));
 sg13g2_nand2_1 _2577_ (.Y(_0636_),
    .A(_0588_),
    .B(_0634_));
 sg13g2_and3_1 _2578_ (.X(_0637_),
    .A(_1035_),
    .B(_0635_),
    .C(_0636_));
 sg13g2_nand3_1 _2579_ (.B(_0635_),
    .C(_0636_),
    .A(_1035_),
    .Y(_0638_));
 sg13g2_nand2_1 _2580_ (.Y(_0639_),
    .A(net732),
    .B(net341));
 sg13g2_xnor2_1 _2581_ (.Y(_0640_),
    .A(\modem.uart.txHdlc.txCrc.crc[15] ),
    .B(_0584_));
 sg13g2_nand2_1 _2582_ (.Y(_0641_),
    .A(net344),
    .B(_0640_));
 sg13g2_nor2_1 _2583_ (.A(net404),
    .B(_0615_),
    .Y(_0642_));
 sg13g2_nand3_1 _2584_ (.B(_0641_),
    .C(net370),
    .A(_0639_),
    .Y(_0177_));
 sg13g2_nand2_1 _2585_ (.Y(_0643_),
    .A(net732),
    .B(net344));
 sg13g2_nand2_1 _2586_ (.Y(_0644_),
    .A(\modem.uart.txHdlc.txCrc.crcNext_2 ),
    .B(net342));
 sg13g2_nand3_1 _2587_ (.B(_0643_),
    .C(_0644_),
    .A(net370),
    .Y(_0178_));
 sg13g2_nand2_1 _2588_ (.Y(_0645_),
    .A(\modem.uart.txHdlc.txCrc.crcNext_3 ),
    .B(net341));
 sg13g2_nand2_1 _2589_ (.Y(_0646_),
    .A(net789),
    .B(net344));
 sg13g2_nand3_1 _2590_ (.B(_0645_),
    .C(_0646_),
    .A(net370),
    .Y(_0179_));
 sg13g2_nand2_1 _2591_ (.Y(_0647_),
    .A(net837),
    .B(net344));
 sg13g2_nand2_1 _2592_ (.Y(_0648_),
    .A(net831),
    .B(net341));
 sg13g2_nand3_1 _2593_ (.B(_0647_),
    .C(_0648_),
    .A(net370),
    .Y(_0180_));
 sg13g2_nand2_1 _2594_ (.Y(_0649_),
    .A(net831),
    .B(net344));
 sg13g2_nand2_1 _2595_ (.Y(_0650_),
    .A(\modem.uart.txHdlc.txCrc.crc[4] ),
    .B(net341));
 sg13g2_nand3_1 _2596_ (.B(_0649_),
    .C(_0650_),
    .A(net370),
    .Y(_0181_));
 sg13g2_xnor2_1 _2597_ (.Y(_0651_),
    .A(\modem.uart.txHdlc.txCrc.crc[4] ),
    .B(_0640_));
 sg13g2_o21ai_1 _2598_ (.B1(net370),
    .Y(_0652_),
    .A1(net341),
    .A2(_0651_));
 sg13g2_a21o_1 _2599_ (.A2(net341),
    .A1(net726),
    .B1(_0652_),
    .X(_0182_));
 sg13g2_nand2_1 _2600_ (.Y(_0653_),
    .A(net731),
    .B(net343));
 sg13g2_nand2_1 _2601_ (.Y(_0654_),
    .A(net726),
    .B(net344));
 sg13g2_nand3_1 _2602_ (.B(_0653_),
    .C(_0654_),
    .A(net371),
    .Y(_0183_));
 sg13g2_nand2_1 _2603_ (.Y(_0655_),
    .A(net754),
    .B(net343));
 sg13g2_nand2_1 _2604_ (.Y(_0656_),
    .A(net731),
    .B(net345));
 sg13g2_nand3_1 _2605_ (.B(_0655_),
    .C(_0656_),
    .A(net371),
    .Y(_0184_));
 sg13g2_nand2_1 _2606_ (.Y(_0657_),
    .A(net754),
    .B(net345));
 sg13g2_nand2_1 _2607_ (.Y(_0658_),
    .A(net744),
    .B(net342));
 sg13g2_nand3_1 _2608_ (.B(_0657_),
    .C(_0658_),
    .A(net371),
    .Y(_0185_));
 sg13g2_nand2_1 _2609_ (.Y(_0659_),
    .A(net744),
    .B(net344));
 sg13g2_nand2_1 _2610_ (.Y(_0660_),
    .A(\modem.uart.txHdlc.txCrc.crcNext_10 ),
    .B(net342));
 sg13g2_nand3_1 _2611_ (.B(_0659_),
    .C(_0660_),
    .A(net371),
    .Y(_0186_));
 sg13g2_nand2_1 _2612_ (.Y(_0661_),
    .A(net791),
    .B(net344));
 sg13g2_nand2_1 _2613_ (.Y(_0662_),
    .A(net782),
    .B(net342));
 sg13g2_nand3_1 _2614_ (.B(_0661_),
    .C(_0662_),
    .A(net370),
    .Y(_0187_));
 sg13g2_nand2_1 _2615_ (.Y(_0663_),
    .A(net782),
    .B(net345));
 sg13g2_nand2_1 _2616_ (.Y(_0664_),
    .A(\modem.uart.txHdlc.txCrc.crc[11] ),
    .B(net342));
 sg13g2_nand3_1 _2617_ (.B(_0663_),
    .C(_0664_),
    .A(net371),
    .Y(_0188_));
 sg13g2_xnor2_1 _2618_ (.Y(_0665_),
    .A(\modem.uart.txHdlc.txCrc.crc[11] ),
    .B(_0640_));
 sg13g2_o21ai_1 _2619_ (.B1(net370),
    .Y(_0666_),
    .A1(net341),
    .A2(_0665_));
 sg13g2_a21o_1 _2620_ (.A2(net341),
    .A1(net738),
    .B1(_0666_),
    .X(_0189_));
 sg13g2_nand2_1 _2621_ (.Y(_0667_),
    .A(net738),
    .B(net345));
 sg13g2_nand2_1 _2622_ (.Y(_0668_),
    .A(net774),
    .B(net343));
 sg13g2_nand3_1 _2623_ (.B(_0667_),
    .C(_0668_),
    .A(_0642_),
    .Y(_0190_));
 sg13g2_nand2_1 _2624_ (.Y(_0669_),
    .A(net774),
    .B(net345));
 sg13g2_nand2_1 _2625_ (.Y(_0670_),
    .A(\modem.uart.txHdlc.txCrc.crcNext_15 ),
    .B(net343));
 sg13g2_nand3_1 _2626_ (.B(_0669_),
    .C(_0670_),
    .A(net371),
    .Y(_0191_));
 sg13g2_nand2_1 _2627_ (.Y(_0671_),
    .A(net830),
    .B(net345));
 sg13g2_nand2_1 _2628_ (.Y(_0672_),
    .A(net750),
    .B(net343));
 sg13g2_nand3_1 _2629_ (.B(_0671_),
    .C(_0672_),
    .A(net371),
    .Y(_0192_));
 sg13g2_nor4_2 _2630_ (.A(net427),
    .B(_1009_),
    .C(_1010_),
    .Y(_0673_),
    .D(net421));
 sg13g2_nand4_1 _2631_ (.B(_0588_),
    .C(_0615_),
    .A(_1033_),
    .Y(_0674_),
    .D(_0673_));
 sg13g2_nor2b_1 _2632_ (.A(net303),
    .B_N(\modem.uart.uart_txCommandDecoder_io_wantTx_regNext ),
    .Y(_0675_));
 sg13g2_o21ai_1 _2633_ (.B1(net444),
    .Y(_0676_),
    .A1(_1034_),
    .A2(_0614_));
 sg13g2_o21ai_1 _2634_ (.B1(_0674_),
    .Y(_0677_),
    .A1(net878),
    .A2(_0675_));
 sg13g2_nor2_1 _2635_ (.A(_0676_),
    .B(net879),
    .Y(_0193_));
 sg13g2_or2_2 _2636_ (.X(_0678_),
    .B(_1144_),
    .A(net815));
 sg13g2_nor3_1 _2637_ (.A(net901),
    .B(_1034_),
    .C(_0613_),
    .Y(_0679_));
 sg13g2_nor2b_1 _2638_ (.A(_0679_),
    .B_N(net875),
    .Y(_0680_));
 sg13g2_and3_1 _2639_ (.X(_0681_),
    .A(net427),
    .B(_1009_),
    .C(_0600_));
 sg13g2_and2_1 _2640_ (.A(\modem.uart.txHdlc.isAbort ),
    .B(net366),
    .X(_0682_));
 sg13g2_and2_1 _2641_ (.A(_0586_),
    .B(_0611_),
    .X(_0683_));
 sg13g2_nand3_1 _2642_ (.B(net421),
    .C(_1036_),
    .A(net422),
    .Y(_0684_));
 sg13g2_nor3_2 _2643_ (.A(_0985_),
    .B(_0683_),
    .C(_0684_),
    .Y(_0685_));
 sg13g2_a21o_1 _2644_ (.A2(_0685_),
    .A1(_1033_),
    .B1(net404),
    .X(_0686_));
 sg13g2_a221oi_1 _2645_ (.B2(_0682_),
    .C1(_0686_),
    .B1(_0681_),
    .A1(_0678_),
    .Y(_0194_),
    .A2(_0680_));
 sg13g2_nor3_1 _2646_ (.A(_1012_),
    .B(net873),
    .C(_0588_),
    .Y(_0687_));
 sg13g2_a21oi_1 _2647_ (.A1(_1033_),
    .A2(_0687_),
    .Y(_0688_),
    .B1(net430));
 sg13g2_nor2_1 _2648_ (.A(_0686_),
    .B(net874),
    .Y(_0195_));
 sg13g2_nand3_1 _2649_ (.B(_1033_),
    .C(_0589_),
    .A(_0985_),
    .Y(_0689_));
 sg13g2_nand3_1 _2650_ (.B(_1144_),
    .C(_0689_),
    .A(net802),
    .Y(_0690_));
 sg13g2_a21oi_1 _2651_ (.A1(_0674_),
    .A2(_0690_),
    .Y(_0196_),
    .B1(net405));
 sg13g2_nor3_2 _2652_ (.A(_1008_),
    .B(\modem.uart.io_isSending ),
    .C(_0673_),
    .Y(_0691_));
 sg13g2_nand2b_1 _2653_ (.Y(_0692_),
    .B(_0691_),
    .A_N(net427));
 sg13g2_and2_1 _2654_ (.A(net427),
    .B(_0678_),
    .X(_0693_));
 sg13g2_mux2_1 _2655_ (.A0(_0056_),
    .A1(_0693_),
    .S(_0634_),
    .X(_0694_));
 sg13g2_nand2b_1 _2656_ (.Y(_0695_),
    .B(\modem.uart.io_isSending ),
    .A_N(_1038_));
 sg13g2_a21oi_1 _2657_ (.A1(_1011_),
    .A2(_0589_),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_o21ai_1 _2658_ (.B1(_0696_),
    .Y(_0697_),
    .A1(_0589_),
    .A2(_0694_));
 sg13g2_a21o_1 _2659_ (.A2(_0697_),
    .A1(_0692_),
    .B1(net429),
    .X(_0698_));
 sg13g2_nor2b_2 _2660_ (.A(_0683_),
    .B_N(_0684_),
    .Y(_0699_));
 sg13g2_mux2_1 _2661_ (.A0(_0693_),
    .A1(net894),
    .S(_0699_),
    .X(_0700_));
 sg13g2_a21oi_1 _2662_ (.A1(net429),
    .A2(_0700_),
    .Y(_0701_),
    .B1(_1034_));
 sg13g2_a21oi_1 _2663_ (.A1(net426),
    .A2(_0682_),
    .Y(_0702_),
    .B1(net404));
 sg13g2_o21ai_1 _2664_ (.B1(_0702_),
    .Y(_0703_),
    .A1(net366),
    .A2(_0693_));
 sg13g2_a21oi_1 _2665_ (.A1(_0698_),
    .A2(net895),
    .Y(_0197_),
    .B1(_0703_));
 sg13g2_xor2_1 _2666_ (.B(net423),
    .A(net427),
    .X(_0704_));
 sg13g2_nor2_1 _2667_ (.A(_0589_),
    .B(_0695_),
    .Y(_0705_));
 sg13g2_and2_1 _2668_ (.A(net423),
    .B(_0678_),
    .X(_0706_));
 sg13g2_mux2_1 _2669_ (.A0(_0704_),
    .A1(_0706_),
    .S(_0634_),
    .X(_0707_));
 sg13g2_a221oi_1 _2670_ (.B2(_0707_),
    .C1(net429),
    .B1(_0705_),
    .A1(_0691_),
    .Y(_0708_),
    .A2(_0704_));
 sg13g2_nand2b_1 _2671_ (.Y(_0709_),
    .B(_0706_),
    .A_N(_0699_));
 sg13g2_nand2b_1 _2672_ (.Y(_0710_),
    .B(_0704_),
    .A_N(_0683_));
 sg13g2_nand3_1 _2673_ (.B(_0709_),
    .C(_0710_),
    .A(net429),
    .Y(_0711_));
 sg13g2_nand3b_1 _2674_ (.B(_0711_),
    .C(_1033_),
    .Y(_0712_),
    .A_N(_0708_));
 sg13g2_nor2b_1 _2675_ (.A(_0681_),
    .B_N(_0682_),
    .Y(_0713_));
 sg13g2_a22oi_1 _2676_ (.Y(_0714_),
    .B1(_0713_),
    .B2(_0704_),
    .A2(_0706_),
    .A1(net368));
 sg13g2_a21oi_1 _2677_ (.A1(_0712_),
    .A2(_0714_),
    .Y(_0198_),
    .B1(net404));
 sg13g2_nor2_1 _2678_ (.A(net900),
    .B(_1037_),
    .Y(_0715_));
 sg13g2_xnor2_1 _2679_ (.Y(_0716_),
    .A(net899),
    .B(_1036_));
 sg13g2_and2_1 _2680_ (.A(net422),
    .B(_0678_),
    .X(_0717_));
 sg13g2_mux2_1 _2681_ (.A0(_0716_),
    .A1(_0717_),
    .S(_0634_),
    .X(_0718_));
 sg13g2_a221oi_1 _2682_ (.B2(_0705_),
    .C1(net429),
    .B1(_0718_),
    .A1(_0691_),
    .Y(_0719_),
    .A2(_0716_));
 sg13g2_nand2b_1 _2683_ (.Y(_0720_),
    .B(_0717_),
    .A_N(_0699_));
 sg13g2_a21oi_1 _2684_ (.A1(_0699_),
    .A2(_0716_),
    .Y(_0721_),
    .B1(_0985_));
 sg13g2_a21oi_1 _2685_ (.A1(_0720_),
    .A2(_0721_),
    .Y(_0722_),
    .B1(_1034_));
 sg13g2_nand2b_1 _2686_ (.Y(_0723_),
    .B(_0722_),
    .A_N(_0719_));
 sg13g2_a22oi_1 _2687_ (.Y(_0724_),
    .B1(_0717_),
    .B2(net368),
    .A2(_0716_),
    .A1(_0713_));
 sg13g2_a21oi_1 _2688_ (.A1(_0723_),
    .A2(_0724_),
    .Y(_0199_),
    .B1(net404));
 sg13g2_nand2_1 _2689_ (.Y(_0725_),
    .A(net421),
    .B(_0678_));
 sg13g2_xnor2_1 _2690_ (.Y(_0726_),
    .A(_1008_),
    .B(_0715_));
 sg13g2_inv_1 _2691_ (.Y(_0727_),
    .A(_0726_));
 sg13g2_o21ai_1 _2692_ (.B1(_0705_),
    .Y(_0728_),
    .A1(_0634_),
    .A2(_0727_));
 sg13g2_a21oi_1 _2693_ (.A1(_0634_),
    .A2(_0725_),
    .Y(_0729_),
    .B1(net429));
 sg13g2_nand2b_1 _2694_ (.Y(_0730_),
    .B(_0729_),
    .A_N(_0728_));
 sg13g2_nand2b_1 _2695_ (.Y(_0731_),
    .B(_0725_),
    .A_N(_0699_));
 sg13g2_a21oi_1 _2696_ (.A1(_0699_),
    .A2(_0726_),
    .Y(_0732_),
    .B1(_0985_));
 sg13g2_a22oi_1 _2697_ (.Y(_0733_),
    .B1(_0731_),
    .B2(_0732_),
    .A2(_0715_),
    .A1(_0616_));
 sg13g2_a21o_1 _2698_ (.A2(_0733_),
    .A1(_0730_),
    .B1(_1034_),
    .X(_0734_));
 sg13g2_nor2_1 _2699_ (.A(net366),
    .B(_0725_),
    .Y(_0735_));
 sg13g2_a21oi_1 _2700_ (.A1(_0713_),
    .A2(_0727_),
    .Y(_0736_),
    .B1(_0735_));
 sg13g2_a21oi_1 _2701_ (.A1(_0734_),
    .A2(_0736_),
    .Y(_0200_),
    .B1(net404));
 sg13g2_nand2_1 _2702_ (.Y(_0737_),
    .A(_0054_),
    .B(_0588_));
 sg13g2_and2_1 _2703_ (.A(_0615_),
    .B(_0737_),
    .X(_0738_));
 sg13g2_o21ai_1 _2704_ (.B1(_0738_),
    .Y(_0739_),
    .A1(_1008_),
    .A2(_0673_));
 sg13g2_nor4_1 _2705_ (.A(\modem.uart.io_isSending ),
    .B(net421),
    .C(_1025_),
    .D(_0673_),
    .Y(_0740_));
 sg13g2_nand4_1 _2706_ (.B(net366),
    .C(_0613_),
    .A(_0059_),
    .Y(_0741_),
    .D(_0739_));
 sg13g2_nor3_2 _2707_ (.A(_0685_),
    .B(_0740_),
    .C(_0741_),
    .Y(_0742_));
 sg13g2_inv_1 _2708_ (.Y(_0743_),
    .A(_0742_));
 sg13g2_o21ai_1 _2709_ (.B1(_0612_),
    .Y(_0744_),
    .A1(_0559_),
    .A2(_0584_));
 sg13g2_nand2_1 _2710_ (.Y(_0745_),
    .A(_0742_),
    .B(_0744_));
 sg13g2_nand2_1 _2711_ (.Y(_0746_),
    .A(net691),
    .B(_0742_));
 sg13g2_nand2_1 _2712_ (.Y(_0747_),
    .A(net444),
    .B(_0746_));
 sg13g2_a21oi_1 _2713_ (.A1(_0984_),
    .A2(_0745_),
    .Y(_0201_),
    .B1(_0747_));
 sg13g2_nand2_1 _2714_ (.Y(_0748_),
    .A(net794),
    .B(net691));
 sg13g2_nand3_1 _2715_ (.B(_0744_),
    .C(_0748_),
    .A(_0585_),
    .Y(_0749_));
 sg13g2_a221oi_1 _2716_ (.B2(_0742_),
    .C1(net404),
    .B1(_0749_),
    .A1(_0983_),
    .Y(_0202_),
    .A2(_0746_));
 sg13g2_nand2_1 _2717_ (.Y(_0750_),
    .A(net462),
    .B(_0743_));
 sg13g2_a21oi_1 _2718_ (.A1(_0053_),
    .A2(_0748_),
    .Y(_0751_),
    .B1(_0743_));
 sg13g2_nand3_1 _2719_ (.B(_0744_),
    .C(_0751_),
    .A(_0585_),
    .Y(_0752_));
 sg13g2_a21oi_1 _2720_ (.A1(_0750_),
    .A2(_0752_),
    .Y(_0203_),
    .B1(net404));
 sg13g2_nand2_1 _2721_ (.Y(_0753_),
    .A(\modem.uart.txFifo.nextIn[0] ),
    .B(_0458_));
 sg13g2_nor2b_1 _2722_ (.A(net439),
    .B_N(\modem.uart.txFifo.nextIn[1] ),
    .Y(_0754_));
 sg13g2_nand3_1 _2723_ (.B(_0458_),
    .C(_0754_),
    .A(\modem.uart.txFifo.nextIn[0] ),
    .Y(_0755_));
 sg13g2_nand2_1 _2724_ (.Y(_0756_),
    .A(net511),
    .B(net357));
 sg13g2_o21ai_1 _2725_ (.B1(_0756_),
    .Y(_0204_),
    .A1(_0980_),
    .A2(net357));
 sg13g2_nand2_1 _2726_ (.Y(_0757_),
    .A(net491),
    .B(net357));
 sg13g2_o21ai_1 _2727_ (.B1(_0757_),
    .Y(_0205_),
    .A1(_0979_),
    .A2(net357));
 sg13g2_nand2_1 _2728_ (.Y(_0758_),
    .A(net525),
    .B(net357));
 sg13g2_o21ai_1 _2729_ (.B1(_0758_),
    .Y(_0206_),
    .A1(_0978_),
    .A2(net357));
 sg13g2_nand2_1 _2730_ (.Y(_0759_),
    .A(net503),
    .B(net358));
 sg13g2_o21ai_1 _2731_ (.B1(_0759_),
    .Y(_0207_),
    .A1(_0977_),
    .A2(net357));
 sg13g2_nand2_1 _2732_ (.Y(_0760_),
    .A(net470),
    .B(net359));
 sg13g2_o21ai_1 _2733_ (.B1(_0760_),
    .Y(_0208_),
    .A1(_0976_),
    .A2(net359));
 sg13g2_nand2_1 _2734_ (.Y(_0761_),
    .A(net464),
    .B(net357));
 sg13g2_o21ai_1 _2735_ (.B1(_0761_),
    .Y(_0209_),
    .A1(_0975_),
    .A2(net358));
 sg13g2_nand2_1 _2736_ (.Y(_0762_),
    .A(net478),
    .B(net358));
 sg13g2_o21ai_1 _2737_ (.B1(_0762_),
    .Y(_0210_),
    .A1(_0974_),
    .A2(net358));
 sg13g2_nand2_1 _2738_ (.Y(_0763_),
    .A(net472),
    .B(net359));
 sg13g2_o21ai_1 _2739_ (.B1(_0763_),
    .Y(_0211_),
    .A1(_0973_),
    .A2(net359));
 sg13g2_o21ai_1 _2740_ (.B1(net452),
    .Y(_0764_),
    .A1(net458),
    .A2(_0459_));
 sg13g2_a21oi_1 _2741_ (.A1(_0982_),
    .A2(_0459_),
    .Y(_0212_),
    .B1(_0764_));
 sg13g2_xor2_1 _2742_ (.B(_0753_),
    .A(net838),
    .X(_0765_));
 sg13g2_nor2_1 _2743_ (.A(net408),
    .B(net839),
    .Y(_0213_));
 sg13g2_o21ai_1 _2744_ (.B1(net452),
    .Y(_0766_),
    .A1(\modem.uart.txFifo.nextOut[0] ),
    .A2(_1206_));
 sg13g2_a21oi_1 _2745_ (.A1(_0981_),
    .A2(_1206_),
    .Y(_0214_),
    .B1(_0766_));
 sg13g2_and3_1 _2746_ (.X(_0767_),
    .A(net420),
    .B(\modem.uart.txFifo.nextOut[0] ),
    .C(_1206_));
 sg13g2_a21oi_1 _2747_ (.A1(net886),
    .A2(_1206_),
    .Y(_0768_),
    .B1(net420));
 sg13g2_nor3_1 _2748_ (.A(net407),
    .B(_0767_),
    .C(net887),
    .Y(_0215_));
 sg13g2_nand3_1 _2749_ (.B(_0458_),
    .C(_0754_),
    .A(_0982_),
    .Y(_0769_));
 sg13g2_nand2_1 _2750_ (.Y(_0770_),
    .A(net468),
    .B(net354));
 sg13g2_o21ai_1 _2751_ (.B1(_0770_),
    .Y(_0216_),
    .A1(_0980_),
    .A2(net354));
 sg13g2_nand2_1 _2752_ (.Y(_0771_),
    .A(net507),
    .B(net354));
 sg13g2_o21ai_1 _2753_ (.B1(_0771_),
    .Y(_0217_),
    .A1(_0979_),
    .A2(net354));
 sg13g2_nand2_1 _2754_ (.Y(_0772_),
    .A(net480),
    .B(net354));
 sg13g2_o21ai_1 _2755_ (.B1(_0772_),
    .Y(_0218_),
    .A1(_0978_),
    .A2(net355));
 sg13g2_nand2_1 _2756_ (.Y(_0773_),
    .A(net532),
    .B(net354));
 sg13g2_o21ai_1 _2757_ (.B1(_0773_),
    .Y(_0219_),
    .A1(_0977_),
    .A2(net355));
 sg13g2_nand2_1 _2758_ (.Y(_0774_),
    .A(net485),
    .B(net356));
 sg13g2_o21ai_1 _2759_ (.B1(_0774_),
    .Y(_0220_),
    .A1(_0976_),
    .A2(net356));
 sg13g2_nand2_1 _2760_ (.Y(_0775_),
    .A(net476),
    .B(net354));
 sg13g2_o21ai_1 _2761_ (.B1(_0775_),
    .Y(_0221_),
    .A1(_0975_),
    .A2(net355));
 sg13g2_nand2_1 _2762_ (.Y(_0776_),
    .A(net483),
    .B(net354));
 sg13g2_o21ai_1 _2763_ (.B1(_0776_),
    .Y(_0222_),
    .A1(_0974_),
    .A2(net355));
 sg13g2_nand2_1 _2764_ (.Y(_0777_),
    .A(net474),
    .B(net356));
 sg13g2_o21ai_1 _2765_ (.B1(_0777_),
    .Y(_0223_),
    .A1(_0973_),
    .A2(net356));
 sg13g2_nor3_1 _2766_ (.A(\modem.uart.txFifo.nextIn[1] ),
    .B(net439),
    .C(_0753_),
    .Y(_0778_));
 sg13g2_nor2_1 _2767_ (.A(net561),
    .B(net349),
    .Y(_0779_));
 sg13g2_a21oi_1 _2768_ (.A1(_0980_),
    .A2(net349),
    .Y(_0224_),
    .B1(_0779_));
 sg13g2_nor2_1 _2769_ (.A(net711),
    .B(net349),
    .Y(_0780_));
 sg13g2_a21oi_1 _2770_ (.A1(_0979_),
    .A2(_0778_),
    .Y(_0225_),
    .B1(_0780_));
 sg13g2_nor2_1 _2771_ (.A(net664),
    .B(net349),
    .Y(_0781_));
 sg13g2_a21oi_1 _2772_ (.A1(_0978_),
    .A2(net349),
    .Y(_0226_),
    .B1(_0781_));
 sg13g2_nor2_1 _2773_ (.A(net595),
    .B(net349),
    .Y(_0782_));
 sg13g2_a21oi_1 _2774_ (.A1(_0977_),
    .A2(net349),
    .Y(_0227_),
    .B1(_0782_));
 sg13g2_nor2_1 _2775_ (.A(net647),
    .B(net350),
    .Y(_0783_));
 sg13g2_a21oi_1 _2776_ (.A1(_0976_),
    .A2(net350),
    .Y(_0228_),
    .B1(_0783_));
 sg13g2_nor2_1 _2777_ (.A(net569),
    .B(net349),
    .Y(_0784_));
 sg13g2_a21oi_1 _2778_ (.A1(_0975_),
    .A2(net350),
    .Y(_0229_),
    .B1(_0784_));
 sg13g2_nor2_1 _2779_ (.A(net581),
    .B(net350),
    .Y(_0785_));
 sg13g2_a21oi_1 _2780_ (.A1(_0974_),
    .A2(net350),
    .Y(_0230_),
    .B1(_0785_));
 sg13g2_nor2_1 _2781_ (.A(net748),
    .B(net350),
    .Y(_0786_));
 sg13g2_a21oi_1 _2782_ (.A1(_0973_),
    .A2(net350),
    .Y(_0231_),
    .B1(_0786_));
 sg13g2_nor3_1 _2783_ (.A(\modem.uart.txFifo.nextIn[1] ),
    .B(\modem.uart.txFifo.nextIn[0] ),
    .C(_0459_),
    .Y(_0787_));
 sg13g2_o21ai_1 _2784_ (.B1(net453),
    .Y(_0788_),
    .A1(net767),
    .A2(net351));
 sg13g2_a21oi_1 _2785_ (.A1(_0980_),
    .A2(net351),
    .Y(_0232_),
    .B1(_0788_));
 sg13g2_o21ai_1 _2786_ (.B1(net453),
    .Y(_0789_),
    .A1(net734),
    .A2(net352));
 sg13g2_a21oi_1 _2787_ (.A1(_0979_),
    .A2(net352),
    .Y(_0233_),
    .B1(_0789_));
 sg13g2_o21ai_1 _2788_ (.B1(net452),
    .Y(_0790_),
    .A1(net708),
    .A2(net351));
 sg13g2_a21oi_1 _2789_ (.A1(_0978_),
    .A2(net351),
    .Y(_0234_),
    .B1(_0790_));
 sg13g2_o21ai_1 _2790_ (.B1(net453),
    .Y(_0791_),
    .A1(net765),
    .A2(net352));
 sg13g2_a21oi_1 _2791_ (.A1(_0977_),
    .A2(net352),
    .Y(_0235_),
    .B1(_0791_));
 sg13g2_o21ai_1 _2792_ (.B1(net453),
    .Y(_0792_),
    .A1(net746),
    .A2(net353));
 sg13g2_a21oi_1 _2793_ (.A1(_0976_),
    .A2(net353),
    .Y(_0236_),
    .B1(_0792_));
 sg13g2_o21ai_1 _2794_ (.B1(net453),
    .Y(_0793_),
    .A1(net792),
    .A2(net351));
 sg13g2_a21oi_1 _2795_ (.A1(_0975_),
    .A2(net351),
    .Y(_0237_),
    .B1(_0793_));
 sg13g2_o21ai_1 _2796_ (.B1(net453),
    .Y(_0794_),
    .A1(net763),
    .A2(net351));
 sg13g2_a21oi_1 _2797_ (.A1(_0974_),
    .A2(net351),
    .Y(_0238_),
    .B1(_0794_));
 sg13g2_o21ai_1 _2798_ (.B1(net452),
    .Y(_0795_),
    .A1(net718),
    .A2(net353));
 sg13g2_a21oi_1 _2799_ (.A1(_0973_),
    .A2(net353),
    .Y(_0239_),
    .B1(_0795_));
 sg13g2_nor2_1 _2800_ (.A(_1206_),
    .B(_0459_),
    .Y(_0796_));
 sg13g2_xnor2_1 _2801_ (.Y(_0797_),
    .A(_1206_),
    .B(_0459_));
 sg13g2_o21ai_1 _2802_ (.B1(net452),
    .Y(_0798_),
    .A1(\modem.uart.txFifo.count[0] ),
    .A2(_0797_));
 sg13g2_a21oi_1 _2803_ (.A1(_0972_),
    .A2(_0797_),
    .Y(_0240_),
    .B1(_0798_));
 sg13g2_nand2_1 _2804_ (.Y(_0799_),
    .A(\modem.uart.txFifo.count[1] ),
    .B(\modem.uart.rxHdlc.io_valid ));
 sg13g2_o21ai_1 _2805_ (.B1(_0799_),
    .Y(_0800_),
    .A1(\modem.uart.txFifo.count[1] ),
    .A2(_0458_));
 sg13g2_xnor2_1 _2806_ (.Y(_0801_),
    .A(_0972_),
    .B(_0800_));
 sg13g2_o21ai_1 _2807_ (.B1(net452),
    .Y(_0802_),
    .A1(net819),
    .A2(_0797_));
 sg13g2_a21oi_1 _2808_ (.A1(_0797_),
    .A2(_0801_),
    .Y(_0241_),
    .B1(_0802_));
 sg13g2_nand3_1 _2809_ (.B(_1206_),
    .C(_0459_),
    .A(_1201_),
    .Y(_0803_));
 sg13g2_nand3_1 _2810_ (.B(\modem.uart.txFifo.count[0] ),
    .C(_0796_),
    .A(\modem.uart.txFifo.count[1] ),
    .Y(_0804_));
 sg13g2_nand2_1 _2811_ (.Y(_0805_),
    .A(_0803_),
    .B(_0804_));
 sg13g2_o21ai_1 _2812_ (.B1(net452),
    .Y(_0806_),
    .A1(net624),
    .A2(_0805_));
 sg13g2_a21oi_1 _2813_ (.A1(net624),
    .A2(_0805_),
    .Y(_0242_),
    .B1(_0806_));
 sg13g2_nor3_1 _2814_ (.A(_1003_),
    .B(_1031_),
    .C(_1213_),
    .Y(_0807_));
 sg13g2_nor3_2 _2815_ (.A(\modem.uart.rxHdlc.fsmHdlcRx_bit[0] ),
    .B(\modem.uart.rxHdlc.fsmHdlcRx_bit[1] ),
    .C(net707),
    .Y(_0808_));
 sg13g2_nand2_1 _2816_ (.Y(_0809_),
    .A(_0807_),
    .B(_0808_));
 sg13g2_mux2_1 _2817_ (.A0(_1208_),
    .A1(net509),
    .S(_0809_),
    .X(_0244_));
 sg13g2_o21ai_1 _2818_ (.B1(\modem.uart.rxHdlc.fsmHdlcRx_bit[2] ),
    .Y(_0810_),
    .A1(\modem.uart.rxHdlc.fsmHdlcRx_bit[0] ),
    .A2(\modem.uart.rxHdlc.fsmHdlcRx_bit[1] ));
 sg13g2_and2_1 _2819_ (.A(_0807_),
    .B(_0810_),
    .X(_0811_));
 sg13g2_nor2b_1 _2820_ (.A(_0808_),
    .B_N(_0811_),
    .Y(_0812_));
 sg13g2_nor2_1 _2821_ (.A(net684),
    .B(_0418_),
    .Y(_0813_));
 sg13g2_nand2_1 _2822_ (.Y(_0814_),
    .A(_0812_),
    .B(_0813_));
 sg13g2_nor2b_2 _2823_ (.A(_0808_),
    .B_N(_1208_),
    .Y(_0815_));
 sg13g2_mux2_1 _2824_ (.A0(_0815_),
    .A1(net620),
    .S(_0814_),
    .X(_0245_));
 sg13g2_nor2b_1 _2825_ (.A(\modem.uart.rxHdlc.fsmHdlcRx_bit[0] ),
    .B_N(\modem.uart.rxHdlc.fsmHdlcRx_bit[1] ),
    .Y(_0816_));
 sg13g2_nand2_1 _2826_ (.Y(_0817_),
    .A(_0811_),
    .B(net686));
 sg13g2_mux2_1 _2827_ (.A0(_0815_),
    .A1(net513),
    .S(_0817_),
    .X(_0246_));
 sg13g2_nand3_1 _2828_ (.B(_0418_),
    .C(_0812_),
    .A(_0997_),
    .Y(_0818_));
 sg13g2_mux2_1 _2829_ (.A0(_0815_),
    .A1(net516),
    .S(_0818_),
    .X(_0247_));
 sg13g2_and2_1 _2830_ (.A(net787),
    .B(_0807_),
    .X(_0819_));
 sg13g2_nand2_1 _2831_ (.Y(_0820_),
    .A(net689),
    .B(_0811_));
 sg13g2_mux2_1 _2832_ (.A0(_1208_),
    .A1(net553),
    .S(_0820_),
    .X(_0248_));
 sg13g2_nand2_1 _2833_ (.Y(_0821_),
    .A(_0813_),
    .B(_0819_));
 sg13g2_mux2_1 _2834_ (.A0(_0815_),
    .A1(net563),
    .S(_0821_),
    .X(_0249_));
 sg13g2_nand2_1 _2835_ (.Y(_0822_),
    .A(net686),
    .B(_0819_));
 sg13g2_mux2_1 _2836_ (.A0(_0815_),
    .A1(net587),
    .S(_0822_),
    .X(_0250_));
 sg13g2_o21ai_1 _2837_ (.B1(_1217_),
    .Y(_0251_),
    .A1(_1026_),
    .A2(net366));
 sg13g2_o21ai_1 _2838_ (.B1(net366),
    .Y(_0823_),
    .A1(_0061_),
    .A2(_1216_));
 sg13g2_a21oi_1 _2839_ (.A1(net431),
    .A2(net321),
    .Y(_0824_),
    .B1(_0823_));
 sg13g2_a21oi_1 _2840_ (.A1(_1007_),
    .A2(net368),
    .Y(_0252_),
    .B1(net322));
 sg13g2_xnor2_1 _2841_ (.Y(_0825_),
    .A(\modem.uart.rxHdlc.oneBitCount[0] ),
    .B(net824));
 sg13g2_nand2_1 _2842_ (.Y(_0826_),
    .A(net824),
    .B(_0823_));
 sg13g2_o21ai_1 _2843_ (.B1(net825),
    .Y(_0253_),
    .A1(_1217_),
    .A2(_0825_));
 sg13g2_nor2_1 _2844_ (.A(_1214_),
    .B(_0823_),
    .Y(_0827_));
 sg13g2_nor2_1 _2845_ (.A(net431),
    .B(_0823_),
    .Y(_0828_));
 sg13g2_xnor2_1 _2846_ (.Y(_0829_),
    .A(net697),
    .B(_0827_));
 sg13g2_nor2_1 _2847_ (.A(_0828_),
    .B(net698),
    .Y(_0254_));
 sg13g2_and3_1 _2848_ (.X(_0830_),
    .A(_0067_),
    .B(net367),
    .C(_1227_));
 sg13g2_nand2_1 _2849_ (.Y(_0831_),
    .A(net509),
    .B(net347));
 sg13g2_o21ai_1 _2850_ (.B1(_0831_),
    .Y(_0255_),
    .A1(_0980_),
    .A2(net348));
 sg13g2_nand2_1 _2851_ (.Y(_0832_),
    .A(net620),
    .B(net347));
 sg13g2_o21ai_1 _2852_ (.B1(_0832_),
    .Y(_0256_),
    .A1(_0979_),
    .A2(net348));
 sg13g2_nand2_1 _2853_ (.Y(_0833_),
    .A(net513),
    .B(net347));
 sg13g2_o21ai_1 _2854_ (.B1(_0833_),
    .Y(_0257_),
    .A1(_0978_),
    .A2(net347));
 sg13g2_nand2_1 _2855_ (.Y(_0834_),
    .A(net516),
    .B(net347));
 sg13g2_o21ai_1 _2856_ (.B1(_0834_),
    .Y(_0258_),
    .A1(_0977_),
    .A2(net347));
 sg13g2_nand2_1 _2857_ (.Y(_0835_),
    .A(net553),
    .B(net348));
 sg13g2_o21ai_1 _2858_ (.B1(_0835_),
    .Y(_0259_),
    .A1(_0976_),
    .A2(net348));
 sg13g2_nand2_1 _2859_ (.Y(_0836_),
    .A(net563),
    .B(net347));
 sg13g2_o21ai_1 _2860_ (.B1(_0836_),
    .Y(_0260_),
    .A1(_0975_),
    .A2(_0830_));
 sg13g2_nand2_1 _2861_ (.Y(_0837_),
    .A(net587),
    .B(net347));
 sg13g2_o21ai_1 _2862_ (.B1(_0837_),
    .Y(_0261_),
    .A1(_0974_),
    .A2(net348));
 sg13g2_nand2_1 _2863_ (.Y(_0838_),
    .A(_1208_),
    .B(net348));
 sg13g2_o21ai_1 _2864_ (.B1(_0838_),
    .Y(_0262_),
    .A1(_0973_),
    .A2(net348));
 sg13g2_nand3_1 _2865_ (.B(net441),
    .C(_0466_),
    .A(\modem.uart.rxFifo.nextIn[2] ),
    .Y(_0839_));
 sg13g2_nand2_1 _2866_ (.Y(_0840_),
    .A(net466),
    .B(net363));
 sg13g2_o21ai_1 _2867_ (.B1(_0840_),
    .Y(_0263_),
    .A1(net409),
    .A2(net363));
 sg13g2_nand2_1 _2868_ (.Y(_0841_),
    .A(net330),
    .B(net362));
 sg13g2_o21ai_1 _2869_ (.B1(_0841_),
    .Y(_0264_),
    .A1(_0992_),
    .A2(net361));
 sg13g2_nand2_1 _2870_ (.Y(_0842_),
    .A(net338),
    .B(net363));
 sg13g2_o21ai_1 _2871_ (.B1(_0842_),
    .Y(_0265_),
    .A1(_0991_),
    .A2(net363));
 sg13g2_nand2_1 _2872_ (.Y(_0843_),
    .A(net460),
    .B(net361));
 sg13g2_o21ai_1 _2873_ (.B1(_0843_),
    .Y(_0266_),
    .A1(net410),
    .A2(net361));
 sg13g2_nand2_1 _2874_ (.Y(_0844_),
    .A(net328),
    .B(net361));
 sg13g2_o21ai_1 _2875_ (.B1(_0844_),
    .Y(_0267_),
    .A1(_0989_),
    .A2(net361));
 sg13g2_nand2_1 _2876_ (.Y(_0845_),
    .A(net326),
    .B(net362));
 sg13g2_o21ai_1 _2877_ (.B1(_0845_),
    .Y(_0268_),
    .A1(_0988_),
    .A2(net362));
 sg13g2_nand2_1 _2878_ (.Y(_0846_),
    .A(net336),
    .B(net361));
 sg13g2_o21ai_1 _2879_ (.B1(_0846_),
    .Y(_0269_),
    .A1(_0987_),
    .A2(net361));
 sg13g2_nand2_1 _2880_ (.Y(_0847_),
    .A(net334),
    .B(net362));
 sg13g2_o21ai_1 _2881_ (.B1(_0847_),
    .Y(_0270_),
    .A1(_0986_),
    .A2(net361));
 sg13g2_a221oi_1 _2882_ (.B2(_1143_),
    .C1(net401),
    .B1(_1133_),
    .A1(_0999_),
    .Y(_0848_),
    .A2(_1000_));
 sg13g2_a21o_1 _2883_ (.A2(_0848_),
    .A1(net442),
    .B1(_1043_),
    .X(_0271_));
 sg13g2_o21ai_1 _2884_ (.B1(\modem.uart.rxUart.fsmUartRx_stateReg[5] ),
    .Y(_0849_),
    .A1(net419),
    .A2(_1162_));
 sg13g2_nand2b_1 _2885_ (.Y(_0850_),
    .B(_0049_),
    .A_N(\modem.uart.rxUart.fsmUartRx_stateReg[1] ));
 sg13g2_and3_2 _2886_ (.X(_0851_),
    .A(_1236_),
    .B(_0849_),
    .C(_0850_));
 sg13g2_nand3_1 _2887_ (.B(net497),
    .C(_0851_),
    .A(\modem.uart.rxUart.fsmUartRx_stateReg[1] ),
    .Y(_0852_));
 sg13g2_o21ai_1 _2888_ (.B1(net498),
    .Y(_0272_),
    .A1(_1005_),
    .A2(_0851_));
 sg13g2_nand3_1 _2889_ (.B(_0440_),
    .C(_0851_),
    .A(net807),
    .Y(_0853_));
 sg13g2_o21ai_1 _2890_ (.B1(_0853_),
    .Y(_0273_),
    .A1(_1020_),
    .A2(_0851_));
 sg13g2_xnor2_1 _2891_ (.Y(_0854_),
    .A(\modem.uart.rxUart.bitId[2] ),
    .B(_1234_));
 sg13g2_nand3_1 _2892_ (.B(_0851_),
    .C(_0854_),
    .A(net807),
    .Y(_0855_));
 sg13g2_o21ai_1 _2893_ (.B1(net808),
    .Y(_0274_),
    .A1(_1021_),
    .A2(_0851_));
 sg13g2_xnor2_1 _2894_ (.Y(_0856_),
    .A(net2),
    .B(\modem.control.zeroCrossDet_7 ));
 sg13g2_xor2_1 _2895_ (.B(\modem.control.zeroCrossDet_7 ),
    .A(net2),
    .X(_0857_));
 sg13g2_o21ai_1 _2896_ (.B1(net451),
    .Y(_0858_),
    .A1(_0036_),
    .A2(_0856_));
 sg13g2_a21oi_1 _2897_ (.A1(_0970_),
    .A2(_0856_),
    .Y(_0275_),
    .B1(_0858_));
 sg13g2_nor2_1 _2898_ (.A(\modem.control.rxAddr[5] ),
    .B(_1028_),
    .Y(_0859_));
 sg13g2_xnor2_1 _2899_ (.Y(_0860_),
    .A(\modem.control.rxAddr[5] ),
    .B(_1028_));
 sg13g2_nor3_1 _2900_ (.A(net827),
    .B(_0856_),
    .C(_0860_),
    .Y(_0861_));
 sg13g2_and3_1 _2901_ (.X(_0862_),
    .A(net827),
    .B(net395),
    .C(_0860_));
 sg13g2_o21ai_1 _2902_ (.B1(net450),
    .Y(_0863_),
    .A1(\modem.control.rxAddr[5] ),
    .A2(net395));
 sg13g2_nor3_1 _2903_ (.A(_0861_),
    .B(_0862_),
    .C(_0863_),
    .Y(_0276_));
 sg13g2_a21oi_1 _2904_ (.A1(\modem.control.rxAddr[5] ),
    .A2(net369),
    .Y(_0864_),
    .B1(net622));
 sg13g2_xnor2_1 _2905_ (.Y(_0865_),
    .A(net796),
    .B(net369));
 sg13g2_nor3_1 _2906_ (.A(_0859_),
    .B(_0864_),
    .C(_0865_),
    .Y(_0866_));
 sg13g2_o21ai_1 _2907_ (.B1(_0865_),
    .Y(_0867_),
    .A1(_0859_),
    .A2(_0864_));
 sg13g2_nand2b_1 _2908_ (.Y(_0868_),
    .B(_0867_),
    .A_N(_0866_));
 sg13g2_o21ai_1 _2909_ (.B1(net450),
    .Y(_0869_),
    .A1(net796),
    .A2(net394));
 sg13g2_a21oi_1 _2910_ (.A1(net394),
    .A2(_0868_),
    .Y(_0277_),
    .B1(_0869_));
 sg13g2_a21oi_1 _2911_ (.A1(_1014_),
    .A2(net369),
    .Y(_0870_),
    .B1(_0866_));
 sg13g2_xnor2_1 _2912_ (.Y(_0871_),
    .A(net804),
    .B(\modem.control.io_upDownOut ));
 sg13g2_nand2b_1 _2913_ (.Y(_0872_),
    .B(_0871_),
    .A_N(_0870_));
 sg13g2_xor2_1 _2914_ (.B(_0871_),
    .A(_0870_),
    .X(_0873_));
 sg13g2_o21ai_1 _2915_ (.B1(net450),
    .Y(_0874_),
    .A1(net804),
    .A2(net395));
 sg13g2_a21oi_1 _2916_ (.A1(net395),
    .A2(_0873_),
    .Y(_0278_),
    .B1(_0874_));
 sg13g2_o21ai_1 _2917_ (.B1(_0872_),
    .Y(_0875_),
    .A1(_0034_),
    .A2(net360));
 sg13g2_xnor2_1 _2918_ (.Y(_0876_),
    .A(net847),
    .B(net360));
 sg13g2_xnor2_1 _2919_ (.Y(_0877_),
    .A(_0875_),
    .B(_0876_));
 sg13g2_o21ai_1 _2920_ (.B1(net450),
    .Y(_0878_),
    .A1(net847),
    .A2(net394));
 sg13g2_a21oi_1 _2921_ (.A1(net394),
    .A2(_0877_),
    .Y(_0279_),
    .B1(_0878_));
 sg13g2_a22oi_1 _2922_ (.Y(_0879_),
    .B1(_0875_),
    .B2(_0876_),
    .A2(net369),
    .A1(_1016_));
 sg13g2_xnor2_1 _2923_ (.Y(_0880_),
    .A(net797),
    .B(net360));
 sg13g2_nor2b_1 _2924_ (.A(_0879_),
    .B_N(_0880_),
    .Y(_0881_));
 sg13g2_xor2_1 _2925_ (.B(_0880_),
    .A(_0879_),
    .X(_0882_));
 sg13g2_o21ai_1 _2926_ (.B1(net447),
    .Y(_0883_),
    .A1(net797),
    .A2(net394));
 sg13g2_a21oi_1 _2927_ (.A1(net394),
    .A2(_0882_),
    .Y(_0280_),
    .B1(_0883_));
 sg13g2_nor2_1 _2928_ (.A(_0032_),
    .B(net360),
    .Y(_0884_));
 sg13g2_xnor2_1 _2929_ (.Y(_0885_),
    .A(\modem.control.rxAddr[10] ),
    .B(net360));
 sg13g2_o21ai_1 _2930_ (.B1(_0885_),
    .Y(_0886_),
    .A1(_0881_),
    .A2(_0884_));
 sg13g2_or3_1 _2931_ (.A(_0881_),
    .B(_0884_),
    .C(_0885_),
    .X(_0887_));
 sg13g2_nand2_1 _2932_ (.Y(_0888_),
    .A(_0886_),
    .B(_0887_));
 sg13g2_o21ai_1 _2933_ (.B1(net450),
    .Y(_0889_),
    .A1(net856),
    .A2(net394));
 sg13g2_a21oi_1 _2934_ (.A1(net394),
    .A2(_0888_),
    .Y(_0281_),
    .B1(_0889_));
 sg13g2_nand3_1 _2935_ (.B(net360),
    .C(_0881_),
    .A(\modem.control.rxAddr[10] ),
    .Y(_0890_));
 sg13g2_nand3_1 _2936_ (.B(net369),
    .C(_0886_),
    .A(_0031_),
    .Y(_0891_));
 sg13g2_a21o_1 _2937_ (.A2(_0891_),
    .A1(_0890_),
    .B1(_0856_),
    .X(_0892_));
 sg13g2_a21oi_1 _2938_ (.A1(net633),
    .A2(_0892_),
    .Y(_0893_),
    .B1(net407));
 sg13g2_o21ai_1 _2939_ (.B1(_0893_),
    .Y(_0282_),
    .A1(net633),
    .A2(_0892_));
 sg13g2_a21oi_1 _2940_ (.A1(_1017_),
    .A2(\latched[3] ),
    .Y(_0894_),
    .B1(\latched[15] ));
 sg13g2_o21ai_1 _2941_ (.B1(_0894_),
    .Y(_0895_),
    .A1(net432),
    .A2(\latched[3] ));
 sg13g2_nor2b_1 _2942_ (.A(\modem.control._zz_txClockInternalFallStb_regNext ),
    .B_N(net318),
    .Y(_0896_));
 sg13g2_xor2_1 _2943_ (.B(_0895_),
    .A(\latched[14] ),
    .X(_0897_));
 sg13g2_o21ai_1 _2944_ (.B1(net446),
    .Y(_0898_),
    .A1(net820),
    .A2(_0896_));
 sg13g2_a21oi_1 _2945_ (.A1(_0896_),
    .A2(_0897_),
    .Y(_0283_),
    .B1(net821));
 sg13g2_o21ai_1 _2946_ (.B1(net449),
    .Y(_0899_),
    .A1(\modem.control.rxAddr[0] ),
    .A2(_0333_));
 sg13g2_a21oi_1 _2947_ (.A1(_0968_),
    .A2(_0333_),
    .Y(_0284_),
    .B1(_0899_));
 sg13g2_a21oi_1 _2948_ (.A1(\modem.control.rxAddr[0] ),
    .A2(_0333_),
    .Y(_0900_),
    .B1(net546));
 sg13g2_nand3_1 _2949_ (.B(net889),
    .C(_0333_),
    .A(net546),
    .Y(_0901_));
 sg13g2_nand2_1 _2950_ (.Y(_0902_),
    .A(net449),
    .B(_0901_));
 sg13g2_nor2_1 _2951_ (.A(net547),
    .B(_0902_),
    .Y(_0285_));
 sg13g2_nor2_1 _2952_ (.A(_0944_),
    .B(_0901_),
    .Y(_0903_));
 sg13g2_a21oi_1 _2953_ (.A1(_0944_),
    .A2(_0901_),
    .Y(_0904_),
    .B1(net407));
 sg13g2_nor2b_1 _2954_ (.A(_0903_),
    .B_N(_0904_),
    .Y(_0286_));
 sg13g2_a21oi_1 _2955_ (.A1(net318),
    .A2(_0903_),
    .Y(_0905_),
    .B1(net407));
 sg13g2_o21ai_1 _2956_ (.B1(_0905_),
    .Y(_0906_),
    .A1(net318),
    .A2(_0903_));
 sg13g2_inv_1 _2957_ (.Y(_0287_),
    .A(_0906_));
 sg13g2_and2_1 _2958_ (.A(net448),
    .B(net304),
    .X(_0288_));
 sg13g2_and3_1 _2959_ (.X(_0289_),
    .A(net450),
    .B(_0332_),
    .C(_0334_));
 sg13g2_nor3_1 _2960_ (.A(net414),
    .B(net412),
    .C(net315),
    .Y(_0907_));
 sg13g2_xnor2_1 _2961_ (.Y(_0908_),
    .A(net315),
    .B(_0330_));
 sg13g2_nor2_1 _2962_ (.A(net407),
    .B(_0908_),
    .Y(_0290_));
 sg13g2_nor2b_1 _2963_ (.A(net713),
    .B_N(_0907_),
    .Y(_0909_));
 sg13g2_xnor2_1 _2964_ (.Y(_0910_),
    .A(net713),
    .B(_0907_));
 sg13g2_nor2_1 _2965_ (.A(net407),
    .B(net714),
    .Y(_0291_));
 sg13g2_xnor2_1 _2966_ (.Y(_0911_),
    .A(net302),
    .B(_0909_));
 sg13g2_nor2_1 _2967_ (.A(net407),
    .B(_0911_),
    .Y(_0292_));
 sg13g2_nand3_1 _2968_ (.B(net309),
    .C(_0909_),
    .A(_1022_),
    .Y(_0912_));
 sg13g2_a21oi_1 _2969_ (.A1(_1022_),
    .A2(_0909_),
    .Y(_0913_),
    .B1(net309));
 sg13g2_nor2_1 _2970_ (.A(net407),
    .B(_0913_),
    .Y(_0914_));
 sg13g2_and2_1 _2971_ (.A(_0912_),
    .B(_0914_),
    .X(_0293_));
 sg13g2_nand2_1 _2972_ (.Y(_0915_),
    .A(\latched[12] ),
    .B(_0330_));
 sg13g2_o21ai_1 _2973_ (.B1(_0915_),
    .Y(_0916_),
    .A1(\latched[12] ),
    .A2(_0334_));
 sg13g2_mux2_1 _2974_ (.A0(net583),
    .A1(\modem.control.rxRcrDacTmp[3] ),
    .S(_0916_),
    .X(_0294_));
 sg13g2_nand2_1 _2975_ (.Y(_0917_),
    .A(\latched[12] ),
    .B(_0333_));
 sg13g2_o21ai_1 _2976_ (.B1(_0917_),
    .Y(_0918_),
    .A1(\latched[12] ),
    .A2(_0332_));
 sg13g2_mux2_1 _2977_ (.A0(net650),
    .A1(net6),
    .S(_0918_),
    .X(_0295_));
 sg13g2_mux2_1 _2978_ (.A0(net2),
    .A1(net618),
    .S(net627),
    .X(_0296_));
 sg13g2_mux2_1 _2979_ (.A0(net618),
    .A1(\modem.control.zeroCrossDet_1 ),
    .S(_1165_),
    .X(_0297_));
 sg13g2_mux2_1 _2980_ (.A0(net646),
    .A1(net639),
    .S(net627),
    .X(_0298_));
 sg13g2_mux2_1 _2981_ (.A0(net639),
    .A1(\modem.control.zeroCrossDet_3 ),
    .S(net627),
    .X(_0299_));
 sg13g2_mux2_1 _2982_ (.A0(net643),
    .A1(net599),
    .S(net627),
    .X(_0300_));
 sg13g2_mux2_1 _2983_ (.A0(net599),
    .A1(\modem.control.zeroCrossDet_5 ),
    .S(_1165_),
    .X(_0301_));
 sg13g2_mux2_1 _2984_ (.A0(net635),
    .A1(\modem.control.zeroCrossDet_5 ),
    .S(\modem.control.io_txClockStb ),
    .X(_0302_));
 sg13g2_nor2b_1 _2985_ (.A(\modem.control._zz_txClockInternalFallStb ),
    .B_N(\modem.control._zz_txClockInternalFallStb_regNext ),
    .Y(_0919_));
 sg13g2_o21ai_1 _2986_ (.B1(net448),
    .Y(_0920_),
    .A1(\modem.control.scrambler_1.io_vecOut[1] ),
    .A2(net392));
 sg13g2_a21oi_1 _2987_ (.A1(_0965_),
    .A2(net392),
    .Y(_0303_),
    .B1(_0920_));
 sg13g2_o21ai_1 _2988_ (.B1(net449),
    .Y(_0921_),
    .A1(net700),
    .A2(net391));
 sg13g2_a21oi_1 _2989_ (.A1(_0964_),
    .A2(net391),
    .Y(_0304_),
    .B1(_0921_));
 sg13g2_o21ai_1 _2990_ (.B1(net449),
    .Y(_0922_),
    .A1(net690),
    .A2(net391));
 sg13g2_a21oi_1 _2991_ (.A1(_0963_),
    .A2(net391),
    .Y(_0305_),
    .B1(_0922_));
 sg13g2_o21ai_1 _2992_ (.B1(net449),
    .Y(_0923_),
    .A1(net670),
    .A2(net391));
 sg13g2_a21oi_1 _2993_ (.A1(_0962_),
    .A2(net391),
    .Y(_0306_),
    .B1(_0923_));
 sg13g2_o21ai_1 _2994_ (.B1(net449),
    .Y(_0924_),
    .A1(net555),
    .A2(net391));
 sg13g2_a21oi_1 _2995_ (.A1(_0961_),
    .A2(net393),
    .Y(_0307_),
    .B1(_0924_));
 sg13g2_o21ai_1 _2996_ (.B1(net448),
    .Y(_0925_),
    .A1(\modem.control.scrambler_1.io_vecOut[6] ),
    .A2(net393));
 sg13g2_a21oi_1 _2997_ (.A1(_0960_),
    .A2(net391),
    .Y(_0308_),
    .B1(_0925_));
 sg13g2_o21ai_1 _2998_ (.B1(net448),
    .Y(_0926_),
    .A1(net655),
    .A2(net392));
 sg13g2_a21oi_1 _2999_ (.A1(_0959_),
    .A2(net392),
    .Y(_0309_),
    .B1(_0926_));
 sg13g2_o21ai_1 _3000_ (.B1(net448),
    .Y(_0927_),
    .A1(net489),
    .A2(net392));
 sg13g2_a21oi_1 _3001_ (.A1(_0958_),
    .A2(net392),
    .Y(_0310_),
    .B1(_0927_));
 sg13g2_o21ai_1 _3002_ (.B1(net448),
    .Y(_0928_),
    .A1(\modem.control.scrambler_1.io_vecOut[9] ),
    .A2(net392));
 sg13g2_a21oi_1 _3003_ (.A1(_0957_),
    .A2(net392),
    .Y(_0311_),
    .B1(_0928_));
 sg13g2_o21ai_1 _3004_ (.B1(net448),
    .Y(_0929_),
    .A1(net324),
    .A2(net390));
 sg13g2_a21oi_1 _3005_ (.A1(_0956_),
    .A2(net390),
    .Y(_0312_),
    .B1(_0929_));
 sg13g2_o21ai_1 _3006_ (.B1(net446),
    .Y(_0930_),
    .A1(\modem.control.scrambler_1.io_vecOut[11] ),
    .A2(net390));
 sg13g2_a21oi_1 _3007_ (.A1(_0955_),
    .A2(net390),
    .Y(_0313_),
    .B1(_0930_));
 sg13g2_o21ai_1 _3008_ (.B1(net446),
    .Y(_0931_),
    .A1(net659),
    .A2(net390));
 sg13g2_a21oi_1 _3009_ (.A1(_0954_),
    .A2(net390),
    .Y(_0314_),
    .B1(_0931_));
 sg13g2_o21ai_1 _3010_ (.B1(net446),
    .Y(_0932_),
    .A1(net521),
    .A2(net389));
 sg13g2_a21oi_1 _3011_ (.A1(_0953_),
    .A2(net389),
    .Y(_0315_),
    .B1(_0932_));
 sg13g2_o21ai_1 _3012_ (.B1(net446),
    .Y(_0933_),
    .A1(\modem.control.scrambler_1.io_vecOut[14] ),
    .A2(net389));
 sg13g2_a21oi_1 _3013_ (.A1(_0952_),
    .A2(net389),
    .Y(_0316_),
    .B1(_0933_));
 sg13g2_o21ai_1 _3014_ (.B1(net446),
    .Y(_0934_),
    .A1(net482),
    .A2(net389));
 sg13g2_a21oi_1 _3015_ (.A1(_0951_),
    .A2(net389),
    .Y(_0317_),
    .B1(_0934_));
 sg13g2_o21ai_1 _3016_ (.B1(net446),
    .Y(_0935_),
    .A1(net332),
    .A2(net389));
 sg13g2_a21oi_1 _3017_ (.A1(_0950_),
    .A2(net389),
    .Y(_0318_),
    .B1(_0935_));
 sg13g2_o21ai_1 _3018_ (.B1(net447),
    .Y(_0936_),
    .A1(net416),
    .A2(\modem.dcdHistory_4 ));
 sg13g2_a21oi_1 _3019_ (.A1(net416),
    .A2(_0949_),
    .Y(_0319_),
    .B1(_0936_));
 sg13g2_o21ai_1 _3020_ (.B1(net447),
    .Y(_0937_),
    .A1(net415),
    .A2(\modem.dcdHistory_3 ));
 sg13g2_a21oi_1 _3021_ (.A1(net415),
    .A2(_0948_),
    .Y(_0320_),
    .B1(_0937_));
 sg13g2_o21ai_1 _3022_ (.B1(net447),
    .Y(_0938_),
    .A1(net415),
    .A2(net776));
 sg13g2_a21oi_1 _3023_ (.A1(net415),
    .A2(_0947_),
    .Y(_0321_),
    .B1(_0938_));
 sg13g2_o21ai_1 _3024_ (.B1(net447),
    .Y(_0939_),
    .A1(net416),
    .A2(net817));
 sg13g2_a21oi_1 _3025_ (.A1(net417),
    .A2(net369),
    .Y(_0322_),
    .B1(_0939_));
 sg13g2_o21ai_1 _3026_ (.B1(net447),
    .Y(_0940_),
    .A1(net415),
    .A2(net841));
 sg13g2_a21oi_1 _3027_ (.A1(net415),
    .A2(_0946_),
    .Y(_0323_),
    .B1(_0940_));
 sg13g2_o21ai_1 _3028_ (.B1(net447),
    .Y(_0941_),
    .A1(net493),
    .A2(net415));
 sg13g2_a21oi_1 _3029_ (.A1(net415),
    .A2(_0945_),
    .Y(_0324_),
    .B1(_0941_));
 sg13g2_o21ai_1 _3030_ (.B1(net447),
    .Y(_0942_),
    .A1(\modem.dcdHistory_7 ),
    .A2(net416));
 sg13g2_a21oi_1 _3031_ (.A1(_0943_),
    .A2(net416),
    .Y(_0325_),
    .B1(_0942_));
 sg13g2_dllrq_1 _3032_ (.D(net2),
    .GATE_N(net450),
    .RESET_B(net15),
    .Q(\latched[0] ));
 sg13g2_dllrq_1 _3033_ (.D(net3),
    .GATE_N(net454),
    .RESET_B(net16),
    .Q(\latched[1] ));
 sg13g2_dllrq_1 _3034_ (.D(net4),
    .GATE_N(net454),
    .RESET_B(net17),
    .Q(\latched[3] ));
 sg13g2_dllrq_1 _3035_ (.D(net5),
    .GATE_N(net454),
    .RESET_B(net18),
    .Q(\latched[5] ));
 sg13g2_dllrq_1 _3036_ (.D(net6),
    .GATE_N(net450),
    .RESET_B(net19),
    .Q(\latched[6] ));
 sg13g2_dllrq_1 _3037_ (.D(net7),
    .GATE_N(net448),
    .RESET_B(net20),
    .Q(\latched[7] ));
 sg13g2_dllrq_1 _3038_ (.D(net9),
    .GATE_N(net454),
    .RESET_B(net21),
    .Q(\latched[12] ));
 sg13g2_dllrq_1 _3039_ (.D(net10),
    .GATE_N(net454),
    .RESET_B(net22),
    .Q(\latched[14] ));
 sg13g2_dllrq_1 _3040_ (.D(net11),
    .GATE_N(net454),
    .RESET_B(net23),
    .Q(\latched[15] ));
 sg13g2_dfrbp_1 _3041_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net26),
    .D(net1),
    .Q_N(_0074_),
    .Q(\modem.control.rst_n ));
 sg13g2_dfrbp_1 _3042_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net27),
    .D(net743),
    .Q_N(_0075_),
    .Q(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[1] ));
 sg13g2_dfrbp_1 _3043_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net28),
    .D(_0017_),
    .Q_N(_1480_),
    .Q(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[2] ));
 sg13g2_dfrbp_1 _3044_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net29),
    .D(net756),
    .Q_N(_0076_),
    .Q(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[3] ));
 sg13g2_dfrbp_1 _3045_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net30),
    .D(net706),
    .Q_N(_1481_),
    .Q(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[4] ));
 sg13g2_dfrbp_1 _3046_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net35),
    .D(net725),
    .Q_N(_1482_),
    .Q(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[5] ));
 sg13g2_dfrbp_1 _3047_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net25),
    .D(net611),
    .Q_N(_1479_),
    .Q(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[6] ));
 sg13g2_dfrbp_1 _3048_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net122),
    .D(net333),
    .Q_N(_1478_),
    .Q(\modem.control.scrambler_1.io_vecOut[0] ));
 sg13g2_dfrbp_1 _3049_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net121),
    .D(net855),
    .Q_N(_0073_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_bit[0] ));
 sg13g2_dfrbp_1 _3050_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net119),
    .D(net850),
    .Q_N(_1477_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_bit[1] ));
 sg13g2_dfrbp_1 _3051_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net36),
    .D(net781),
    .Q_N(_0077_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_bit[2] ));
 sg13g2_dfrbp_1 _3052_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net37),
    .D(_0008_),
    .Q_N(_1483_),
    .Q(\modem.uart.tx.fsmUartTx_stateReg[1] ));
 sg13g2_dfrbp_1 _3053_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net38),
    .D(_0009_),
    .Q_N(_0078_),
    .Q(\modem.uart.tx.fsmUartTx_stateReg[2] ));
 sg13g2_dfrbp_1 _3054_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net39),
    .D(net773),
    .Q_N(_1484_),
    .Q(\modem.uart.tx.fsmUartTx_stateReg[3] ));
 sg13g2_dfrbp_1 _3055_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net40),
    .D(net694),
    .Q_N(_0079_),
    .Q(\modem.uart.tx.fsmUartTx_stateReg[4] ));
 sg13g2_dfrbp_1 _3056_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net41),
    .D(net801),
    .Q_N(_0080_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[1] ));
 sg13g2_dfrbp_1 _3057_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net42),
    .D(net877),
    .Q_N(_1485_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[2] ));
 sg13g2_dfrbp_1 _3058_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net43),
    .D(net702),
    .Q_N(_1486_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[3] ));
 sg13g2_dfrbp_1 _3059_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net44),
    .D(net786),
    .Q_N(_0081_),
    .Q(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[1] ));
 sg13g2_dfrbp_1 _3060_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net45),
    .D(net519),
    .Q_N(_1487_),
    .Q(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[2] ));
 sg13g2_dfrbp_1 _3061_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net46),
    .D(_0014_),
    .Q_N(_1488_),
    .Q(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[3] ));
 sg13g2_dfrbp_1 _3062_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net47),
    .D(_0015_),
    .Q_N(_1489_),
    .Q(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[4] ));
 sg13g2_dfrbp_1 _3063_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net48),
    .D(\modem.uart.txPacketUpper.io_ready ),
    .Q_N(_1490_),
    .Q(\modem.uart.uart_txPacketUpper_io_ready_regNext ));
 sg13g2_dfrbp_1 _3064_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net49),
    .D(net303),
    .Q_N(_1491_),
    .Q(\modem.uart.uart_txCommandDecoder_io_wantTx_regNext ));
 sg13g2_dfrbp_1 _3065_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net51),
    .D(net301),
    .Q_N(_1492_),
    .Q(\modem.uart.rxUart.io_uartRxIn_buffercc.buffers_1 ));
 sg13g2_dfrbp_1 _3066_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net117),
    .D(net7),
    .Q_N(_1476_),
    .Q(\modem.uart.rxUart.io_uartRxIn_buffercc.buffers_0 ));
 sg13g2_dfrbp_1 _3067_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net52),
    .D(net496),
    .Q_N(_0082_),
    .Q(\modem.uart.rxUart.samples_5 ));
 sg13g2_dfrbp_1 _3068_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net53),
    .D(net859),
    .Q_N(_1493_),
    .Q(\modem.uart.rxUart.sampleTimer_counter[0] ));
 sg13g2_dfrbp_1 _3069_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net207),
    .D(net753),
    .Q_N(_1494_),
    .Q(\modem.uart.rxUart.sampleTimer_counter[1] ));
 sg13g2_dfrbp_1 _3070_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net115),
    .D(net502),
    .Q_N(_0072_),
    .Q(\modem.uart.rxUart.sampleTimer_counter[2] ));
 sg13g2_dfrbp_1 _3071_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net114),
    .D(_0091_),
    .Q_N(_1475_),
    .Q(\modem.uart.rxUart.samples_6 ));
 sg13g2_dfrbp_1 _3072_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net113),
    .D(net312),
    .Q_N(_0071_),
    .Q(\modem.uart.tx.bitId[0] ));
 sg13g2_dfrbp_1 _3073_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net111),
    .D(_0093_),
    .Q_N(_1474_),
    .Q(\modem.uart.tx.bitId[1] ));
 sg13g2_dfrbp_1 _3074_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net109),
    .D(_0094_),
    .Q_N(_0070_),
    .Q(\modem.uart.tx.bitId[2] ));
 sg13g2_dfrbp_1 _3075_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net107),
    .D(net543),
    .Q_N(_1473_),
    .Q(\modem.uart.rxFifo.io_dataIn[0] ));
 sg13g2_dfrbp_1 _3076_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net106),
    .D(net845),
    .Q_N(_1472_),
    .Q(\modem.uart.rxFifo.io_dataIn[1] ));
 sg13g2_dfrbp_1 _3077_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net105),
    .D(net722),
    .Q_N(_1471_),
    .Q(\modem.uart.rxFifo.io_dataIn[2] ));
 sg13g2_dfrbp_1 _3078_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net104),
    .D(net865),
    .Q_N(_1470_),
    .Q(\modem.uart.rxFifo.io_dataIn[3] ));
 sg13g2_dfrbp_1 _3079_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net103),
    .D(net771),
    .Q_N(_1469_),
    .Q(\modem.uart.rxFifo.io_dataIn[4] ));
 sg13g2_dfrbp_1 _3080_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net102),
    .D(net759),
    .Q_N(_1468_),
    .Q(\modem.uart.rxFifo.io_dataIn[5] ));
 sg13g2_dfrbp_1 _3081_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net101),
    .D(net730),
    .Q_N(_1467_),
    .Q(\modem.uart.rxFifo.io_dataIn[6] ));
 sg13g2_dfrbp_1 _3082_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net100),
    .D(net717),
    .Q_N(_1466_),
    .Q(\modem.uart.rxFifo.io_dataIn[7] ));
 sg13g2_dfrbp_1 _3083_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net99),
    .D(net762),
    .Q_N(_1465_),
    .Q(\modem.uart.rxUart._zz_sampleValue_29 ));
 sg13g2_dfrbp_1 _3084_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net98),
    .D(_0104_),
    .Q_N(_1464_),
    .Q(\modem.uart.rxUart.samples_2 ));
 sg13g2_dfrbp_1 _3085_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net97),
    .D(_0105_),
    .Q_N(_0069_),
    .Q(\modem.uart.rxUart.samples_3 ));
 sg13g2_dfrbp_1 _3086_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net96),
    .D(net737),
    .Q_N(_0068_),
    .Q(\modem.uart.rxUart.samples_4 ));
 sg13g2_dfrbp_1 _3087_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net95),
    .D(net882),
    .Q_N(_0067_),
    .Q(\modem.uart.rxHdlc.io_valid ));
 sg13g2_dfrbp_1 _3088_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net94),
    .D(net314),
    .Q_N(_0066_),
    .Q(\modem.uart.rxFifo.nextIn[0] ));
 sg13g2_dfrbp_1 _3089_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net92),
    .D(_0109_),
    .Q_N(_1463_),
    .Q(\modem.uart.rxFifo.nextIn[1] ));
 sg13g2_dfrbp_1 _3090_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net90),
    .D(_0110_),
    .Q_N(_0065_),
    .Q(\modem.uart.rxFifo.nextIn[2] ));
 sg13g2_dfrbp_1 _3091_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net88),
    .D(net320),
    .Q_N(_0064_),
    .Q(\modem.uart.rxFifo.nextOut[0] ));
 sg13g2_dfrbp_1 _3092_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net86),
    .D(_0112_),
    .Q_N(_1462_),
    .Q(\modem.uart.rxFifo.nextOut[1] ));
 sg13g2_dfrbp_1 _3093_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net84),
    .D(_0113_),
    .Q_N(_0063_),
    .Q(\modem.uart.rxFifo.nextOut[2] ));
 sg13g2_dfrbp_1 _3094_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net82),
    .D(_0114_),
    .Q_N(_1461_),
    .Q(\modem.uart.rxFifo.fifo_6[0] ));
 sg13g2_dfrbp_1 _3095_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net81),
    .D(net541),
    .Q_N(_1460_),
    .Q(\modem.uart.rxFifo.fifo_6[1] ));
 sg13g2_dfrbp_1 _3096_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net80),
    .D(net586),
    .Q_N(_1459_),
    .Q(\modem.uart.rxFifo.fifo_6[2] ));
 sg13g2_dfrbp_1 _3097_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net79),
    .D(net598),
    .Q_N(_1458_),
    .Q(\modem.uart.rxFifo.fifo_6[3] ));
 sg13g2_dfrbp_1 _3098_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net78),
    .D(net602),
    .Q_N(_1457_),
    .Q(\modem.uart.rxFifo.fifo_6[4] ));
 sg13g2_dfrbp_1 _3099_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net77),
    .D(net524),
    .Q_N(_1456_),
    .Q(\modem.uart.rxFifo.fifo_6[5] ));
 sg13g2_dfrbp_1 _3100_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net76),
    .D(net578),
    .Q_N(_1455_),
    .Q(\modem.uart.rxFifo.fifo_6[6] ));
 sg13g2_dfrbp_1 _3101_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net75),
    .D(net535),
    .Q_N(_1454_),
    .Q(\modem.uart.rxFifo.fifo_6[7] ));
 sg13g2_dfrbp_1 _3102_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net74),
    .D(_0122_),
    .Q_N(_1453_),
    .Q(\modem.uart.rxFifo.fifo_5[0] ));
 sg13g2_dfrbp_1 _3103_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net73),
    .D(net568),
    .Q_N(_1452_),
    .Q(\modem.uart.rxFifo.fifo_5[1] ));
 sg13g2_dfrbp_1 _3104_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net72),
    .D(net673),
    .Q_N(_1451_),
    .Q(\modem.uart.rxFifo.fifo_5[2] ));
 sg13g2_dfrbp_1 _3105_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net71),
    .D(_0125_),
    .Q_N(_1450_),
    .Q(\modem.uart.rxFifo.fifo_5[3] ));
 sg13g2_dfrbp_1 _3106_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net70),
    .D(net572),
    .Q_N(_1449_),
    .Q(\modem.uart.rxFifo.fifo_5[4] ));
 sg13g2_dfrbp_1 _3107_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net69),
    .D(net537),
    .Q_N(_1448_),
    .Q(\modem.uart.rxFifo.fifo_5[5] ));
 sg13g2_dfrbp_1 _3108_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net68),
    .D(net574),
    .Q_N(_1447_),
    .Q(\modem.uart.rxFifo.fifo_5[6] ));
 sg13g2_dfrbp_1 _3109_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net67),
    .D(net669),
    .Q_N(_1446_),
    .Q(\modem.uart.rxFifo.fifo_5[7] ));
 sg13g2_dfrbp_1 _3110_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net66),
    .D(_0130_),
    .Q_N(_1445_),
    .Q(\modem.uart.rxFifo.fifo_4[0] ));
 sg13g2_dfrbp_1 _3111_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net65),
    .D(net580),
    .Q_N(_1444_),
    .Q(\modem.uart.rxFifo.fifo_4[1] ));
 sg13g2_dfrbp_1 _3112_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net64),
    .D(net594),
    .Q_N(_1443_),
    .Q(\modem.uart.rxFifo.fifo_4[2] ));
 sg13g2_dfrbp_1 _3113_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net63),
    .D(_0133_),
    .Q_N(_1442_),
    .Q(\modem.uart.rxFifo.fifo_4[3] ));
 sg13g2_dfrbp_1 _3114_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net62),
    .D(net638),
    .Q_N(_1441_),
    .Q(\modem.uart.rxFifo.fifo_4[4] ));
 sg13g2_dfrbp_1 _3115_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net61),
    .D(net558),
    .Q_N(_1440_),
    .Q(\modem.uart.rxFifo.fifo_4[5] ));
 sg13g2_dfrbp_1 _3116_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net60),
    .D(net545),
    .Q_N(_1439_),
    .Q(\modem.uart.rxFifo.fifo_4[6] ));
 sg13g2_dfrbp_1 _3117_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net59),
    .D(net657),
    .Q_N(_1438_),
    .Q(\modem.uart.rxFifo.fifo_4[7] ));
 sg13g2_dfrbp_1 _3118_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net58),
    .D(_0138_),
    .Q_N(_1437_),
    .Q(\modem.uart.rxFifo.fifo_3[0] ));
 sg13g2_dfrbp_1 _3119_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net57),
    .D(net741),
    .Q_N(_1436_),
    .Q(\modem.uart.rxFifo.fifo_3[1] ));
 sg13g2_dfrbp_1 _3120_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net56),
    .D(net629),
    .Q_N(_1435_),
    .Q(\modem.uart.rxFifo.fifo_3[2] ));
 sg13g2_dfrbp_1 _3121_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net55),
    .D(net607),
    .Q_N(_1434_),
    .Q(\modem.uart.rxFifo.fifo_3[3] ));
 sg13g2_dfrbp_1 _3122_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net54),
    .D(net609),
    .Q_N(_1433_),
    .Q(\modem.uart.rxFifo.fifo_3[4] ));
 sg13g2_dfrbp_1 _3123_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net50),
    .D(net652),
    .Q_N(_1432_),
    .Q(\modem.uart.rxFifo.fifo_3[5] ));
 sg13g2_dfrbp_1 _3124_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net34),
    .D(net645),
    .Q_N(_1431_),
    .Q(\modem.uart.rxFifo.fifo_3[6] ));
 sg13g2_dfrbp_1 _3125_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net33),
    .D(net696),
    .Q_N(_1430_),
    .Q(\modem.uart.rxFifo.fifo_3[7] ));
 sg13g2_dfrbp_1 _3126_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net32),
    .D(_0146_),
    .Q_N(_1429_),
    .Q(\modem.uart.rxFifo.fifo_2[0] ));
 sg13g2_dfrbp_1 _3127_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net31),
    .D(net550),
    .Q_N(_1428_),
    .Q(\modem.uart.rxFifo.fifo_2[1] ));
 sg13g2_dfrbp_1 _3128_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net24),
    .D(net528),
    .Q_N(_1427_),
    .Q(\modem.uart.rxFifo.fifo_2[2] ));
 sg13g2_dfrbp_1 _3129_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net300),
    .D(_0149_),
    .Q_N(_1426_),
    .Q(\modem.uart.rxFifo.fifo_2[3] ));
 sg13g2_dfrbp_1 _3130_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net299),
    .D(net539),
    .Q_N(_1425_),
    .Q(\modem.uart.rxFifo.fifo_2[4] ));
 sg13g2_dfrbp_1 _3131_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net298),
    .D(net576),
    .Q_N(_1424_),
    .Q(\modem.uart.rxFifo.fifo_2[5] ));
 sg13g2_dfrbp_1 _3132_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net297),
    .D(net617),
    .Q_N(_1423_),
    .Q(\modem.uart.rxFifo.fifo_2[6] ));
 sg13g2_dfrbp_1 _3133_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net296),
    .D(net592),
    .Q_N(_1422_),
    .Q(\modem.uart.rxFifo.fifo_2[7] ));
 sg13g2_dfrbp_1 _3134_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net295),
    .D(_0154_),
    .Q_N(_1421_),
    .Q(\modem.uart.rxFifo.fifo_1[0] ));
 sg13g2_dfrbp_1 _3135_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net294),
    .D(net683),
    .Q_N(_1420_),
    .Q(\modem.uart.rxFifo.fifo_1[1] ));
 sg13g2_dfrbp_1 _3136_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net293),
    .D(net530),
    .Q_N(_1419_),
    .Q(\modem.uart.rxFifo.fifo_1[2] ));
 sg13g2_dfrbp_1 _3137_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net292),
    .D(net560),
    .Q_N(_1418_),
    .Q(\modem.uart.rxFifo.fifo_1[3] ));
 sg13g2_dfrbp_1 _3138_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net291),
    .D(net642),
    .Q_N(_1417_),
    .Q(\modem.uart.rxFifo.fifo_1[4] ));
 sg13g2_dfrbp_1 _3139_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net290),
    .D(net552),
    .Q_N(_1416_),
    .Q(\modem.uart.rxFifo.fifo_1[5] ));
 sg13g2_dfrbp_1 _3140_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net289),
    .D(net615),
    .Q_N(_1415_),
    .Q(\modem.uart.rxFifo.fifo_1[6] ));
 sg13g2_dfrbp_1 _3141_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net288),
    .D(net613),
    .Q_N(_1414_),
    .Q(\modem.uart.rxFifo.fifo_1[7] ));
 sg13g2_dfrbp_1 _3142_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net287),
    .D(net661),
    .Q_N(_1413_),
    .Q(\modem.control.zeroCrossDet_7 ));
 sg13g2_dfrbp_1 _3143_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net286),
    .D(_0163_),
    .Q_N(_1412_),
    .Q(\modem.uart.rxFifo.fifo_0[0] ));
 sg13g2_dfrbp_1 _3144_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net284),
    .D(net811),
    .Q_N(_1411_),
    .Q(\modem.uart.rxFifo.fifo_0[1] ));
 sg13g2_dfrbp_1 _3145_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net282),
    .D(_0165_),
    .Q_N(_1410_),
    .Q(\modem.uart.rxFifo.fifo_0[2] ));
 sg13g2_dfrbp_1 _3146_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net280),
    .D(_0166_),
    .Q_N(_1409_),
    .Q(\modem.uart.rxFifo.fifo_0[3] ));
 sg13g2_dfrbp_1 _3147_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net278),
    .D(_0167_),
    .Q_N(_1408_),
    .Q(\modem.uart.rxFifo.fifo_0[4] ));
 sg13g2_dfrbp_1 _3148_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net276),
    .D(_0168_),
    .Q_N(_1407_),
    .Q(\modem.uart.rxFifo.fifo_0[5] ));
 sg13g2_dfrbp_1 _3149_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net274),
    .D(_0169_),
    .Q_N(_1406_),
    .Q(\modem.uart.rxFifo.fifo_0[6] ));
 sg13g2_dfrbp_1 _3150_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net272),
    .D(_0170_),
    .Q_N(_1405_),
    .Q(\modem.uart.rxFifo.fifo_0[7] ));
 sg13g2_dfrbp_1 _3151_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net270),
    .D(net488),
    .Q_N(_0062_),
    .Q(\modem.uart.rxFifo.count[0] ));
 sg13g2_dfrbp_1 _3152_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net268),
    .D(_0172_),
    .Q_N(_1404_),
    .Q(\modem.uart.rxFifo.count[1] ));
 sg13g2_dfrbp_1 _3153_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net266),
    .D(_0173_),
    .Q_N(_1403_),
    .Q(\modem.uart.rxFifo.count[2] ));
 sg13g2_dfrbp_1 _3154_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net264),
    .D(net663),
    .Q_N(_1402_),
    .Q(\modem.uart.rxFifo.count[3] ));
 sg13g2_dfrbp_1 _3155_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net261),
    .D(net869),
    .Q_N(_0061_),
    .Q(\modem.uart.descram.io_dataIn ));
 sg13g2_dfrbp_1 _3156_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net260),
    .D(net317),
    .Q_N(_1401_),
    .Q(\modem.uart.txCommandDecoder.io_wantTx ));
 sg13g2_dfrbp_1 _3157_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net258),
    .D(_0177_),
    .Q_N(_1400_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_1 ));
 sg13g2_dfrbp_1 _3158_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net252),
    .D(net733),
    .Q_N(_1399_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_2 ));
 sg13g2_dfrbp_1 _3159_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net250),
    .D(net790),
    .Q_N(_1398_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_3 ));
 sg13g2_dfrbp_1 _3160_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net248),
    .D(_0180_),
    .Q_N(_1397_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_4 ));
 sg13g2_dfrbp_1 _3161_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net246),
    .D(net832),
    .Q_N(_1396_),
    .Q(\modem.uart.txHdlc.txCrc.crc[4] ));
 sg13g2_dfrbp_1 _3162_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net244),
    .D(net727),
    .Q_N(_1395_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_6 ));
 sg13g2_dfrbp_1 _3163_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net242),
    .D(_0183_),
    .Q_N(_1394_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_7 ));
 sg13g2_dfrbp_1 _3164_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net240),
    .D(_0184_),
    .Q_N(_1393_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_8 ));
 sg13g2_dfrbp_1 _3165_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net238),
    .D(_0185_),
    .Q_N(_1392_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_9 ));
 sg13g2_dfrbp_1 _3166_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net236),
    .D(net745),
    .Q_N(_1391_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_10 ));
 sg13g2_dfrbp_1 _3167_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net234),
    .D(_0187_),
    .Q_N(_1390_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_11 ));
 sg13g2_dfrbp_1 _3168_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net232),
    .D(net783),
    .Q_N(_1389_),
    .Q(\modem.uart.txHdlc.txCrc.crc[11] ));
 sg13g2_dfrbp_1 _3169_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net230),
    .D(net739),
    .Q_N(_1388_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_13 ));
 sg13g2_dfrbp_1 _3170_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net228),
    .D(_0190_),
    .Q_N(_1387_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_14 ));
 sg13g2_dfrbp_1 _3171_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net226),
    .D(net775),
    .Q_N(_1386_),
    .Q(\modem.uart.txHdlc.txCrc.crcNext_15 ));
 sg13g2_dfrbp_1 _3172_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net223),
    .D(_0192_),
    .Q_N(_1385_),
    .Q(\modem.uart.txHdlc.txCrc.crc[15] ));
 sg13g2_dfrbp_1 _3173_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net221),
    .D(_0193_),
    .Q_N(_0060_),
    .Q(\modem.uart.txHdlc.wantFrameEnd ));
 sg13g2_dfrbp_1 _3174_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net220),
    .D(_0194_),
    .Q_N(_0059_),
    .Q(\modem.uart.txHdlc.isAbort ));
 sg13g2_dfrbp_1 _3175_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net219),
    .D(_0195_),
    .Q_N(_0058_),
    .Q(\modem.uart.txHdlc.isCRC ));
 sg13g2_dfrbp_1 _3176_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net217),
    .D(_0196_),
    .Q_N(_0057_),
    .Q(\modem.uart.io_isSending ));
 sg13g2_dfrbp_1 _3177_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net216),
    .D(net896),
    .Q_N(_0056_),
    .Q(\modem.uart.txHdlc.bit8[0] ));
 sg13g2_dfrbp_1 _3178_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net215),
    .D(_0198_),
    .Q_N(_1384_),
    .Q(\modem.uart.txHdlc.bit8[1] ));
 sg13g2_dfrbp_1 _3179_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net214),
    .D(_0199_),
    .Q_N(_0055_),
    .Q(\modem.uart.txHdlc.bit8[2] ));
 sg13g2_dfrbp_1 _3180_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net213),
    .D(_0200_),
    .Q_N(_0054_),
    .Q(\modem.uart.txHdlc.when_ModemTop_l593 ));
 sg13g2_dfrbp_1 _3181_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net206),
    .D(net692),
    .Q_N(_1383_),
    .Q(\modem.uart.txHdlc.bitstuffCnt[0] ));
 sg13g2_dfrbp_1 _3182_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net204),
    .D(net795),
    .Q_N(_1382_),
    .Q(\modem.uart.txHdlc.bitstuffCnt[1] ));
 sg13g2_dfrbp_1 _3183_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net202),
    .D(net463),
    .Q_N(_0053_),
    .Q(\modem.uart.txHdlc.bitstuffCnt[2] ));
 sg13g2_dfrbp_1 _3184_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net200),
    .D(net512),
    .Q_N(_1381_),
    .Q(\modem.uart.txFifo.fifo_3[0] ));
 sg13g2_dfrbp_1 _3185_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net199),
    .D(net492),
    .Q_N(_1380_),
    .Q(\modem.uart.txFifo.fifo_3[1] ));
 sg13g2_dfrbp_1 _3186_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net198),
    .D(net526),
    .Q_N(_1379_),
    .Q(\modem.uart.txFifo.fifo_3[2] ));
 sg13g2_dfrbp_1 _3187_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net197),
    .D(net504),
    .Q_N(_1378_),
    .Q(\modem.uart.txFifo.fifo_3[3] ));
 sg13g2_dfrbp_1 _3188_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net196),
    .D(net471),
    .Q_N(_1377_),
    .Q(\modem.uart.txFifo.fifo_3[4] ));
 sg13g2_dfrbp_1 _3189_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net195),
    .D(net465),
    .Q_N(_1376_),
    .Q(\modem.uart.txFifo.fifo_3[5] ));
 sg13g2_dfrbp_1 _3190_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net194),
    .D(net479),
    .Q_N(_1375_),
    .Q(\modem.uart.txFifo.fifo_3[6] ));
 sg13g2_dfrbp_1 _3191_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net193),
    .D(net473),
    .Q_N(_1374_),
    .Q(\modem.uart.txFifo.fifo_3[7] ));
 sg13g2_dfrbp_1 _3192_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net192),
    .D(net459),
    .Q_N(_0052_),
    .Q(\modem.uart.txFifo.nextIn[0] ));
 sg13g2_dfrbp_1 _3193_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net190),
    .D(_0213_),
    .Q_N(_1373_),
    .Q(\modem.uart.txFifo.nextIn[1] ));
 sg13g2_dfrbp_1 _3194_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net188),
    .D(net306),
    .Q_N(_0051_),
    .Q(\modem.uart.txFifo.nextOut[0] ));
 sg13g2_dfrbp_1 _3195_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net186),
    .D(net888),
    .Q_N(_1372_),
    .Q(\modem.uart.txFifo.nextOut[1] ));
 sg13g2_dfrbp_1 _3196_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net184),
    .D(net469),
    .Q_N(_1371_),
    .Q(\modem.uart.txFifo.fifo_2[0] ));
 sg13g2_dfrbp_1 _3197_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net183),
    .D(net508),
    .Q_N(_1370_),
    .Q(\modem.uart.txFifo.fifo_2[1] ));
 sg13g2_dfrbp_1 _3198_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net182),
    .D(net481),
    .Q_N(_1369_),
    .Q(\modem.uart.txFifo.fifo_2[2] ));
 sg13g2_dfrbp_1 _3199_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net181),
    .D(net533),
    .Q_N(_1368_),
    .Q(\modem.uart.txFifo.fifo_2[3] ));
 sg13g2_dfrbp_1 _3200_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net180),
    .D(net486),
    .Q_N(_1367_),
    .Q(\modem.uart.txFifo.fifo_2[4] ));
 sg13g2_dfrbp_1 _3201_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net179),
    .D(net477),
    .Q_N(_1366_),
    .Q(\modem.uart.txFifo.fifo_2[5] ));
 sg13g2_dfrbp_1 _3202_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net178),
    .D(net484),
    .Q_N(_1365_),
    .Q(\modem.uart.txFifo.fifo_2[6] ));
 sg13g2_dfrbp_1 _3203_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net177),
    .D(net475),
    .Q_N(_1364_),
    .Q(\modem.uart.txFifo.fifo_2[7] ));
 sg13g2_dfrbp_1 _3204_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net176),
    .D(net562),
    .Q_N(_1363_),
    .Q(\modem.uart.txFifo.fifo_1[0] ));
 sg13g2_dfrbp_1 _3205_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net175),
    .D(net712),
    .Q_N(_1362_),
    .Q(\modem.uart.txFifo.fifo_1[1] ));
 sg13g2_dfrbp_1 _3206_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net174),
    .D(net665),
    .Q_N(_1361_),
    .Q(\modem.uart.txFifo.fifo_1[2] ));
 sg13g2_dfrbp_1 _3207_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net173),
    .D(net596),
    .Q_N(_1360_),
    .Q(\modem.uart.txFifo.fifo_1[3] ));
 sg13g2_dfrbp_1 _3208_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net172),
    .D(net648),
    .Q_N(_1359_),
    .Q(\modem.uart.txFifo.fifo_1[4] ));
 sg13g2_dfrbp_1 _3209_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net171),
    .D(net570),
    .Q_N(_1358_),
    .Q(\modem.uart.txFifo.fifo_1[5] ));
 sg13g2_dfrbp_1 _3210_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net170),
    .D(net582),
    .Q_N(_1357_),
    .Q(\modem.uart.txFifo.fifo_1[6] ));
 sg13g2_dfrbp_1 _3211_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net169),
    .D(net749),
    .Q_N(_1356_),
    .Q(\modem.uart.txFifo.fifo_1[7] ));
 sg13g2_dfrbp_1 _3212_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net168),
    .D(net768),
    .Q_N(_1355_),
    .Q(\modem.uart.txFifo.fifo_0[0] ));
 sg13g2_dfrbp_1 _3213_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net166),
    .D(net735),
    .Q_N(_1354_),
    .Q(\modem.uart.txFifo.fifo_0[1] ));
 sg13g2_dfrbp_1 _3214_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net164),
    .D(net709),
    .Q_N(_1353_),
    .Q(\modem.uart.txFifo.fifo_0[2] ));
 sg13g2_dfrbp_1 _3215_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net162),
    .D(net766),
    .Q_N(_1352_),
    .Q(\modem.uart.txFifo.fifo_0[3] ));
 sg13g2_dfrbp_1 _3216_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net160),
    .D(net747),
    .Q_N(_1351_),
    .Q(\modem.uart.txFifo.fifo_0[4] ));
 sg13g2_dfrbp_1 _3217_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net158),
    .D(net793),
    .Q_N(_1350_),
    .Q(\modem.uart.txFifo.fifo_0[5] ));
 sg13g2_dfrbp_1 _3218_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net156),
    .D(net764),
    .Q_N(_1349_),
    .Q(\modem.uart.txFifo.fifo_0[6] ));
 sg13g2_dfrbp_1 _3219_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net154),
    .D(net719),
    .Q_N(_1348_),
    .Q(\modem.uart.txFifo.fifo_0[7] ));
 sg13g2_dfrbp_1 _3220_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net152),
    .D(net457),
    .Q_N(_0050_),
    .Q(\modem.uart.txFifo.count[0] ));
 sg13g2_dfrbp_1 _3221_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net150),
    .D(_0241_),
    .Q_N(_1347_),
    .Q(\modem.uart.txFifo.count[1] ));
 sg13g2_dfrbp_1 _3222_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net148),
    .D(net625),
    .Q_N(_1346_),
    .Q(\modem.uart.txFifo.count[2] ));
 sg13g2_dfrbp_1 _3223_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net208),
    .D(_0243_),
    .Q_N(_0083_),
    .Q(\modem.uart.rxFifo.io_dataInEn ));
 sg13g2_dfrbp_1 _3224_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net209),
    .D(net439),
    .Q_N(_1495_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[0] ));
 sg13g2_dfrbp_1 _3225_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net210),
    .D(net506),
    .Q_N(_0084_),
    .Q(\modem.uart.rxUart.fsmUartRx_stateReg[1] ));
 sg13g2_dfrbp_1 _3226_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net211),
    .D(_0004_),
    .Q_N(_1496_),
    .Q(\modem.uart.rxUart.fsmUartRx_stateReg[2] ));
 sg13g2_dfrbp_1 _3227_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net212),
    .D(net680),
    .Q_N(_1497_),
    .Q(\modem.uart.rxUart.fsmUartRx_stateReg[3] ));
 sg13g2_dfrbp_1 _3228_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net224),
    .D(net813),
    .Q_N(_1498_),
    .Q(\modem.uart.rxUart.fsmUartRx_stateReg[4] ));
 sg13g2_dfrbp_1 _3229_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net146),
    .D(_0007_),
    .Q_N(_0049_),
    .Q(\modem.uart.rxUart.fsmUartRx_stateReg[5] ));
 sg13g2_dfrbp_1 _3230_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net145),
    .D(_0244_),
    .Q_N(_1345_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[0] ));
 sg13g2_dfrbp_1 _3231_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net144),
    .D(_0245_),
    .Q_N(_1344_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[1] ));
 sg13g2_dfrbp_1 _3232_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net143),
    .D(_0246_),
    .Q_N(_1343_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[2] ));
 sg13g2_dfrbp_1 _3233_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net142),
    .D(_0247_),
    .Q_N(_1342_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[3] ));
 sg13g2_dfrbp_1 _3234_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net141),
    .D(_0248_),
    .Q_N(_1341_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[4] ));
 sg13g2_dfrbp_1 _3235_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net140),
    .D(_0249_),
    .Q_N(_1340_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[5] ));
 sg13g2_dfrbp_1 _3236_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net139),
    .D(_0250_),
    .Q_N(_1339_),
    .Q(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[6] ));
 sg13g2_dfrbp_1 _3237_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net138),
    .D(_0251_),
    .Q_N(_1338_),
    .Q(\modem.uart.rxHdlc.regNextRxDataIn ));
 sg13g2_dfrbp_1 _3238_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net137),
    .D(net323),
    .Q_N(_0048_),
    .Q(\modem.uart.rxHdlc.oneBitCount[0] ));
 sg13g2_dfrbp_1 _3239_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net135),
    .D(net826),
    .Q_N(_1337_),
    .Q(\modem.uart.rxHdlc.oneBitCount[1] ));
 sg13g2_dfrbp_1 _3240_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net254),
    .D(net699),
    .Q_N(_0085_),
    .Q(\modem.uart.rxHdlc.oneBitCount[2] ));
 sg13g2_dfrbp_1 _3241_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net133),
    .D(_0022_),
    .Q_N(_0047_),
    .Q(\modem.uart.rxHdlc.canInhibit ));
 sg13g2_dfrbp_1 _3242_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net131),
    .D(net510),
    .Q_N(_1336_),
    .Q(\modem.uart.rxHdlc.io_payload[0] ));
 sg13g2_dfrbp_1 _3243_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net130),
    .D(net621),
    .Q_N(_1335_),
    .Q(\modem.uart.rxHdlc.io_payload[1] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net129),
    .D(net514),
    .Q_N(_1334_),
    .Q(\modem.uart.rxHdlc.io_payload[2] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net128),
    .D(net517),
    .Q_N(_1333_),
    .Q(\modem.uart.rxHdlc.io_payload[3] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net127),
    .D(net554),
    .Q_N(_1332_),
    .Q(\modem.uart.rxHdlc.io_payload[4] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net126),
    .D(net564),
    .Q_N(_1331_),
    .Q(\modem.uart.rxHdlc.io_payload[5] ));
 sg13g2_dfrbp_1 _3248_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net125),
    .D(net588),
    .Q_N(_1330_),
    .Q(\modem.uart.rxHdlc.io_payload[6] ));
 sg13g2_dfrbp_1 _3249_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net124),
    .D(_0262_),
    .Q_N(_1329_),
    .Q(\modem.uart.rxHdlc.io_payload[7] ));
 sg13g2_dfrbp_1 _3250_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net123),
    .D(net467),
    .Q_N(_0046_),
    .Q(\modem.uart.rxFifo.fifo_7[0] ));
 sg13g2_dfrbp_1 _3251_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net120),
    .D(net331),
    .Q_N(_0045_),
    .Q(\modem.uart.rxFifo.fifo_7[1] ));
 sg13g2_dfrbp_1 _3252_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net118),
    .D(net339),
    .Q_N(_0044_),
    .Q(\modem.uart.rxFifo.fifo_7[2] ));
 sg13g2_dfrbp_1 _3253_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net116),
    .D(net461),
    .Q_N(_0043_),
    .Q(\modem.uart.rxFifo.fifo_7[3] ));
 sg13g2_dfrbp_1 _3254_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net112),
    .D(net329),
    .Q_N(_0042_),
    .Q(\modem.uart.rxFifo.fifo_7[4] ));
 sg13g2_dfrbp_1 _3255_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net110),
    .D(net327),
    .Q_N(_0041_),
    .Q(\modem.uart.rxFifo.fifo_7[5] ));
 sg13g2_dfrbp_1 _3256_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net108),
    .D(net337),
    .Q_N(_0040_),
    .Q(\modem.uart.rxFifo.fifo_7[6] ));
 sg13g2_dfrbp_1 _3257_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net93),
    .D(net335),
    .Q_N(_0039_),
    .Q(\modem.uart.rxFifo.fifo_7[7] ));
 sg13g2_dfrbp_1 _3258_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net91),
    .D(net898),
    .Q_N(_1328_),
    .Q(\modem.uart.txCommandDecoder.io_valid ));
 sg13g2_dfrbp_1 _3259_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net89),
    .D(net499),
    .Q_N(_0038_),
    .Q(\modem.uart.rxUart.bitId[0] ));
 sg13g2_dfrbp_1 _3260_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net85),
    .D(net853),
    .Q_N(_1327_),
    .Q(\modem.uart.rxUart.bitId[1] ));
 sg13g2_dfrbp_1 _3261_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net285),
    .D(net809),
    .Q_N(_0037_),
    .Q(\modem.uart.rxUart.bitId[2] ));
 sg13g2_dfrbp_1 _3262_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net281),
    .D(net623),
    .Q_N(_0036_),
    .Q(\modem.control.rxAddr[4] ));
 sg13g2_dfrbp_1 _3263_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net277),
    .D(net828),
    .Q_N(_1326_),
    .Q(\modem.control.rxAddr[5] ));
 sg13g2_dfrbp_1 _3264_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net273),
    .D(_0277_),
    .Q_N(_0035_),
    .Q(\modem.control.rxAddr[6] ));
 sg13g2_dfrbp_1 _3265_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net269),
    .D(net805),
    .Q_N(_0034_),
    .Q(\modem.control.rxAddr[7] ));
 sg13g2_dfrbp_1 _3266_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net265),
    .D(net848),
    .Q_N(_0033_),
    .Q(\modem.control.rxAddr[8] ));
 sg13g2_dfrbp_1 _3267_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net259),
    .D(_0280_),
    .Q_N(_0032_),
    .Q(\modem.control.rxAddr[9] ));
 sg13g2_dfrbp_1 _3268_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net251),
    .D(net857),
    .Q_N(_0031_),
    .Q(\modem.control.rxAddr[10] ));
 sg13g2_dfrbp_1 _3269_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net247),
    .D(net634),
    .Q_N(_1325_),
    .Q(\modem.control.rxAddr[11] ));
 sg13g2_dfrbp_1 _3270_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net255),
    .D(net822),
    .Q_N(_1499_),
    .Q(\modem.control.scrambler_1.io_dataIn ));
 sg13g2_dfrbp_1 _3271_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net256),
    .D(net315),
    .Q_N(_1500_),
    .Q(\modem.control._zz__3_regNext ));
 sg13g2_dfrbp_1 _3272_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net257),
    .D(net302),
    .Q_N(_1501_),
    .Q(\modem.control._zz__regNext ));
 sg13g2_dfrbp_1 _3273_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net262),
    .D(net309),
    .Q_N(_1502_),
    .Q(\modem.control._zz__1_regNext ));
 sg13g2_dfrbp_1 _3274_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net243),
    .D(net412),
    .Q_N(_1324_),
    .Q(\modem.control._zz__2_regNext ));
 sg13g2_dfrbp_1 _3275_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net239),
    .D(net308),
    .Q_N(_0030_),
    .Q(\modem.control.rxAddr[0] ));
 sg13g2_dfrbp_1 _3276_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net235),
    .D(net548),
    .Q_N(_1323_),
    .Q(\modem.control.rxAddr[1] ));
 sg13g2_dfrbp_1 _3277_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net231),
    .D(_0286_),
    .Q_N(_1322_),
    .Q(\modem.control.io_rxClock ));
 sg13g2_dfrbp_1 _3278_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net263),
    .D(_0287_),
    .Q_N(_1503_),
    .Q(\modem.control._zz_txClockInternalFallStb ));
 sg13g2_dfrbp_1 _3279_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net227),
    .D(net318),
    .Q_N(_1321_),
    .Q(\modem.control._zz_txClockInternalFallStb_regNext ));
 sg13g2_dfrbp_1 _3280_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net222),
    .D(_0288_),
    .Q_N(_0029_),
    .Q(\modem.control.phase[0] ));
 sg13g2_dfrbp_1 _3281_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net218),
    .D(_0289_),
    .Q_N(_1320_),
    .Q(\modem.control._zz__2 ));
 sg13g2_dfrbp_1 _3282_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net205),
    .D(_0290_),
    .Q_N(_1319_),
    .Q(\modem.control._zz__3 ));
 sg13g2_dfrbp_1 _3283_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net203),
    .D(_0291_),
    .Q_N(_1318_),
    .Q(\modem.control.tablePhase[3] ));
 sg13g2_dfrbp_1 _3284_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net201),
    .D(_0292_),
    .Q_N(_1317_),
    .Q(\modem.control._zz_ ));
 sg13g2_dfrbp_1 _3285_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net191),
    .D(_0293_),
    .Q_N(_1316_),
    .Q(\modem.control._zz__1 ));
 sg13g2_dfrbp_1 _3286_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net189),
    .D(net584),
    .Q_N(_1315_),
    .Q(\modem.analog_rxDac8[7] ));
 sg13g2_dfrbp_1 _3287_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net187),
    .D(_0295_),
    .Q_N(_1314_),
    .Q(\modem.control.rxRcrDacTmp[3] ));
 sg13g2_dfrbp_1 _3288_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net185),
    .D(_0296_),
    .Q_N(_1313_),
    .Q(\modem.control.zeroCrossDet_0 ));
 sg13g2_dfrbp_1 _3289_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net167),
    .D(net619),
    .Q_N(_1312_),
    .Q(\modem.control.zeroCrossDet_1 ));
 sg13g2_dfrbp_1 _3290_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net165),
    .D(_0298_),
    .Q_N(_1311_),
    .Q(\modem.control.zeroCrossDet_2 ));
 sg13g2_dfrbp_1 _3291_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net163),
    .D(net640),
    .Q_N(_1310_),
    .Q(\modem.control.zeroCrossDet_3 ));
 sg13g2_dfrbp_1 _3292_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net161),
    .D(_0300_),
    .Q_N(_1309_),
    .Q(\modem.control.zeroCrossDet_4 ));
 sg13g2_dfrbp_1 _3293_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net159),
    .D(net600),
    .Q_N(_1308_),
    .Q(\modem.control.zeroCrossDet_5 ));
 sg13g2_dfrbp_1 _3294_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net157),
    .D(net636),
    .Q_N(_1307_),
    .Q(\modem.control.zeroCrossDet_6 ));
 sg13g2_dfrbp_1 _3295_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net155),
    .D(net704),
    .Q_N(_1306_),
    .Q(\modem.control.scrambler_1.io_vecOut[1] ));
 sg13g2_dfrbp_1 _3296_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net151),
    .D(_0304_),
    .Q_N(_1305_),
    .Q(\modem.control.scrambler_1.io_vecOut[2] ));
 sg13g2_dfrbp_1 _3297_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net147),
    .D(_0305_),
    .Q_N(_1304_),
    .Q(\modem.control.scrambler_1.io_vecOut[3] ));
 sg13g2_dfrbp_1 _3298_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net134),
    .D(_0306_),
    .Q_N(_1303_),
    .Q(\modem.control.scrambler_1.io_vecOut[4] ));
 sg13g2_dfrbp_1 _3299_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net87),
    .D(net671),
    .Q_N(_1302_),
    .Q(\modem.control.scrambler_1.io_vecOut[5] ));
 sg13g2_dfrbp_1 _3300_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net283),
    .D(net556),
    .Q_N(_1301_),
    .Q(\modem.control.scrambler_1.io_vecOut[6] ));
 sg13g2_dfrbp_1 _3301_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net275),
    .D(_0309_),
    .Q_N(_1300_),
    .Q(\modem.control.scrambler_1.io_vecOut[7] ));
 sg13g2_dfrbp_1 _3302_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net267),
    .D(_0310_),
    .Q_N(_1299_),
    .Q(\modem.control.scrambler_1.io_vecOut[8] ));
 sg13g2_dfrbp_1 _3303_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net253),
    .D(net490),
    .Q_N(_1298_),
    .Q(\modem.control.scrambler_1.io_vecOut[9] ));
 sg13g2_dfrbp_1 _3304_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net245),
    .D(_0312_),
    .Q_N(_1297_),
    .Q(\modem.control.scrambler_1.io_vecOut[10] ));
 sg13g2_dfrbp_1 _3305_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net237),
    .D(net325),
    .Q_N(_1296_),
    .Q(\modem.control.scrambler_1.io_vecOut[11] ));
 sg13g2_dfrbp_1 _3306_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net229),
    .D(_0314_),
    .Q_N(_1295_),
    .Q(\modem.control.scrambler_1.io_vecOut[12] ));
 sg13g2_dfrbp_1 _3307_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net153),
    .D(_0315_),
    .Q_N(_1294_),
    .Q(\modem.control.scrambler_1.io_vecOut[13] ));
 sg13g2_dfrbp_1 _3308_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net136),
    .D(net522),
    .Q_N(_1293_),
    .Q(\modem.control.scrambler_1.io_vecOut[14] ));
 sg13g2_dfrbp_1 _3309_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net83),
    .D(_0317_),
    .Q_N(_1292_),
    .Q(\modem.control.scrambler_1.io_vecOut[15] ));
 sg13g2_dfrbp_1 _3310_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net271),
    .D(_0318_),
    .Q_N(_1291_),
    .Q(\modem.control.scrambler_1.io_vecOut[16] ));
 sg13g2_dfrbp_1 _3311_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net249),
    .D(net867),
    .Q_N(_1290_),
    .Q(\modem.dcdHistory_4 ));
 sg13g2_dfrbp_1 _3312_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net233),
    .D(net777),
    .Q_N(_1289_),
    .Q(\modem.dcdHistory_3 ));
 sg13g2_dfrbp_1 _3313_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net149),
    .D(_0321_),
    .Q_N(_0028_),
    .Q(\modem.dcdHistory_2 ));
 sg13g2_dfrbp_1 _3314_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net279),
    .D(_0322_),
    .Q_N(_0027_),
    .Q(\modem.dcdHistory_1 ));
 sg13g2_dfrbp_1 _3315_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net241),
    .D(net842),
    .Q_N(_0026_),
    .Q(\modem.dcdHistory_5 ));
 sg13g2_dfrbp_1 _3316_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net132),
    .D(_0324_),
    .Q_N(_1288_),
    .Q(\modem.dcdHistory_6 ));
 sg13g2_dfrbp_1 _3317_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net225),
    .D(net494),
    .Q_N(_1287_),
    .Q(\modem.dcdHistory_7 ));
 sg13g2_tiehi _3033__16 (.L_HI(net16));
 sg13g2_tiehi _3034__17 (.L_HI(net17));
 sg13g2_tiehi _3035__18 (.L_HI(net18));
 sg13g2_tiehi _3036__19 (.L_HI(net19));
 sg13g2_tiehi _3037__20 (.L_HI(net20));
 sg13g2_tiehi _3038__21 (.L_HI(net21));
 sg13g2_tiehi _3039__22 (.L_HI(net22));
 sg13g2_tiehi _3040__23 (.L_HI(net23));
 sg13g2_tiehi _3128__24 (.L_HI(net24));
 sg13g2_tiehi _3047__25 (.L_HI(net25));
 sg13g2_tiehi _3041__26 (.L_HI(net26));
 sg13g2_tiehi _3042__27 (.L_HI(net27));
 sg13g2_tiehi _3043__28 (.L_HI(net28));
 sg13g2_tiehi _3044__29 (.L_HI(net29));
 sg13g2_tiehi _3045__30 (.L_HI(net30));
 sg13g2_tiehi _3127__31 (.L_HI(net31));
 sg13g2_tiehi _3126__32 (.L_HI(net32));
 sg13g2_tiehi _3125__33 (.L_HI(net33));
 sg13g2_tiehi _3124__34 (.L_HI(net34));
 sg13g2_tiehi _3046__35 (.L_HI(net35));
 sg13g2_tiehi _3051__36 (.L_HI(net36));
 sg13g2_tiehi _3052__37 (.L_HI(net37));
 sg13g2_tiehi _3053__38 (.L_HI(net38));
 sg13g2_tiehi _3054__39 (.L_HI(net39));
 sg13g2_tiehi _3055__40 (.L_HI(net40));
 sg13g2_tiehi _3056__41 (.L_HI(net41));
 sg13g2_tiehi _3057__42 (.L_HI(net42));
 sg13g2_tiehi _3058__43 (.L_HI(net43));
 sg13g2_tiehi _3059__44 (.L_HI(net44));
 sg13g2_tiehi _3060__45 (.L_HI(net45));
 sg13g2_tiehi _3061__46 (.L_HI(net46));
 sg13g2_tiehi _3062__47 (.L_HI(net47));
 sg13g2_tiehi _3063__48 (.L_HI(net48));
 sg13g2_tiehi _3064__49 (.L_HI(net49));
 sg13g2_tiehi _3123__50 (.L_HI(net50));
 sg13g2_tiehi _3065__51 (.L_HI(net51));
 sg13g2_tiehi _3067__52 (.L_HI(net52));
 sg13g2_tiehi _3068__53 (.L_HI(net53));
 sg13g2_tiehi _3122__54 (.L_HI(net54));
 sg13g2_tiehi _3121__55 (.L_HI(net55));
 sg13g2_tiehi _3120__56 (.L_HI(net56));
 sg13g2_tiehi _3119__57 (.L_HI(net57));
 sg13g2_tiehi _3118__58 (.L_HI(net58));
 sg13g2_tiehi _3117__59 (.L_HI(net59));
 sg13g2_tiehi _3116__60 (.L_HI(net60));
 sg13g2_tiehi _3115__61 (.L_HI(net61));
 sg13g2_tiehi _3114__62 (.L_HI(net62));
 sg13g2_tiehi _3113__63 (.L_HI(net63));
 sg13g2_tiehi _3112__64 (.L_HI(net64));
 sg13g2_tiehi _3111__65 (.L_HI(net65));
 sg13g2_tiehi _3110__66 (.L_HI(net66));
 sg13g2_tiehi _3109__67 (.L_HI(net67));
 sg13g2_tiehi _3108__68 (.L_HI(net68));
 sg13g2_tiehi _3107__69 (.L_HI(net69));
 sg13g2_tiehi _3106__70 (.L_HI(net70));
 sg13g2_tiehi _3105__71 (.L_HI(net71));
 sg13g2_tiehi _3104__72 (.L_HI(net72));
 sg13g2_tiehi _3103__73 (.L_HI(net73));
 sg13g2_tiehi _3102__74 (.L_HI(net74));
 sg13g2_tiehi _3101__75 (.L_HI(net75));
 sg13g2_tiehi _3100__76 (.L_HI(net76));
 sg13g2_tiehi _3099__77 (.L_HI(net77));
 sg13g2_tiehi _3098__78 (.L_HI(net78));
 sg13g2_tiehi _3097__79 (.L_HI(net79));
 sg13g2_tiehi _3096__80 (.L_HI(net80));
 sg13g2_tiehi _3095__81 (.L_HI(net81));
 sg13g2_tiehi _3094__82 (.L_HI(net82));
 sg13g2_tiehi _3309__83 (.L_HI(net83));
 sg13g2_tiehi _3093__84 (.L_HI(net84));
 sg13g2_tiehi _3260__85 (.L_HI(net85));
 sg13g2_tiehi _3092__86 (.L_HI(net86));
 sg13g2_tiehi _3299__87 (.L_HI(net87));
 sg13g2_tiehi _3091__88 (.L_HI(net88));
 sg13g2_tiehi _3259__89 (.L_HI(net89));
 sg13g2_tiehi _3090__90 (.L_HI(net90));
 sg13g2_tiehi _3258__91 (.L_HI(net91));
 sg13g2_tiehi _3089__92 (.L_HI(net92));
 sg13g2_tiehi _3257__93 (.L_HI(net93));
 sg13g2_tiehi _3088__94 (.L_HI(net94));
 sg13g2_tiehi _3087__95 (.L_HI(net95));
 sg13g2_tiehi _3086__96 (.L_HI(net96));
 sg13g2_tiehi _3085__97 (.L_HI(net97));
 sg13g2_tiehi _3084__98 (.L_HI(net98));
 sg13g2_tiehi _3083__99 (.L_HI(net99));
 sg13g2_tiehi _3082__100 (.L_HI(net100));
 sg13g2_tiehi _3081__101 (.L_HI(net101));
 sg13g2_tiehi _3080__102 (.L_HI(net102));
 sg13g2_tiehi _3079__103 (.L_HI(net103));
 sg13g2_tiehi _3078__104 (.L_HI(net104));
 sg13g2_tiehi _3077__105 (.L_HI(net105));
 sg13g2_tiehi _3076__106 (.L_HI(net106));
 sg13g2_tiehi _3075__107 (.L_HI(net107));
 sg13g2_tiehi _3256__108 (.L_HI(net108));
 sg13g2_tiehi _3074__109 (.L_HI(net109));
 sg13g2_tiehi _3255__110 (.L_HI(net110));
 sg13g2_tiehi _3073__111 (.L_HI(net111));
 sg13g2_tiehi _3254__112 (.L_HI(net112));
 sg13g2_tiehi _3072__113 (.L_HI(net113));
 sg13g2_tiehi _3071__114 (.L_HI(net114));
 sg13g2_tiehi _3070__115 (.L_HI(net115));
 sg13g2_tiehi _3253__116 (.L_HI(net116));
 sg13g2_tiehi _3066__117 (.L_HI(net117));
 sg13g2_tiehi _3252__118 (.L_HI(net118));
 sg13g2_tiehi _3050__119 (.L_HI(net119));
 sg13g2_tiehi _3251__120 (.L_HI(net120));
 sg13g2_tiehi _3049__121 (.L_HI(net121));
 sg13g2_tiehi _3048__122 (.L_HI(net122));
 sg13g2_tiehi _3250__123 (.L_HI(net123));
 sg13g2_tiehi _3249__124 (.L_HI(net124));
 sg13g2_tiehi _3248__125 (.L_HI(net125));
 sg13g2_tiehi _3247__126 (.L_HI(net126));
 sg13g2_tiehi _3246__127 (.L_HI(net127));
 sg13g2_tiehi _3245__128 (.L_HI(net128));
 sg13g2_tiehi _3244__129 (.L_HI(net129));
 sg13g2_tiehi _3243__130 (.L_HI(net130));
 sg13g2_tiehi _3242__131 (.L_HI(net131));
 sg13g2_tiehi _3316__132 (.L_HI(net132));
 sg13g2_tiehi _3241__133 (.L_HI(net133));
 sg13g2_tiehi _3298__134 (.L_HI(net134));
 sg13g2_tiehi _3239__135 (.L_HI(net135));
 sg13g2_tiehi _3308__136 (.L_HI(net136));
 sg13g2_tiehi _3238__137 (.L_HI(net137));
 sg13g2_tiehi _3237__138 (.L_HI(net138));
 sg13g2_tiehi _3236__139 (.L_HI(net139));
 sg13g2_tiehi _3235__140 (.L_HI(net140));
 sg13g2_tiehi _3234__141 (.L_HI(net141));
 sg13g2_tiehi _3233__142 (.L_HI(net142));
 sg13g2_tiehi _3232__143 (.L_HI(net143));
 sg13g2_tiehi _3231__144 (.L_HI(net144));
 sg13g2_tiehi _3230__145 (.L_HI(net145));
 sg13g2_tiehi _3229__146 (.L_HI(net146));
 sg13g2_tiehi _3297__147 (.L_HI(net147));
 sg13g2_tiehi _3222__148 (.L_HI(net148));
 sg13g2_tiehi _3313__149 (.L_HI(net149));
 sg13g2_tiehi _3221__150 (.L_HI(net150));
 sg13g2_tiehi _3296__151 (.L_HI(net151));
 sg13g2_tiehi _3220__152 (.L_HI(net152));
 sg13g2_tiehi _3307__153 (.L_HI(net153));
 sg13g2_tiehi _3219__154 (.L_HI(net154));
 sg13g2_tiehi _3295__155 (.L_HI(net155));
 sg13g2_tiehi _3218__156 (.L_HI(net156));
 sg13g2_tiehi _3294__157 (.L_HI(net157));
 sg13g2_tiehi _3217__158 (.L_HI(net158));
 sg13g2_tiehi _3293__159 (.L_HI(net159));
 sg13g2_tiehi _3216__160 (.L_HI(net160));
 sg13g2_tiehi _3292__161 (.L_HI(net161));
 sg13g2_tiehi _3215__162 (.L_HI(net162));
 sg13g2_tiehi _3291__163 (.L_HI(net163));
 sg13g2_tiehi _3214__164 (.L_HI(net164));
 sg13g2_tiehi _3290__165 (.L_HI(net165));
 sg13g2_tiehi _3213__166 (.L_HI(net166));
 sg13g2_tiehi _3289__167 (.L_HI(net167));
 sg13g2_tiehi _3212__168 (.L_HI(net168));
 sg13g2_tiehi _3211__169 (.L_HI(net169));
 sg13g2_tiehi _3210__170 (.L_HI(net170));
 sg13g2_tiehi _3209__171 (.L_HI(net171));
 sg13g2_tiehi _3208__172 (.L_HI(net172));
 sg13g2_tiehi _3207__173 (.L_HI(net173));
 sg13g2_tiehi _3206__174 (.L_HI(net174));
 sg13g2_tiehi _3205__175 (.L_HI(net175));
 sg13g2_tiehi _3204__176 (.L_HI(net176));
 sg13g2_tiehi _3203__177 (.L_HI(net177));
 sg13g2_tiehi _3202__178 (.L_HI(net178));
 sg13g2_tiehi _3201__179 (.L_HI(net179));
 sg13g2_tiehi _3200__180 (.L_HI(net180));
 sg13g2_tiehi _3199__181 (.L_HI(net181));
 sg13g2_tiehi _3198__182 (.L_HI(net182));
 sg13g2_tiehi _3197__183 (.L_HI(net183));
 sg13g2_tiehi _3196__184 (.L_HI(net184));
 sg13g2_tiehi _3288__185 (.L_HI(net185));
 sg13g2_tiehi _3195__186 (.L_HI(net186));
 sg13g2_tiehi _3287__187 (.L_HI(net187));
 sg13g2_tiehi _3194__188 (.L_HI(net188));
 sg13g2_tiehi _3286__189 (.L_HI(net189));
 sg13g2_tiehi _3193__190 (.L_HI(net190));
 sg13g2_tiehi _3285__191 (.L_HI(net191));
 sg13g2_tiehi _3192__192 (.L_HI(net192));
 sg13g2_tiehi _3191__193 (.L_HI(net193));
 sg13g2_tiehi _3190__194 (.L_HI(net194));
 sg13g2_tiehi _3189__195 (.L_HI(net195));
 sg13g2_tiehi _3188__196 (.L_HI(net196));
 sg13g2_tiehi _3187__197 (.L_HI(net197));
 sg13g2_tiehi _3186__198 (.L_HI(net198));
 sg13g2_tiehi _3185__199 (.L_HI(net199));
 sg13g2_tiehi _3184__200 (.L_HI(net200));
 sg13g2_tiehi _3284__201 (.L_HI(net201));
 sg13g2_tiehi _3183__202 (.L_HI(net202));
 sg13g2_tiehi _3283__203 (.L_HI(net203));
 sg13g2_tiehi _3182__204 (.L_HI(net204));
 sg13g2_tiehi _3282__205 (.L_HI(net205));
 sg13g2_tiehi _3181__206 (.L_HI(net206));
 sg13g2_tiehi _3069__207 (.L_HI(net207));
 sg13g2_tiehi _3223__208 (.L_HI(net208));
 sg13g2_tiehi _3224__209 (.L_HI(net209));
 sg13g2_tiehi _3225__210 (.L_HI(net210));
 sg13g2_tiehi _3226__211 (.L_HI(net211));
 sg13g2_tiehi _3227__212 (.L_HI(net212));
 sg13g2_tiehi _3180__213 (.L_HI(net213));
 sg13g2_tiehi _3179__214 (.L_HI(net214));
 sg13g2_tiehi _3178__215 (.L_HI(net215));
 sg13g2_tiehi _3177__216 (.L_HI(net216));
 sg13g2_tiehi _3176__217 (.L_HI(net217));
 sg13g2_tiehi _3281__218 (.L_HI(net218));
 sg13g2_tiehi _3175__219 (.L_HI(net219));
 sg13g2_tiehi _3174__220 (.L_HI(net220));
 sg13g2_tiehi _3173__221 (.L_HI(net221));
 sg13g2_tiehi _3280__222 (.L_HI(net222));
 sg13g2_tiehi _3172__223 (.L_HI(net223));
 sg13g2_tiehi _3228__224 (.L_HI(net224));
 sg13g2_tiehi _3317__225 (.L_HI(net225));
 sg13g2_tiehi _3171__226 (.L_HI(net226));
 sg13g2_tiehi _3279__227 (.L_HI(net227));
 sg13g2_tiehi _3170__228 (.L_HI(net228));
 sg13g2_tiehi _3306__229 (.L_HI(net229));
 sg13g2_tiehi _3169__230 (.L_HI(net230));
 sg13g2_tiehi _3277__231 (.L_HI(net231));
 sg13g2_tiehi _3168__232 (.L_HI(net232));
 sg13g2_tiehi _3312__233 (.L_HI(net233));
 sg13g2_tiehi _3167__234 (.L_HI(net234));
 sg13g2_tiehi _3276__235 (.L_HI(net235));
 sg13g2_tiehi _3166__236 (.L_HI(net236));
 sg13g2_tiehi _3305__237 (.L_HI(net237));
 sg13g2_tiehi _3165__238 (.L_HI(net238));
 sg13g2_tiehi _3275__239 (.L_HI(net239));
 sg13g2_tiehi _3164__240 (.L_HI(net240));
 sg13g2_tiehi _3315__241 (.L_HI(net241));
 sg13g2_tiehi _3163__242 (.L_HI(net242));
 sg13g2_tiehi _3274__243 (.L_HI(net243));
 sg13g2_tiehi _3162__244 (.L_HI(net244));
 sg13g2_tiehi _3304__245 (.L_HI(net245));
 sg13g2_tiehi _3161__246 (.L_HI(net246));
 sg13g2_tiehi _3269__247 (.L_HI(net247));
 sg13g2_tiehi _3160__248 (.L_HI(net248));
 sg13g2_tiehi _3311__249 (.L_HI(net249));
 sg13g2_tiehi _3159__250 (.L_HI(net250));
 sg13g2_tiehi _3268__251 (.L_HI(net251));
 sg13g2_tiehi _3158__252 (.L_HI(net252));
 sg13g2_tiehi _3303__253 (.L_HI(net253));
 sg13g2_tiehi _3240__254 (.L_HI(net254));
 sg13g2_tiehi _3270__255 (.L_HI(net255));
 sg13g2_tiehi _3271__256 (.L_HI(net256));
 sg13g2_tiehi _3272__257 (.L_HI(net257));
 sg13g2_tiehi _3157__258 (.L_HI(net258));
 sg13g2_tiehi _3267__259 (.L_HI(net259));
 sg13g2_tiehi _3156__260 (.L_HI(net260));
 sg13g2_tiehi _3155__261 (.L_HI(net261));
 sg13g2_tiehi _3273__262 (.L_HI(net262));
 sg13g2_tiehi _3278__263 (.L_HI(net263));
 sg13g2_tiehi _3154__264 (.L_HI(net264));
 sg13g2_tiehi _3266__265 (.L_HI(net265));
 sg13g2_tiehi _3153__266 (.L_HI(net266));
 sg13g2_tiehi _3302__267 (.L_HI(net267));
 sg13g2_tiehi _3152__268 (.L_HI(net268));
 sg13g2_tiehi _3265__269 (.L_HI(net269));
 sg13g2_tiehi _3151__270 (.L_HI(net270));
 sg13g2_tiehi _3310__271 (.L_HI(net271));
 sg13g2_tiehi _3150__272 (.L_HI(net272));
 sg13g2_tiehi _3264__273 (.L_HI(net273));
 sg13g2_tiehi _3149__274 (.L_HI(net274));
 sg13g2_tiehi _3301__275 (.L_HI(net275));
 sg13g2_tiehi _3148__276 (.L_HI(net276));
 sg13g2_tiehi _3263__277 (.L_HI(net277));
 sg13g2_tiehi _3147__278 (.L_HI(net278));
 sg13g2_tiehi _3314__279 (.L_HI(net279));
 sg13g2_tiehi _3146__280 (.L_HI(net280));
 sg13g2_tiehi _3262__281 (.L_HI(net281));
 sg13g2_tiehi _3145__282 (.L_HI(net282));
 sg13g2_tiehi _3300__283 (.L_HI(net283));
 sg13g2_tiehi _3144__284 (.L_HI(net284));
 sg13g2_tiehi _3261__285 (.L_HI(net285));
 sg13g2_tiehi _3143__286 (.L_HI(net286));
 sg13g2_tiehi _3142__287 (.L_HI(net287));
 sg13g2_tiehi _3141__288 (.L_HI(net288));
 sg13g2_tiehi _3140__289 (.L_HI(net289));
 sg13g2_tiehi _3139__290 (.L_HI(net290));
 sg13g2_tiehi _3138__291 (.L_HI(net291));
 sg13g2_tiehi _3137__292 (.L_HI(net292));
 sg13g2_tiehi _3136__293 (.L_HI(net293));
 sg13g2_tiehi _3135__294 (.L_HI(net294));
 sg13g2_tiehi _3134__295 (.L_HI(net295));
 sg13g2_tiehi _3133__296 (.L_HI(net296));
 sg13g2_tiehi _3132__297 (.L_HI(net297));
 sg13g2_tiehi _3131__298 (.L_HI(net298));
 sg13g2_tiehi _3130__299 (.L_HI(net299));
 sg13g2_tiehi _3129__300 (.L_HI(net300));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_dlmiles_poc_fskmodem_hdlctrx_13 (.L_LO(net13));
 sg13g2_tielo tt_um_dlmiles_poc_fskmodem_hdlctrx_14 (.L_LO(net14));
 sg13g2_tiehi _3032__15 (.L_HI(net15));
 sg13g2_buf_2 _3607_ (.A(\modem.cfgRxClockDirection ),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3608_ (.A(\modem.cfgUpDownSource ),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3609_ (.A(\modem.cfgAddrDirection ),
    .X(uio_oe[2]));
 sg13g2_buf_2 _3610_ (.A(\modem.cfgAddrDirection ),
    .X(uio_oe[3]));
 sg13g2_buf_2 _3611_ (.A(\modem.cfgAddrDirection ),
    .X(uio_oe[4]));
 sg13g2_buf_2 _3612_ (.A(\modem.cfgAddrDirection ),
    .X(uio_oe[5]));
 sg13g2_buf_2 _3613_ (.A(\modem.cfgAddrDirection ),
    .X(uio_oe[6]));
 sg13g2_buf_2 _3614_ (.A(\modem.cfgAddrDirection ),
    .X(uio_oe[7]));
 sg13g2_buf_2 _3615_ (.A(net417),
    .X(uio_out[0]));
 sg13g2_buf_1 _3616_ (.A(\modem.control.io_upDownOut ),
    .X(uio_out[1]));
 sg13g2_buf_1 _3617_ (.A(\modem.uart.io_uartTxOut ),
    .X(uo_out[0]));
 sg13g2_buf_2 _3618_ (.A(\modem.uart.io_uartCtsOut ),
    .X(uo_out[1]));
 sg13g2_buf_1 _3619_ (.A(\modem.dcd ),
    .X(uo_out[2]));
 sg13g2_buf_4 _3620_ (.X(uo_out[5]),
    .A(\modem.uart.io_isSending ));
 sg13g2_buf_1 _3621_ (.A(\modem.control.io_txClockStb ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout341 (.A(net343),
    .X(net341));
 sg13g2_buf_1 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_0638_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_0637_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_0468_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_0830_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(net350),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_0778_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net353),
    .X(net351));
 sg13g2_buf_1 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_0787_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(net355),
    .X(net354));
 sg13g2_buf_1 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_0769_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_1 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_1 fanout359 (.A(_0755_),
    .X(net359));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(\modem.control.io_upDownOut ));
 sg13g2_buf_2 fanout361 (.A(net363),
    .X(net361));
 sg13g2_buf_1 fanout362 (.A(net363),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_0839_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(net365),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_1166_),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(net367));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(_1032_));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(_1031_));
 sg13g2_buf_2 fanout369 (.A(_1028_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(net371),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_0642_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_0532_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_0532_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_0523_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(net379),
    .X(net377));
 sg13g2_buf_1 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_0514_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(net381),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_0505_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(net383),
    .X(net382));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(_0495_));
 sg13g2_buf_2 fanout384 (.A(net385),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_0486_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_0476_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_0476_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_1057_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(net393),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(net393),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(net393),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_0919_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_0857_),
    .X(net394));
 sg13g2_buf_1 fanout395 (.A(_0857_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_1056_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_1053_),
    .X(net397));
 sg13g2_buf_1 fanout398 (.A(_1053_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_1046_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_1046_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_1044_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_1023_),
    .X(net402));
 sg13g2_buf_1 fanout403 (.A(_1023_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(net405),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_1001_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_1001_),
    .X(net408));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(_0993_));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(_0990_));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(\modem.control._zz__2 ));
 sg13g2_buf_1 fanout412 (.A(net675),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(net788),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(net416),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(net818),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(net419),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(\modem.uart.rxFifo.io_dataInEn ),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(\modem.uart.txFifo.nextOut[1] ),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(\modem.uart.txHdlc.when_ModemTop_l593 ),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(\modem.uart.txHdlc.bit8[2] ),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(\modem.uart.txHdlc.bit8[1] ),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(\modem.uart.txHdlc.bit8[1] ),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(net428),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(net428),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(\modem.uart.txHdlc.bit8[0] ),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(\modem.uart.txHdlc.isCRC ),
    .X(net429));
 sg13g2_buf_1 fanout430 (.A(\modem.uart.txHdlc.isCRC ),
    .X(net430));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(net432));
 sg13g2_buf_2 fanout432 (.A(\modem.uart.descram.io_dataIn ),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_0063_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(net436),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(\modem.uart.rxFifo.nextOut[2] ),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(net890),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(\modem.uart.tx.bitId[0] ),
    .X(net438));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(net515));
 sg13g2_buf_2 fanout440 (.A(net515),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(net442),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_4 fanout443 (.X(net443),
    .A(net456));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(net456));
 sg13g2_buf_1 fanout445 (.A(net456),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(net455),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net455),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net451),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net451),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(net451),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net455),
    .X(net451));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net454));
 sg13g2_buf_2 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(net456),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net851),
    .X(net456));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[4]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[6]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[7]),
    .X(net11));
 sg13g2_tielo tt_um_dlmiles_poc_fskmodem_hdlctrx_12 (.L_LO(net12));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_35_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_30_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_12_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\modem.uart.rxUart.io_uartRxIn_buffercc.buffers_0 ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold2 (.A(\modem.control._zz_ ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold3 (.A(\modem.uart.txCommandDecoder.io_wantTx ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0029_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0051_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0214_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0030_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0284_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold9 (.A(\modem.control._zz__1 ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0071_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0425_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0092_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0066_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0108_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold15 (.A(\modem.control._zz__3 ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0081_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0176_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold18 (.A(\modem.control._zz_txClockInternalFallStb ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0064_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0111_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0048_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0824_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0252_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold24 (.A(\modem.control.scrambler_1.io_vecOut[10] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0313_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold26 (.A(\modem.uart.rxFifo.fifo_7[5] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0268_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold28 (.A(\modem.uart.rxFifo.fifo_7[4] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0267_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold30 (.A(\modem.uart.rxFifo.fifo_7[1] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0264_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold32 (.A(\modem.control.scrambler_1.io_vecOut[16] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0086_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold34 (.A(\modem.uart.rxFifo.fifo_7[7] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0270_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold36 (.A(\modem.uart.rxFifo.fifo_7[6] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0269_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold38 (.A(\modem.uart.rxFifo.fifo_7[2] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0265_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0050_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0240_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0052_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0212_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold44 (.A(\modem.uart.rxFifo.fifo_7[3] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0266_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold46 (.A(\modem.uart.txHdlc.bitstuffCnt[2] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0203_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold48 (.A(\modem.uart.txFifo.fifo_3[5] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0209_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold50 (.A(\modem.uart.rxFifo.fifo_7[0] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0263_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold52 (.A(\modem.uart.txFifo.fifo_2[0] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0216_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold54 (.A(\modem.uart.txFifo.fifo_3[4] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0208_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold56 (.A(\modem.uart.txFifo.fifo_3[7] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0211_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold58 (.A(\modem.uart.txFifo.fifo_2[7] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0223_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold60 (.A(\modem.uart.txFifo.fifo_2[5] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0221_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold62 (.A(\modem.uart.txFifo.fifo_3[6] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0210_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold64 (.A(\modem.uart.txFifo.fifo_2[2] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0218_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold66 (.A(\modem.control.scrambler_1.io_vecOut[15] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold67 (.A(\modem.uart.txFifo.fifo_2[6] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0222_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold69 (.A(\modem.uart.txFifo.fifo_2[4] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0220_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0062_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0171_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold73 (.A(\modem.control.scrambler_1.io_vecOut[8] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0311_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold75 (.A(\modem.uart.txFifo.fifo_3[1] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0205_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold77 (.A(\modem.dcdHistory_6 ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0325_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold79 (.A(\modem.uart.rxUart.samples_5 ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0090_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0038_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0852_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0272_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0072_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0326_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0025_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold87 (.A(\modem.uart.txFifo.fifo_3[3] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0207_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0083_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0003_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold91 (.A(\modem.uart.txFifo.fifo_2[1] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0217_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold93 (.A(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[0] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0255_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold95 (.A(\modem.uart.txFifo.fifo_3[0] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0204_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold97 (.A(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[2] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0257_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0074_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold100 (.A(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[3] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0258_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold102 (.A(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[2] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0013_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold104 (.A(\modem.control.scrambler_1.io_vecOut[9] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold105 (.A(\modem.control.scrambler_1.io_vecOut[13] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0316_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold107 (.A(\modem.uart.rxFifo.fifo_6[5] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0119_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold109 (.A(\modem.uart.txFifo.fifo_3[2] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0206_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold111 (.A(\modem.uart.rxFifo.fifo_2[2] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0148_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold113 (.A(\modem.uart.rxFifo.fifo_1[2] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0156_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold115 (.A(\modem.control.scrambler_1.io_vecOut[14] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold116 (.A(\modem.uart.txFifo.fifo_2[3] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0219_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold118 (.A(\modem.uart.rxFifo.fifo_6[7] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0121_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold120 (.A(\modem.uart.rxFifo.fifo_5[5] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0127_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold122 (.A(\modem.uart.rxFifo.fifo_2[4] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0150_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold124 (.A(\modem.uart.rxFifo.fifo_6[1] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0115_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold126 (.A(\modem.uart.rxFifo.io_dataIn[0] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0095_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold128 (.A(\modem.uart.rxFifo.fifo_4[6] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0136_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold130 (.A(\modem.control.rxAddr[1] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0900_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0285_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold133 (.A(\modem.uart.rxFifo.fifo_2[1] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0147_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold135 (.A(\modem.uart.rxFifo.fifo_1[5] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0159_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold137 (.A(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[4] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0259_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold139 (.A(\modem.control.scrambler_1.io_vecOut[5] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0308_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold141 (.A(\modem.uart.rxFifo.fifo_4[5] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0135_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold143 (.A(\modem.uart.rxFifo.fifo_1[3] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0157_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold145 (.A(\modem.uart.txFifo.fifo_1[0] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0224_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold147 (.A(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[5] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0260_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0047_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0329_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold151 (.A(\modem.uart.rxFifo.fifo_5[1] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0123_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold153 (.A(\modem.uart.txFifo.fifo_1[5] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0229_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold155 (.A(\modem.uart.rxFifo.fifo_5[4] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0126_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold157 (.A(\modem.uart.rxFifo.fifo_5[6] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0128_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold159 (.A(\modem.uart.rxFifo.fifo_2[5] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0151_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold161 (.A(\modem.uart.rxFifo.fifo_6[6] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0120_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold163 (.A(\modem.uart.rxFifo.fifo_4[1] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0131_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold165 (.A(\modem.uart.txFifo.fifo_1[6] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0230_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold167 (.A(\modem.analog_rxDac8[7] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0294_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold169 (.A(\modem.uart.rxFifo.fifo_6[2] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0116_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold171 (.A(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[6] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0261_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold173 (.A(\modem.uart.rxFifo.fifo_6[0] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold174 (.A(\modem.uart.rxFifo.fifo_2[0] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold175 (.A(\modem.uart.rxFifo.fifo_2[7] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0153_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold177 (.A(\modem.uart.rxFifo.fifo_4[2] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0132_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold179 (.A(\modem.uart.txFifo.fifo_1[3] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0227_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold181 (.A(\modem.uart.rxFifo.fifo_6[3] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0117_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold183 (.A(\modem.control.zeroCrossDet_4 ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0301_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold185 (.A(\modem.uart.rxFifo.fifo_6[4] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0118_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold187 (.A(\modem.uart.rxFifo.fifo_1[0] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold188 (.A(\modem.uart.tx.fsmUartTx_stateReg[1] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1207_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold190 (.A(\modem.uart.rxFifo.io_dataIn[3] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0141_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold192 (.A(\modem.uart.rxFifo.fifo_3[4] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0142_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold194 (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[6] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0021_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold196 (.A(\modem.uart.rxFifo.fifo_1[7] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0161_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold198 (.A(\modem.uart.rxFifo.fifo_1[6] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0160_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold200 (.A(\modem.uart.rxFifo.fifo_2[6] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0152_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold202 (.A(\modem.control.zeroCrossDet_0 ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0297_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold204 (.A(\modem.uart.rxHdlc.fsmHdlcRx_rxByte[1] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0256_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold206 (.A(\modem.control.rxAddr[4] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0275_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold208 (.A(\modem.uart.txFifo.count[2] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0242_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold210 (.A(\modem.control._zz__3 ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold211 (.A(_1165_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold212 (.A(\modem.uart.rxFifo.fifo_3[2] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0140_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold214 (.A(\modem.uart.rxHdlc.regNextRxDataIn ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold215 (.A(\modem.uart.rxFifo.fifo_5[3] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold216 (.A(\modem.uart.rxFifo.fifo_5[0] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold217 (.A(\modem.control.rxAddr[11] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0282_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold219 (.A(\modem.control.zeroCrossDet_6 ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0302_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold221 (.A(\modem.uart.rxFifo.fifo_4[4] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0134_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold223 (.A(\modem.control.zeroCrossDet_2 ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0299_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold225 (.A(\modem.uart.rxFifo.fifo_1[4] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0158_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold227 (.A(\modem.control.zeroCrossDet_3 ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold228 (.A(\modem.uart.rxFifo.fifo_3[6] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0144_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold230 (.A(\modem.control.zeroCrossDet_1 ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold231 (.A(\modem.uart.txFifo.fifo_1[4] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0228_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold233 (.A(\modem.uart.rxFifo.fifo_4[3] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold234 (.A(\modem.control.rxRcrDacTmp[3] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold235 (.A(\modem.uart.rxFifo.fifo_3[5] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0143_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold237 (.A(\modem.uart.rxUart.fsmUartRx_stateReg[5] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold238 (.A(_1176_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold239 (.A(\modem.control.scrambler_1.io_vecOut[7] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold240 (.A(\modem.uart.rxFifo.fifo_4[7] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0137_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold242 (.A(\modem.uart.rxUart.fsmUartRx_stateReg[4] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold243 (.A(\modem.control.scrambler_1.io_vecOut[12] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold244 (.A(\modem.control.zeroCrossDet_7 ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0162_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold246 (.A(\modem.uart.rxFifo.count[3] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0174_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold248 (.A(\modem.uart.txFifo.fifo_1[2] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0226_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold250 (.A(\modem.uart.rxFifo.fifo_2[3] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold251 (.A(\modem.uart.rxFifo.fifo_5[7] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0494_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0129_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold254 (.A(\modem.control.scrambler_1.io_vecOut[4] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0307_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold256 (.A(\modem.uart.rxFifo.fifo_5[2] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0124_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold258 (.A(\modem.control.scrambler_1.io_vecOut[6] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold259 (.A(\modem.control._zz__2 ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold260 (.A(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[1] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold261 (.A(\modem.uart.rxFifo.fifo_3[0] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold262 (.A(\modem.uart.rxUart.fsmUartRx_stateReg[3] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold263 (.A(_1238_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0005_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold265 (.A(\modem.control.scrambler_1.io_vecOut[11] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold266 (.A(\modem.uart.rxFifo.fifo_1[1] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0155_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0073_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold269 (.A(\modem.uart.rxHdlc.fsmHdlcRx_bit[0] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0816_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold271 (.A(\modem.uart.rxFifo.fifo_4[0] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold272 (.A(\modem.uart.rxUart.samples_6 ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold273 (.A(\modem.uart.rxHdlc.fsmHdlcRx_bit[2] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold274 (.A(\modem.control.scrambler_1.io_vecOut[3] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold275 (.A(\modem.uart.txHdlc.bitstuffCnt[0] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0201_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold277 (.A(\modem.uart.tx.fsmUartTx_stateReg[2] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0011_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold279 (.A(\modem.uart.rxFifo.fifo_3[7] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0145_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold281 (.A(\modem.uart.rxHdlc.oneBitCount[2] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0829_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0254_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold284 (.A(\modem.control.scrambler_1.io_vecOut[2] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold285 (.A(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[3] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0002_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold287 (.A(\modem.control.scrambler_1.io_vecOut[0] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0303_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold289 (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[4] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0019_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold291 (.A(\modem.uart.rxHdlc.fsmHdlcRx_bit[2] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold292 (.A(\modem.uart.txFifo.fifo_0[2] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0234_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold294 (.A(\modem.uart.tx.fsmUartTx_stateReg[3] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold295 (.A(\modem.uart.txFifo.fifo_1[1] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0225_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold297 (.A(\modem.control.tablePhase[3] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0910_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold299 (.A(\modem.uart.rxFifo.io_dataIn[7] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0454_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0102_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold302 (.A(\modem.uart.txFifo.fifo_0[7] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0239_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold304 (.A(\modem.uart.rxFifo.io_dataIn[2] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0444_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0097_),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold307 (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[5] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold308 (.A(_1139_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0020_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold310 (.A(\modem.uart.txHdlc.txCrc.crcNext_6 ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0182_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold312 (.A(\modem.uart.rxFifo.io_dataIn[6] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0453_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0101_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold315 (.A(\modem.uart.txHdlc.txCrc.crcNext_7 ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold316 (.A(\modem.uart.txHdlc.txCrc.crcNext_1 ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0178_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold318 (.A(\modem.uart.txFifo.fifo_0[1] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0233_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold320 (.A(\modem.uart.rxUart.samples_3 ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0106_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold322 (.A(\modem.uart.txHdlc.txCrc.crcNext_13 ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0189_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold324 (.A(\modem.uart.rxFifo.fifo_3[1] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0139_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold326 (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[1] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0016_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold328 (.A(\modem.uart.txHdlc.txCrc.crcNext_9 ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0186_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold330 (.A(\modem.uart.txFifo.fifo_0[4] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0236_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold332 (.A(\modem.uart.txFifo.fifo_1[7] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0231_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold334 (.A(\modem.uart.txHdlc.txCrc.crc[15] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold335 (.A(\modem.uart.rxUart.sampleTimer_counter[1] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold336 (.A(_1286_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0024_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold338 (.A(\modem.uart.txHdlc.txCrc.crcNext_8 ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold339 (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[3] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0018_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold341 (.A(\modem.uart.rxFifo.io_dataIn[5] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0451_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0100_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold344 (.A(\modem.control.scrambler_1.io_vecOut[1] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold345 (.A(\modem.uart.rxUart.io_uartRxIn_buffercc.buffers_1 ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0103_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold347 (.A(\modem.uart.txFifo.fifo_0[6] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0238_),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold349 (.A(\modem.uart.txFifo.fifo_0[3] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0235_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold351 (.A(\modem.uart.txFifo.fifo_0[0] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0232_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold353 (.A(\modem.uart.rxFifo.io_dataIn[4] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0449_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0099_),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold356 (.A(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[0] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0010_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold358 (.A(\modem.uart.txHdlc.txCrc.crcNext_14 ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0191_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold360 (.A(\modem.dcdHistory_2 ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0320_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0080_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0421_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0422_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0089_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold366 (.A(\modem.uart.txHdlc.txCrc.crcNext_11 ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0188_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold368 (.A(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[1] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold369 (.A(_1193_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0012_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold371 (.A(\modem.uart.rxHdlc.fsmHdlcRx_bit[2] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold372 (.A(\modem.control.phase[0] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold373 (.A(\modem.uart.txHdlc.txCrc.crcNext_2 ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0179_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold375 (.A(\modem.uart.txHdlc.txCrc.crcNext_10 ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold376 (.A(\modem.uart.txFifo.fifo_0[5] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0237_),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold378 (.A(\modem.uart.txHdlc.bitstuffCnt[1] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0202_),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold380 (.A(\modem.control.rxAddr[6] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold381 (.A(\modem.control.rxAddr[9] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold382 (.A(\modem.uart.rxFifo.fifo_0[3] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold383 (.A(\modem.uart.rxHdlc.fsmHdlcRx_stateReg[2] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold384 (.A(_1229_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0000_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold386 (.A(\modem.uart.io_isSending ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold387 (.A(\modem.uart.rxFifo.fifo_0[7] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold388 (.A(\modem.control.rxAddr[7] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0278_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold390 (.A(\modem.uart.rxFifo.fifo_0[0] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold391 (.A(\modem.uart.rxUart.fsmUartRx_stateReg[1] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0855_),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0274_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold394 (.A(\modem.uart.rxFifo.fifo_0[1] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0164_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0037_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0006_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold398 (.A(\modem.uart.rxFifo.fifo_0[5] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0057_),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold400 (.A(_1035_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold401 (.A(\modem.dcdHistory_1 ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold402 (.A(\modem.control.io_rxClock ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold403 (.A(\modem.uart.txFifo.count[1] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold404 (.A(\modem.control.scrambler_1.io_dataIn ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0898_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0283_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold407 (.A(\modem.uart.rxUart.samples_2 ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold408 (.A(\modem.uart.rxHdlc.oneBitCount[1] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0826_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0253_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0036_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0276_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold413 (.A(\modem.uart.rxFifo.fifo_0[4] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold414 (.A(\modem.uart.txHdlc.txCrc.crcNext_15 ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold415 (.A(\modem.uart.txHdlc.txCrc.crcNext_4 ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0181_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold417 (.A(\modem.uart.rxFifo.nextOut[1] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0470_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold419 (.A(\modem.uart.rxHdlc.io_payload[7] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold420 (.A(\modem.uart.rxUart._zz_sampleValue_29 ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold421 (.A(\modem.uart.txHdlc.txCrc.crcNext_3 ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold422 (.A(\modem.uart.txFifo.nextIn[1] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0765_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold424 (.A(\modem.uart.rxFifo.fifo_0[2] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold425 (.A(\modem.dcdHistory_5 ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0323_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold427 (.A(\modem.uart.rxFifo.io_dataIn[1] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0442_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0096_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold430 (.A(\modem.uart.rxFifo.fifo_0[6] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold431 (.A(\modem.control.rxAddr[8] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0279_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold433 (.A(\modem.uart.rxHdlc.fsmHdlcRx_bit[1] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0088_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold435 (.A(\modem.control.rst_n ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold436 (.A(\modem.uart.rxUart.bitId[1] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0273_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0077_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0087_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold440 (.A(\modem.control.rxAddr[10] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0281_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold442 (.A(\modem.uart.rxUart.sampleTimer_counter[0] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0023_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold444 (.A(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[3] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold445 (.A(_0403_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold446 (.A(\modem.uart.rxFifo.nextIn[1] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0464_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0084_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0098_),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold450 (.A(\modem.dcdHistory_3 ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0319_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0061_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold453 (.A(_0175_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold454 (.A(\modem.uart.tx.bitId[2] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold455 (.A(_0430_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold456 (.A(\modem.uart.rxFifo.nextIn[2] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0060_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0688_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold459 (.A(_0059_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0085_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0001_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold462 (.A(\modem.uart.txHdlc.wantFrameEnd ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0677_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold464 (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[2] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0067_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0107_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold467 (.A(\modem.uart.rxFifo.count[2] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold468 (.A(\modem.uart.txCommandDecoder.fsmCmdDecoder_stateReg[4] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold469 (.A(\modem.uart.txHdlc.isAbort ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold470 (.A(\modem.uart.txFifo.nextOut[0] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0768_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0215_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold473 (.A(\modem.control.rxAddr[0] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold474 (.A(\modem.uart.tx.bitId[1] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0428_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold476 (.A(\modem.uart.rxUart.fsmUartRx_stateReg[2] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold477 (.A(\modem.uart.rxFifo.count[1] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0056_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0701_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0197_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold481 (.A(\modem.uart.txPacketUpper.fsmKissDecoder_stateReg[2] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0271_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0055_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0055_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold485 (.A(\modem.uart.txHdlc.wantFrameEnd ),
    .X(net901));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_4 FILLER_0_91 ();
 sg13g2_fill_2 FILLER_0_95 ();
 sg13g2_decap_8 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_141 ();
 sg13g2_decap_8 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_155 ();
 sg13g2_decap_8 FILLER_0_162 ();
 sg13g2_decap_8 FILLER_0_169 ();
 sg13g2_decap_8 FILLER_0_176 ();
 sg13g2_decap_8 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_197 ();
 sg13g2_decap_8 FILLER_0_204 ();
 sg13g2_decap_8 FILLER_0_211 ();
 sg13g2_decap_8 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_253 ();
 sg13g2_decap_8 FILLER_0_260 ();
 sg13g2_decap_8 FILLER_0_267 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_fill_2 FILLER_1_77 ();
 sg13g2_fill_2 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_142 ();
 sg13g2_decap_8 FILLER_1_149 ();
 sg13g2_decap_8 FILLER_1_156 ();
 sg13g2_decap_8 FILLER_1_163 ();
 sg13g2_decap_8 FILLER_1_170 ();
 sg13g2_decap_8 FILLER_1_177 ();
 sg13g2_decap_8 FILLER_1_184 ();
 sg13g2_decap_8 FILLER_1_191 ();
 sg13g2_decap_8 FILLER_1_198 ();
 sg13g2_decap_8 FILLER_1_205 ();
 sg13g2_decap_8 FILLER_1_212 ();
 sg13g2_decap_8 FILLER_1_219 ();
 sg13g2_decap_8 FILLER_1_226 ();
 sg13g2_decap_8 FILLER_1_233 ();
 sg13g2_decap_8 FILLER_1_240 ();
 sg13g2_decap_8 FILLER_1_247 ();
 sg13g2_decap_8 FILLER_1_254 ();
 sg13g2_decap_4 FILLER_1_261 ();
 sg13g2_fill_1 FILLER_1_265 ();
 sg13g2_fill_2 FILLER_1_296 ();
 sg13g2_fill_1 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_325 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_4 FILLER_2_70 ();
 sg13g2_fill_2 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_150 ();
 sg13g2_decap_8 FILLER_2_157 ();
 sg13g2_decap_8 FILLER_2_164 ();
 sg13g2_decap_8 FILLER_2_171 ();
 sg13g2_decap_8 FILLER_2_178 ();
 sg13g2_decap_8 FILLER_2_185 ();
 sg13g2_decap_8 FILLER_2_192 ();
 sg13g2_decap_8 FILLER_2_199 ();
 sg13g2_decap_8 FILLER_2_206 ();
 sg13g2_decap_8 FILLER_2_213 ();
 sg13g2_decap_8 FILLER_2_220 ();
 sg13g2_decap_8 FILLER_2_227 ();
 sg13g2_decap_8 FILLER_2_234 ();
 sg13g2_decap_8 FILLER_2_241 ();
 sg13g2_decap_8 FILLER_2_248 ();
 sg13g2_decap_4 FILLER_2_255 ();
 sg13g2_fill_1 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_fill_2 FILLER_3_70 ();
 sg13g2_fill_2 FILLER_3_131 ();
 sg13g2_fill_1 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_160 ();
 sg13g2_decap_8 FILLER_3_167 ();
 sg13g2_decap_8 FILLER_3_174 ();
 sg13g2_decap_8 FILLER_3_181 ();
 sg13g2_decap_8 FILLER_3_188 ();
 sg13g2_decap_8 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_3_202 ();
 sg13g2_decap_8 FILLER_3_209 ();
 sg13g2_decap_8 FILLER_3_216 ();
 sg13g2_decap_8 FILLER_3_223 ();
 sg13g2_decap_8 FILLER_3_230 ();
 sg13g2_decap_8 FILLER_3_237 ();
 sg13g2_decap_8 FILLER_3_244 ();
 sg13g2_decap_4 FILLER_3_251 ();
 sg13g2_decap_8 FILLER_3_328 ();
 sg13g2_decap_8 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_342 ();
 sg13g2_decap_8 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_fill_1 FILLER_4_70 ();
 sg13g2_fill_1 FILLER_4_93 ();
 sg13g2_fill_1 FILLER_4_122 ();
 sg13g2_fill_2 FILLER_4_149 ();
 sg13g2_fill_1 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_170 ();
 sg13g2_decap_8 FILLER_4_177 ();
 sg13g2_decap_8 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_decap_8 FILLER_4_219 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_decap_8 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_240 ();
 sg13g2_fill_1 FILLER_4_247 ();
 sg13g2_fill_2 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_fill_2 FILLER_5_70 ();
 sg13g2_fill_1 FILLER_5_108 ();
 sg13g2_fill_1 FILLER_5_143 ();
 sg13g2_fill_1 FILLER_5_148 ();
 sg13g2_decap_8 FILLER_5_181 ();
 sg13g2_decap_8 FILLER_5_188 ();
 sg13g2_decap_8 FILLER_5_195 ();
 sg13g2_decap_8 FILLER_5_202 ();
 sg13g2_decap_8 FILLER_5_209 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_8 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_4 FILLER_5_251 ();
 sg13g2_fill_1 FILLER_5_255 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_fill_2 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_298 ();
 sg13g2_fill_2 FILLER_5_308 ();
 sg13g2_fill_1 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_4 FILLER_6_56 ();
 sg13g2_fill_1 FILLER_6_60 ();
 sg13g2_fill_2 FILLER_6_153 ();
 sg13g2_decap_8 FILLER_6_194 ();
 sg13g2_decap_8 FILLER_6_201 ();
 sg13g2_decap_8 FILLER_6_208 ();
 sg13g2_decap_8 FILLER_6_215 ();
 sg13g2_decap_8 FILLER_6_222 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_decap_8 FILLER_6_236 ();
 sg13g2_fill_2 FILLER_6_243 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_fill_1 FILLER_6_272 ();
 sg13g2_fill_2 FILLER_6_294 ();
 sg13g2_fill_1 FILLER_6_296 ();
 sg13g2_fill_2 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_4 FILLER_7_63 ();
 sg13g2_fill_1 FILLER_7_67 ();
 sg13g2_fill_1 FILLER_7_138 ();
 sg13g2_decap_8 FILLER_7_183 ();
 sg13g2_decap_8 FILLER_7_190 ();
 sg13g2_decap_8 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_211 ();
 sg13g2_decap_8 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_225 ();
 sg13g2_decap_8 FILLER_7_232 ();
 sg13g2_fill_2 FILLER_7_239 ();
 sg13g2_fill_1 FILLER_7_241 ();
 sg13g2_fill_2 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_288 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_fill_2 FILLER_8_63 ();
 sg13g2_fill_1 FILLER_8_65 ();
 sg13g2_fill_1 FILLER_8_167 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_4 FILLER_8_245 ();
 sg13g2_fill_1 FILLER_8_249 ();
 sg13g2_fill_2 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_4 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_101 ();
 sg13g2_fill_1 FILLER_9_160 ();
 sg13g2_fill_2 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_201 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_229 ();
 sg13g2_decap_8 FILLER_9_236 ();
 sg13g2_decap_8 FILLER_9_243 ();
 sg13g2_decap_4 FILLER_9_250 ();
 sg13g2_fill_2 FILLER_9_254 ();
 sg13g2_fill_2 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_fill_2 FILLER_9_285 ();
 sg13g2_fill_2 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_4 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_74 ();
 sg13g2_fill_2 FILLER_10_136 ();
 sg13g2_fill_1 FILLER_10_138 ();
 sg13g2_decap_8 FILLER_10_192 ();
 sg13g2_decap_8 FILLER_10_199 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_213 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_decap_8 FILLER_10_227 ();
 sg13g2_decap_8 FILLER_10_234 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_fill_2 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_4 FILLER_11_63 ();
 sg13g2_fill_1 FILLER_11_125 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_275 ();
 sg13g2_fill_1 FILLER_11_277 ();
 sg13g2_fill_1 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_decap_8 FILLER_11_344 ();
 sg13g2_decap_8 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_358 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_94 ();
 sg13g2_fill_1 FILLER_12_101 ();
 sg13g2_fill_2 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_113 ();
 sg13g2_fill_2 FILLER_12_128 ();
 sg13g2_fill_1 FILLER_12_130 ();
 sg13g2_fill_1 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_fill_2 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_fill_1 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_4 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_53 ();
 sg13g2_decap_4 FILLER_13_187 ();
 sg13g2_fill_2 FILLER_13_191 ();
 sg13g2_decap_8 FILLER_13_223 ();
 sg13g2_decap_4 FILLER_13_230 ();
 sg13g2_fill_2 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_293 ();
 sg13g2_fill_1 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_fill_2 FILLER_14_114 ();
 sg13g2_fill_2 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_4 FILLER_14_240 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_fill_2 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_4 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_60 ();
 sg13g2_fill_2 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_160 ();
 sg13g2_fill_1 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_243 ();
 sg13g2_decap_4 FILLER_15_250 ();
 sg13g2_fill_2 FILLER_15_254 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_fill_2 FILLER_16_217 ();
 sg13g2_fill_2 FILLER_16_247 ();
 sg13g2_fill_1 FILLER_16_249 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_51 ();
 sg13g2_fill_1 FILLER_17_86 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_167 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_fill_2 FILLER_17_254 ();
 sg13g2_fill_2 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_fill_2 FILLER_17_281 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_93 ();
 sg13g2_fill_1 FILLER_18_99 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_146 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_fill_1 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_2 FILLER_18_205 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_fill_1 FILLER_18_237 ();
 sg13g2_fill_1 FILLER_18_244 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_331 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_decap_4 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_240 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_271 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_decap_4 FILLER_19_299 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_4 FILLER_20_56 ();
 sg13g2_fill_1 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_2 FILLER_20_116 ();
 sg13g2_fill_1 FILLER_20_196 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_decap_4 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_229 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_decap_4 FILLER_20_243 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_263 ();
 sg13g2_decap_4 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_206 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_4 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_fill_2 FILLER_22_99 ();
 sg13g2_fill_2 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_fill_1 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_202 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_decap_4 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_337 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_fill_1 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_195 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_152 ();
 sg13g2_decap_4 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_251 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_2 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_276 ();
 sg13g2_decap_8 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_313 ();
 sg13g2_decap_8 FILLER_25_320 ();
 sg13g2_decap_8 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_2 FILLER_26_136 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_260 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_352 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_180 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_337 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_fill_1 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_decap_4 FILLER_28_154 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_185 ();
 sg13g2_fill_2 FILLER_28_189 ();
 sg13g2_fill_2 FILLER_28_208 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_257 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_decap_8 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_60 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_decap_4 FILLER_29_179 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_107 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_120 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_decap_4 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_decap_4 FILLER_30_188 ();
 sg13g2_fill_2 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_4 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_31_114 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_136 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_182 ();
 sg13g2_decap_4 FILLER_31_193 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_decap_4 FILLER_31_206 ();
 sg13g2_fill_2 FILLER_31_250 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_314 ();
 sg13g2_decap_8 FILLER_31_321 ();
 sg13g2_decap_8 FILLER_31_328 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_decap_8 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_4 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_320 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_132 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_decap_8 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_334 ();
 sg13g2_decap_8 FILLER_33_341 ();
 sg13g2_decap_8 FILLER_33_348 ();
 sg13g2_decap_8 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_33_362 ();
 sg13g2_decap_8 FILLER_33_369 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_383 ();
 sg13g2_decap_8 FILLER_33_390 ();
 sg13g2_decap_8 FILLER_33_397 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_72 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_fill_2 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_decap_8 FILLER_34_339 ();
 sg13g2_decap_8 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_70 ();
 sg13g2_fill_2 FILLER_35_90 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_143 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_fill_1 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_decap_8 FILLER_35_319 ();
 sg13g2_decap_8 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_361 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_4 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_decap_4 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_311 ();
 sg13g2_decap_8 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_77 ();
 sg13g2_fill_1 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_117 ();
 sg13g2_fill_2 FILLER_37_169 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_decap_4 FILLER_37_180 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_201 ();
 sg13g2_decap_4 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_283 ();
 sg13g2_fill_2 FILLER_37_289 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_88 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_fill_2 FILLER_38_213 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_decap_8 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_decap_8 FILLER_38_319 ();
 sg13g2_decap_8 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_4 FILLER_39_77 ();
 sg13g2_fill_1 FILLER_39_81 ();
 sg13g2_fill_2 FILLER_39_100 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_fill_2 FILLER_39_117 ();
 sg13g2_fill_1 FILLER_39_133 ();
 sg13g2_fill_2 FILLER_39_149 ();
 sg13g2_fill_1 FILLER_39_189 ();
 sg13g2_fill_2 FILLER_39_226 ();
 sg13g2_fill_1 FILLER_39_228 ();
 sg13g2_fill_2 FILLER_39_242 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_fill_2 FILLER_39_272 ();
 sg13g2_decap_8 FILLER_39_300 ();
 sg13g2_decap_8 FILLER_39_307 ();
 sg13g2_decap_8 FILLER_39_314 ();
 sg13g2_decap_8 FILLER_39_321 ();
 sg13g2_decap_8 FILLER_39_328 ();
 sg13g2_decap_8 FILLER_39_335 ();
 sg13g2_decap_8 FILLER_39_342 ();
 sg13g2_decap_8 FILLER_39_349 ();
 sg13g2_decap_8 FILLER_39_356 ();
 sg13g2_decap_8 FILLER_39_363 ();
 sg13g2_decap_8 FILLER_39_370 ();
 sg13g2_decap_8 FILLER_39_377 ();
 sg13g2_decap_8 FILLER_39_384 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_4 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_60 ();
 sg13g2_fill_2 FILLER_40_103 ();
 sg13g2_fill_1 FILLER_40_155 ();
 sg13g2_fill_2 FILLER_40_187 ();
 sg13g2_fill_1 FILLER_40_189 ();
 sg13g2_fill_1 FILLER_40_242 ();
 sg13g2_fill_1 FILLER_40_252 ();
 sg13g2_fill_1 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_310 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_324 ();
 sg13g2_decap_8 FILLER_40_331 ();
 sg13g2_decap_8 FILLER_40_338 ();
 sg13g2_decap_8 FILLER_40_345 ();
 sg13g2_decap_8 FILLER_40_352 ();
 sg13g2_decap_8 FILLER_40_359 ();
 sg13g2_decap_8 FILLER_40_366 ();
 sg13g2_decap_8 FILLER_40_373 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_4 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_60 ();
 sg13g2_fill_2 FILLER_41_88 ();
 sg13g2_decap_4 FILLER_41_175 ();
 sg13g2_decap_4 FILLER_41_224 ();
 sg13g2_fill_1 FILLER_41_276 ();
 sg13g2_fill_1 FILLER_41_303 ();
 sg13g2_fill_2 FILLER_41_307 ();
 sg13g2_fill_1 FILLER_41_309 ();
 sg13g2_decap_8 FILLER_41_327 ();
 sg13g2_decap_8 FILLER_41_334 ();
 sg13g2_decap_8 FILLER_41_341 ();
 sg13g2_decap_8 FILLER_41_348 ();
 sg13g2_decap_8 FILLER_41_355 ();
 sg13g2_decap_8 FILLER_41_362 ();
 sg13g2_decap_8 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_376 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_56 ();
 sg13g2_fill_1 FILLER_42_60 ();
 sg13g2_fill_2 FILLER_42_82 ();
 sg13g2_fill_2 FILLER_42_128 ();
 sg13g2_fill_2 FILLER_42_174 ();
 sg13g2_fill_2 FILLER_42_196 ();
 sg13g2_fill_1 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_233 ();
 sg13g2_fill_1 FILLER_42_261 ();
 sg13g2_fill_1 FILLER_42_296 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_decap_8 FILLER_42_356 ();
 sg13g2_decap_8 FILLER_42_363 ();
 sg13g2_decap_8 FILLER_42_370 ();
 sg13g2_decap_8 FILLER_42_377 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_4 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_fill_1 FILLER_43_63 ();
 sg13g2_fill_2 FILLER_43_101 ();
 sg13g2_fill_2 FILLER_43_117 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_fill_2 FILLER_43_140 ();
 sg13g2_fill_1 FILLER_43_142 ();
 sg13g2_fill_1 FILLER_43_197 ();
 sg13g2_decap_4 FILLER_43_203 ();
 sg13g2_fill_2 FILLER_43_207 ();
 sg13g2_decap_4 FILLER_43_222 ();
 sg13g2_fill_2 FILLER_43_226 ();
 sg13g2_fill_2 FILLER_43_232 ();
 sg13g2_fill_1 FILLER_43_234 ();
 sg13g2_fill_1 FILLER_43_274 ();
 sg13g2_fill_2 FILLER_43_292 ();
 sg13g2_fill_2 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_fill_1 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_201 ();
 sg13g2_decap_8 FILLER_44_208 ();
 sg13g2_decap_8 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_decap_8 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_335 ();
 sg13g2_decap_8 FILLER_44_362 ();
 sg13g2_decap_8 FILLER_44_369 ();
 sg13g2_decap_8 FILLER_44_376 ();
 sg13g2_decap_8 FILLER_44_383 ();
 sg13g2_decap_8 FILLER_44_390 ();
 sg13g2_decap_8 FILLER_44_397 ();
 sg13g2_decap_4 FILLER_44_404 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_fill_1 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_148 ();
 sg13g2_decap_8 FILLER_45_155 ();
 sg13g2_decap_8 FILLER_45_162 ();
 sg13g2_fill_2 FILLER_45_169 ();
 sg13g2_fill_1 FILLER_45_171 ();
 sg13g2_fill_1 FILLER_45_207 ();
 sg13g2_decap_8 FILLER_45_211 ();
 sg13g2_fill_2 FILLER_45_244 ();
 sg13g2_fill_1 FILLER_45_250 ();
 sg13g2_fill_1 FILLER_45_259 ();
 sg13g2_fill_1 FILLER_45_283 ();
 sg13g2_fill_2 FILLER_45_325 ();
 sg13g2_decap_8 FILLER_45_363 ();
 sg13g2_decap_8 FILLER_45_370 ();
 sg13g2_decap_8 FILLER_45_377 ();
 sg13g2_decap_8 FILLER_45_384 ();
 sg13g2_decap_8 FILLER_45_391 ();
 sg13g2_decap_8 FILLER_45_398 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_fill_2 FILLER_46_56 ();
 sg13g2_fill_2 FILLER_46_120 ();
 sg13g2_fill_2 FILLER_46_136 ();
 sg13g2_decap_4 FILLER_46_169 ();
 sg13g2_fill_1 FILLER_46_181 ();
 sg13g2_decap_8 FILLER_46_246 ();
 sg13g2_fill_2 FILLER_46_253 ();
 sg13g2_decap_4 FILLER_46_263 ();
 sg13g2_fill_1 FILLER_46_267 ();
 sg13g2_fill_2 FILLER_46_273 ();
 sg13g2_fill_1 FILLER_46_284 ();
 sg13g2_decap_8 FILLER_46_372 ();
 sg13g2_decap_8 FILLER_46_379 ();
 sg13g2_decap_8 FILLER_46_386 ();
 sg13g2_decap_8 FILLER_46_393 ();
 sg13g2_decap_8 FILLER_46_400 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_4 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_60 ();
 sg13g2_fill_2 FILLER_47_121 ();
 sg13g2_fill_1 FILLER_47_123 ();
 sg13g2_fill_2 FILLER_47_163 ();
 sg13g2_fill_2 FILLER_47_183 ();
 sg13g2_fill_2 FILLER_47_199 ();
 sg13g2_fill_2 FILLER_47_252 ();
 sg13g2_fill_2 FILLER_47_263 ();
 sg13g2_fill_2 FILLER_47_270 ();
 sg13g2_fill_1 FILLER_47_298 ();
 sg13g2_fill_2 FILLER_47_328 ();
 sg13g2_fill_1 FILLER_47_330 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_decap_8 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_47_388 ();
 sg13g2_decap_8 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_86 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_fill_1 FILLER_48_123 ();
 sg13g2_fill_1 FILLER_48_139 ();
 sg13g2_fill_1 FILLER_48_178 ();
 sg13g2_fill_2 FILLER_48_225 ();
 sg13g2_fill_1 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_4 FILLER_49_56 ();
 sg13g2_fill_2 FILLER_49_60 ();
 sg13g2_fill_2 FILLER_49_86 ();
 sg13g2_fill_1 FILLER_49_93 ();
 sg13g2_fill_1 FILLER_49_139 ();
 sg13g2_fill_2 FILLER_49_152 ();
 sg13g2_fill_1 FILLER_49_154 ();
 sg13g2_fill_1 FILLER_49_217 ();
 sg13g2_fill_2 FILLER_49_227 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_1 FILLER_49_344 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_fill_2 FILLER_50_63 ();
 sg13g2_fill_1 FILLER_50_65 ();
 sg13g2_fill_1 FILLER_50_134 ();
 sg13g2_fill_1 FILLER_50_154 ();
 sg13g2_fill_1 FILLER_50_178 ();
 sg13g2_decap_4 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_221 ();
 sg13g2_fill_1 FILLER_50_267 ();
 sg13g2_fill_1 FILLER_50_292 ();
 sg13g2_fill_1 FILLER_50_348 ();
 sg13g2_decap_8 FILLER_50_384 ();
 sg13g2_decap_8 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_398 ();
 sg13g2_decap_4 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_fill_1 FILLER_51_70 ();
 sg13g2_fill_1 FILLER_51_102 ();
 sg13g2_fill_1 FILLER_51_188 ();
 sg13g2_fill_2 FILLER_51_214 ();
 sg13g2_fill_1 FILLER_51_216 ();
 sg13g2_fill_2 FILLER_51_243 ();
 sg13g2_fill_1 FILLER_51_306 ();
 sg13g2_fill_2 FILLER_51_343 ();
 sg13g2_fill_1 FILLER_51_345 ();
 sg13g2_fill_2 FILLER_51_351 ();
 sg13g2_fill_1 FILLER_51_353 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_386 ();
 sg13g2_decap_8 FILLER_51_393 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_4 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_decap_8 FILLER_52_218 ();
 sg13g2_fill_2 FILLER_52_225 ();
 sg13g2_fill_1 FILLER_52_236 ();
 sg13g2_fill_1 FILLER_52_252 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_fill_1 FILLER_52_333 ();
 sg13g2_decap_8 FILLER_52_390 ();
 sg13g2_decap_8 FILLER_52_397 ();
 sg13g2_decap_4 FILLER_52_404 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_fill_2 FILLER_53_70 ();
 sg13g2_fill_2 FILLER_53_88 ();
 sg13g2_fill_1 FILLER_53_105 ();
 sg13g2_fill_1 FILLER_53_171 ();
 sg13g2_decap_4 FILLER_53_208 ();
 sg13g2_fill_1 FILLER_53_212 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_226 ();
 sg13g2_decap_4 FILLER_53_244 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_decap_4 FILLER_53_253 ();
 sg13g2_fill_1 FILLER_53_257 ();
 sg13g2_fill_2 FILLER_53_263 ();
 sg13g2_decap_8 FILLER_53_270 ();
 sg13g2_fill_2 FILLER_53_277 ();
 sg13g2_fill_2 FILLER_53_284 ();
 sg13g2_fill_1 FILLER_53_286 ();
 sg13g2_decap_8 FILLER_53_386 ();
 sg13g2_decap_8 FILLER_53_393 ();
 sg13g2_decap_8 FILLER_53_400 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_fill_1 FILLER_54_63 ();
 sg13g2_fill_2 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_110 ();
 sg13g2_fill_1 FILLER_54_210 ();
 sg13g2_fill_2 FILLER_54_250 ();
 sg13g2_fill_1 FILLER_54_252 ();
 sg13g2_fill_2 FILLER_54_287 ();
 sg13g2_fill_1 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_386 ();
 sg13g2_decap_8 FILLER_54_393 ();
 sg13g2_decap_8 FILLER_54_400 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_fill_2 FILLER_55_122 ();
 sg13g2_fill_1 FILLER_55_179 ();
 sg13g2_fill_2 FILLER_55_214 ();
 sg13g2_fill_1 FILLER_55_216 ();
 sg13g2_fill_2 FILLER_55_227 ();
 sg13g2_fill_1 FILLER_55_229 ();
 sg13g2_fill_2 FILLER_55_289 ();
 sg13g2_fill_1 FILLER_55_305 ();
 sg13g2_fill_1 FILLER_55_319 ();
 sg13g2_fill_1 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_348 ();
 sg13g2_decap_8 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_4 FILLER_56_63 ();
 sg13g2_fill_2 FILLER_56_67 ();
 sg13g2_fill_1 FILLER_56_95 ();
 sg13g2_fill_1 FILLER_56_122 ();
 sg13g2_fill_2 FILLER_56_176 ();
 sg13g2_decap_8 FILLER_56_220 ();
 sg13g2_decap_8 FILLER_56_227 ();
 sg13g2_fill_1 FILLER_56_234 ();
 sg13g2_fill_1 FILLER_56_270 ();
 sg13g2_fill_1 FILLER_56_319 ();
 sg13g2_fill_2 FILLER_56_362 ();
 sg13g2_decap_8 FILLER_56_390 ();
 sg13g2_decap_8 FILLER_56_397 ();
 sg13g2_decap_4 FILLER_56_404 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_4 FILLER_57_70 ();
 sg13g2_fill_2 FILLER_57_74 ();
 sg13g2_fill_2 FILLER_57_94 ();
 sg13g2_fill_2 FILLER_57_105 ();
 sg13g2_fill_1 FILLER_57_135 ();
 sg13g2_fill_1 FILLER_57_158 ();
 sg13g2_fill_2 FILLER_57_176 ();
 sg13g2_fill_1 FILLER_57_187 ();
 sg13g2_fill_2 FILLER_57_202 ();
 sg13g2_fill_1 FILLER_57_204 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_fill_2 FILLER_57_283 ();
 sg13g2_fill_1 FILLER_57_293 ();
 sg13g2_fill_2 FILLER_57_303 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_fill_1 FILLER_58_63 ();
 sg13g2_fill_2 FILLER_58_104 ();
 sg13g2_fill_2 FILLER_58_164 ();
 sg13g2_fill_2 FILLER_58_269 ();
 sg13g2_fill_1 FILLER_58_271 ();
 sg13g2_fill_2 FILLER_58_277 ();
 sg13g2_fill_1 FILLER_58_279 ();
 sg13g2_fill_1 FILLER_58_303 ();
 sg13g2_fill_2 FILLER_58_356 ();
 sg13g2_fill_1 FILLER_58_358 ();
 sg13g2_fill_1 FILLER_58_377 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_4 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_78 ();
 sg13g2_fill_1 FILLER_59_106 ();
 sg13g2_fill_2 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_157 ();
 sg13g2_fill_1 FILLER_59_189 ();
 sg13g2_fill_2 FILLER_59_231 ();
 sg13g2_fill_1 FILLER_59_233 ();
 sg13g2_fill_2 FILLER_59_275 ();
 sg13g2_fill_1 FILLER_59_277 ();
 sg13g2_fill_2 FILLER_59_327 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_405 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_fill_2 FILLER_60_77 ();
 sg13g2_fill_1 FILLER_60_79 ();
 sg13g2_decap_8 FILLER_60_216 ();
 sg13g2_decap_8 FILLER_60_223 ();
 sg13g2_fill_2 FILLER_60_282 ();
 sg13g2_fill_1 FILLER_60_284 ();
 sg13g2_fill_1 FILLER_60_317 ();
 sg13g2_fill_1 FILLER_60_331 ();
 sg13g2_fill_1 FILLER_60_341 ();
 sg13g2_fill_2 FILLER_60_384 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_4 FILLER_61_63 ();
 sg13g2_fill_2 FILLER_61_197 ();
 sg13g2_fill_2 FILLER_61_203 ();
 sg13g2_fill_1 FILLER_61_214 ();
 sg13g2_fill_2 FILLER_61_239 ();
 sg13g2_fill_2 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_322 ();
 sg13g2_decap_4 FILLER_61_403 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_4 FILLER_62_70 ();
 sg13g2_fill_1 FILLER_62_74 ();
 sg13g2_fill_1 FILLER_62_107 ();
 sg13g2_fill_2 FILLER_62_141 ();
 sg13g2_decap_4 FILLER_62_171 ();
 sg13g2_fill_1 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_fill_2 FILLER_62_217 ();
 sg13g2_fill_2 FILLER_62_249 ();
 sg13g2_fill_2 FILLER_62_260 ();
 sg13g2_fill_2 FILLER_62_296 ();
 sg13g2_fill_1 FILLER_62_303 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_fill_1 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_118 ();
 sg13g2_decap_8 FILLER_63_145 ();
 sg13g2_fill_1 FILLER_63_152 ();
 sg13g2_decap_8 FILLER_63_157 ();
 sg13g2_decap_4 FILLER_63_164 ();
 sg13g2_fill_1 FILLER_63_178 ();
 sg13g2_fill_1 FILLER_63_189 ();
 sg13g2_fill_2 FILLER_63_219 ();
 sg13g2_fill_1 FILLER_63_221 ();
 sg13g2_fill_1 FILLER_63_287 ();
 sg13g2_fill_2 FILLER_63_349 ();
 sg13g2_fill_2 FILLER_63_391 ();
 sg13g2_fill_1 FILLER_63_393 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_4 FILLER_64_70 ();
 sg13g2_fill_2 FILLER_64_74 ();
 sg13g2_fill_2 FILLER_64_231 ();
 sg13g2_fill_1 FILLER_64_254 ();
 sg13g2_decap_4 FILLER_64_261 ();
 sg13g2_fill_1 FILLER_64_265 ();
 sg13g2_decap_4 FILLER_64_291 ();
 sg13g2_fill_1 FILLER_64_295 ();
 sg13g2_fill_2 FILLER_64_301 ();
 sg13g2_fill_1 FILLER_64_317 ();
 sg13g2_fill_2 FILLER_64_332 ();
 sg13g2_fill_2 FILLER_64_355 ();
 sg13g2_fill_1 FILLER_64_357 ();
 sg13g2_fill_1 FILLER_64_378 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_fill_2 FILLER_65_84 ();
 sg13g2_fill_1 FILLER_65_86 ();
 sg13g2_fill_2 FILLER_65_101 ();
 sg13g2_fill_1 FILLER_65_103 ();
 sg13g2_fill_1 FILLER_65_127 ();
 sg13g2_decap_8 FILLER_65_145 ();
 sg13g2_decap_8 FILLER_65_152 ();
 sg13g2_fill_2 FILLER_65_159 ();
 sg13g2_fill_1 FILLER_65_161 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_fill_1 FILLER_65_203 ();
 sg13g2_fill_1 FILLER_65_216 ();
 sg13g2_fill_1 FILLER_65_222 ();
 sg13g2_decap_8 FILLER_65_232 ();
 sg13g2_fill_2 FILLER_65_239 ();
 sg13g2_decap_8 FILLER_65_244 ();
 sg13g2_fill_1 FILLER_65_251 ();
 sg13g2_decap_4 FILLER_65_256 ();
 sg13g2_fill_1 FILLER_65_260 ();
 sg13g2_decap_4 FILLER_65_268 ();
 sg13g2_fill_2 FILLER_65_298 ();
 sg13g2_fill_1 FILLER_65_300 ();
 sg13g2_fill_2 FILLER_65_330 ();
 sg13g2_fill_1 FILLER_65_332 ();
 sg13g2_fill_2 FILLER_65_362 ();
 sg13g2_fill_1 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_101 ();
 sg13g2_fill_1 FILLER_66_108 ();
 sg13g2_fill_1 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_118 ();
 sg13g2_fill_2 FILLER_66_145 ();
 sg13g2_fill_1 FILLER_66_151 ();
 sg13g2_fill_2 FILLER_66_159 ();
 sg13g2_decap_4 FILLER_66_176 ();
 sg13g2_fill_1 FILLER_66_180 ();
 sg13g2_decap_8 FILLER_66_216 ();
 sg13g2_decap_4 FILLER_66_223 ();
 sg13g2_fill_2 FILLER_66_231 ();
 sg13g2_fill_2 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_398 ();
 sg13g2_decap_4 FILLER_66_405 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_110 ();
 sg13g2_fill_2 FILLER_67_117 ();
 sg13g2_decap_4 FILLER_67_187 ();
 sg13g2_fill_1 FILLER_67_191 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_4 FILLER_67_210 ();
 sg13g2_fill_2 FILLER_67_218 ();
 sg13g2_fill_1 FILLER_67_220 ();
 sg13g2_fill_1 FILLER_67_261 ();
 sg13g2_fill_2 FILLER_67_308 ();
 sg13g2_fill_2 FILLER_67_315 ();
 sg13g2_fill_1 FILLER_67_317 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_fill_2 FILLER_68_87 ();
 sg13g2_fill_2 FILLER_68_129 ();
 sg13g2_fill_1 FILLER_68_136 ();
 sg13g2_fill_2 FILLER_68_160 ();
 sg13g2_decap_8 FILLER_68_190 ();
 sg13g2_decap_8 FILLER_68_197 ();
 sg13g2_decap_4 FILLER_68_204 ();
 sg13g2_fill_1 FILLER_68_208 ();
 sg13g2_fill_1 FILLER_68_253 ();
 sg13g2_fill_1 FILLER_68_279 ();
 sg13g2_fill_2 FILLER_68_299 ();
 sg13g2_fill_1 FILLER_68_301 ();
 sg13g2_fill_2 FILLER_68_321 ();
 sg13g2_fill_2 FILLER_68_355 ();
 sg13g2_fill_1 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_fill_2 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_121 ();
 sg13g2_decap_4 FILLER_69_128 ();
 sg13g2_fill_1 FILLER_69_132 ();
 sg13g2_fill_2 FILLER_69_189 ();
 sg13g2_fill_2 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_271 ();
 sg13g2_fill_2 FILLER_69_355 ();
 sg13g2_decap_8 FILLER_69_401 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_fill_2 FILLER_70_70 ();
 sg13g2_fill_2 FILLER_70_105 ();
 sg13g2_fill_1 FILLER_70_133 ();
 sg13g2_fill_2 FILLER_70_167 ();
 sg13g2_fill_2 FILLER_70_218 ();
 sg13g2_fill_1 FILLER_70_224 ();
 sg13g2_fill_2 FILLER_70_238 ();
 sg13g2_fill_1 FILLER_70_240 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_fill_2 FILLER_71_84 ();
 sg13g2_fill_2 FILLER_71_113 ();
 sg13g2_fill_1 FILLER_71_115 ();
 sg13g2_fill_2 FILLER_71_153 ();
 sg13g2_fill_1 FILLER_71_167 ();
 sg13g2_fill_2 FILLER_71_178 ();
 sg13g2_fill_2 FILLER_71_203 ();
 sg13g2_fill_1 FILLER_71_205 ();
 sg13g2_decap_8 FILLER_71_215 ();
 sg13g2_decap_8 FILLER_71_222 ();
 sg13g2_fill_2 FILLER_71_229 ();
 sg13g2_fill_1 FILLER_71_231 ();
 sg13g2_fill_2 FILLER_71_236 ();
 sg13g2_decap_4 FILLER_71_247 ();
 sg13g2_fill_2 FILLER_71_268 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_fill_1 FILLER_71_329 ();
 sg13g2_fill_1 FILLER_71_365 ();
 sg13g2_decap_8 FILLER_71_396 ();
 sg13g2_decap_4 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_4 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_98 ();
 sg13g2_fill_1 FILLER_72_110 ();
 sg13g2_fill_2 FILLER_72_116 ();
 sg13g2_fill_2 FILLER_72_127 ();
 sg13g2_fill_1 FILLER_72_145 ();
 sg13g2_fill_1 FILLER_72_159 ();
 sg13g2_fill_1 FILLER_72_207 ();
 sg13g2_decap_8 FILLER_72_241 ();
 sg13g2_fill_2 FILLER_72_248 ();
 sg13g2_fill_1 FILLER_72_250 ();
 sg13g2_decap_8 FILLER_72_256 ();
 sg13g2_decap_4 FILLER_72_263 ();
 sg13g2_fill_2 FILLER_72_267 ();
 sg13g2_fill_2 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_323 ();
 sg13g2_fill_2 FILLER_72_332 ();
 sg13g2_fill_1 FILLER_72_348 ();
 sg13g2_decap_8 FILLER_72_393 ();
 sg13g2_decap_8 FILLER_72_400 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_fill_1 FILLER_73_147 ();
 sg13g2_fill_2 FILLER_73_182 ();
 sg13g2_fill_1 FILLER_73_241 ();
 sg13g2_decap_8 FILLER_73_272 ();
 sg13g2_fill_2 FILLER_73_279 ();
 sg13g2_fill_1 FILLER_73_281 ();
 sg13g2_fill_1 FILLER_73_294 ();
 sg13g2_fill_2 FILLER_73_335 ();
 sg13g2_fill_1 FILLER_73_337 ();
 sg13g2_fill_1 FILLER_73_347 ();
 sg13g2_fill_1 FILLER_73_352 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_fill_1 FILLER_74_84 ();
 sg13g2_fill_1 FILLER_74_133 ();
 sg13g2_fill_2 FILLER_74_146 ();
 sg13g2_fill_1 FILLER_74_160 ();
 sg13g2_fill_1 FILLER_74_170 ();
 sg13g2_fill_2 FILLER_74_190 ();
 sg13g2_fill_1 FILLER_74_192 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_fill_2 FILLER_74_280 ();
 sg13g2_fill_2 FILLER_74_312 ();
 sg13g2_fill_1 FILLER_74_314 ();
 sg13g2_fill_2 FILLER_74_351 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_4 FILLER_75_84 ();
 sg13g2_fill_2 FILLER_75_88 ();
 sg13g2_fill_2 FILLER_75_117 ();
 sg13g2_decap_8 FILLER_75_197 ();
 sg13g2_decap_8 FILLER_75_208 ();
 sg13g2_decap_4 FILLER_75_215 ();
 sg13g2_fill_2 FILLER_75_231 ();
 sg13g2_fill_1 FILLER_75_233 ();
 sg13g2_fill_1 FILLER_75_258 ();
 sg13g2_fill_1 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_4 FILLER_76_77 ();
 sg13g2_fill_2 FILLER_76_190 ();
 sg13g2_decap_4 FILLER_76_215 ();
 sg13g2_fill_2 FILLER_76_219 ();
 sg13g2_fill_1 FILLER_76_256 ();
 sg13g2_fill_1 FILLER_76_299 ();
 sg13g2_fill_1 FILLER_76_353 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_fill_1 FILLER_77_77 ();
 sg13g2_fill_1 FILLER_77_163 ();
 sg13g2_fill_1 FILLER_77_265 ();
 sg13g2_fill_2 FILLER_77_297 ();
 sg13g2_fill_1 FILLER_77_348 ();
 sg13g2_fill_1 FILLER_77_381 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_84 ();
 sg13g2_fill_2 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_165 ();
 sg13g2_fill_2 FILLER_78_175 ();
 sg13g2_fill_2 FILLER_78_282 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_88 ();
 sg13g2_fill_2 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_260 ();
 sg13g2_fill_1 FILLER_79_265 ();
 sg13g2_fill_2 FILLER_79_292 ();
 sg13g2_fill_1 FILLER_79_294 ();
 sg13g2_fill_2 FILLER_79_352 ();
 sg13g2_fill_1 FILLER_79_354 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_decap_8 FILLER_80_84 ();
 sg13g2_decap_8 FILLER_80_91 ();
 sg13g2_fill_2 FILLER_80_98 ();
 sg13g2_fill_1 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_122 ();
 sg13g2_fill_2 FILLER_80_138 ();
 sg13g2_fill_1 FILLER_80_140 ();
 sg13g2_fill_2 FILLER_80_163 ();
 sg13g2_fill_1 FILLER_80_165 ();
 sg13g2_decap_8 FILLER_80_184 ();
 sg13g2_fill_1 FILLER_80_191 ();
 sg13g2_fill_2 FILLER_80_196 ();
 sg13g2_fill_1 FILLER_80_207 ();
 sg13g2_fill_1 FILLER_80_229 ();
 sg13g2_fill_2 FILLER_80_310 ();
 sg13g2_fill_2 FILLER_80_317 ();
 sg13g2_fill_1 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uo_out[3] = net12;
 assign uo_out[4] = net13;
 assign uo_out[6] = net14;
endmodule

module tt_um_ultra_tiny_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \ACC[0] ;
 wire \ACC[1] ;
 wire \ACC[2] ;
 wire \ACC[3] ;
 wire \ACC[4] ;
 wire \ACC[5] ;
 wire \ACC[6] ;
 wire \ACC[7] ;
 wire \B[0] ;
 wire \B[1] ;
 wire \B[2] ;
 wire \B[3] ;
 wire \B[4] ;
 wire \B[5] ;
 wire \B[6] ;
 wire \B[7] ;
 wire \IR[0] ;
 wire \IR[1] ;
 wire \IR[2] ;
 wire \IR[4] ;
 wire \IR[5] ;
 wire \IR[6] ;
 wire \IR[7] ;
 wire \PC[0] ;
 wire \PC[1] ;
 wire \PC[2] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire clknet_0_clk;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;

 sg13g2_inv_1 _0644_ (.Y(_0107_),
    .A(net128));
 sg13g2_inv_1 _0645_ (.Y(_0108_),
    .A(net129));
 sg13g2_inv_1 _0646_ (.Y(_0109_),
    .A(_0004_));
 sg13g2_inv_1 _0647_ (.Y(_0110_),
    .A(net97));
 sg13g2_inv_1 _0648_ (.Y(_0111_),
    .A(net93));
 sg13g2_inv_1 _0649_ (.Y(_0112_),
    .A(net94));
 sg13g2_inv_1 _0650_ (.Y(_0113_),
    .A(net95));
 sg13g2_inv_1 _0651_ (.Y(_0114_),
    .A(net229));
 sg13g2_nor2_2 _0652_ (.A(net127),
    .B(net129),
    .Y(_0115_));
 sg13g2_nor2_2 _0653_ (.A(net122),
    .B(net129),
    .Y(_0116_));
 sg13g2_inv_1 _0654_ (.Y(_0117_),
    .A(_0116_));
 sg13g2_a21oi_1 _0655_ (.A1(net130),
    .A2(net147),
    .Y(_0118_),
    .B1(_0116_));
 sg13g2_and2_1 _0656_ (.A(net1),
    .B(_0118_),
    .X(_0016_));
 sg13g2_nor2_2 _0657_ (.A(\IR[7] ),
    .B(\IR[6] ),
    .Y(_0119_));
 sg13g2_nor2b_2 _0658_ (.A(\IR[5] ),
    .B_N(\IR[4] ),
    .Y(_0120_));
 sg13g2_nand2_1 _0659_ (.Y(_0121_),
    .A(_0119_),
    .B(_0120_));
 sg13g2_nor2_2 _0660_ (.A(\IR[4] ),
    .B(\IR[5] ),
    .Y(_0122_));
 sg13g2_nor2b_2 _0661_ (.A(\IR[6] ),
    .B_N(\IR[7] ),
    .Y(_0123_));
 sg13g2_a22oi_1 _0662_ (.Y(_0124_),
    .B1(_0122_),
    .B2(_0123_),
    .A2(_0120_),
    .A1(_0119_));
 sg13g2_nor2b_2 _0663_ (.A(net131),
    .B_N(net1),
    .Y(_0125_));
 sg13g2_nand2_1 _0664_ (.Y(_0126_),
    .A(net167),
    .B(_0125_));
 sg13g2_nand3_1 _0665_ (.B(_0124_),
    .C(_0125_),
    .A(net167),
    .Y(_0127_));
 sg13g2_nand2_1 _0666_ (.Y(_0128_),
    .A(net217),
    .B(_0125_));
 sg13g2_nand3_1 _0667_ (.B(net127),
    .C(net131),
    .A(net1),
    .Y(_0129_));
 sg13g2_nand3_1 _0668_ (.B(_0128_),
    .C(_0129_),
    .A(_0127_),
    .Y(_0000_));
 sg13g2_nand2_1 _0669_ (.Y(_0130_),
    .A(net147),
    .B(_0125_));
 sg13g2_nand3_1 _0670_ (.B(net131),
    .C(net167),
    .A(net1),
    .Y(_0131_));
 sg13g2_nand2_1 _0671_ (.Y(_0001_),
    .A(net120),
    .B(_0131_));
 sg13g2_nand3_1 _0672_ (.B(net131),
    .C(\state[3] ),
    .A(net1),
    .Y(_0132_));
 sg13g2_o21ai_1 _0673_ (.B1(_0132_),
    .Y(_0002_),
    .A1(_0124_),
    .A2(_0126_));
 sg13g2_a21o_1 _0674_ (.A2(_0123_),
    .A1(_0120_),
    .B1(_0117_),
    .X(_0133_));
 sg13g2_nand3_1 _0675_ (.B(net1),
    .C(_0133_),
    .A(net137),
    .Y(_0134_));
 sg13g2_a21oi_1 _0676_ (.A1(_0108_),
    .A2(_0004_),
    .Y(_0135_),
    .B1(_0134_));
 sg13g2_nand2_1 _0677_ (.Y(_0136_),
    .A(\IR[1] ),
    .B(\IR[0] ));
 sg13g2_nor2_1 _0678_ (.A(_0003_),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_inv_1 _0679_ (.Y(_0138_),
    .A(_0137_));
 sg13g2_nand2_1 _0680_ (.Y(_0139_),
    .A(net3),
    .B(net2));
 sg13g2_nand3_1 _0681_ (.B(net2),
    .C(net4),
    .A(net3),
    .Y(_0140_));
 sg13g2_a22oi_1 _0682_ (.Y(_0141_),
    .B1(_0140_),
    .B2(net130),
    .A2(_0138_),
    .A1(_0116_));
 sg13g2_nand2_2 _0683_ (.Y(_0142_),
    .A(_0135_),
    .B(_0141_));
 sg13g2_mux2_2 _0684_ (.A0(\ACC[0] ),
    .A1(net5),
    .S(net132),
    .X(_0143_));
 sg13g2_mux2_1 _0685_ (.A0(_0143_),
    .A1(net197),
    .S(_0142_),
    .X(_0017_));
 sg13g2_nand2_1 _0686_ (.Y(_0144_),
    .A(net132),
    .B(net6));
 sg13g2_o21ai_1 _0687_ (.B1(_0144_),
    .Y(_0145_),
    .A1(net132),
    .A2(_0110_));
 sg13g2_mux2_1 _0688_ (.A0(_0145_),
    .A1(net185),
    .S(_0142_),
    .X(_0018_));
 sg13g2_nand2_1 _0689_ (.Y(_0146_),
    .A(net133),
    .B(net7));
 sg13g2_o21ai_1 _0690_ (.B1(_0146_),
    .Y(_0147_),
    .A1(net133),
    .A2(_0111_));
 sg13g2_mux2_1 _0691_ (.A0(_0147_),
    .A1(net165),
    .S(_0142_),
    .X(_0019_));
 sg13g2_mux2_2 _0692_ (.A0(net126),
    .A1(net8),
    .S(net132),
    .X(_0148_));
 sg13g2_mux2_1 _0693_ (.A0(_0148_),
    .A1(net191),
    .S(_0142_),
    .X(_0020_));
 sg13g2_nand2_1 _0694_ (.Y(_0149_),
    .A(net133),
    .B(net9));
 sg13g2_o21ai_1 _0695_ (.B1(_0149_),
    .Y(_0150_),
    .A1(net133),
    .A2(_0112_));
 sg13g2_mux2_1 _0696_ (.A0(_0150_),
    .A1(net189),
    .S(_0142_),
    .X(_0021_));
 sg13g2_mux2_2 _0697_ (.A0(net125),
    .A1(net10),
    .S(net133),
    .X(_0151_));
 sg13g2_mux2_1 _0698_ (.A0(_0151_),
    .A1(net190),
    .S(_0142_),
    .X(_0022_));
 sg13g2_nand2_1 _0699_ (.Y(_0152_),
    .A(net133),
    .B(net11));
 sg13g2_o21ai_1 _0700_ (.B1(_0152_),
    .Y(_0153_),
    .A1(net133),
    .A2(_0113_));
 sg13g2_mux2_1 _0701_ (.A0(_0153_),
    .A1(net181),
    .S(_0142_),
    .X(_0023_));
 sg13g2_mux2_2 _0702_ (.A0(\ACC[7] ),
    .A1(net12),
    .S(net133),
    .X(_0154_));
 sg13g2_mux2_1 _0703_ (.A0(_0154_),
    .A1(net195),
    .S(_0142_),
    .X(_0024_));
 sg13g2_nand3_1 _0704_ (.B(_0123_),
    .C(_0125_),
    .A(_0122_),
    .Y(_0155_));
 sg13g2_nor2_1 _0705_ (.A(net102),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_nor2_1 _0706_ (.A(\B[0] ),
    .B(_0156_),
    .Y(_0157_));
 sg13g2_o21ai_1 _0707_ (.B1(net123),
    .Y(_0158_),
    .A1(\PC[2] ),
    .A2(_0007_));
 sg13g2_o21ai_1 _0708_ (.B1(_0158_),
    .Y(_0159_),
    .A1(net123),
    .A2(_0007_));
 sg13g2_nor2_2 _0709_ (.A(net124),
    .B(_0159_),
    .Y(_0160_));
 sg13g2_or2_2 _0710_ (.X(_0161_),
    .B(_0159_),
    .A(net124));
 sg13g2_nor2b_1 _0711_ (.A(net124),
    .B_N(net123),
    .Y(_0162_));
 sg13g2_and2_2 _0712_ (.A(\PC[2] ),
    .B(_0162_),
    .X(_0163_));
 sg13g2_and3_1 _0713_ (.X(_0164_),
    .A(net124),
    .B(net123),
    .C(\PC[2] ));
 sg13g2_a22oi_1 _0714_ (.Y(_0165_),
    .B1(net117),
    .B2(\mem[7][0] ),
    .A2(_0163_),
    .A1(\mem[6][0] ));
 sg13g2_and2_2 _0715_ (.A(_0007_),
    .B(_0162_),
    .X(_0166_));
 sg13g2_nand2_1 _0716_ (.Y(_0167_),
    .A(\mem[2][0] ),
    .B(_0166_));
 sg13g2_nor2b_1 _0717_ (.A(net123),
    .B_N(net124),
    .Y(_0168_));
 sg13g2_and2_2 _0718_ (.A(_0007_),
    .B(_0168_),
    .X(_0169_));
 sg13g2_nor2b_2 _0719_ (.A(_0007_),
    .B_N(_0168_),
    .Y(_0170_));
 sg13g2_and3_2 _0720_ (.X(_0171_),
    .A(net124),
    .B(net123),
    .C(_0114_));
 sg13g2_nor3_2 _0721_ (.A(net124),
    .B(net123),
    .C(_0007_),
    .Y(_0172_));
 sg13g2_a22oi_1 _0722_ (.Y(_0173_),
    .B1(_0172_),
    .B2(\mem[4][0] ),
    .A2(_0169_),
    .A1(\mem[1][0] ));
 sg13g2_a22oi_1 _0723_ (.Y(_0174_),
    .B1(_0171_),
    .B2(\mem[3][0] ),
    .A2(_0170_),
    .A1(\mem[5][0] ));
 sg13g2_nand4_1 _0724_ (.B(_0167_),
    .C(_0173_),
    .A(_0165_),
    .Y(_0175_),
    .D(_0174_));
 sg13g2_a21oi_2 _0725_ (.B1(_0175_),
    .Y(_0176_),
    .A2(_0160_),
    .A1(net212));
 sg13g2_a21oi_1 _0726_ (.A1(net109),
    .A2(_0176_),
    .Y(_0025_),
    .B1(net103));
 sg13g2_a22oi_1 _0727_ (.Y(_0177_),
    .B1(_0170_),
    .B2(\mem[5][1] ),
    .A2(_0163_),
    .A1(\mem[6][1] ));
 sg13g2_a22oi_1 _0728_ (.Y(_0178_),
    .B1(_0166_),
    .B2(\mem[2][1] ),
    .A2(net117),
    .A1(\mem[7][1] ));
 sg13g2_and2_1 _0729_ (.A(_0177_),
    .B(_0178_),
    .X(_0179_));
 sg13g2_a21oi_1 _0730_ (.A1(\mem[4][1] ),
    .A2(_0172_),
    .Y(_0180_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0731_ (.Y(_0181_),
    .B1(_0171_),
    .B2(\mem[3][1] ),
    .A2(_0169_),
    .A1(\mem[1][1] ));
 sg13g2_nand3_1 _0732_ (.B(_0180_),
    .C(_0181_),
    .A(_0179_),
    .Y(_0182_));
 sg13g2_o21ai_1 _0733_ (.B1(_0182_),
    .Y(_0183_),
    .A1(\mem[0][1] ),
    .A2(_0161_));
 sg13g2_nor2_1 _0734_ (.A(net228),
    .B(net109),
    .Y(_0184_));
 sg13g2_a21oi_1 _0735_ (.A1(net109),
    .A2(_0183_),
    .Y(_0026_),
    .B1(_0184_));
 sg13g2_nor2_1 _0736_ (.A(net223),
    .B(net109),
    .Y(_0185_));
 sg13g2_a22oi_1 _0737_ (.Y(_0186_),
    .B1(_0171_),
    .B2(\mem[3][2] ),
    .A2(_0163_),
    .A1(\mem[6][2] ));
 sg13g2_a22oi_1 _0738_ (.Y(_0187_),
    .B1(_0172_),
    .B2(\mem[4][2] ),
    .A2(_0169_),
    .A1(\mem[1][2] ));
 sg13g2_and2_1 _0739_ (.A(_0186_),
    .B(_0187_),
    .X(_0188_));
 sg13g2_a21oi_1 _0740_ (.A1(\mem[2][2] ),
    .A2(_0166_),
    .Y(_0189_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0741_ (.Y(_0190_),
    .B1(_0170_),
    .B2(\mem[5][2] ),
    .A2(net117),
    .A1(\mem[7][2] ));
 sg13g2_nand3_1 _0742_ (.B(_0189_),
    .C(_0190_),
    .A(_0188_),
    .Y(_0191_));
 sg13g2_o21ai_1 _0743_ (.B1(_0191_),
    .Y(_0192_),
    .A1(net198),
    .A2(_0161_));
 sg13g2_a21oi_1 _0744_ (.A1(net109),
    .A2(_0192_),
    .Y(_0027_),
    .B1(_0185_));
 sg13g2_nor2_1 _0745_ (.A(net216),
    .B(net109),
    .Y(_0193_));
 sg13g2_nand2b_1 _0746_ (.Y(_0194_),
    .B(_0160_),
    .A_N(net199));
 sg13g2_a22oi_1 _0747_ (.Y(_0195_),
    .B1(_0169_),
    .B2(\mem[1][3] ),
    .A2(_0163_),
    .A1(\mem[6][3] ));
 sg13g2_a22oi_1 _0748_ (.Y(_0196_),
    .B1(_0166_),
    .B2(\mem[2][3] ),
    .A2(net117),
    .A1(\mem[7][3] ));
 sg13g2_nand2_1 _0749_ (.Y(_0197_),
    .A(_0195_),
    .B(_0196_));
 sg13g2_nand2_1 _0750_ (.Y(_0198_),
    .A(\mem[4][3] ),
    .B(_0172_));
 sg13g2_a22oi_1 _0751_ (.Y(_0199_),
    .B1(_0171_),
    .B2(\mem[3][3] ),
    .A2(_0170_),
    .A1(\mem[5][3] ));
 sg13g2_nand3_1 _0752_ (.B(_0198_),
    .C(_0199_),
    .A(_0161_),
    .Y(_0200_));
 sg13g2_o21ai_1 _0753_ (.B1(_0194_),
    .Y(_0201_),
    .A1(_0197_),
    .A2(_0200_));
 sg13g2_a21oi_1 _0754_ (.A1(net109),
    .A2(_0201_),
    .Y(_0028_),
    .B1(_0193_));
 sg13g2_nor2_1 _0755_ (.A(net221),
    .B(net108),
    .Y(_0202_));
 sg13g2_a22oi_1 _0756_ (.Y(_0203_),
    .B1(_0172_),
    .B2(\mem[4][4] ),
    .A2(_0163_),
    .A1(\mem[6][4] ));
 sg13g2_a22oi_1 _0757_ (.Y(_0204_),
    .B1(_0170_),
    .B2(\mem[5][4] ),
    .A2(_0169_),
    .A1(\mem[1][4] ));
 sg13g2_and2_1 _0758_ (.A(_0203_),
    .B(_0204_),
    .X(_0205_));
 sg13g2_a21oi_1 _0759_ (.A1(\mem[7][4] ),
    .A2(net117),
    .Y(_0206_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0760_ (.Y(_0207_),
    .B1(_0171_),
    .B2(\mem[3][4] ),
    .A2(_0166_),
    .A1(\mem[2][4] ));
 sg13g2_nand3_1 _0761_ (.B(_0206_),
    .C(_0207_),
    .A(_0205_),
    .Y(_0208_));
 sg13g2_o21ai_1 _0762_ (.B1(_0208_),
    .Y(_0209_),
    .A1(\mem[0][4] ),
    .A2(_0161_));
 sg13g2_a21oi_1 _0763_ (.A1(net108),
    .A2(_0209_),
    .Y(_0029_),
    .B1(_0202_));
 sg13g2_a22oi_1 _0764_ (.Y(_0210_),
    .B1(net117),
    .B2(\mem[7][5] ),
    .A2(_0163_),
    .A1(\mem[6][5] ));
 sg13g2_a22oi_1 _0765_ (.Y(_0211_),
    .B1(_0170_),
    .B2(\mem[5][5] ),
    .A2(_0166_),
    .A1(\mem[2][5] ));
 sg13g2_a22oi_1 _0766_ (.Y(_0212_),
    .B1(_0171_),
    .B2(\mem[3][5] ),
    .A2(_0169_),
    .A1(\mem[1][5] ));
 sg13g2_and2_1 _0767_ (.A(_0211_),
    .B(_0212_),
    .X(_0213_));
 sg13g2_a21oi_1 _0768_ (.A1(\mem[4][5] ),
    .A2(_0172_),
    .Y(_0214_),
    .B1(_0160_));
 sg13g2_nand3_1 _0769_ (.B(_0213_),
    .C(_0214_),
    .A(_0210_),
    .Y(_0215_));
 sg13g2_o21ai_1 _0770_ (.B1(_0215_),
    .Y(_0216_),
    .A1(\mem[0][5] ),
    .A2(_0161_));
 sg13g2_nor2_1 _0771_ (.A(net207),
    .B(net108),
    .Y(_0217_));
 sg13g2_a21oi_1 _0772_ (.A1(net108),
    .A2(_0216_),
    .Y(_0030_),
    .B1(_0217_));
 sg13g2_a22oi_1 _0773_ (.Y(_0218_),
    .B1(_0172_),
    .B2(\mem[4][6] ),
    .A2(_0169_),
    .A1(\mem[1][6] ));
 sg13g2_a22oi_1 _0774_ (.Y(_0219_),
    .B1(_0170_),
    .B2(\mem[5][6] ),
    .A2(net117),
    .A1(\mem[7][6] ));
 sg13g2_and2_1 _0775_ (.A(_0218_),
    .B(_0219_),
    .X(_0220_));
 sg13g2_a21oi_1 _0776_ (.A1(\mem[2][6] ),
    .A2(_0166_),
    .Y(_0221_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0777_ (.Y(_0222_),
    .B1(_0171_),
    .B2(\mem[3][6] ),
    .A2(_0163_),
    .A1(\mem[6][6] ));
 sg13g2_nand3_1 _0778_ (.B(_0221_),
    .C(_0222_),
    .A(_0220_),
    .Y(_0223_));
 sg13g2_o21ai_1 _0779_ (.B1(_0223_),
    .Y(_0224_),
    .A1(net200),
    .A2(_0161_));
 sg13g2_nor2_1 _0780_ (.A(net215),
    .B(net108),
    .Y(_0225_));
 sg13g2_a21oi_1 _0781_ (.A1(net108),
    .A2(_0224_),
    .Y(_0031_),
    .B1(_0225_));
 sg13g2_a22oi_1 _0782_ (.Y(_0226_),
    .B1(_0172_),
    .B2(\mem[4][7] ),
    .A2(_0169_),
    .A1(\mem[1][7] ));
 sg13g2_a22oi_1 _0783_ (.Y(_0227_),
    .B1(_0171_),
    .B2(\mem[3][7] ),
    .A2(_0163_),
    .A1(\mem[6][7] ));
 sg13g2_a21o_1 _0784_ (.A2(_0170_),
    .A1(\mem[5][7] ),
    .B1(_0160_),
    .X(_0228_));
 sg13g2_a221oi_1 _0785_ (.B2(\mem[2][7] ),
    .C1(_0228_),
    .B1(_0166_),
    .A1(\mem[7][7] ),
    .Y(_0229_),
    .A2(net117));
 sg13g2_nand3_1 _0786_ (.B(_0227_),
    .C(_0229_),
    .A(_0226_),
    .Y(_0230_));
 sg13g2_o21ai_1 _0787_ (.B1(_0230_),
    .Y(_0231_),
    .A1(net231),
    .A2(_0161_));
 sg13g2_nor2_1 _0788_ (.A(net176),
    .B(net108),
    .Y(_0232_));
 sg13g2_a21oi_1 _0789_ (.A1(net108),
    .A2(_0231_),
    .Y(_0032_),
    .B1(_0232_));
 sg13g2_nor2b_2 _0790_ (.A(\IR[7] ),
    .B_N(\IR[6] ),
    .Y(_0233_));
 sg13g2_nor2b_1 _0791_ (.A(\IR[4] ),
    .B_N(\IR[5] ),
    .Y(_0234_));
 sg13g2_and2_1 _0792_ (.A(_0123_),
    .B(_0234_),
    .X(_0235_));
 sg13g2_nor2_1 _0793_ (.A(_0233_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_a21oi_1 _0794_ (.A1(\IR[5] ),
    .A2(_0119_),
    .Y(_0237_),
    .B1(net122));
 sg13g2_nand2_1 _0795_ (.Y(_0238_),
    .A(net107),
    .B(_0237_));
 sg13g2_o21ai_1 _0796_ (.B1(_0125_),
    .Y(_0239_),
    .A1(net127),
    .A2(\state[3] ));
 sg13g2_a21oi_1 _0797_ (.A1(\state[3] ),
    .A2(_0121_),
    .Y(_0240_),
    .B1(_0239_));
 sg13g2_nand2_1 _0798_ (.Y(_0241_),
    .A(_0238_),
    .B(_0240_));
 sg13g2_nand2b_1 _0799_ (.Y(_0242_),
    .B(\IR[0] ),
    .A_N(\IR[1] ));
 sg13g2_nor2_1 _0800_ (.A(_0003_),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_inv_1 _0801_ (.Y(_0244_),
    .A(_0243_));
 sg13g2_a22oi_1 _0802_ (.Y(_0245_),
    .B1(net114),
    .B2(\mem[5][0] ),
    .A2(net116),
    .A1(\mem[7][0] ));
 sg13g2_nor2_1 _0803_ (.A(\IR[2] ),
    .B(_0242_),
    .Y(_0246_));
 sg13g2_nor2_2 _0804_ (.A(\IR[1] ),
    .B(\IR[0] ),
    .Y(_0247_));
 sg13g2_nor2_1 _0805_ (.A(\IR[2] ),
    .B(_0247_),
    .Y(_0248_));
 sg13g2_nor2b_2 _0806_ (.A(_0248_),
    .B_N(_0003_),
    .Y(_0249_));
 sg13g2_o21ai_1 _0807_ (.B1(_0003_),
    .Y(_0250_),
    .A1(\IR[2] ),
    .A2(_0247_));
 sg13g2_nand2b_1 _0808_ (.Y(_0251_),
    .B(\IR[1] ),
    .A_N(\IR[0] ));
 sg13g2_nor2_1 _0809_ (.A(\IR[2] ),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_nor2_1 _0810_ (.A(\IR[2] ),
    .B(_0136_),
    .Y(_0253_));
 sg13g2_a22oi_1 _0811_ (.Y(_0254_),
    .B1(_0253_),
    .B2(\mem[3][0] ),
    .A2(net112),
    .A1(\mem[2][0] ));
 sg13g2_nor3_2 _0812_ (.A(\IR[1] ),
    .B(\IR[0] ),
    .C(_0003_),
    .Y(_0255_));
 sg13g2_inv_1 _0813_ (.Y(_0256_),
    .A(_0255_));
 sg13g2_nor2_1 _0814_ (.A(_0003_),
    .B(_0251_),
    .Y(_0257_));
 sg13g2_a22oi_1 _0815_ (.Y(_0258_),
    .B1(_0255_),
    .B2(\mem[4][0] ),
    .A2(net113),
    .A1(\mem[1][0] ));
 sg13g2_nand3_1 _0816_ (.B(_0254_),
    .C(_0258_),
    .A(_0245_),
    .Y(_0259_));
 sg13g2_a22oi_1 _0817_ (.Y(_0260_),
    .B1(_0257_),
    .B2(\mem[6][0] ),
    .A2(_0249_),
    .A1(\mem[0][0] ));
 sg13g2_nand2b_1 _0818_ (.Y(_0261_),
    .B(_0260_),
    .A_N(_0259_));
 sg13g2_nand2_2 _0819_ (.Y(_0262_),
    .A(_0120_),
    .B(_0233_));
 sg13g2_and2_1 _0820_ (.A(\ACC[0] ),
    .B(\B[0] ),
    .X(_0263_));
 sg13g2_nand3b_1 _0821_ (.B(\IR[5] ),
    .C(_0233_),
    .Y(_0264_),
    .A_N(\IR[4] ));
 sg13g2_nor2b_1 _0822_ (.A(net107),
    .B_N(_0264_),
    .Y(_0265_));
 sg13g2_o21ai_1 _0823_ (.B1(_0262_),
    .Y(_0266_),
    .A1(_0263_),
    .A2(_0265_));
 sg13g2_o21ai_1 _0824_ (.B1(_0266_),
    .Y(_0267_),
    .A1(\ACC[0] ),
    .A2(\B[0] ));
 sg13g2_and2_2 _0825_ (.A(_0122_),
    .B(_0233_),
    .X(_0268_));
 sg13g2_and2_2 _0826_ (.A(\IR[4] ),
    .B(\IR[5] ),
    .X(_0269_));
 sg13g2_nand2_2 _0827_ (.Y(_0270_),
    .A(_0233_),
    .B(_0269_));
 sg13g2_o21ai_1 _0828_ (.B1(net127),
    .Y(_0271_),
    .A1(\ACC[0] ),
    .A2(_0270_));
 sg13g2_a221oi_1 _0829_ (.B2(_0268_),
    .C1(_0271_),
    .B1(_0263_),
    .A1(net115),
    .Y(_0272_),
    .A2(_0261_));
 sg13g2_a221oi_1 _0830_ (.B2(_0272_),
    .C1(_0241_),
    .B1(_0267_),
    .A1(net122),
    .Y(_0273_),
    .A2(_0176_));
 sg13g2_a21o_1 _0831_ (.A2(net105),
    .A1(net96),
    .B1(_0273_),
    .X(_0033_));
 sg13g2_nor2b_1 _0832_ (.A(\ACC[0] ),
    .B_N(\B[0] ),
    .Y(_0274_));
 sg13g2_and2_2 _0833_ (.A(_0119_),
    .B(_0269_),
    .X(_0275_));
 sg13g2_nand2_2 _0834_ (.Y(_0276_),
    .A(_0119_),
    .B(_0269_));
 sg13g2_nor2_1 _0835_ (.A(\B[0] ),
    .B(\B[1] ),
    .Y(_0277_));
 sg13g2_xnor2_1 _0836_ (.Y(_0278_),
    .A(\B[0] ),
    .B(\B[1] ));
 sg13g2_nand3b_1 _0837_ (.B(_0119_),
    .C(_0269_),
    .Y(_0279_),
    .A_N(_0008_));
 sg13g2_a21o_1 _0838_ (.A2(_0269_),
    .A1(_0119_),
    .B1(_0278_),
    .X(_0280_));
 sg13g2_and3_1 _0839_ (.X(_0281_),
    .A(\ACC[1] ),
    .B(_0279_),
    .C(_0280_));
 sg13g2_nand3_1 _0840_ (.B(_0279_),
    .C(_0280_),
    .A(\ACC[1] ),
    .Y(_0282_));
 sg13g2_a21oi_1 _0841_ (.A1(_0279_),
    .A2(_0280_),
    .Y(_0283_),
    .B1(\ACC[1] ));
 sg13g2_nor2_1 _0842_ (.A(_0281_),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_xnor2_1 _0843_ (.Y(_0285_),
    .A(_0274_),
    .B(_0284_));
 sg13g2_a22oi_1 _0844_ (.Y(_0286_),
    .B1(_0255_),
    .B2(\mem[4][1] ),
    .A2(net113),
    .A1(\mem[1][1] ));
 sg13g2_a22oi_1 _0845_ (.Y(_0287_),
    .B1(net111),
    .B2(\mem[3][1] ),
    .A2(net116),
    .A1(\mem[7][1] ));
 sg13g2_a22oi_1 _0846_ (.Y(_0288_),
    .B1(net110),
    .B2(\mem[6][1] ),
    .A2(net112),
    .A1(\mem[2][1] ));
 sg13g2_nand3_1 _0847_ (.B(_0287_),
    .C(_0288_),
    .A(_0286_),
    .Y(_0289_));
 sg13g2_a22oi_1 _0848_ (.Y(_0290_),
    .B1(_0249_),
    .B2(\mem[0][1] ),
    .A2(net114),
    .A1(\mem[5][1] ));
 sg13g2_nand2b_1 _0849_ (.Y(_0291_),
    .B(_0290_),
    .A_N(_0289_));
 sg13g2_and2_1 _0850_ (.A(\ACC[1] ),
    .B(\B[1] ),
    .X(_0292_));
 sg13g2_o21ai_1 _0851_ (.B1(_0262_),
    .Y(_0293_),
    .A1(_0264_),
    .A2(_0292_));
 sg13g2_o21ai_1 _0852_ (.B1(_0293_),
    .Y(_0294_),
    .A1(\ACC[1] ),
    .A2(\B[1] ));
 sg13g2_nand2_1 _0853_ (.Y(_0295_),
    .A(_0268_),
    .B(_0292_));
 sg13g2_nand3_1 _0854_ (.B(_0233_),
    .C(_0269_),
    .A(_0110_),
    .Y(_0296_));
 sg13g2_nand2b_1 _0855_ (.Y(_0297_),
    .B(net122),
    .A_N(_0183_));
 sg13g2_a22oi_1 _0856_ (.Y(_0298_),
    .B1(_0291_),
    .B2(net115),
    .A2(_0285_),
    .A1(net107));
 sg13g2_nand4_1 _0857_ (.B(_0295_),
    .C(_0296_),
    .A(_0294_),
    .Y(_0299_),
    .D(_0298_));
 sg13g2_a21oi_1 _0858_ (.A1(net214),
    .A2(_0299_),
    .Y(_0300_),
    .B1(net105));
 sg13g2_a22oi_1 _0859_ (.Y(_0034_),
    .B1(_0297_),
    .B2(_0300_),
    .A2(net105),
    .A1(_0110_));
 sg13g2_nor3_1 _0860_ (.A(\B[0] ),
    .B(\B[1] ),
    .C(\B[2] ),
    .Y(_0301_));
 sg13g2_xor2_1 _0861_ (.B(_0277_),
    .A(\B[2] ),
    .X(_0302_));
 sg13g2_mux2_1 _0862_ (.A0(_0009_),
    .A1(_0302_),
    .S(_0276_),
    .X(_0303_));
 sg13g2_and2_1 _0863_ (.A(\ACC[2] ),
    .B(_0303_),
    .X(_0304_));
 sg13g2_xnor2_1 _0864_ (.Y(_0305_),
    .A(_0111_),
    .B(_0303_));
 sg13g2_o21ai_1 _0865_ (.B1(_0282_),
    .Y(_0306_),
    .A1(_0274_),
    .A2(_0283_));
 sg13g2_xnor2_1 _0866_ (.Y(_0307_),
    .A(_0305_),
    .B(_0306_));
 sg13g2_a22oi_1 _0867_ (.Y(_0308_),
    .B1(net110),
    .B2(\mem[6][2] ),
    .A2(net111),
    .A1(\mem[3][2] ));
 sg13g2_a22oi_1 _0868_ (.Y(_0309_),
    .B1(net113),
    .B2(\mem[1][2] ),
    .A2(net114),
    .A1(\mem[5][2] ));
 sg13g2_a21oi_1 _0869_ (.A1(\mem[4][2] ),
    .A2(_0247_),
    .Y(_0310_),
    .B1(_0249_));
 sg13g2_a22oi_1 _0870_ (.Y(_0311_),
    .B1(net112),
    .B2(\mem[2][2] ),
    .A2(net116),
    .A1(\mem[7][2] ));
 sg13g2_nand4_1 _0871_ (.B(_0309_),
    .C(_0310_),
    .A(_0308_),
    .Y(_0312_),
    .D(_0311_));
 sg13g2_o21ai_1 _0872_ (.B1(net115),
    .Y(_0313_),
    .A1(\mem[0][2] ),
    .A2(_0250_));
 sg13g2_nor2b_1 _0873_ (.A(_0313_),
    .B_N(_0312_),
    .Y(_0314_));
 sg13g2_and2_1 _0874_ (.A(\ACC[2] ),
    .B(\B[2] ),
    .X(_0315_));
 sg13g2_o21ai_1 _0875_ (.B1(_0262_),
    .Y(_0316_),
    .A1(_0264_),
    .A2(_0315_));
 sg13g2_o21ai_1 _0876_ (.B1(_0316_),
    .Y(_0317_),
    .A1(\ACC[2] ),
    .A2(\B[2] ));
 sg13g2_nand2_1 _0877_ (.Y(_0318_),
    .A(_0268_),
    .B(_0315_));
 sg13g2_o21ai_1 _0878_ (.B1(_0318_),
    .Y(_0319_),
    .A1(\ACC[2] ),
    .A2(_0270_));
 sg13g2_nor3_1 _0879_ (.A(net106),
    .B(_0314_),
    .C(_0319_),
    .Y(_0320_));
 sg13g2_a22oi_1 _0880_ (.Y(_0321_),
    .B1(_0317_),
    .B2(_0320_),
    .A2(_0307_),
    .A1(net107));
 sg13g2_nand2b_1 _0881_ (.Y(_0322_),
    .B(net121),
    .A_N(_0192_));
 sg13g2_a21oi_1 _0882_ (.A1(net128),
    .A2(_0321_),
    .Y(_0323_),
    .B1(net104));
 sg13g2_a22oi_1 _0883_ (.Y(_0035_),
    .B1(_0322_),
    .B2(_0323_),
    .A2(net104),
    .A1(_0111_));
 sg13g2_nand2_1 _0884_ (.Y(_0324_),
    .A(_0010_),
    .B(_0275_));
 sg13g2_or4_2 _0885_ (.A(\B[0] ),
    .B(\B[1] ),
    .C(\B[2] ),
    .D(\B[3] ),
    .X(_0325_));
 sg13g2_xnor2_1 _0886_ (.Y(_0326_),
    .A(\B[3] ),
    .B(_0301_));
 sg13g2_o21ai_1 _0887_ (.B1(_0324_),
    .Y(_0327_),
    .A1(_0275_),
    .A2(_0326_));
 sg13g2_nand2_1 _0888_ (.Y(_0328_),
    .A(\ACC[3] ),
    .B(_0327_));
 sg13g2_nor2_1 _0889_ (.A(\ACC[3] ),
    .B(_0327_),
    .Y(_0329_));
 sg13g2_xnor2_1 _0890_ (.Y(_0330_),
    .A(net126),
    .B(_0327_));
 sg13g2_a21oi_2 _0891_ (.B1(_0304_),
    .Y(_0331_),
    .A2(_0306_),
    .A1(_0305_));
 sg13g2_o21ai_1 _0892_ (.B1(net106),
    .Y(_0332_),
    .A1(_0330_),
    .A2(_0331_));
 sg13g2_a21o_1 _0893_ (.A2(_0331_),
    .A1(_0330_),
    .B1(_0332_),
    .X(_0333_));
 sg13g2_a22oi_1 _0894_ (.Y(_0334_),
    .B1(_0252_),
    .B2(\mem[2][3] ),
    .A2(net116),
    .A1(\mem[7][3] ));
 sg13g2_a22oi_1 _0895_ (.Y(_0335_),
    .B1(net110),
    .B2(\mem[6][3] ),
    .A2(net114),
    .A1(\mem[5][3] ));
 sg13g2_a22oi_1 _0896_ (.Y(_0336_),
    .B1(net111),
    .B2(\mem[3][3] ),
    .A2(net113),
    .A1(\mem[1][3] ));
 sg13g2_a22oi_1 _0897_ (.Y(_0337_),
    .B1(_0255_),
    .B2(\mem[4][3] ),
    .A2(_0249_),
    .A1(\mem[0][3] ));
 sg13g2_nand4_1 _0898_ (.B(_0335_),
    .C(_0336_),
    .A(_0334_),
    .Y(_0338_),
    .D(_0337_));
 sg13g2_and2_1 _0899_ (.A(net126),
    .B(\B[3] ),
    .X(_0339_));
 sg13g2_o21ai_1 _0900_ (.B1(_0262_),
    .Y(_0340_),
    .A1(_0264_),
    .A2(_0339_));
 sg13g2_o21ai_1 _0901_ (.B1(_0340_),
    .Y(_0341_),
    .A1(net126),
    .A2(\B[3] ));
 sg13g2_o21ai_1 _0902_ (.B1(net127),
    .Y(_0342_),
    .A1(net126),
    .A2(_0270_));
 sg13g2_a21oi_1 _0903_ (.A1(_0268_),
    .A2(_0339_),
    .Y(_0343_),
    .B1(_0342_));
 sg13g2_nand2_1 _0904_ (.Y(_0344_),
    .A(_0341_),
    .B(_0343_));
 sg13g2_a21oi_1 _0905_ (.A1(net115),
    .A2(_0338_),
    .Y(_0345_),
    .B1(_0344_));
 sg13g2_a221oi_1 _0906_ (.B2(_0345_),
    .C1(net105),
    .B1(_0333_),
    .A1(net122),
    .Y(_0346_),
    .A2(_0201_));
 sg13g2_a21o_1 _0907_ (.A2(net105),
    .A1(net126),
    .B1(_0346_),
    .X(_0036_));
 sg13g2_xnor2_1 _0908_ (.Y(_0347_),
    .A(\B[4] ),
    .B(_0325_));
 sg13g2_mux2_1 _0909_ (.A0(_0011_),
    .A1(_0347_),
    .S(_0276_),
    .X(_0348_));
 sg13g2_nand2_1 _0910_ (.Y(_0349_),
    .A(\ACC[4] ),
    .B(_0348_));
 sg13g2_inv_1 _0911_ (.Y(_0350_),
    .A(_0349_));
 sg13g2_xnor2_1 _0912_ (.Y(_0351_),
    .A(_0112_),
    .B(_0348_));
 sg13g2_inv_1 _0913_ (.Y(_0352_),
    .A(_0351_));
 sg13g2_o21ai_1 _0914_ (.B1(_0328_),
    .Y(_0353_),
    .A1(_0329_),
    .A2(_0331_));
 sg13g2_a22oi_1 _0915_ (.Y(_0354_),
    .B1(net111),
    .B2(\mem[3][4] ),
    .A2(_0247_),
    .A1(\mem[4][4] ));
 sg13g2_a21oi_1 _0916_ (.A1(\mem[5][4] ),
    .A2(net114),
    .Y(_0355_),
    .B1(_0249_));
 sg13g2_a22oi_1 _0917_ (.Y(_0356_),
    .B1(net112),
    .B2(\mem[2][4] ),
    .A2(net113),
    .A1(\mem[1][4] ));
 sg13g2_a22oi_1 _0918_ (.Y(_0357_),
    .B1(net110),
    .B2(\mem[6][4] ),
    .A2(net116),
    .A1(\mem[7][4] ));
 sg13g2_nand4_1 _0919_ (.B(_0355_),
    .C(_0356_),
    .A(_0354_),
    .Y(_0358_),
    .D(_0357_));
 sg13g2_o21ai_1 _0920_ (.B1(net115),
    .Y(_0359_),
    .A1(\mem[0][4] ),
    .A2(_0250_));
 sg13g2_nor2b_1 _0921_ (.A(_0359_),
    .B_N(_0358_),
    .Y(_0360_));
 sg13g2_and2_1 _0922_ (.A(\ACC[4] ),
    .B(\B[4] ),
    .X(_0361_));
 sg13g2_o21ai_1 _0923_ (.B1(_0262_),
    .Y(_0362_),
    .A1(_0264_),
    .A2(_0361_));
 sg13g2_o21ai_1 _0924_ (.B1(_0362_),
    .Y(_0363_),
    .A1(\ACC[4] ),
    .A2(\B[4] ));
 sg13g2_nand2_1 _0925_ (.Y(_0364_),
    .A(_0268_),
    .B(_0361_));
 sg13g2_o21ai_1 _0926_ (.B1(_0364_),
    .Y(_0365_),
    .A1(\ACC[4] ),
    .A2(_0270_));
 sg13g2_nand2b_1 _0927_ (.Y(_0366_),
    .B(net121),
    .A_N(_0209_));
 sg13g2_xnor2_1 _0928_ (.Y(_0367_),
    .A(_0351_),
    .B(_0353_));
 sg13g2_nor3_1 _0929_ (.A(net106),
    .B(_0360_),
    .C(_0365_),
    .Y(_0368_));
 sg13g2_a22oi_1 _0930_ (.Y(_0369_),
    .B1(_0368_),
    .B2(_0363_),
    .A2(_0367_),
    .A1(net106));
 sg13g2_a21oi_1 _0931_ (.A1(net128),
    .A2(_0369_),
    .Y(_0370_),
    .B1(net105));
 sg13g2_a22oi_1 _0932_ (.Y(_0037_),
    .B1(_0366_),
    .B2(_0370_),
    .A2(net105),
    .A1(_0112_));
 sg13g2_a21oi_1 _0933_ (.A1(_0351_),
    .A2(_0353_),
    .Y(_0371_),
    .B1(_0350_));
 sg13g2_o21ai_1 _0934_ (.B1(\B[5] ),
    .Y(_0372_),
    .A1(\B[4] ),
    .A2(_0325_));
 sg13g2_or3_1 _0935_ (.A(\B[4] ),
    .B(\B[5] ),
    .C(_0325_),
    .X(_0373_));
 sg13g2_a21oi_1 _0936_ (.A1(_0372_),
    .A2(_0373_),
    .Y(_0374_),
    .B1(_0275_));
 sg13g2_a21o_1 _0937_ (.A2(_0275_),
    .A1(_0012_),
    .B1(_0374_),
    .X(_0375_));
 sg13g2_nor2_1 _0938_ (.A(net125),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_xnor2_1 _0939_ (.Y(_0377_),
    .A(net125),
    .B(_0375_));
 sg13g2_o21ai_1 _0940_ (.B1(net106),
    .Y(_0378_),
    .A1(_0371_),
    .A2(_0377_));
 sg13g2_a21o_1 _0941_ (.A2(_0377_),
    .A1(_0371_),
    .B1(_0378_),
    .X(_0379_));
 sg13g2_a22oi_1 _0942_ (.Y(_0380_),
    .B1(net110),
    .B2(\mem[6][5] ),
    .A2(net116),
    .A1(\mem[7][5] ));
 sg13g2_a22oi_1 _0943_ (.Y(_0381_),
    .B1(net111),
    .B2(\mem[3][5] ),
    .A2(net113),
    .A1(\mem[1][5] ));
 sg13g2_a22oi_1 _0944_ (.Y(_0382_),
    .B1(_0255_),
    .B2(\mem[4][5] ),
    .A2(net112),
    .A1(\mem[2][5] ));
 sg13g2_a22oi_1 _0945_ (.Y(_0383_),
    .B1(_0249_),
    .B2(\mem[0][5] ),
    .A2(net114),
    .A1(\mem[5][5] ));
 sg13g2_nand4_1 _0946_ (.B(_0381_),
    .C(_0382_),
    .A(_0380_),
    .Y(_0384_),
    .D(_0383_));
 sg13g2_and2_1 _0947_ (.A(\ACC[5] ),
    .B(\B[5] ),
    .X(_0385_));
 sg13g2_o21ai_1 _0948_ (.B1(_0262_),
    .Y(_0386_),
    .A1(_0264_),
    .A2(_0385_));
 sg13g2_o21ai_1 _0949_ (.B1(_0386_),
    .Y(_0387_),
    .A1(net125),
    .A2(\B[5] ));
 sg13g2_o21ai_1 _0950_ (.B1(net128),
    .Y(_0388_),
    .A1(net125),
    .A2(_0270_));
 sg13g2_a21oi_1 _0951_ (.A1(_0268_),
    .A2(_0385_),
    .Y(_0389_),
    .B1(_0388_));
 sg13g2_nand2_1 _0952_ (.Y(_0390_),
    .A(_0387_),
    .B(_0389_));
 sg13g2_a21oi_1 _0953_ (.A1(net115),
    .A2(_0384_),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_a221oi_1 _0954_ (.B2(_0391_),
    .C1(net104),
    .B1(_0379_),
    .A1(net121),
    .Y(_0392_),
    .A2(_0216_));
 sg13g2_a21o_1 _0955_ (.A2(net104),
    .A1(net125),
    .B1(_0392_),
    .X(_0038_));
 sg13g2_nor2_1 _0956_ (.A(_0352_),
    .B(_0377_),
    .Y(_0393_));
 sg13g2_nor2_1 _0957_ (.A(_0349_),
    .B(_0376_),
    .Y(_0394_));
 sg13g2_a221oi_1 _0958_ (.B2(_0353_),
    .C1(_0394_),
    .B1(_0393_),
    .A1(\ACC[5] ),
    .Y(_0395_),
    .A2(_0375_));
 sg13g2_nand2_1 _0959_ (.Y(_0396_),
    .A(_0013_),
    .B(_0275_));
 sg13g2_nor2_1 _0960_ (.A(\B[6] ),
    .B(_0373_),
    .Y(_0397_));
 sg13g2_xor2_1 _0961_ (.B(_0373_),
    .A(\B[6] ),
    .X(_0398_));
 sg13g2_o21ai_1 _0962_ (.B1(_0396_),
    .Y(_0399_),
    .A1(_0275_),
    .A2(_0398_));
 sg13g2_nand2_1 _0963_ (.Y(_0400_),
    .A(\ACC[6] ),
    .B(_0399_));
 sg13g2_xnor2_1 _0964_ (.Y(_0401_),
    .A(_0113_),
    .B(_0399_));
 sg13g2_inv_1 _0965_ (.Y(_0402_),
    .A(_0401_));
 sg13g2_xnor2_1 _0966_ (.Y(_0403_),
    .A(_0395_),
    .B(_0402_));
 sg13g2_a22oi_1 _0967_ (.Y(_0404_),
    .B1(net110),
    .B2(\mem[6][6] ),
    .A2(net116),
    .A1(\mem[7][6] ));
 sg13g2_a21oi_1 _0968_ (.A1(\mem[4][6] ),
    .A2(_0247_),
    .Y(_0405_),
    .B1(_0249_));
 sg13g2_a22oi_1 _0969_ (.Y(_0406_),
    .B1(net113),
    .B2(\mem[1][6] ),
    .A2(net114),
    .A1(\mem[5][6] ));
 sg13g2_a22oi_1 _0970_ (.Y(_0407_),
    .B1(net111),
    .B2(\mem[3][6] ),
    .A2(net112),
    .A1(\mem[2][6] ));
 sg13g2_nand4_1 _0971_ (.B(_0405_),
    .C(_0406_),
    .A(_0404_),
    .Y(_0408_),
    .D(_0407_));
 sg13g2_o21ai_1 _0972_ (.B1(net115),
    .Y(_0409_),
    .A1(\mem[0][6] ),
    .A2(_0250_));
 sg13g2_nor2b_1 _0973_ (.A(_0409_),
    .B_N(_0408_),
    .Y(_0410_));
 sg13g2_and2_1 _0974_ (.A(\ACC[6] ),
    .B(\B[6] ),
    .X(_0411_));
 sg13g2_o21ai_1 _0975_ (.B1(_0262_),
    .Y(_0412_),
    .A1(_0264_),
    .A2(_0411_));
 sg13g2_o21ai_1 _0976_ (.B1(_0412_),
    .Y(_0413_),
    .A1(\ACC[6] ),
    .A2(\B[6] ));
 sg13g2_nand2_1 _0977_ (.Y(_0414_),
    .A(_0268_),
    .B(_0411_));
 sg13g2_o21ai_1 _0978_ (.B1(_0414_),
    .Y(_0415_),
    .A1(\ACC[6] ),
    .A2(_0270_));
 sg13g2_nor3_1 _0979_ (.A(net106),
    .B(_0410_),
    .C(_0415_),
    .Y(_0416_));
 sg13g2_a22oi_1 _0980_ (.Y(_0417_),
    .B1(_0413_),
    .B2(_0416_),
    .A2(_0403_),
    .A1(net106));
 sg13g2_nand2b_1 _0981_ (.Y(_0418_),
    .B(net121),
    .A_N(_0224_));
 sg13g2_a21oi_1 _0982_ (.A1(net128),
    .A2(_0417_),
    .Y(_0419_),
    .B1(net104));
 sg13g2_a22oi_1 _0983_ (.Y(_0039_),
    .B1(_0418_),
    .B2(_0419_),
    .A2(net104),
    .A1(_0113_));
 sg13g2_o21ai_1 _0984_ (.B1(_0400_),
    .Y(_0420_),
    .A1(_0395_),
    .A2(_0402_));
 sg13g2_xor2_1 _0985_ (.B(_0397_),
    .A(_0014_),
    .X(_0421_));
 sg13g2_mux2_1 _0986_ (.A0(\B[7] ),
    .A1(_0421_),
    .S(_0276_),
    .X(_0422_));
 sg13g2_xor2_1 _0987_ (.B(_0422_),
    .A(\ACC[7] ),
    .X(_0423_));
 sg13g2_xnor2_1 _0988_ (.Y(_0424_),
    .A(_0420_),
    .B(_0423_));
 sg13g2_a22oi_1 _0989_ (.Y(_0425_),
    .B1(net111),
    .B2(\mem[3][7] ),
    .A2(net114),
    .A1(\mem[5][7] ));
 sg13g2_a22oi_1 _0990_ (.Y(_0426_),
    .B1(_0255_),
    .B2(\mem[4][7] ),
    .A2(net113),
    .A1(\mem[1][7] ));
 sg13g2_a22oi_1 _0991_ (.Y(_0427_),
    .B1(net110),
    .B2(\mem[6][7] ),
    .A2(net112),
    .A1(\mem[2][7] ));
 sg13g2_a22oi_1 _0992_ (.Y(_0428_),
    .B1(_0249_),
    .B2(\mem[0][7] ),
    .A2(net116),
    .A1(\mem[7][7] ));
 sg13g2_nand4_1 _0993_ (.B(_0426_),
    .C(_0427_),
    .A(_0425_),
    .Y(_0429_),
    .D(_0428_));
 sg13g2_and2_1 _0994_ (.A(\ACC[7] ),
    .B(\B[7] ),
    .X(_0430_));
 sg13g2_o21ai_1 _0995_ (.B1(_0262_),
    .Y(_0431_),
    .A1(_0264_),
    .A2(_0430_));
 sg13g2_o21ai_1 _0996_ (.B1(_0431_),
    .Y(_0432_),
    .A1(\ACC[7] ),
    .A2(\B[7] ));
 sg13g2_o21ai_1 _0997_ (.B1(net128),
    .Y(_0433_),
    .A1(\ACC[7] ),
    .A2(_0270_));
 sg13g2_a21oi_1 _0998_ (.A1(_0268_),
    .A2(_0430_),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_nand2_1 _0999_ (.Y(_0435_),
    .A(_0432_),
    .B(_0434_));
 sg13g2_a221oi_1 _1000_ (.B2(net115),
    .C1(_0435_),
    .B1(_0429_),
    .A1(net106),
    .Y(_0436_),
    .A2(_0424_));
 sg13g2_a21o_1 _1001_ (.A2(_0231_),
    .A1(net121),
    .B1(net104),
    .X(_0437_));
 sg13g2_nand2_1 _1002_ (.Y(_0438_),
    .A(net100),
    .B(net104));
 sg13g2_o21ai_1 _1003_ (.B1(_0438_),
    .Y(_0040_),
    .A1(_0436_),
    .A2(_0437_));
 sg13g2_nor4_1 _1004_ (.A(net125),
    .B(\ACC[4] ),
    .C(\ACC[7] ),
    .D(\ACC[6] ),
    .Y(_0439_));
 sg13g2_nor4_1 _1005_ (.A(\ACC[1] ),
    .B(\ACC[0] ),
    .C(net126),
    .D(\ACC[2] ),
    .Y(_0440_));
 sg13g2_and3_1 _1006_ (.X(_0441_),
    .A(\IR[7] ),
    .B(\IR[6] ),
    .C(_0122_));
 sg13g2_a21oi_1 _1007_ (.A1(_0439_),
    .A2(_0440_),
    .Y(_0442_),
    .B1(_0004_));
 sg13g2_a21o_1 _1008_ (.A2(_0269_),
    .A1(_0123_),
    .B1(net121),
    .X(_0443_));
 sg13g2_o21ai_1 _1009_ (.B1(_0125_),
    .Y(_0444_),
    .A1(_0109_),
    .A2(\state[3] ));
 sg13g2_a22oi_1 _1010_ (.Y(_0445_),
    .B1(_0444_),
    .B2(net120),
    .A2(_0442_),
    .A1(_0441_));
 sg13g2_o21ai_1 _1011_ (.B1(_0445_),
    .Y(_0446_),
    .A1(_0441_),
    .A2(_0443_));
 sg13g2_nor2b_1 _1012_ (.A(net127),
    .B_N(_0006_),
    .Y(_0447_));
 sg13g2_a21oi_1 _1013_ (.A1(net127),
    .A2(\IR[0] ),
    .Y(_0448_),
    .B1(_0447_));
 sg13g2_nand2_1 _1014_ (.Y(_0449_),
    .A(net98),
    .B(_0446_));
 sg13g2_o21ai_1 _1015_ (.B1(_0449_),
    .Y(_0041_),
    .A1(_0446_),
    .A2(_0448_));
 sg13g2_o21ai_1 _1016_ (.B1(net121),
    .Y(_0450_),
    .A1(_0162_),
    .A2(_0168_));
 sg13g2_nand2_1 _1017_ (.Y(_0451_),
    .A(net127),
    .B(net230));
 sg13g2_a21oi_1 _1018_ (.A1(_0450_),
    .A2(_0451_),
    .Y(_0452_),
    .B1(_0446_));
 sg13g2_a21o_1 _1019_ (.A2(_0446_),
    .A1(net101),
    .B1(_0452_),
    .X(_0042_));
 sg13g2_a21oi_1 _1020_ (.A1(net124),
    .A2(net123),
    .Y(_0453_),
    .B1(net128));
 sg13g2_o21ai_1 _1021_ (.B1(_0114_),
    .Y(_0454_),
    .A1(_0446_),
    .A2(_0453_));
 sg13g2_nand2_1 _1022_ (.Y(_0455_),
    .A(net122),
    .B(_0164_));
 sg13g2_o21ai_1 _1023_ (.B1(_0455_),
    .Y(_0456_),
    .A1(net121),
    .A2(\IR[2] ));
 sg13g2_nand2b_1 _1024_ (.Y(_0457_),
    .B(_0456_),
    .A_N(_0446_));
 sg13g2_and2_1 _1025_ (.A(_0454_),
    .B(_0457_),
    .X(_0043_));
 sg13g2_nand2_1 _1026_ (.Y(_0458_),
    .A(net227),
    .B(net120));
 sg13g2_o21ai_1 _1027_ (.B1(_0458_),
    .Y(_0044_),
    .A1(net120),
    .A2(_0176_));
 sg13g2_nand2_1 _1028_ (.Y(_0459_),
    .A(net222),
    .B(net119));
 sg13g2_o21ai_1 _1029_ (.B1(_0459_),
    .Y(_0045_),
    .A1(net119),
    .A2(_0183_));
 sg13g2_nand2_1 _1030_ (.Y(_0460_),
    .A(net226),
    .B(net118));
 sg13g2_o21ai_1 _1031_ (.B1(_0460_),
    .Y(_0046_),
    .A1(net118),
    .A2(_0192_));
 sg13g2_nand2_1 _1032_ (.Y(_0461_),
    .A(net204),
    .B(net119));
 sg13g2_o21ai_1 _1033_ (.B1(_0461_),
    .Y(_0047_),
    .A1(net119),
    .A2(_0209_));
 sg13g2_nand2_1 _1034_ (.Y(_0462_),
    .A(net224),
    .B(net118));
 sg13g2_o21ai_1 _1035_ (.B1(_0462_),
    .Y(_0048_),
    .A1(net118),
    .A2(_0216_));
 sg13g2_nand2_1 _1036_ (.Y(_0463_),
    .A(net211),
    .B(net118));
 sg13g2_o21ai_1 _1037_ (.B1(_0463_),
    .Y(_0049_),
    .A1(net118),
    .A2(_0224_));
 sg13g2_nand2_1 _1038_ (.Y(_0464_),
    .A(net210),
    .B(net118));
 sg13g2_o21ai_1 _1039_ (.B1(_0464_),
    .Y(_0050_),
    .A1(net118),
    .A2(_0231_));
 sg13g2_nor2_2 _1040_ (.A(_0115_),
    .B(_0134_),
    .Y(_0465_));
 sg13g2_nand2b_1 _1041_ (.Y(_0466_),
    .B(_0247_),
    .A_N(\IR[2] ));
 sg13g2_nor2_1 _1042_ (.A(net3),
    .B(net2),
    .Y(_0467_));
 sg13g2_nand2b_1 _1043_ (.Y(_0468_),
    .B(_0467_),
    .A_N(net4));
 sg13g2_a22oi_1 _1044_ (.Y(_0469_),
    .B1(_0468_),
    .B2(net129),
    .A2(_0466_),
    .A1(_0116_));
 sg13g2_nand2_2 _1045_ (.Y(_0470_),
    .A(_0465_),
    .B(_0469_));
 sg13g2_mux2_1 _1046_ (.A0(_0143_),
    .A1(net212),
    .S(_0470_),
    .X(_0051_));
 sg13g2_mux2_1 _1047_ (.A0(_0145_),
    .A1(net196),
    .S(_0470_),
    .X(_0052_));
 sg13g2_mux2_1 _1048_ (.A0(_0147_),
    .A1(net198),
    .S(_0470_),
    .X(_0053_));
 sg13g2_mux2_1 _1049_ (.A0(_0148_),
    .A1(net199),
    .S(_0470_),
    .X(_0054_));
 sg13g2_mux2_1 _1050_ (.A0(_0150_),
    .A1(net193),
    .S(_0470_),
    .X(_0055_));
 sg13g2_mux2_1 _1051_ (.A0(_0151_),
    .A1(net208),
    .S(_0470_),
    .X(_0056_));
 sg13g2_mux2_1 _1052_ (.A0(_0153_),
    .A1(net200),
    .S(_0470_),
    .X(_0057_));
 sg13g2_mux2_1 _1053_ (.A0(_0154_),
    .A1(net218),
    .S(_0470_),
    .X(_0058_));
 sg13g2_nand2b_1 _1054_ (.Y(_0471_),
    .B(net2),
    .A_N(net3));
 sg13g2_o21ai_1 _1055_ (.B1(net129),
    .Y(_0472_),
    .A1(net4),
    .A2(_0471_));
 sg13g2_o21ai_1 _1056_ (.B1(_0472_),
    .Y(_0473_),
    .A1(_0117_),
    .A2(_0246_));
 sg13g2_nor3_2 _1057_ (.A(_0115_),
    .B(_0134_),
    .C(_0473_),
    .Y(_0474_));
 sg13g2_mux2_1 _1058_ (.A0(net154),
    .A1(_0143_),
    .S(_0474_),
    .X(_0059_));
 sg13g2_mux2_1 _1059_ (.A0(net152),
    .A1(_0145_),
    .S(_0474_),
    .X(_0060_));
 sg13g2_mux2_1 _1060_ (.A0(net163),
    .A1(_0147_),
    .S(_0474_),
    .X(_0061_));
 sg13g2_mux2_1 _1061_ (.A0(net162),
    .A1(_0148_),
    .S(_0474_),
    .X(_0062_));
 sg13g2_mux2_1 _1062_ (.A0(net160),
    .A1(_0150_),
    .S(_0474_),
    .X(_0063_));
 sg13g2_mux2_1 _1063_ (.A0(net142),
    .A1(_0151_),
    .S(_0474_),
    .X(_0064_));
 sg13g2_mux2_1 _1064_ (.A0(net153),
    .A1(_0153_),
    .S(_0474_),
    .X(_0065_));
 sg13g2_mux2_1 _1065_ (.A0(net144),
    .A1(_0154_),
    .S(_0474_),
    .X(_0066_));
 sg13g2_nand2b_1 _1066_ (.Y(_0475_),
    .B(net3),
    .A_N(net2));
 sg13g2_o21ai_1 _1067_ (.B1(net130),
    .Y(_0476_),
    .A1(net4),
    .A2(_0475_));
 sg13g2_o21ai_1 _1068_ (.B1(_0476_),
    .Y(_0477_),
    .A1(_0117_),
    .A2(net112));
 sg13g2_nor3_2 _1069_ (.A(_0115_),
    .B(_0134_),
    .C(_0477_),
    .Y(_0478_));
 sg13g2_mux2_1 _1070_ (.A0(net172),
    .A1(_0143_),
    .S(_0478_),
    .X(_0067_));
 sg13g2_mux2_1 _1071_ (.A0(net157),
    .A1(_0145_),
    .S(_0478_),
    .X(_0068_));
 sg13g2_mux2_1 _1072_ (.A0(net166),
    .A1(_0147_),
    .S(_0478_),
    .X(_0069_));
 sg13g2_mux2_1 _1073_ (.A0(net158),
    .A1(_0148_),
    .S(_0478_),
    .X(_0070_));
 sg13g2_mux2_1 _1074_ (.A0(net171),
    .A1(_0150_),
    .S(_0478_),
    .X(_0071_));
 sg13g2_mux2_1 _1075_ (.A0(net146),
    .A1(_0151_),
    .S(_0478_),
    .X(_0072_));
 sg13g2_mux2_1 _1076_ (.A0(net164),
    .A1(_0153_),
    .S(_0478_),
    .X(_0073_));
 sg13g2_mux2_1 _1077_ (.A0(net159),
    .A1(_0154_),
    .S(_0478_),
    .X(_0074_));
 sg13g2_nand2b_1 _1078_ (.Y(_0479_),
    .B(_0116_),
    .A_N(net111));
 sg13g2_o21ai_1 _1079_ (.B1(net129),
    .Y(_0480_),
    .A1(net4),
    .A2(_0139_));
 sg13g2_nand3_1 _1080_ (.B(_0479_),
    .C(_0480_),
    .A(_0465_),
    .Y(_0481_));
 sg13g2_mux2_1 _1081_ (.A0(_0143_),
    .A1(net184),
    .S(_0481_),
    .X(_0075_));
 sg13g2_mux2_1 _1082_ (.A0(_0145_),
    .A1(net187),
    .S(_0481_),
    .X(_0076_));
 sg13g2_mux2_1 _1083_ (.A0(_0147_),
    .A1(net182),
    .S(_0481_),
    .X(_0077_));
 sg13g2_mux2_1 _1084_ (.A0(_0148_),
    .A1(net186),
    .S(_0481_),
    .X(_0078_));
 sg13g2_mux2_1 _1085_ (.A0(_0150_),
    .A1(net178),
    .S(_0481_),
    .X(_0079_));
 sg13g2_mux2_1 _1086_ (.A0(_0151_),
    .A1(net179),
    .S(_0481_),
    .X(_0080_));
 sg13g2_mux2_1 _1087_ (.A0(_0153_),
    .A1(net192),
    .S(_0481_),
    .X(_0081_));
 sg13g2_mux2_1 _1088_ (.A0(_0154_),
    .A1(net180),
    .S(_0481_),
    .X(_0082_));
 sg13g2_nand2_1 _1089_ (.Y(_0482_),
    .A(net4),
    .B(_0467_));
 sg13g2_a22oi_1 _1090_ (.Y(_0483_),
    .B1(_0482_),
    .B2(net129),
    .A2(_0256_),
    .A1(_0116_));
 sg13g2_nand2_2 _1091_ (.Y(_0484_),
    .A(_0465_),
    .B(_0483_));
 sg13g2_mux2_1 _1092_ (.A0(_0143_),
    .A1(net206),
    .S(_0484_),
    .X(_0083_));
 sg13g2_mux2_1 _1093_ (.A0(_0145_),
    .A1(net209),
    .S(_0484_),
    .X(_0084_));
 sg13g2_mux2_1 _1094_ (.A0(_0147_),
    .A1(net213),
    .S(_0484_),
    .X(_0085_));
 sg13g2_mux2_1 _1095_ (.A0(_0148_),
    .A1(net203),
    .S(_0484_),
    .X(_0086_));
 sg13g2_mux2_1 _1096_ (.A0(_0150_),
    .A1(net201),
    .S(_0484_),
    .X(_0087_));
 sg13g2_mux2_1 _1097_ (.A0(_0151_),
    .A1(net194),
    .S(_0484_),
    .X(_0088_));
 sg13g2_mux2_1 _1098_ (.A0(_0153_),
    .A1(net202),
    .S(_0484_),
    .X(_0089_));
 sg13g2_mux2_1 _1099_ (.A0(_0154_),
    .A1(net188),
    .S(_0484_),
    .X(_0090_));
 sg13g2_nand3b_1 _1100_ (.B(net2),
    .C(net4),
    .Y(_0485_),
    .A_N(net3));
 sg13g2_a22oi_1 _1101_ (.Y(_0486_),
    .B1(_0485_),
    .B2(net129),
    .A2(_0244_),
    .A1(_0116_));
 sg13g2_and2_2 _1102_ (.A(_0465_),
    .B(_0486_),
    .X(_0487_));
 sg13g2_mux2_1 _1103_ (.A0(net161),
    .A1(_0143_),
    .S(_0487_),
    .X(_0091_));
 sg13g2_mux2_1 _1104_ (.A0(net175),
    .A1(_0145_),
    .S(_0487_),
    .X(_0092_));
 sg13g2_mux2_1 _1105_ (.A0(net169),
    .A1(_0147_),
    .S(_0487_),
    .X(_0093_));
 sg13g2_mux2_1 _1106_ (.A0(net143),
    .A1(_0148_),
    .S(_0487_),
    .X(_0094_));
 sg13g2_mux2_1 _1107_ (.A0(net183),
    .A1(_0150_),
    .S(_0487_),
    .X(_0095_));
 sg13g2_mux2_1 _1108_ (.A0(net174),
    .A1(_0151_),
    .S(_0487_),
    .X(_0096_));
 sg13g2_mux2_1 _1109_ (.A0(net173),
    .A1(_0153_),
    .S(_0487_),
    .X(_0097_));
 sg13g2_mux2_1 _1110_ (.A0(net177),
    .A1(_0154_),
    .S(_0487_),
    .X(_0098_));
 sg13g2_nand3b_1 _1111_ (.B(net4),
    .C(net3),
    .Y(_0488_),
    .A_N(net2));
 sg13g2_o21ai_1 _1112_ (.B1(_0135_),
    .Y(_0489_),
    .A1(_0117_),
    .A2(net110));
 sg13g2_a21oi_2 _1113_ (.B1(_0489_),
    .Y(_0490_),
    .A2(_0488_),
    .A1(net130));
 sg13g2_mux2_1 _1114_ (.A0(net155),
    .A1(_0143_),
    .S(_0490_),
    .X(_0099_));
 sg13g2_mux2_1 _1115_ (.A0(net156),
    .A1(_0145_),
    .S(_0490_),
    .X(_0100_));
 sg13g2_mux2_1 _1116_ (.A0(net148),
    .A1(_0147_),
    .S(_0490_),
    .X(_0101_));
 sg13g2_mux2_1 _1117_ (.A0(net170),
    .A1(_0148_),
    .S(_0490_),
    .X(_0102_));
 sg13g2_mux2_1 _1118_ (.A0(net145),
    .A1(_0150_),
    .S(_0490_),
    .X(_0103_));
 sg13g2_mux2_1 _1119_ (.A0(net149),
    .A1(_0151_),
    .S(_0490_),
    .X(_0104_));
 sg13g2_mux2_1 _1120_ (.A0(net150),
    .A1(_0153_),
    .S(_0490_),
    .X(_0105_));
 sg13g2_mux2_1 _1121_ (.A0(net151),
    .A1(_0154_),
    .S(_0490_),
    .X(_0106_));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net137),
    .D(_0016_),
    .Q_N(\state[0] ),
    .Q(_0015_));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net137),
    .D(_0000_),
    .Q_N(_0004_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net137),
    .D(_0001_),
    .Q_N(_0571_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net137),
    .D(net168),
    .Q_N(_0005_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net36),
    .D(_0017_),
    .Q_N(_0570_),
    .Q(\mem[7][0] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net35),
    .D(_0018_),
    .Q_N(_0569_),
    .Q(\mem[7][1] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net34),
    .D(_0019_),
    .Q_N(_0568_),
    .Q(\mem[7][2] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net33),
    .D(_0020_),
    .Q_N(_0567_),
    .Q(\mem[7][3] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net32),
    .D(_0021_),
    .Q_N(_0566_),
    .Q(\mem[7][4] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net31),
    .D(_0022_),
    .Q_N(_0565_),
    .Q(\mem[7][5] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net30),
    .D(_0023_),
    .Q_N(_0564_),
    .Q(\mem[7][6] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net29),
    .D(_0024_),
    .Q_N(_0572_),
    .Q(\mem[7][7] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net138),
    .D(net96),
    .Q_N(_0573_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net138),
    .D(net97),
    .Q_N(_0574_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net135),
    .D(net93),
    .Q_N(_0575_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net139),
    .D(net126),
    .Q_N(_0576_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net135),
    .D(net94),
    .Q_N(_0577_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(net125),
    .Q_N(_0578_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(net95),
    .Q_N(_0579_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net134),
    .D(net100),
    .Q_N(_0563_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net137),
    .D(net141),
    .Q_N(_0562_),
    .Q(\B[0] ));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net138),
    .D(_0026_),
    .Q_N(_0008_),
    .Q(\B[1] ));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net136),
    .D(_0027_),
    .Q_N(_0009_),
    .Q(\B[2] ));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net136),
    .D(_0028_),
    .Q_N(_0010_),
    .Q(\B[3] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net140),
    .D(_0029_),
    .Q_N(_0011_),
    .Q(\B[4] ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net135),
    .D(_0030_),
    .Q_N(_0012_),
    .Q(\B[5] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_0031_),
    .Q_N(_0013_),
    .Q(\B[6] ));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_0032_),
    .Q_N(_0014_),
    .Q(\B[7] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net137),
    .D(_0033_),
    .Q_N(_0561_),
    .Q(\ACC[0] ));
 sg13g2_dfrbp_1 _1151_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net138),
    .D(_0034_),
    .Q_N(_0560_),
    .Q(\ACC[1] ));
 sg13g2_dfrbp_1 _1152_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net136),
    .D(_0035_),
    .Q_N(_0559_),
    .Q(\ACC[2] ));
 sg13g2_dfrbp_1 _1153_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net138),
    .D(_0036_),
    .Q_N(_0558_),
    .Q(\ACC[3] ));
 sg13g2_dfrbp_1 _1154_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net140),
    .D(_0037_),
    .Q_N(_0557_),
    .Q(\ACC[4] ));
 sg13g2_dfrbp_1 _1155_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_0038_),
    .Q_N(_0556_),
    .Q(\ACC[5] ));
 sg13g2_dfrbp_1 _1156_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_0039_),
    .Q_N(_0555_),
    .Q(\ACC[6] ));
 sg13g2_dfrbp_1 _1157_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net134),
    .D(_0040_),
    .Q_N(_0554_),
    .Q(\ACC[7] ));
 sg13g2_dfrbp_1 _1158_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net136),
    .D(net99),
    .Q_N(_0006_),
    .Q(\PC[0] ));
 sg13g2_dfrbp_1 _1159_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(_0042_),
    .Q_N(_0553_),
    .Q(\PC[1] ));
 sg13g2_dfrbp_1 _1160_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net135),
    .D(_0043_),
    .Q_N(_0007_),
    .Q(\PC[2] ));
 sg13g2_dfrbp_1 _1161_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net137),
    .D(_0044_),
    .Q_N(_0552_),
    .Q(\IR[0] ));
 sg13g2_dfrbp_1 _1162_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net136),
    .D(_0045_),
    .Q_N(_0551_),
    .Q(\IR[1] ));
 sg13g2_dfrbp_1 _1163_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net136),
    .D(_0046_),
    .Q_N(_0003_),
    .Q(\IR[2] ));
 sg13g2_dfrbp_1 _1164_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net136),
    .D(net205),
    .Q_N(_0550_),
    .Q(\IR[4] ));
 sg13g2_dfrbp_1 _1165_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net136),
    .D(net225),
    .Q_N(_0549_),
    .Q(\IR[5] ));
 sg13g2_dfrbp_1 _1166_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(_0049_),
    .Q_N(_0548_),
    .Q(\IR[6] ));
 sg13g2_dfrbp_1 _1167_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net135),
    .D(_0050_),
    .Q_N(_0547_),
    .Q(\IR[7] ));
 sg13g2_dfrbp_1 _1168_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net92),
    .D(_0051_),
    .Q_N(_0546_),
    .Q(\mem[0][0] ));
 sg13g2_dfrbp_1 _1169_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net91),
    .D(_0052_),
    .Q_N(_0545_),
    .Q(\mem[0][1] ));
 sg13g2_dfrbp_1 _1170_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net90),
    .D(_0053_),
    .Q_N(_0544_),
    .Q(\mem[0][2] ));
 sg13g2_dfrbp_1 _1171_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net89),
    .D(_0054_),
    .Q_N(_0543_),
    .Q(\mem[0][3] ));
 sg13g2_dfrbp_1 _1172_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net88),
    .D(_0055_),
    .Q_N(_0542_),
    .Q(\mem[0][4] ));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net87),
    .D(_0056_),
    .Q_N(_0541_),
    .Q(\mem[0][5] ));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net86),
    .D(_0057_),
    .Q_N(_0540_),
    .Q(\mem[0][6] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net85),
    .D(_0058_),
    .Q_N(_0539_),
    .Q(\mem[0][7] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net84),
    .D(_0059_),
    .Q_N(_0538_),
    .Q(\mem[1][0] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net83),
    .D(_0060_),
    .Q_N(_0537_),
    .Q(\mem[1][1] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(_0061_),
    .Q_N(_0536_),
    .Q(\mem[1][2] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net81),
    .D(_0062_),
    .Q_N(_0535_),
    .Q(\mem[1][3] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net80),
    .D(_0063_),
    .Q_N(_0534_),
    .Q(\mem[1][4] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net79),
    .D(_0064_),
    .Q_N(_0533_),
    .Q(\mem[1][5] ));
 sg13g2_dfrbp_1 _1182_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net78),
    .D(_0065_),
    .Q_N(_0532_),
    .Q(\mem[1][6] ));
 sg13g2_dfrbp_1 _1183_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net77),
    .D(_0066_),
    .Q_N(_0531_),
    .Q(\mem[1][7] ));
 sg13g2_dfrbp_1 _1184_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net76),
    .D(_0067_),
    .Q_N(_0530_),
    .Q(\mem[2][0] ));
 sg13g2_dfrbp_1 _1185_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net75),
    .D(_0068_),
    .Q_N(_0529_),
    .Q(\mem[2][1] ));
 sg13g2_dfrbp_1 _1186_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net74),
    .D(_0069_),
    .Q_N(_0528_),
    .Q(\mem[2][2] ));
 sg13g2_dfrbp_1 _1187_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net73),
    .D(_0070_),
    .Q_N(_0527_),
    .Q(\mem[2][3] ));
 sg13g2_dfrbp_1 _1188_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net72),
    .D(_0071_),
    .Q_N(_0526_),
    .Q(\mem[2][4] ));
 sg13g2_dfrbp_1 _1189_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net71),
    .D(_0072_),
    .Q_N(_0525_),
    .Q(\mem[2][5] ));
 sg13g2_dfrbp_1 _1190_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net70),
    .D(_0073_),
    .Q_N(_0524_),
    .Q(\mem[2][6] ));
 sg13g2_dfrbp_1 _1191_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net69),
    .D(_0074_),
    .Q_N(_0523_),
    .Q(\mem[2][7] ));
 sg13g2_dfrbp_1 _1192_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net68),
    .D(_0075_),
    .Q_N(_0522_),
    .Q(\mem[3][0] ));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net67),
    .D(_0076_),
    .Q_N(_0521_),
    .Q(\mem[3][1] ));
 sg13g2_dfrbp_1 _1194_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net66),
    .D(_0077_),
    .Q_N(_0520_),
    .Q(\mem[3][2] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net65),
    .D(_0078_),
    .Q_N(_0519_),
    .Q(\mem[3][3] ));
 sg13g2_dfrbp_1 _1196_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net64),
    .D(_0079_),
    .Q_N(_0518_),
    .Q(\mem[3][4] ));
 sg13g2_dfrbp_1 _1197_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net63),
    .D(_0080_),
    .Q_N(_0517_),
    .Q(\mem[3][5] ));
 sg13g2_dfrbp_1 _1198_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net62),
    .D(_0081_),
    .Q_N(_0516_),
    .Q(\mem[3][6] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net61),
    .D(_0082_),
    .Q_N(_0515_),
    .Q(\mem[3][7] ));
 sg13g2_dfrbp_1 _1200_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net60),
    .D(_0083_),
    .Q_N(_0514_),
    .Q(\mem[4][0] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net59),
    .D(_0084_),
    .Q_N(_0513_),
    .Q(\mem[4][1] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net58),
    .D(_0085_),
    .Q_N(_0512_),
    .Q(\mem[4][2] ));
 sg13g2_dfrbp_1 _1203_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net57),
    .D(_0086_),
    .Q_N(_0511_),
    .Q(\mem[4][3] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net56),
    .D(_0087_),
    .Q_N(_0510_),
    .Q(\mem[4][4] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net55),
    .D(_0088_),
    .Q_N(_0509_),
    .Q(\mem[4][5] ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net54),
    .D(_0089_),
    .Q_N(_0508_),
    .Q(\mem[4][6] ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net53),
    .D(_0090_),
    .Q_N(_0507_),
    .Q(\mem[4][7] ));
 sg13g2_dfrbp_1 _1208_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net52),
    .D(_0091_),
    .Q_N(_0506_),
    .Q(\mem[5][0] ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net51),
    .D(_0092_),
    .Q_N(_0505_),
    .Q(\mem[5][1] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net50),
    .D(_0093_),
    .Q_N(_0504_),
    .Q(\mem[5][2] ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net49),
    .D(_0094_),
    .Q_N(_0503_),
    .Q(\mem[5][3] ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net48),
    .D(_0095_),
    .Q_N(_0502_),
    .Q(\mem[5][4] ));
 sg13g2_dfrbp_1 _1213_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net47),
    .D(_0096_),
    .Q_N(_0501_),
    .Q(\mem[5][5] ));
 sg13g2_dfrbp_1 _1214_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net46),
    .D(_0097_),
    .Q_N(_0500_),
    .Q(\mem[5][6] ));
 sg13g2_dfrbp_1 _1215_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net45),
    .D(_0098_),
    .Q_N(_0499_),
    .Q(\mem[5][7] ));
 sg13g2_dfrbp_1 _1216_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net44),
    .D(_0099_),
    .Q_N(_0498_),
    .Q(\mem[6][0] ));
 sg13g2_dfrbp_1 _1217_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net43),
    .D(_0100_),
    .Q_N(_0497_),
    .Q(\mem[6][1] ));
 sg13g2_dfrbp_1 _1218_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net42),
    .D(_0101_),
    .Q_N(_0496_),
    .Q(\mem[6][2] ));
 sg13g2_dfrbp_1 _1219_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net41),
    .D(_0102_),
    .Q_N(_0495_),
    .Q(\mem[6][3] ));
 sg13g2_dfrbp_1 _1220_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net40),
    .D(_0103_),
    .Q_N(_0494_),
    .Q(\mem[6][4] ));
 sg13g2_dfrbp_1 _1221_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net39),
    .D(_0104_),
    .Q_N(_0493_),
    .Q(\mem[6][5] ));
 sg13g2_dfrbp_1 _1222_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net38),
    .D(_0105_),
    .Q_N(_0492_),
    .Q(\mem[6][6] ));
 sg13g2_dfrbp_1 _1223_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net37),
    .D(_0106_),
    .Q_N(_0491_),
    .Q(\mem[6][7] ));
 sg13g2_tiehi _1132__30 (.L_HI(net30));
 sg13g2_tiehi _1131__31 (.L_HI(net31));
 sg13g2_tiehi _1130__32 (.L_HI(net32));
 sg13g2_tiehi _1129__33 (.L_HI(net33));
 sg13g2_tiehi _1128__34 (.L_HI(net34));
 sg13g2_tiehi _1127__35 (.L_HI(net35));
 sg13g2_tiehi _1126__36 (.L_HI(net36));
 sg13g2_tiehi _1223__37 (.L_HI(net37));
 sg13g2_tiehi _1222__38 (.L_HI(net38));
 sg13g2_tiehi _1221__39 (.L_HI(net39));
 sg13g2_tiehi _1220__40 (.L_HI(net40));
 sg13g2_tiehi _1219__41 (.L_HI(net41));
 sg13g2_tiehi _1218__42 (.L_HI(net42));
 sg13g2_tiehi _1217__43 (.L_HI(net43));
 sg13g2_tiehi _1216__44 (.L_HI(net44));
 sg13g2_tiehi _1215__45 (.L_HI(net45));
 sg13g2_tiehi _1214__46 (.L_HI(net46));
 sg13g2_tiehi _1213__47 (.L_HI(net47));
 sg13g2_tiehi _1212__48 (.L_HI(net48));
 sg13g2_tiehi _1211__49 (.L_HI(net49));
 sg13g2_tiehi _1210__50 (.L_HI(net50));
 sg13g2_tiehi _1209__51 (.L_HI(net51));
 sg13g2_tiehi _1208__52 (.L_HI(net52));
 sg13g2_tiehi _1207__53 (.L_HI(net53));
 sg13g2_tiehi _1206__54 (.L_HI(net54));
 sg13g2_tiehi _1205__55 (.L_HI(net55));
 sg13g2_tiehi _1204__56 (.L_HI(net56));
 sg13g2_tiehi _1203__57 (.L_HI(net57));
 sg13g2_tiehi _1202__58 (.L_HI(net58));
 sg13g2_tiehi _1201__59 (.L_HI(net59));
 sg13g2_tiehi _1200__60 (.L_HI(net60));
 sg13g2_tiehi _1199__61 (.L_HI(net61));
 sg13g2_tiehi _1198__62 (.L_HI(net62));
 sg13g2_tiehi _1197__63 (.L_HI(net63));
 sg13g2_tiehi _1196__64 (.L_HI(net64));
 sg13g2_tiehi _1195__65 (.L_HI(net65));
 sg13g2_tiehi _1194__66 (.L_HI(net66));
 sg13g2_tiehi _1193__67 (.L_HI(net67));
 sg13g2_tiehi _1192__68 (.L_HI(net68));
 sg13g2_tiehi _1191__69 (.L_HI(net69));
 sg13g2_tiehi _1190__70 (.L_HI(net70));
 sg13g2_tiehi _1189__71 (.L_HI(net71));
 sg13g2_tiehi _1188__72 (.L_HI(net72));
 sg13g2_tiehi _1187__73 (.L_HI(net73));
 sg13g2_tiehi _1186__74 (.L_HI(net74));
 sg13g2_tiehi _1185__75 (.L_HI(net75));
 sg13g2_tiehi _1184__76 (.L_HI(net76));
 sg13g2_tiehi _1183__77 (.L_HI(net77));
 sg13g2_tiehi _1182__78 (.L_HI(net78));
 sg13g2_tiehi _1181__79 (.L_HI(net79));
 sg13g2_tiehi _1180__80 (.L_HI(net80));
 sg13g2_tiehi _1179__81 (.L_HI(net81));
 sg13g2_tiehi _1178__82 (.L_HI(net82));
 sg13g2_tiehi _1177__83 (.L_HI(net83));
 sg13g2_tiehi _1176__84 (.L_HI(net84));
 sg13g2_tiehi _1175__85 (.L_HI(net85));
 sg13g2_tiehi _1174__86 (.L_HI(net86));
 sg13g2_tiehi _1173__87 (.L_HI(net87));
 sg13g2_tiehi _1172__88 (.L_HI(net88));
 sg13g2_tiehi _1171__89 (.L_HI(net89));
 sg13g2_tiehi _1170__90 (.L_HI(net90));
 sg13g2_tiehi _1169__91 (.L_HI(net91));
 sg13g2_tiehi _1168__92 (.L_HI(net92));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_ultra_tiny_cpu_14 (.L_LO(net14));
 sg13g2_tielo tt_um_ultra_tiny_cpu_15 (.L_LO(net15));
 sg13g2_tielo tt_um_ultra_tiny_cpu_16 (.L_LO(net16));
 sg13g2_tielo tt_um_ultra_tiny_cpu_17 (.L_LO(net17));
 sg13g2_tielo tt_um_ultra_tiny_cpu_18 (.L_LO(net18));
 sg13g2_tielo tt_um_ultra_tiny_cpu_19 (.L_LO(net19));
 sg13g2_tielo tt_um_ultra_tiny_cpu_20 (.L_LO(net20));
 sg13g2_tielo tt_um_ultra_tiny_cpu_21 (.L_LO(net21));
 sg13g2_tielo tt_um_ultra_tiny_cpu_22 (.L_LO(net22));
 sg13g2_tielo tt_um_ultra_tiny_cpu_23 (.L_LO(net23));
 sg13g2_tielo tt_um_ultra_tiny_cpu_24 (.L_LO(net24));
 sg13g2_tielo tt_um_ultra_tiny_cpu_25 (.L_LO(net25));
 sg13g2_tielo tt_um_ultra_tiny_cpu_26 (.L_LO(net26));
 sg13g2_tielo tt_um_ultra_tiny_cpu_27 (.L_LO(net27));
 sg13g2_tielo tt_um_ultra_tiny_cpu_28 (.L_LO(net28));
 sg13g2_tiehi _1133__29 (.L_HI(net29));
 sg13g2_buf_2 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0241_),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_0236_));
 sg13g2_buf_1 fanout107 (.A(_0236_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0156_),
    .X(net109));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_0257_));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_0253_));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(_0252_));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(_0246_));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(_0243_));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(_0235_));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_0137_));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(_0164_));
 sg13g2_buf_2 fanout118 (.A(net120),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0130_),
    .X(net120));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(_0107_));
 sg13g2_buf_2 fanout122 (.A(_0107_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(\PC[1] ),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(\PC[0] ),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(net219),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net220),
    .X(net126));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(net128));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(net214));
 sg13g2_buf_2 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(ui_in[7]),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(ui_in[7]),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net135));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net140));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net139));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net139));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(rst_n),
    .X(net140));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[0]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[3]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[4]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[5]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[6]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[7]),
    .X(net12));
 sg13g2_tielo tt_um_ultra_tiny_cpu_13 (.L_LO(net13));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ACC[2] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ACC[4] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ACC[6] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold4 (.A(\ACC[0] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ACC[1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold6 (.A(\PC[0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0041_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold8 (.A(\ACC[7] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold9 (.A(\PC[1] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0005_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0157_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0025_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mem[1][5] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mem[5][3] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mem[1][7] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mem[6][4] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mem[2][5] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold18 (.A(\state[0] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mem[6][2] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mem[6][5] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mem[6][6] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mem[6][7] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mem[1][1] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mem[1][6] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mem[1][0] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mem[6][0] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mem[6][1] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mem[2][1] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mem[2][3] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mem[2][7] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mem[1][4] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mem[5][0] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mem[1][3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mem[1][2] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mem[2][6] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mem[7][2] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mem[2][2] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold38 (.A(\state[2] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0002_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mem[5][2] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mem[6][3] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mem[2][4] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mem[2][0] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mem[5][6] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mem[5][5] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mem[5][1] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold47 (.A(\B[7] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mem[5][7] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mem[3][4] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mem[3][5] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mem[3][7] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mem[7][6] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mem[3][2] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mem[5][4] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mem[3][0] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mem[7][1] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mem[3][3] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mem[3][1] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mem[4][7] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mem[7][4] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mem[7][5] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mem[7][3] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mem[3][6] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mem[0][4] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mem[4][5] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mem[7][7] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mem[0][1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mem[7][0] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mem[0][2] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mem[0][3] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mem[0][6] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mem[4][4] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mem[4][6] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mem[4][3] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold75 (.A(\IR[4] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0047_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mem[4][0] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold78 (.A(\B[5] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mem[0][5] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mem[4][1] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold81 (.A(\IR[7] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold82 (.A(\IR[6] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mem[0][0] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mem[4][2] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold85 (.A(\state[1] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold86 (.A(\B[6] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold87 (.A(\B[3] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold88 (.A(\state[3] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mem[0][7] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold90 (.A(\ACC[5] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ACC[3] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold92 (.A(\B[4] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold93 (.A(\IR[1] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold94 (.A(\B[2] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold95 (.A(\IR[5] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0048_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold97 (.A(\IR[2] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold98 (.A(\IR[0] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold99 (.A(\B[1] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold100 (.A(\PC[2] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold101 (.A(\IR[1] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mem[0][7] ),
    .X(net231));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_173 ();
 sg13g2_fill_2 FILLER_11_187 ();
 sg13g2_decap_4 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_213 ();
 sg13g2_decap_8 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_227 ();
 sg13g2_decap_4 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_fill_2 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_327 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_161 ();
 sg13g2_fill_2 FILLER_12_215 ();
 sg13g2_fill_1 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_4 FILLER_13_140 ();
 sg13g2_fill_2 FILLER_13_177 ();
 sg13g2_fill_1 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_208 ();
 sg13g2_fill_1 FILLER_13_215 ();
 sg13g2_fill_2 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_228 ();
 sg13g2_fill_1 FILLER_13_257 ();
 sg13g2_fill_2 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_decap_4 FILLER_13_313 ();
 sg13g2_fill_1 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_fill_2 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_decap_4 FILLER_14_124 ();
 sg13g2_fill_2 FILLER_14_128 ();
 sg13g2_fill_1 FILLER_14_143 ();
 sg13g2_fill_2 FILLER_14_170 ();
 sg13g2_fill_2 FILLER_14_198 ();
 sg13g2_fill_1 FILLER_14_200 ();
 sg13g2_fill_1 FILLER_14_227 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_2 FILLER_14_312 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_fill_2 FILLER_14_325 ();
 sg13g2_fill_1 FILLER_14_327 ();
 sg13g2_fill_1 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_fill_1 FILLER_15_109 ();
 sg13g2_fill_2 FILLER_15_146 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_fill_1 FILLER_15_164 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_1 FILLER_15_177 ();
 sg13g2_fill_2 FILLER_15_191 ();
 sg13g2_decap_4 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_decap_4 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_328 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_fill_1 FILLER_15_354 ();
 sg13g2_fill_2 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_93 ();
 sg13g2_decap_8 FILLER_16_120 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_decap_4 FILLER_16_164 ();
 sg13g2_decap_8 FILLER_16_225 ();
 sg13g2_fill_2 FILLER_16_232 ();
 sg13g2_fill_2 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_decap_4 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_335 ();
 sg13g2_fill_2 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_4 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_decap_4 FILLER_17_100 ();
 sg13g2_decap_4 FILLER_17_144 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_decap_4 FILLER_17_153 ();
 sg13g2_fill_2 FILLER_17_157 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_4 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_decap_4 FILLER_17_208 ();
 sg13g2_decap_4 FILLER_17_268 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_decap_4 FILLER_17_331 ();
 sg13g2_fill_1 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_146 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_decap_4 FILLER_18_177 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_decap_4 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_363 ();
 sg13g2_fill_1 FILLER_18_383 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_fill_2 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_2 FILLER_19_196 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_decap_4 FILLER_19_335 ();
 sg13g2_decap_4 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_fill_2 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_185 ();
 sg13g2_decap_4 FILLER_20_192 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_decap_4 FILLER_20_212 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_decap_4 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_4 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_decap_4 FILLER_20_298 ();
 sg13g2_decap_4 FILLER_20_310 ();
 sg13g2_fill_2 FILLER_20_314 ();
 sg13g2_decap_4 FILLER_20_327 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_4 FILLER_21_100 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_fill_2 FILLER_21_115 ();
 sg13g2_fill_2 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_fill_1 FILLER_21_306 ();
 sg13g2_decap_4 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_156 ();
 sg13g2_fill_2 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_decap_4 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_227 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_2 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_4 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_130 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_decap_4 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_178 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_decap_8 FILLER_23_212 ();
 sg13g2_decap_4 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_275 ();
 sg13g2_fill_2 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_362 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_fill_2 FILLER_24_97 ();
 sg13g2_fill_2 FILLER_24_162 ();
 sg13g2_fill_1 FILLER_24_164 ();
 sg13g2_fill_1 FILLER_24_171 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_284 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_310 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_318 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_349 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_decap_4 FILLER_24_367 ();
 sg13g2_fill_2 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_100 ();
 sg13g2_fill_1 FILLER_25_104 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_fill_1 FILLER_25_173 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_4 FILLER_25_295 ();
 sg13g2_decap_4 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_fill_2 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_228 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_348 ();
 sg13g2_fill_2 FILLER_26_370 ();
 sg13g2_fill_1 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_110 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_decap_4 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_decap_4 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_227 ();
 sg13g2_decap_4 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_115 ();
 sg13g2_fill_2 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_decap_4 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_240 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_decap_4 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_4 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_349 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_127 ();
 sg13g2_decap_4 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_205 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_decap_4 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_354 ();
 sg13g2_fill_1 FILLER_29_356 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_4 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_decap_4 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_decap_4 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_fill_1 FILLER_30_342 ();
 sg13g2_decap_4 FILLER_30_348 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_125 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_260 ();
 sg13g2_decap_4 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_315 ();
 sg13g2_fill_1 FILLER_31_368 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_93 ();
 sg13g2_decap_4 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_245 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_decap_4 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_decap_4 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_116 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_decap_4 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_188 ();
 sg13g2_decap_8 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_decap_4 FILLER_33_268 ();
 sg13g2_decap_8 FILLER_33_278 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_fill_2 FILLER_33_315 ();
 sg13g2_fill_2 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_324 ();
 sg13g2_decap_4 FILLER_33_346 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_4 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_109 ();
 sg13g2_fill_2 FILLER_34_137 ();
 sg13g2_fill_2 FILLER_34_153 ();
 sg13g2_decap_4 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_decap_4 FILLER_34_273 ();
 sg13g2_decap_4 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_1 FILLER_34_309 ();
 sg13g2_fill_2 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_331 ();
 sg13g2_decap_8 FILLER_34_337 ();
 sg13g2_fill_2 FILLER_34_344 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_decap_4 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_fill_2 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_186 ();
 sg13g2_fill_2 FILLER_35_212 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_fill_2 FILLER_35_308 ();
 sg13g2_fill_2 FILLER_35_319 ();
 sg13g2_fill_1 FILLER_35_321 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_4 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_232 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_decap_4 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_146 ();
 sg13g2_fill_2 FILLER_37_170 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_205 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_decap_4 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_fill_1 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_4 FILLER_37_323 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_fill_1 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_fill_2 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_fill_2 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_311 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
 assign uio_out[4] = net25;
 assign uio_out[5] = net26;
 assign uio_out[6] = net27;
 assign uio_out[7] = net28;
endmodule

module tt_um_dlmiles_dffram32x8_2r1w (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire clknet_leaf_0_clk;
 wire addrhi;
 wire \mem[100] ;
 wire \mem[101] ;
 wire \mem[102] ;
 wire \mem[103] ;
 wire \mem[104] ;
 wire \mem[105] ;
 wire \mem[106] ;
 wire \mem[107] ;
 wire \mem[108] ;
 wire \mem[109] ;
 wire \mem[110] ;
 wire \mem[111] ;
 wire \mem[112] ;
 wire \mem[113] ;
 wire \mem[114] ;
 wire \mem[115] ;
 wire \mem[116] ;
 wire \mem[117] ;
 wire \mem[118] ;
 wire \mem[119] ;
 wire \mem[120] ;
 wire \mem[121] ;
 wire \mem[122] ;
 wire \mem[123] ;
 wire \mem[124] ;
 wire \mem[125] ;
 wire \mem[126] ;
 wire \mem[127] ;
 wire \mem[128] ;
 wire \mem[129] ;
 wire \mem[130] ;
 wire \mem[131] ;
 wire \mem[132] ;
 wire \mem[133] ;
 wire \mem[134] ;
 wire \mem[135] ;
 wire \mem[136] ;
 wire \mem[137] ;
 wire \mem[138] ;
 wire \mem[139] ;
 wire \mem[140] ;
 wire \mem[141] ;
 wire \mem[142] ;
 wire \mem[143] ;
 wire \mem[144] ;
 wire \mem[145] ;
 wire \mem[146] ;
 wire \mem[147] ;
 wire \mem[148] ;
 wire \mem[149] ;
 wire \mem[150] ;
 wire \mem[151] ;
 wire \mem[152] ;
 wire \mem[153] ;
 wire \mem[154] ;
 wire \mem[155] ;
 wire \mem[156] ;
 wire \mem[157] ;
 wire \mem[158] ;
 wire \mem[159] ;
 wire \mem[160] ;
 wire \mem[161] ;
 wire \mem[162] ;
 wire \mem[163] ;
 wire \mem[164] ;
 wire \mem[165] ;
 wire \mem[166] ;
 wire \mem[167] ;
 wire \mem[168] ;
 wire \mem[169] ;
 wire \mem[170] ;
 wire \mem[171] ;
 wire \mem[172] ;
 wire \mem[173] ;
 wire \mem[174] ;
 wire \mem[175] ;
 wire \mem[176] ;
 wire \mem[177] ;
 wire \mem[178] ;
 wire \mem[179] ;
 wire \mem[180] ;
 wire \mem[181] ;
 wire \mem[182] ;
 wire \mem[183] ;
 wire \mem[184] ;
 wire \mem[185] ;
 wire \mem[186] ;
 wire \mem[187] ;
 wire \mem[188] ;
 wire \mem[189] ;
 wire \mem[190] ;
 wire \mem[191] ;
 wire \mem[192] ;
 wire \mem[193] ;
 wire \mem[194] ;
 wire \mem[195] ;
 wire \mem[196] ;
 wire \mem[197] ;
 wire \mem[198] ;
 wire \mem[199] ;
 wire \mem[200] ;
 wire \mem[201] ;
 wire \mem[202] ;
 wire \mem[203] ;
 wire \mem[204] ;
 wire \mem[205] ;
 wire \mem[206] ;
 wire \mem[207] ;
 wire \mem[208] ;
 wire \mem[209] ;
 wire \mem[210] ;
 wire \mem[211] ;
 wire \mem[212] ;
 wire \mem[213] ;
 wire \mem[214] ;
 wire \mem[215] ;
 wire \mem[216] ;
 wire \mem[217] ;
 wire \mem[218] ;
 wire \mem[219] ;
 wire \mem[220] ;
 wire \mem[221] ;
 wire \mem[222] ;
 wire \mem[223] ;
 wire \mem[224] ;
 wire \mem[225] ;
 wire \mem[226] ;
 wire \mem[227] ;
 wire \mem[228] ;
 wire \mem[229] ;
 wire \mem[230] ;
 wire \mem[231] ;
 wire \mem[232] ;
 wire \mem[233] ;
 wire \mem[234] ;
 wire \mem[235] ;
 wire \mem[236] ;
 wire \mem[237] ;
 wire \mem[238] ;
 wire \mem[239] ;
 wire \mem[240] ;
 wire \mem[241] ;
 wire \mem[242] ;
 wire \mem[243] ;
 wire \mem[244] ;
 wire \mem[245] ;
 wire \mem[246] ;
 wire \mem[247] ;
 wire \mem[248] ;
 wire \mem[249] ;
 wire \mem[250] ;
 wire \mem[251] ;
 wire \mem[252] ;
 wire \mem[253] ;
 wire \mem[254] ;
 wire \mem[255] ;
 wire \mem[64] ;
 wire \mem[65] ;
 wire \mem[66] ;
 wire \mem[67] ;
 wire \mem[68] ;
 wire \mem[69] ;
 wire \mem[70] ;
 wire \mem[71] ;
 wire \mem[72] ;
 wire \mem[73] ;
 wire \mem[74] ;
 wire \mem[75] ;
 wire \mem[76] ;
 wire \mem[77] ;
 wire \mem[78] ;
 wire \mem[79] ;
 wire \mem[80] ;
 wire \mem[81] ;
 wire \mem[82] ;
 wire \mem[83] ;
 wire \mem[84] ;
 wire \mem[85] ;
 wire \mem[86] ;
 wire \mem[87] ;
 wire \mem[88] ;
 wire \mem[89] ;
 wire \mem[90] ;
 wire \mem[91] ;
 wire \mem[92] ;
 wire \mem[93] ;
 wire \mem[94] ;
 wire \mem[95] ;
 wire \mem[96] ;
 wire \mem[97] ;
 wire \mem[98] ;
 wire \mem[99] ;
 wire \rdata_buff_a[0] ;
 wire \rdata_buff_a[1] ;
 wire \rdata_buff_a[2] ;
 wire \rdata_buff_a[3] ;
 wire \rdata_buff_a[4] ;
 wire \rdata_buff_a[5] ;
 wire \rdata_buff_a[6] ;
 wire \rdata_buff_a[7] ;
 wire \rdata_buff_b[0] ;
 wire \rdata_buff_b[1] ;
 wire \rdata_buff_b[2] ;
 wire \rdata_buff_b[3] ;
 wire \rdata_buff_b[4] ;
 wire \rdata_buff_b[5] ;
 wire \rdata_buff_b[6] ;
 wire \rdata_buff_b[7] ;
 wire \rdata_curr_a[0] ;
 wire \rdata_curr_a[1] ;
 wire \rdata_curr_a[2] ;
 wire \rdata_curr_a[3] ;
 wire \rdata_curr_a[4] ;
 wire \rdata_curr_a[5] ;
 wire \rdata_curr_a[6] ;
 wire \rdata_curr_a[7] ;
 wire \rdata_curr_b[0] ;
 wire \rdata_curr_b[1] ;
 wire \rdata_curr_b[2] ;
 wire \rdata_curr_b[3] ;
 wire \rdata_curr_b[4] ;
 wire \rdata_curr_b[5] ;
 wire \rdata_curr_b[6] ;
 wire \rdata_curr_b[7] ;
 wire read_buffer_a;
 wire read_buffer_b;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire write_through;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;

 sg13g2_inv_1 _1264_ (.Y(_0430_),
    .A(net589));
 sg13g2_inv_1 _1265_ (.Y(_0431_),
    .A(net2));
 sg13g2_inv_1 _1266_ (.Y(_0432_),
    .A(net3));
 sg13g2_inv_1 _1267_ (.Y(_0433_),
    .A(\mem[231] ));
 sg13g2_inv_1 _1268_ (.Y(_0434_),
    .A(\mem[199] ));
 sg13g2_inv_1 _1269_ (.Y(_0435_),
    .A(\mem[207] ));
 sg13g2_inv_1 _1270_ (.Y(_0436_),
    .A(net267));
 sg13g2_inv_1 _1271_ (.Y(_0437_),
    .A(net285));
 sg13g2_inv_1 _1272_ (.Y(_0438_),
    .A(\mem[143] ));
 sg13g2_inv_1 _1273_ (.Y(_0439_),
    .A(net264));
 sg13g2_inv_1 _1274_ (.Y(_0440_),
    .A(net257));
 sg13g2_inv_1 _1275_ (.Y(_0441_),
    .A(net306));
 sg13g2_inv_1 _1276_ (.Y(_0442_),
    .A(\mem[230] ));
 sg13g2_inv_1 _1277_ (.Y(_0443_),
    .A(\mem[198] ));
 sg13g2_inv_2 _1278_ (.Y(_0444_),
    .A(\mem[206] ));
 sg13g2_inv_2 _1279_ (.Y(_0445_),
    .A(net315));
 sg13g2_inv_2 _1280_ (.Y(_0446_),
    .A(net294));
 sg13g2_inv_1 _1281_ (.Y(_0447_),
    .A(\mem[142] ));
 sg13g2_inv_1 _1282_ (.Y(_0448_),
    .A(net244));
 sg13g2_inv_1 _1283_ (.Y(_0449_),
    .A(net286));
 sg13g2_inv_1 _1284_ (.Y(_0450_),
    .A(\mem[229] ));
 sg13g2_inv_1 _1285_ (.Y(_0451_),
    .A(\mem[197] ));
 sg13g2_inv_1 _1286_ (.Y(_0452_),
    .A(\mem[205] ));
 sg13g2_inv_2 _1287_ (.Y(_0453_),
    .A(net325));
 sg13g2_inv_2 _1288_ (.Y(_0454_),
    .A(net293));
 sg13g2_inv_1 _1289_ (.Y(_0455_),
    .A(\mem[141] ));
 sg13g2_inv_1 _1290_ (.Y(_0456_),
    .A(net248));
 sg13g2_inv_1 _1291_ (.Y(_0457_),
    .A(net252));
 sg13g2_inv_1 _1292_ (.Y(_0458_),
    .A(\mem[228] ));
 sg13g2_inv_1 _1293_ (.Y(_0459_),
    .A(\mem[196] ));
 sg13g2_inv_1 _1294_ (.Y(_0460_),
    .A(\mem[204] ));
 sg13g2_inv_1 _1295_ (.Y(_0461_),
    .A(net283));
 sg13g2_inv_1 _1296_ (.Y(_0462_),
    .A(net290));
 sg13g2_inv_1 _1297_ (.Y(_0463_),
    .A(\mem[140] ));
 sg13g2_inv_1 _1298_ (.Y(_0464_),
    .A(net266));
 sg13g2_inv_1 _1299_ (.Y(_0465_),
    .A(net259));
 sg13g2_inv_1 _1300_ (.Y(_0466_),
    .A(\mem[227] ));
 sg13g2_inv_1 _1301_ (.Y(_0467_),
    .A(\mem[195] ));
 sg13g2_inv_1 _1302_ (.Y(_0468_),
    .A(\mem[203] ));
 sg13g2_inv_1 _1303_ (.Y(_0469_),
    .A(net353));
 sg13g2_inv_1 _1304_ (.Y(_0470_),
    .A(net270));
 sg13g2_inv_1 _1305_ (.Y(_0471_),
    .A(\mem[139] ));
 sg13g2_inv_1 _1306_ (.Y(_0472_),
    .A(net268));
 sg13g2_inv_1 _1307_ (.Y(_0473_),
    .A(net277));
 sg13g2_inv_1 _1308_ (.Y(_0474_),
    .A(\mem[226] ));
 sg13g2_inv_1 _1309_ (.Y(_0475_),
    .A(\mem[194] ));
 sg13g2_inv_1 _1310_ (.Y(_0476_),
    .A(\mem[202] ));
 sg13g2_inv_1 _1311_ (.Y(_0477_),
    .A(net253));
 sg13g2_inv_1 _1312_ (.Y(_0478_),
    .A(net282));
 sg13g2_inv_1 _1313_ (.Y(_0479_),
    .A(\mem[138] ));
 sg13g2_inv_1 _1314_ (.Y(_0480_),
    .A(net272));
 sg13g2_inv_1 _1315_ (.Y(_0481_),
    .A(net260));
 sg13g2_inv_1 _1316_ (.Y(_0482_),
    .A(\mem[225] ));
 sg13g2_inv_1 _1317_ (.Y(_0483_),
    .A(\mem[193] ));
 sg13g2_inv_1 _1318_ (.Y(_0484_),
    .A(\mem[201] ));
 sg13g2_inv_1 _1319_ (.Y(_0485_),
    .A(net317));
 sg13g2_inv_1 _1320_ (.Y(_0486_),
    .A(net298));
 sg13g2_inv_1 _1321_ (.Y(_0487_),
    .A(\mem[137] ));
 sg13g2_inv_1 _1322_ (.Y(_0488_),
    .A(net249));
 sg13g2_inv_1 _1323_ (.Y(_0489_),
    .A(net284));
 sg13g2_inv_1 _1324_ (.Y(_0490_),
    .A(\mem[224] ));
 sg13g2_inv_1 _1325_ (.Y(_0491_),
    .A(\mem[192] ));
 sg13g2_inv_1 _1326_ (.Y(_0492_),
    .A(\mem[200] ));
 sg13g2_inv_1 _1327_ (.Y(_0493_),
    .A(net364));
 sg13g2_inv_1 _1328_ (.Y(_0494_),
    .A(net305));
 sg13g2_inv_1 _1329_ (.Y(_0495_),
    .A(\mem[136] ));
 sg13g2_inv_1 _1330_ (.Y(_0496_),
    .A(net261));
 sg13g2_inv_1 _1331_ (.Y(_0497_),
    .A(net275));
 sg13g2_inv_2 _1332_ (.Y(_0498_),
    .A(read_buffer_a));
 sg13g2_inv_1 _1333_ (.Y(_0499_),
    .A(\rdata_buff_a[4] ));
 sg13g2_inv_1 _1334_ (.Y(_0500_),
    .A(\rdata_buff_a[5] ));
 sg13g2_inv_1 _1335_ (.Y(_0501_),
    .A(\rdata_buff_a[6] ));
 sg13g2_inv_1 _1336_ (.Y(_0502_),
    .A(\rdata_buff_a[7] ));
 sg13g2_inv_1 _1337_ (.Y(_0503_),
    .A(net580));
 sg13g2_and2_1 _1338_ (.A(net4),
    .B(net566),
    .X(_0504_));
 sg13g2_nand2_1 _1339_ (.Y(_0505_),
    .A(net585),
    .B(net567));
 sg13g2_nor2b_2 _1340_ (.A(net585),
    .B_N(net567),
    .Y(_0506_));
 sg13g2_nand2_1 _1341_ (.Y(_0507_),
    .A(net567),
    .B(net557));
 sg13g2_nor2_2 _1342_ (.A(net576),
    .B(net564),
    .Y(_0508_));
 sg13g2_nand2_1 _1343_ (.Y(_0509_),
    .A(net588),
    .B(net554));
 sg13g2_nor3_1 _1344_ (.A(_0431_),
    .B(net3),
    .C(net561),
    .Y(_0510_));
 sg13g2_nand3_1 _1345_ (.B(_0432_),
    .C(net555),
    .A(net2),
    .Y(_0511_));
 sg13g2_nor3_1 _1346_ (.A(_0431_),
    .B(_0432_),
    .C(net561),
    .Y(_0512_));
 sg13g2_nand3_1 _1347_ (.B(net3),
    .C(net556),
    .A(net2),
    .Y(_0513_));
 sg13g2_o21ai_1 _1348_ (.B1(net555),
    .Y(_0514_),
    .A1(net2),
    .A2(net3));
 sg13g2_a21oi_2 _1349_ (.B1(net561),
    .Y(_0515_),
    .A2(_0432_),
    .A1(_0431_));
 sg13g2_a21oi_1 _1350_ (.A1(_0439_),
    .A2(net539),
    .Y(_0516_),
    .B1(net515));
 sg13g2_o21ai_1 _1351_ (.B1(_0516_),
    .Y(_0517_),
    .A1(\mem[119] ),
    .A2(net539));
 sg13g2_a21oi_1 _1352_ (.A1(net590),
    .A2(net557),
    .Y(_0518_),
    .B1(\mem[95] ));
 sg13g2_nor3_1 _1353_ (.A(net2),
    .B(_0432_),
    .C(net561),
    .Y(_0519_));
 sg13g2_nand3_1 _1354_ (.B(net3),
    .C(net554),
    .A(_0431_),
    .Y(_0520_));
 sg13g2_nor3_1 _1355_ (.A(net576),
    .B(\mem[87] ),
    .C(net564),
    .Y(_0521_));
 sg13g2_nor3_1 _1356_ (.A(_0518_),
    .B(_0520_),
    .C(_0521_),
    .Y(_0522_));
 sg13g2_mux2_1 _1357_ (.A0(\mem[103] ),
    .A1(\mem[111] ),
    .S(net539),
    .X(_0523_));
 sg13g2_mux2_1 _1358_ (.A0(\mem[71] ),
    .A1(\mem[79] ),
    .S(net539),
    .X(_0524_));
 sg13g2_a221oi_1 _1359_ (.B2(net524),
    .C1(_0522_),
    .B1(_0524_),
    .A1(net529),
    .Y(_0525_),
    .A2(_0523_));
 sg13g2_a21oi_1 _1360_ (.A1(_0517_),
    .A2(_0525_),
    .Y(_0526_),
    .B1(net544));
 sg13g2_nor2b_1 _1361_ (.A(net567),
    .B_N(net585),
    .Y(_0527_));
 sg13g2_nand2_2 _1362_ (.Y(_0528_),
    .A(net585),
    .B(net553));
 sg13g2_nor2_1 _1363_ (.A(_0506_),
    .B(_0527_),
    .Y(_0529_));
 sg13g2_nand2_2 _1364_ (.Y(_0530_),
    .A(net543),
    .B(_0528_));
 sg13g2_mux2_2 _1365_ (.A0(\mem[231] ),
    .A1(\mem[239] ),
    .S(net531),
    .X(_0531_));
 sg13g2_mux2_1 _1366_ (.A0(\mem[247] ),
    .A1(\mem[255] ),
    .S(net537),
    .X(_0532_));
 sg13g2_a22oi_1 _1367_ (.Y(_0533_),
    .B1(_0532_),
    .B2(net517),
    .A2(_0531_),
    .A1(net525));
 sg13g2_mux2_1 _1368_ (.A0(\mem[215] ),
    .A1(\mem[223] ),
    .S(net533),
    .X(_0534_));
 sg13g2_mux2_1 _1369_ (.A0(\mem[199] ),
    .A1(\mem[207] ),
    .S(net531),
    .X(_0535_));
 sg13g2_a22oi_1 _1370_ (.Y(_0536_),
    .B1(_0535_),
    .B2(net521),
    .A2(_0534_),
    .A1(net511));
 sg13g2_a21oi_2 _1371_ (.B1(_0530_),
    .Y(_0537_),
    .A2(_0536_),
    .A1(_0533_));
 sg13g2_mux2_1 _1372_ (.A0(\mem[135] ),
    .A1(\mem[143] ),
    .S(net534),
    .X(_0538_));
 sg13g2_mux2_1 _1373_ (.A0(\mem[151] ),
    .A1(\mem[159] ),
    .S(net534),
    .X(_0539_));
 sg13g2_a22oi_1 _1374_ (.Y(_0540_),
    .B1(_0539_),
    .B2(net512),
    .A2(_0538_),
    .A1(net522));
 sg13g2_mux2_2 _1375_ (.A0(\mem[167] ),
    .A1(\mem[175] ),
    .S(net534),
    .X(_0541_));
 sg13g2_mux2_2 _1376_ (.A0(\mem[183] ),
    .A1(\mem[191] ),
    .S(net541),
    .X(_0542_));
 sg13g2_a22oi_1 _1377_ (.Y(_0543_),
    .B1(_0542_),
    .B2(net518),
    .A2(_0541_),
    .A1(net526));
 sg13g2_a21oi_2 _1378_ (.B1(_0528_),
    .Y(_0544_),
    .A2(_0543_),
    .A1(_0540_));
 sg13g2_or3_1 _1379_ (.A(_0526_),
    .B(_0537_),
    .C(_0544_),
    .X(\rdata_curr_a[0] ));
 sg13g2_nand3_1 _1380_ (.B(_0442_),
    .C(net552),
    .A(net586),
    .Y(_0545_));
 sg13g2_a21oi_1 _1381_ (.A1(net586),
    .A2(net552),
    .Y(_0546_),
    .B1(\mem[238] ));
 sg13g2_nand3b_1 _1382_ (.B(net525),
    .C(_0545_),
    .Y(_0547_),
    .A_N(_0546_));
 sg13g2_nand3_1 _1383_ (.B(_0443_),
    .C(net552),
    .A(net586),
    .Y(_0548_));
 sg13g2_o21ai_1 _1384_ (.B1(_0444_),
    .Y(_0549_),
    .A1(net572),
    .A2(net559));
 sg13g2_nand3_1 _1385_ (.B(_0548_),
    .C(_0549_),
    .A(net521),
    .Y(_0550_));
 sg13g2_a21oi_1 _1386_ (.A1(net590),
    .A2(net557),
    .Y(_0551_),
    .B1(\mem[254] ));
 sg13g2_nor3_1 _1387_ (.A(net576),
    .B(\mem[246] ),
    .C(net564),
    .Y(_0552_));
 sg13g2_or3_2 _1388_ (.A(net515),
    .B(_0551_),
    .C(_0552_),
    .X(_0553_));
 sg13g2_nor3_1 _1389_ (.A(net573),
    .B(\mem[214] ),
    .C(net560),
    .Y(_0554_));
 sg13g2_a21oi_1 _1390_ (.A1(net587),
    .A2(net553),
    .Y(_0555_),
    .B1(\mem[222] ));
 sg13g2_or3_1 _1391_ (.A(net510),
    .B(_0554_),
    .C(_0555_),
    .X(_0556_));
 sg13g2_nand4_1 _1392_ (.B(_0550_),
    .C(_0553_),
    .A(_0547_),
    .Y(_0557_),
    .D(_0556_));
 sg13g2_mux2_1 _1393_ (.A0(\mem[102] ),
    .A1(\mem[110] ),
    .S(net538),
    .X(_0558_));
 sg13g2_mux2_1 _1394_ (.A0(\mem[70] ),
    .A1(\mem[78] ),
    .S(net538),
    .X(_0559_));
 sg13g2_a22oi_1 _1395_ (.Y(_0560_),
    .B1(_0559_),
    .B2(net524),
    .A2(_0558_),
    .A1(net529));
 sg13g2_mux2_1 _1396_ (.A0(\mem[118] ),
    .A1(\mem[126] ),
    .S(net538),
    .X(_0561_));
 sg13g2_mux2_1 _1397_ (.A0(\mem[86] ),
    .A1(\mem[94] ),
    .S(net538),
    .X(_0562_));
 sg13g2_a22oi_1 _1398_ (.Y(_0563_),
    .B1(_0562_),
    .B2(net513),
    .A2(_0561_),
    .A1(net517));
 sg13g2_a21o_1 _1399_ (.A2(_0563_),
    .A1(_0560_),
    .B1(net544),
    .X(_0564_));
 sg13g2_nor3_1 _1400_ (.A(net576),
    .B(\mem[182] ),
    .C(net564),
    .Y(_0565_));
 sg13g2_a21oi_1 _1401_ (.A1(net590),
    .A2(net557),
    .Y(_0566_),
    .B1(\mem[190] ));
 sg13g2_or3_2 _1402_ (.A(_0515_),
    .B(_0565_),
    .C(_0566_),
    .X(_0567_));
 sg13g2_nor3_1 _1403_ (.A(net573),
    .B(\mem[150] ),
    .C(net560),
    .Y(_0568_));
 sg13g2_a21oi_1 _1404_ (.A1(net587),
    .A2(net553),
    .Y(_0569_),
    .B1(\mem[158] ));
 sg13g2_or3_1 _1405_ (.A(net510),
    .B(_0568_),
    .C(_0569_),
    .X(_0570_));
 sg13g2_nand3_1 _1406_ (.B(_0445_),
    .C(net553),
    .A(net587),
    .Y(_0571_));
 sg13g2_o21ai_1 _1407_ (.B1(_0446_),
    .Y(_0572_),
    .A1(net572),
    .A2(net559));
 sg13g2_nand3_1 _1408_ (.B(_0571_),
    .C(_0572_),
    .A(net526),
    .Y(_0573_));
 sg13g2_o21ai_1 _1409_ (.B1(_0447_),
    .Y(_0574_),
    .A1(net572),
    .A2(net559));
 sg13g2_nor3_1 _1410_ (.A(net572),
    .B(\mem[134] ),
    .C(net559),
    .Y(_0575_));
 sg13g2_nand3b_1 _1411_ (.B(net522),
    .C(_0574_),
    .Y(_0576_),
    .A_N(_0575_));
 sg13g2_nand4_1 _1412_ (.B(_0570_),
    .C(_0573_),
    .A(_0567_),
    .Y(_0577_),
    .D(_0576_));
 sg13g2_a22oi_1 _1413_ (.Y(_0578_),
    .B1(_0577_),
    .B2(net551),
    .A2(_0557_),
    .A1(net508));
 sg13g2_nand2_1 _1414_ (.Y(\rdata_curr_a[1] ),
    .A(_0564_),
    .B(_0578_));
 sg13g2_nor3_1 _1415_ (.A(net572),
    .B(\mem[133] ),
    .C(net559),
    .Y(_0579_));
 sg13g2_a21oi_1 _1416_ (.A1(net586),
    .A2(net552),
    .Y(_0580_),
    .B1(\mem[141] ));
 sg13g2_or3_1 _1417_ (.A(_0513_),
    .B(_0579_),
    .C(_0580_),
    .X(_0581_));
 sg13g2_a21oi_1 _1418_ (.A1(net587),
    .A2(net553),
    .Y(_0582_),
    .B1(\mem[157] ));
 sg13g2_nor3_1 _1419_ (.A(net573),
    .B(\mem[149] ),
    .C(net560),
    .Y(_0583_));
 sg13g2_or3_1 _1420_ (.A(net510),
    .B(_0582_),
    .C(_0583_),
    .X(_0584_));
 sg13g2_nand3_1 _1421_ (.B(_0453_),
    .C(net552),
    .A(net586),
    .Y(_0585_));
 sg13g2_o21ai_1 _1422_ (.B1(_0454_),
    .Y(_0586_),
    .A1(net572),
    .A2(net559));
 sg13g2_nand3_1 _1423_ (.B(_0585_),
    .C(_0586_),
    .A(net526),
    .Y(_0587_));
 sg13g2_nor3_1 _1424_ (.A(net576),
    .B(\mem[181] ),
    .C(net564),
    .Y(_0588_));
 sg13g2_a21oi_1 _1425_ (.A1(net590),
    .A2(net557),
    .Y(_0589_),
    .B1(\mem[189] ));
 sg13g2_or3_2 _1426_ (.A(net515),
    .B(_0588_),
    .C(_0589_),
    .X(_0590_));
 sg13g2_nand4_1 _1427_ (.B(_0584_),
    .C(_0587_),
    .A(_0581_),
    .Y(_0591_),
    .D(_0590_));
 sg13g2_mux2_1 _1428_ (.A0(\mem[101] ),
    .A1(\mem[109] ),
    .S(net538),
    .X(_0592_));
 sg13g2_mux2_1 _1429_ (.A0(\mem[85] ),
    .A1(\mem[93] ),
    .S(net538),
    .X(_0593_));
 sg13g2_a22oi_1 _1430_ (.Y(_0594_),
    .B1(_0593_),
    .B2(net513),
    .A2(_0592_),
    .A1(net529));
 sg13g2_mux2_1 _1431_ (.A0(\mem[69] ),
    .A1(\mem[77] ),
    .S(net538),
    .X(_0595_));
 sg13g2_mux2_1 _1432_ (.A0(\mem[117] ),
    .A1(\mem[125] ),
    .S(net538),
    .X(_0596_));
 sg13g2_a22oi_1 _1433_ (.Y(_0597_),
    .B1(_0596_),
    .B2(net517),
    .A2(_0595_),
    .A1(net524));
 sg13g2_a21o_1 _1434_ (.A2(_0597_),
    .A1(_0594_),
    .B1(net544),
    .X(_0598_));
 sg13g2_nand3_1 _1435_ (.B(_0450_),
    .C(net552),
    .A(net586),
    .Y(_0599_));
 sg13g2_a21oi_1 _1436_ (.A1(net586),
    .A2(net552),
    .Y(_0600_),
    .B1(\mem[237] ));
 sg13g2_nand3b_1 _1437_ (.B(net525),
    .C(_0599_),
    .Y(_0601_),
    .A_N(_0600_));
 sg13g2_nor3_1 _1438_ (.A(net576),
    .B(\mem[245] ),
    .C(net564),
    .Y(_0602_));
 sg13g2_a21oi_1 _1439_ (.A1(net590),
    .A2(net557),
    .Y(_0603_),
    .B1(\mem[253] ));
 sg13g2_or3_2 _1440_ (.A(net515),
    .B(_0602_),
    .C(_0603_),
    .X(_0604_));
 sg13g2_a21oi_1 _1441_ (.A1(net587),
    .A2(net553),
    .Y(_0605_),
    .B1(\mem[221] ));
 sg13g2_nor3_1 _1442_ (.A(net572),
    .B(\mem[213] ),
    .C(net559),
    .Y(_0606_));
 sg13g2_or3_1 _1443_ (.A(net510),
    .B(_0605_),
    .C(_0606_),
    .X(_0607_));
 sg13g2_nand3_1 _1444_ (.B(_0451_),
    .C(net552),
    .A(net586),
    .Y(_0608_));
 sg13g2_o21ai_1 _1445_ (.B1(_0452_),
    .Y(_0609_),
    .A1(net572),
    .A2(net559));
 sg13g2_nand3_1 _1446_ (.B(_0608_),
    .C(_0609_),
    .A(net521),
    .Y(_0610_));
 sg13g2_nand4_1 _1447_ (.B(_0604_),
    .C(_0607_),
    .A(_0601_),
    .Y(_0611_),
    .D(_0610_));
 sg13g2_a22oi_1 _1448_ (.Y(_0612_),
    .B1(_0611_),
    .B2(net508),
    .A2(_0591_),
    .A1(net551));
 sg13g2_nand2_1 _1449_ (.Y(\rdata_curr_a[2] ),
    .A(_0598_),
    .B(_0612_));
 sg13g2_mux2_1 _1450_ (.A0(\mem[100] ),
    .A1(\mem[108] ),
    .S(net536),
    .X(_0613_));
 sg13g2_mux2_1 _1451_ (.A0(\mem[84] ),
    .A1(\mem[92] ),
    .S(net536),
    .X(_0614_));
 sg13g2_a22oi_1 _1452_ (.Y(_0615_),
    .B1(_0614_),
    .B2(net513),
    .A2(_0613_),
    .A1(net529));
 sg13g2_mux2_1 _1453_ (.A0(\mem[68] ),
    .A1(\mem[76] ),
    .S(net536),
    .X(_0616_));
 sg13g2_mux2_1 _1454_ (.A0(\mem[116] ),
    .A1(\mem[124] ),
    .S(net536),
    .X(_0617_));
 sg13g2_a22oi_1 _1455_ (.Y(_0618_),
    .B1(_0617_),
    .B2(net517),
    .A2(_0616_),
    .A1(net524));
 sg13g2_a21oi_1 _1456_ (.A1(_0615_),
    .A2(_0618_),
    .Y(_0619_),
    .B1(net544));
 sg13g2_mux2_1 _1457_ (.A0(\mem[132] ),
    .A1(\mem[140] ),
    .S(net530),
    .X(_0620_));
 sg13g2_mux2_1 _1458_ (.A0(\mem[148] ),
    .A1(\mem[156] ),
    .S(net534),
    .X(_0621_));
 sg13g2_a22oi_1 _1459_ (.Y(_0622_),
    .B1(_0621_),
    .B2(net512),
    .A2(_0620_),
    .A1(net522));
 sg13g2_mux2_2 _1460_ (.A0(\mem[164] ),
    .A1(\mem[172] ),
    .S(net534),
    .X(_0623_));
 sg13g2_mux2_1 _1461_ (.A0(\mem[180] ),
    .A1(\mem[188] ),
    .S(net537),
    .X(_0624_));
 sg13g2_a22oi_1 _1462_ (.Y(_0625_),
    .B1(_0624_),
    .B2(net518),
    .A2(_0623_),
    .A1(net526));
 sg13g2_a21oi_1 _1463_ (.A1(_0622_),
    .A2(_0625_),
    .Y(_0626_),
    .B1(_0528_));
 sg13g2_mux2_2 _1464_ (.A0(\mem[228] ),
    .A1(\mem[236] ),
    .S(net531),
    .X(_0627_));
 sg13g2_mux2_1 _1465_ (.A0(\mem[244] ),
    .A1(\mem[252] ),
    .S(net537),
    .X(_0628_));
 sg13g2_a22oi_1 _1466_ (.Y(_0629_),
    .B1(_0628_),
    .B2(net516),
    .A2(_0627_),
    .A1(net525));
 sg13g2_mux2_1 _1467_ (.A0(\mem[212] ),
    .A1(\mem[220] ),
    .S(net532),
    .X(_0630_));
 sg13g2_mux2_1 _1468_ (.A0(\mem[196] ),
    .A1(\mem[204] ),
    .S(net531),
    .X(_0631_));
 sg13g2_a22oi_1 _1469_ (.Y(_0632_),
    .B1(_0631_),
    .B2(net521),
    .A2(_0630_),
    .A1(net511));
 sg13g2_a21oi_1 _1470_ (.A1(_0629_),
    .A2(_0632_),
    .Y(_0633_),
    .B1(_0530_));
 sg13g2_or3_2 _1471_ (.A(_0619_),
    .B(_0626_),
    .C(_0633_),
    .X(\rdata_curr_a[3] ));
 sg13g2_a21oi_1 _1472_ (.A1(net588),
    .A2(net555),
    .Y(_0634_),
    .B1(\mem[251] ));
 sg13g2_nor3_1 _1473_ (.A(net575),
    .B(\mem[243] ),
    .C(net562),
    .Y(_0635_));
 sg13g2_nor3_1 _1474_ (.A(_0515_),
    .B(_0634_),
    .C(_0635_),
    .Y(_0636_));
 sg13g2_a21oi_1 _1475_ (.A1(net589),
    .A2(net556),
    .Y(_0637_),
    .B1(\mem[235] ));
 sg13g2_nor3_1 _1476_ (.A(net574),
    .B(\mem[227] ),
    .C(net563),
    .Y(_0638_));
 sg13g2_nor3_1 _1477_ (.A(_0511_),
    .B(_0637_),
    .C(_0638_),
    .Y(_0639_));
 sg13g2_nor3_1 _1478_ (.A(net575),
    .B(\mem[211] ),
    .C(net561),
    .Y(_0640_));
 sg13g2_a21oi_1 _1479_ (.A1(net590),
    .A2(net554),
    .Y(_0641_),
    .B1(\mem[219] ));
 sg13g2_nor3_1 _1480_ (.A(net510),
    .B(_0640_),
    .C(_0641_),
    .Y(_0642_));
 sg13g2_nor3_1 _1481_ (.A(net574),
    .B(\mem[195] ),
    .C(net563),
    .Y(_0643_));
 sg13g2_a21oi_1 _1482_ (.A1(net589),
    .A2(net556),
    .Y(_0644_),
    .B1(\mem[203] ));
 sg13g2_nor3_1 _1483_ (.A(_0513_),
    .B(_0643_),
    .C(_0644_),
    .Y(_0645_));
 sg13g2_or4_1 _1484_ (.A(_0636_),
    .B(_0639_),
    .C(_0642_),
    .D(_0645_),
    .X(_0646_));
 sg13g2_mux2_1 _1485_ (.A0(\mem[99] ),
    .A1(\mem[107] ),
    .S(net532),
    .X(_0647_));
 sg13g2_mux2_1 _1486_ (.A0(\mem[83] ),
    .A1(\mem[91] ),
    .S(net532),
    .X(_0648_));
 sg13g2_a22oi_1 _1487_ (.Y(_0649_),
    .B1(_0648_),
    .B2(net511),
    .A2(_0647_),
    .A1(net528));
 sg13g2_mux2_1 _1488_ (.A0(\mem[115] ),
    .A1(\mem[123] ),
    .S(net532),
    .X(_0650_));
 sg13g2_mux2_1 _1489_ (.A0(\mem[67] ),
    .A1(\mem[75] ),
    .S(net530),
    .X(_0651_));
 sg13g2_a22oi_1 _1490_ (.Y(_0652_),
    .B1(_0651_),
    .B2(net523),
    .A2(_0650_),
    .A1(net516));
 sg13g2_a21o_2 _1491_ (.A2(_0652_),
    .A1(_0649_),
    .B1(net543),
    .X(_0653_));
 sg13g2_nor3_1 _1492_ (.A(net575),
    .B(\mem[179] ),
    .C(net562),
    .Y(_0654_));
 sg13g2_a21oi_1 _1493_ (.A1(net588),
    .A2(net554),
    .Y(_0655_),
    .B1(\mem[187] ));
 sg13g2_nor3_1 _1494_ (.A(_0515_),
    .B(_0654_),
    .C(_0655_),
    .Y(_0656_));
 sg13g2_nor3_1 _1495_ (.A(net574),
    .B(\mem[131] ),
    .C(net563),
    .Y(_0657_));
 sg13g2_a21oi_1 _1496_ (.A1(net589),
    .A2(net556),
    .Y(_0658_),
    .B1(\mem[139] ));
 sg13g2_nor3_1 _1497_ (.A(_0513_),
    .B(_0657_),
    .C(_0658_),
    .Y(_0659_));
 sg13g2_nor3_1 _1498_ (.A(net574),
    .B(\mem[163] ),
    .C(net563),
    .Y(_0660_));
 sg13g2_a21oi_1 _1499_ (.A1(net589),
    .A2(net556),
    .Y(_0661_),
    .B1(\mem[171] ));
 sg13g2_nor3_1 _1500_ (.A(_0511_),
    .B(_0660_),
    .C(_0661_),
    .Y(_0662_));
 sg13g2_a21oi_1 _1501_ (.A1(net588),
    .A2(net555),
    .Y(_0663_),
    .B1(\mem[155] ));
 sg13g2_nor3_1 _1502_ (.A(net575),
    .B(\mem[147] ),
    .C(net562),
    .Y(_0664_));
 sg13g2_nor3_1 _1503_ (.A(net510),
    .B(_0663_),
    .C(_0664_),
    .Y(_0665_));
 sg13g2_or4_1 _1504_ (.A(_0656_),
    .B(_0659_),
    .C(_0662_),
    .D(_0665_),
    .X(_0666_));
 sg13g2_a22oi_1 _1505_ (.Y(_0667_),
    .B1(_0666_),
    .B2(net551),
    .A2(_0646_),
    .A1(net509));
 sg13g2_nand2_1 _1506_ (.Y(\rdata_curr_a[4] ),
    .A(_0653_),
    .B(_0667_));
 sg13g2_mux2_1 _1507_ (.A0(\mem[66] ),
    .A1(\mem[74] ),
    .S(net530),
    .X(_0668_));
 sg13g2_mux2_1 _1508_ (.A0(\mem[98] ),
    .A1(\mem[106] ),
    .S(net530),
    .X(_0669_));
 sg13g2_mux2_1 _1509_ (.A0(\mem[114] ),
    .A1(\mem[122] ),
    .S(net532),
    .X(_0670_));
 sg13g2_mux2_1 _1510_ (.A0(\mem[82] ),
    .A1(\mem[90] ),
    .S(net532),
    .X(_0671_));
 sg13g2_a22oi_1 _1511_ (.Y(_0672_),
    .B1(_0671_),
    .B2(net511),
    .A2(_0668_),
    .A1(net521));
 sg13g2_a22oi_1 _1512_ (.Y(_0673_),
    .B1(_0670_),
    .B2(net516),
    .A2(_0669_),
    .A1(net525));
 sg13g2_a21oi_1 _1513_ (.A1(_0672_),
    .A2(_0673_),
    .Y(_0674_),
    .B1(net543));
 sg13g2_mux2_1 _1514_ (.A0(\mem[194] ),
    .A1(\mem[202] ),
    .S(net535),
    .X(_0675_));
 sg13g2_mux2_2 _1515_ (.A0(\mem[210] ),
    .A1(\mem[218] ),
    .S(net541),
    .X(_0676_));
 sg13g2_a22oi_1 _1516_ (.Y(_0677_),
    .B1(_0676_),
    .B2(net512),
    .A2(_0675_),
    .A1(net522));
 sg13g2_mux2_2 _1517_ (.A0(\mem[242] ),
    .A1(\mem[250] ),
    .S(net541),
    .X(_0678_));
 sg13g2_mux2_1 _1518_ (.A0(\mem[226] ),
    .A1(\mem[234] ),
    .S(net535),
    .X(_0679_));
 sg13g2_a22oi_1 _1519_ (.Y(_0680_),
    .B1(_0679_),
    .B2(net527),
    .A2(_0678_),
    .A1(net518));
 sg13g2_a21oi_1 _1520_ (.A1(_0677_),
    .A2(_0680_),
    .Y(_0681_),
    .B1(_0530_));
 sg13g2_mux2_1 _1521_ (.A0(\mem[162] ),
    .A1(\mem[170] ),
    .S(net535),
    .X(_0682_));
 sg13g2_mux2_2 _1522_ (.A0(\mem[146] ),
    .A1(\mem[154] ),
    .S(net542),
    .X(_0683_));
 sg13g2_a22oi_1 _1523_ (.Y(_0684_),
    .B1(_0683_),
    .B2(net512),
    .A2(_0682_),
    .A1(net526));
 sg13g2_mux2_1 _1524_ (.A0(\mem[130] ),
    .A1(\mem[138] ),
    .S(net535),
    .X(_0685_));
 sg13g2_mux2_2 _1525_ (.A0(\mem[178] ),
    .A1(\mem[186] ),
    .S(net541),
    .X(_0686_));
 sg13g2_a22oi_1 _1526_ (.Y(_0687_),
    .B1(_0686_),
    .B2(net518),
    .A2(_0685_),
    .A1(net522));
 sg13g2_a21oi_1 _1527_ (.A1(_0684_),
    .A2(_0687_),
    .Y(_0688_),
    .B1(_0528_));
 sg13g2_or3_2 _1528_ (.A(_0674_),
    .B(_0681_),
    .C(_0688_),
    .X(\rdata_curr_a[5] ));
 sg13g2_mux2_1 _1529_ (.A0(\mem[241] ),
    .A1(\mem[249] ),
    .S(net541),
    .X(_0689_));
 sg13g2_mux2_1 _1530_ (.A0(\mem[225] ),
    .A1(\mem[233] ),
    .S(net535),
    .X(_0690_));
 sg13g2_mux2_1 _1531_ (.A0(\mem[193] ),
    .A1(\mem[201] ),
    .S(net534),
    .X(_0691_));
 sg13g2_mux2_1 _1532_ (.A0(\mem[209] ),
    .A1(\mem[217] ),
    .S(net541),
    .X(_0692_));
 sg13g2_a22oi_1 _1533_ (.Y(_0693_),
    .B1(_0691_),
    .B2(net522),
    .A2(_0690_),
    .A1(net526));
 sg13g2_a22oi_1 _1534_ (.Y(_0694_),
    .B1(_0692_),
    .B2(net514),
    .A2(_0689_),
    .A1(net519));
 sg13g2_a21oi_1 _1535_ (.A1(_0693_),
    .A2(_0694_),
    .Y(_0695_),
    .B1(_0530_));
 sg13g2_mux2_1 _1536_ (.A0(\mem[97] ),
    .A1(\mem[105] ),
    .S(net530),
    .X(_0696_));
 sg13g2_mux2_1 _1537_ (.A0(\mem[81] ),
    .A1(\mem[89] ),
    .S(net532),
    .X(_0697_));
 sg13g2_a22oi_1 _1538_ (.Y(_0698_),
    .B1(_0697_),
    .B2(net511),
    .A2(_0696_),
    .A1(net525));
 sg13g2_mux2_1 _1539_ (.A0(\mem[113] ),
    .A1(\mem[121] ),
    .S(net532),
    .X(_0699_));
 sg13g2_mux2_1 _1540_ (.A0(\mem[65] ),
    .A1(\mem[73] ),
    .S(net530),
    .X(_0700_));
 sg13g2_a22oi_1 _1541_ (.Y(_0701_),
    .B1(_0700_),
    .B2(net521),
    .A2(_0699_),
    .A1(net516));
 sg13g2_a21oi_1 _1542_ (.A1(_0698_),
    .A2(_0701_),
    .Y(_0702_),
    .B1(net543));
 sg13g2_mux2_1 _1543_ (.A0(\mem[177] ),
    .A1(\mem[185] ),
    .S(net541),
    .X(_0703_));
 sg13g2_mux2_1 _1544_ (.A0(\mem[145] ),
    .A1(\mem[153] ),
    .S(net541),
    .X(_0704_));
 sg13g2_a22oi_1 _1545_ (.Y(_0705_),
    .B1(_0704_),
    .B2(net514),
    .A2(_0703_),
    .A1(net518));
 sg13g2_mux2_1 _1546_ (.A0(\mem[161] ),
    .A1(\mem[169] ),
    .S(net534),
    .X(_0706_));
 sg13g2_mux2_1 _1547_ (.A0(\mem[129] ),
    .A1(\mem[137] ),
    .S(net534),
    .X(_0707_));
 sg13g2_a22oi_1 _1548_ (.Y(_0708_),
    .B1(_0707_),
    .B2(net522),
    .A2(_0706_),
    .A1(net526));
 sg13g2_a21oi_1 _1549_ (.A1(_0705_),
    .A2(_0708_),
    .Y(_0709_),
    .B1(_0528_));
 sg13g2_or3_2 _1550_ (.A(_0695_),
    .B(_0702_),
    .C(_0709_),
    .X(\rdata_curr_a[6] ));
 sg13g2_a21oi_1 _1551_ (.A1(net588),
    .A2(net554),
    .Y(_0710_),
    .B1(\mem[248] ));
 sg13g2_nor3_1 _1552_ (.A(net575),
    .B(\mem[240] ),
    .C(net561),
    .Y(_0711_));
 sg13g2_nor3_1 _1553_ (.A(net515),
    .B(_0710_),
    .C(_0711_),
    .Y(_0712_));
 sg13g2_a21oi_1 _1554_ (.A1(net591),
    .A2(net558),
    .Y(_0713_),
    .B1(\mem[200] ));
 sg13g2_nor3_1 _1555_ (.A(net573),
    .B(\mem[192] ),
    .C(net560),
    .Y(_0714_));
 sg13g2_nor3_2 _1556_ (.A(net520),
    .B(_0713_),
    .C(_0714_),
    .Y(_0715_));
 sg13g2_nor3_1 _1557_ (.A(net574),
    .B(\mem[224] ),
    .C(net563),
    .Y(_0716_));
 sg13g2_a21oi_1 _1558_ (.A1(net589),
    .A2(net556),
    .Y(_0717_),
    .B1(\mem[232] ));
 sg13g2_nor3_1 _1559_ (.A(_0511_),
    .B(_0716_),
    .C(_0717_),
    .Y(_0718_));
 sg13g2_nor3_1 _1560_ (.A(net574),
    .B(\mem[208] ),
    .C(net561),
    .Y(_0719_));
 sg13g2_a21oi_1 _1561_ (.A1(net588),
    .A2(net554),
    .Y(_0720_),
    .B1(\mem[216] ));
 sg13g2_nor3_1 _1562_ (.A(net510),
    .B(_0719_),
    .C(_0720_),
    .Y(_0721_));
 sg13g2_or4_1 _1563_ (.A(_0712_),
    .B(_0715_),
    .C(_0718_),
    .D(_0721_),
    .X(_0722_));
 sg13g2_mux2_2 _1564_ (.A0(\mem[96] ),
    .A1(\mem[104] ),
    .S(net530),
    .X(_0723_));
 sg13g2_mux2_1 _1565_ (.A0(\mem[80] ),
    .A1(\mem[88] ),
    .S(net536),
    .X(_0724_));
 sg13g2_a22oi_1 _1566_ (.Y(_0725_),
    .B1(_0724_),
    .B2(net511),
    .A2(_0723_),
    .A1(net528));
 sg13g2_mux2_1 _1567_ (.A0(\mem[112] ),
    .A1(\mem[120] ),
    .S(net536),
    .X(_0726_));
 sg13g2_mux2_2 _1568_ (.A0(\mem[64] ),
    .A1(\mem[72] ),
    .S(net530),
    .X(_0727_));
 sg13g2_a22oi_1 _1569_ (.Y(_0728_),
    .B1(_0727_),
    .B2(net521),
    .A2(_0726_),
    .A1(net516));
 sg13g2_a21o_2 _1570_ (.A2(_0728_),
    .A1(_0725_),
    .B1(net543),
    .X(_0729_));
 sg13g2_nor3_1 _1571_ (.A(net574),
    .B(\mem[160] ),
    .C(net563),
    .Y(_0730_));
 sg13g2_a21oi_1 _1572_ (.A1(net589),
    .A2(net556),
    .Y(_0731_),
    .B1(\mem[168] ));
 sg13g2_nor3_1 _1573_ (.A(_0511_),
    .B(_0730_),
    .C(_0731_),
    .Y(_0732_));
 sg13g2_nor3_1 _1574_ (.A(net575),
    .B(\mem[144] ),
    .C(net561),
    .Y(_0733_));
 sg13g2_a21oi_1 _1575_ (.A1(net588),
    .A2(net554),
    .Y(_0734_),
    .B1(\mem[152] ));
 sg13g2_nor3_1 _1576_ (.A(net510),
    .B(_0733_),
    .C(_0734_),
    .Y(_0735_));
 sg13g2_nor3_1 _1577_ (.A(net573),
    .B(\mem[128] ),
    .C(net560),
    .Y(_0736_));
 sg13g2_a21oi_1 _1578_ (.A1(net591),
    .A2(net558),
    .Y(_0737_),
    .B1(\mem[136] ));
 sg13g2_nor3_2 _1579_ (.A(net520),
    .B(_0736_),
    .C(_0737_),
    .Y(_0738_));
 sg13g2_a21oi_1 _1580_ (.A1(net588),
    .A2(net554),
    .Y(_0739_),
    .B1(\mem[184] ));
 sg13g2_nor3_1 _1581_ (.A(net574),
    .B(\mem[176] ),
    .C(net562),
    .Y(_0740_));
 sg13g2_nor3_1 _1582_ (.A(net515),
    .B(_0739_),
    .C(_0740_),
    .Y(_0741_));
 sg13g2_or4_1 _1583_ (.A(_0732_),
    .B(_0735_),
    .C(_0738_),
    .D(_0741_),
    .X(_0742_));
 sg13g2_a22oi_1 _1584_ (.Y(_0743_),
    .B1(_0742_),
    .B2(net551),
    .A2(_0722_),
    .A1(net509));
 sg13g2_nand2_1 _1585_ (.Y(\rdata_curr_a[7] ),
    .A(_0729_),
    .B(_0743_));
 sg13g2_a21oi_1 _1586_ (.A1(_0653_),
    .A2(_0667_),
    .Y(_0744_),
    .B1(net565));
 sg13g2_o21ai_1 _1587_ (.B1(net577),
    .Y(_0745_),
    .A1(_0498_),
    .A2(_0499_));
 sg13g2_a21o_1 _1588_ (.A2(net565),
    .A1(\rdata_buff_a[0] ),
    .B1(net577),
    .X(_0746_));
 sg13g2_a21oi_1 _1589_ (.A1(_0498_),
    .A2(\rdata_curr_a[0] ),
    .Y(_0747_),
    .B1(_0746_));
 sg13g2_nand2_2 _1590_ (.Y(_0748_),
    .A(write_through),
    .B(net11));
 sg13g2_o21ai_1 _1591_ (.B1(_0748_),
    .Y(_0749_),
    .A1(_0744_),
    .A2(_0745_));
 sg13g2_nand3_1 _1592_ (.B(net11),
    .C(net623),
    .A(write_through),
    .Y(_0750_));
 sg13g2_o21ai_1 _1593_ (.B1(_0750_),
    .Y(uo_out[0]),
    .A1(_0747_),
    .A2(_0749_));
 sg13g2_o21ai_1 _1594_ (.B1(net577),
    .Y(_0751_),
    .A1(_0498_),
    .A2(_0500_));
 sg13g2_a21oi_1 _1595_ (.A1(_0498_),
    .A2(\rdata_curr_a[5] ),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_a21oi_1 _1596_ (.A1(_0564_),
    .A2(_0578_),
    .Y(_0753_),
    .B1(net565));
 sg13g2_a21o_1 _1597_ (.A2(\rdata_buff_a[1] ),
    .A1(net565),
    .B1(net577),
    .X(_0754_));
 sg13g2_o21ai_1 _1598_ (.B1(_0748_),
    .Y(_0755_),
    .A1(_0753_),
    .A2(_0754_));
 sg13g2_nand3_1 _1599_ (.B(net11),
    .C(net617),
    .A(write_through),
    .Y(_0756_));
 sg13g2_o21ai_1 _1600_ (.B1(_0756_),
    .Y(uo_out[1]),
    .A1(_0752_),
    .A2(_0755_));
 sg13g2_o21ai_1 _1601_ (.B1(net8),
    .Y(_0757_),
    .A1(_0498_),
    .A2(_0501_));
 sg13g2_a21oi_1 _1602_ (.A1(_0498_),
    .A2(\rdata_curr_a[6] ),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_a21oi_1 _1603_ (.A1(_0598_),
    .A2(_0612_),
    .Y(_0759_),
    .B1(net565));
 sg13g2_a21o_1 _1604_ (.A2(\rdata_buff_a[2] ),
    .A1(net565),
    .B1(net577),
    .X(_0760_));
 sg13g2_o21ai_1 _1605_ (.B1(_0748_),
    .Y(_0761_),
    .A1(_0759_),
    .A2(_0760_));
 sg13g2_nand3_1 _1606_ (.B(net11),
    .C(net607),
    .A(write_through),
    .Y(_0762_));
 sg13g2_o21ai_1 _1607_ (.B1(_0762_),
    .Y(uo_out[2]),
    .A1(_0758_),
    .A2(_0761_));
 sg13g2_a21oi_1 _1608_ (.A1(_0729_),
    .A2(_0743_),
    .Y(_0763_),
    .B1(net565));
 sg13g2_o21ai_1 _1609_ (.B1(net577),
    .Y(_0764_),
    .A1(_0498_),
    .A2(_0502_));
 sg13g2_a21o_1 _1610_ (.A2(\rdata_buff_a[3] ),
    .A1(net565),
    .B1(net8),
    .X(_0765_));
 sg13g2_a21oi_1 _1611_ (.A1(_0498_),
    .A2(\rdata_curr_a[3] ),
    .Y(_0766_),
    .B1(_0765_));
 sg13g2_o21ai_1 _1612_ (.B1(_0748_),
    .Y(_0767_),
    .A1(_0763_),
    .A2(_0764_));
 sg13g2_nand3_1 _1613_ (.B(net11),
    .C(net600),
    .A(write_through),
    .Y(_0768_));
 sg13g2_o21ai_1 _1614_ (.B1(_0768_),
    .Y(uo_out[3]),
    .A1(_0766_),
    .A2(_0767_));
 sg13g2_nand2_2 _1615_ (.Y(_0769_),
    .A(net566),
    .B(net7));
 sg13g2_and2_1 _1616_ (.A(net584),
    .B(_0769_),
    .X(_0770_));
 sg13g2_nand2_1 _1617_ (.Y(_0771_),
    .A(net584),
    .B(_0769_));
 sg13g2_and2_1 _1618_ (.A(net6),
    .B(_0769_),
    .X(_0772_));
 sg13g2_nand2_1 _1619_ (.Y(_0773_),
    .A(net6),
    .B(_0769_));
 sg13g2_a21oi_1 _1620_ (.A1(_0440_),
    .A2(net583),
    .Y(_0774_),
    .B1(net488));
 sg13g2_o21ai_1 _1621_ (.B1(_0774_),
    .Y(_0775_),
    .A1(\mem[111] ),
    .A2(net507));
 sg13g2_a21oi_1 _1622_ (.A1(_0441_),
    .A2(net583),
    .Y(_0776_),
    .B1(net481));
 sg13g2_o21ai_1 _1623_ (.B1(_0776_),
    .Y(_0777_),
    .A1(\mem[79] ),
    .A2(net507));
 sg13g2_and2_1 _1624_ (.A(net5),
    .B(_0769_),
    .X(_0778_));
 sg13g2_nand2_2 _1625_ (.Y(_0779_),
    .A(net5),
    .B(_0769_));
 sg13g2_nand3_1 _1626_ (.B(_0777_),
    .C(net476),
    .A(_0775_),
    .Y(_0780_));
 sg13g2_nor2b_1 _1627_ (.A(net7),
    .B_N(net566),
    .Y(_0781_));
 sg13g2_mux4_1 _1628_ (.S0(net496),
    .A0(\mem[119] ),
    .A1(\mem[127] ),
    .A2(\mem[87] ),
    .A3(\mem[95] ),
    .S1(net488),
    .X(_0782_));
 sg13g2_nand2_1 _1629_ (.Y(_0783_),
    .A(\mem[255] ),
    .B(net493));
 sg13g2_nor2b_1 _1630_ (.A(net566),
    .B_N(net7),
    .Y(_0784_));
 sg13g2_nand2_1 _1631_ (.Y(_0785_),
    .A(net7),
    .B(_0769_));
 sg13g2_a21oi_1 _1632_ (.A1(\mem[247] ),
    .A2(net502),
    .Y(_0786_),
    .B1(net546));
 sg13g2_nand2_1 _1633_ (.Y(_0787_),
    .A(\mem[191] ),
    .B(net494));
 sg13g2_a21oi_1 _1634_ (.A1(\mem[183] ),
    .A2(net503),
    .Y(_0788_),
    .B1(net472));
 sg13g2_a221oi_1 _1635_ (.B2(_0788_),
    .C1(net487),
    .B1(_0787_),
    .A1(_0783_),
    .Y(_0789_),
    .A2(_0786_));
 sg13g2_a221oi_1 _1636_ (.B2(\mem[215] ),
    .C1(net548),
    .B1(net500),
    .A1(\mem[223] ),
    .Y(_0790_),
    .A2(net569));
 sg13g2_a221oi_1 _1637_ (.B2(\mem[151] ),
    .C1(net471),
    .B1(net501),
    .A1(\mem[159] ),
    .Y(_0791_),
    .A2(net569));
 sg13g2_nor3_2 _1638_ (.A(net480),
    .B(_0790_),
    .C(_0791_),
    .Y(_0792_));
 sg13g2_o21ai_1 _1639_ (.B1(_0779_),
    .Y(_0793_),
    .A1(_0789_),
    .A2(_0792_));
 sg13g2_a22oi_1 _1640_ (.Y(_0794_),
    .B1(net490),
    .B2(_0437_),
    .A2(net580),
    .A1(_0436_));
 sg13g2_a22oi_1 _1641_ (.Y(_0795_),
    .B1(net492),
    .B2(_0435_),
    .A2(net579),
    .A1(_0434_));
 sg13g2_a21oi_1 _1642_ (.A1(_0438_),
    .A2(net568),
    .Y(_0796_),
    .B1(net478));
 sg13g2_o21ai_1 _1643_ (.B1(_0796_),
    .Y(_0797_),
    .A1(\mem[135] ),
    .A2(net490));
 sg13g2_a21oi_1 _1644_ (.A1(net478),
    .A2(_0794_),
    .Y(_0798_),
    .B1(net470));
 sg13g2_a21oi_1 _1645_ (.A1(_0433_),
    .A2(net579),
    .Y(_0799_),
    .B1(net484));
 sg13g2_o21ai_1 _1646_ (.B1(_0799_),
    .Y(_0800_),
    .A1(\mem[239] ),
    .A2(net499));
 sg13g2_a21oi_1 _1647_ (.A1(net484),
    .A2(_0795_),
    .Y(_0801_),
    .B1(net545));
 sg13g2_a22oi_1 _1648_ (.Y(_0802_),
    .B1(_0800_),
    .B2(_0801_),
    .A2(_0798_),
    .A1(_0797_));
 sg13g2_o21ai_1 _1649_ (.B1(_0780_),
    .Y(_0803_),
    .A1(net475),
    .A2(_0782_));
 sg13g2_a21oi_1 _1650_ (.A1(net475),
    .A2(_0802_),
    .Y(_0804_),
    .B1(net550));
 sg13g2_a22oi_1 _1651_ (.Y(\rdata_curr_b[0] ),
    .B1(_0804_),
    .B2(_0793_),
    .A2(_0803_),
    .A1(net550));
 sg13g2_a21oi_1 _1652_ (.A1(_0448_),
    .A2(net583),
    .Y(_0805_),
    .B1(net488));
 sg13g2_o21ai_1 _1653_ (.B1(_0805_),
    .Y(_0806_),
    .A1(\mem[110] ),
    .A2(net507));
 sg13g2_a21oi_1 _1654_ (.A1(_0449_),
    .A2(net583),
    .Y(_0807_),
    .B1(net481));
 sg13g2_o21ai_1 _1655_ (.B1(_0807_),
    .Y(_0808_),
    .A1(\mem[78] ),
    .A2(net502));
 sg13g2_nand3_1 _1656_ (.B(_0806_),
    .C(_0808_),
    .A(net476),
    .Y(_0809_));
 sg13g2_mux4_1 _1657_ (.S0(net496),
    .A0(\mem[118] ),
    .A1(\mem[126] ),
    .A2(\mem[86] ),
    .A3(\mem[94] ),
    .S1(net487),
    .X(_0810_));
 sg13g2_nand2_1 _1658_ (.Y(_0811_),
    .A(\mem[254] ),
    .B(net493));
 sg13g2_a21oi_1 _1659_ (.A1(\mem[246] ),
    .A2(net503),
    .Y(_0812_),
    .B1(net546));
 sg13g2_nand2_1 _1660_ (.Y(_0813_),
    .A(\mem[190] ),
    .B(net494));
 sg13g2_a21oi_1 _1661_ (.A1(\mem[182] ),
    .A2(net503),
    .Y(_0814_),
    .B1(net472));
 sg13g2_a221oi_1 _1662_ (.B2(_0814_),
    .C1(net489),
    .B1(_0813_),
    .A1(_0811_),
    .Y(_0815_),
    .A2(_0812_));
 sg13g2_a221oi_1 _1663_ (.B2(\mem[214] ),
    .C1(net548),
    .B1(net500),
    .A1(\mem[222] ),
    .Y(_0816_),
    .A2(net569));
 sg13g2_a221oi_1 _1664_ (.B2(\mem[150] ),
    .C1(net470),
    .B1(net501),
    .A1(\mem[158] ),
    .Y(_0817_),
    .A2(net569));
 sg13g2_nor3_2 _1665_ (.A(net479),
    .B(_0816_),
    .C(_0817_),
    .Y(_0818_));
 sg13g2_o21ai_1 _1666_ (.B1(_0779_),
    .Y(_0819_),
    .A1(_0815_),
    .A2(_0818_));
 sg13g2_a22oi_1 _1667_ (.Y(_0820_),
    .B1(net490),
    .B2(_0446_),
    .A2(net580),
    .A1(_0445_));
 sg13g2_a22oi_1 _1668_ (.Y(_0821_),
    .B1(net492),
    .B2(_0444_),
    .A2(net579),
    .A1(_0443_));
 sg13g2_a21oi_1 _1669_ (.A1(_0447_),
    .A2(net568),
    .Y(_0822_),
    .B1(net478));
 sg13g2_o21ai_1 _1670_ (.B1(_0822_),
    .Y(_0823_),
    .A1(\mem[134] ),
    .A2(net490));
 sg13g2_a21oi_1 _1671_ (.A1(net478),
    .A2(_0820_),
    .Y(_0824_),
    .B1(net470));
 sg13g2_a21oi_1 _1672_ (.A1(_0442_),
    .A2(net579),
    .Y(_0825_),
    .B1(net483));
 sg13g2_o21ai_1 _1673_ (.B1(_0825_),
    .Y(_0826_),
    .A1(\mem[238] ),
    .A2(net499));
 sg13g2_a21oi_1 _1674_ (.A1(net483),
    .A2(_0821_),
    .Y(_0827_),
    .B1(net545));
 sg13g2_a22oi_1 _1675_ (.Y(_0828_),
    .B1(_0826_),
    .B2(_0827_),
    .A2(_0824_),
    .A1(_0823_));
 sg13g2_o21ai_1 _1676_ (.B1(_0809_),
    .Y(_0829_),
    .A1(net476),
    .A2(_0810_));
 sg13g2_a21oi_1 _1677_ (.A1(_0778_),
    .A2(_0828_),
    .Y(_0830_),
    .B1(net550));
 sg13g2_a22oi_1 _1678_ (.Y(\rdata_curr_b[1] ),
    .B1(_0830_),
    .B2(_0819_),
    .A2(_0829_),
    .A1(net550));
 sg13g2_a21oi_1 _1679_ (.A1(_0456_),
    .A2(net583),
    .Y(_0831_),
    .B1(net487));
 sg13g2_o21ai_1 _1680_ (.B1(_0831_),
    .Y(_0832_),
    .A1(\mem[109] ),
    .A2(net502));
 sg13g2_a21oi_1 _1681_ (.A1(_0457_),
    .A2(net583),
    .Y(_0833_),
    .B1(net481));
 sg13g2_o21ai_1 _1682_ (.B1(_0833_),
    .Y(_0834_),
    .A1(\mem[77] ),
    .A2(net502));
 sg13g2_nand3_1 _1683_ (.B(_0832_),
    .C(_0834_),
    .A(net476),
    .Y(_0835_));
 sg13g2_mux4_1 _1684_ (.S0(net493),
    .A0(\mem[117] ),
    .A1(\mem[125] ),
    .A2(\mem[85] ),
    .A3(\mem[93] ),
    .S1(net487),
    .X(_0836_));
 sg13g2_nand2_1 _1685_ (.Y(_0837_),
    .A(\mem[253] ),
    .B(net493));
 sg13g2_a21oi_1 _1686_ (.A1(\mem[245] ),
    .A2(net503),
    .Y(_0838_),
    .B1(net546));
 sg13g2_nand2_1 _1687_ (.Y(_0839_),
    .A(\mem[189] ),
    .B(net494));
 sg13g2_a21oi_1 _1688_ (.A1(\mem[181] ),
    .A2(net503),
    .Y(_0840_),
    .B1(net472));
 sg13g2_a221oi_1 _1689_ (.B2(_0840_),
    .C1(net489),
    .B1(_0839_),
    .A1(_0837_),
    .Y(_0841_),
    .A2(_0838_));
 sg13g2_a221oi_1 _1690_ (.B2(\mem[213] ),
    .C1(net545),
    .B1(net500),
    .A1(\mem[221] ),
    .Y(_0842_),
    .A2(net569));
 sg13g2_a221oi_1 _1691_ (.B2(\mem[149] ),
    .C1(net470),
    .B1(net501),
    .A1(\mem[157] ),
    .Y(_0843_),
    .A2(net568));
 sg13g2_nor3_2 _1692_ (.A(net479),
    .B(_0842_),
    .C(_0843_),
    .Y(_0192_));
 sg13g2_o21ai_1 _1693_ (.B1(_0779_),
    .Y(_0193_),
    .A1(_0841_),
    .A2(_0192_));
 sg13g2_a22oi_1 _1694_ (.Y(_0194_),
    .B1(net490),
    .B2(_0454_),
    .A2(net580),
    .A1(_0453_));
 sg13g2_a22oi_1 _1695_ (.Y(_0195_),
    .B1(net492),
    .B2(_0452_),
    .A2(net579),
    .A1(_0451_));
 sg13g2_a21oi_1 _1696_ (.A1(_0455_),
    .A2(net568),
    .Y(_0196_),
    .B1(net478));
 sg13g2_o21ai_1 _1697_ (.B1(_0196_),
    .Y(_0197_),
    .A1(\mem[133] ),
    .A2(net490));
 sg13g2_a21oi_1 _1698_ (.A1(net478),
    .A2(_0194_),
    .Y(_0198_),
    .B1(net470));
 sg13g2_a21oi_1 _1699_ (.A1(_0450_),
    .A2(net579),
    .Y(_0199_),
    .B1(net483));
 sg13g2_o21ai_1 _1700_ (.B1(_0199_),
    .Y(_0200_),
    .A1(\mem[237] ),
    .A2(net499));
 sg13g2_a21oi_1 _1701_ (.A1(net483),
    .A2(_0195_),
    .Y(_0201_),
    .B1(net545));
 sg13g2_a22oi_1 _1702_ (.Y(_0202_),
    .B1(_0200_),
    .B2(_0201_),
    .A2(_0198_),
    .A1(_0197_));
 sg13g2_o21ai_1 _1703_ (.B1(_0835_),
    .Y(_0203_),
    .A1(net476),
    .A2(_0836_));
 sg13g2_a21oi_1 _1704_ (.A1(net475),
    .A2(_0202_),
    .Y(_0204_),
    .B1(net550));
 sg13g2_a22oi_1 _1705_ (.Y(\rdata_curr_b[2] ),
    .B1(_0204_),
    .B2(_0193_),
    .A2(_0203_),
    .A1(net550));
 sg13g2_a21oi_1 _1706_ (.A1(_0464_),
    .A2(net583),
    .Y(_0205_),
    .B1(net487));
 sg13g2_o21ai_1 _1707_ (.B1(_0205_),
    .Y(_0206_),
    .A1(\mem[108] ),
    .A2(net502));
 sg13g2_a21oi_1 _1708_ (.A1(_0465_),
    .A2(net583),
    .Y(_0207_),
    .B1(net481));
 sg13g2_o21ai_1 _1709_ (.B1(_0207_),
    .Y(_0208_),
    .A1(\mem[76] ),
    .A2(net502));
 sg13g2_nand3_1 _1710_ (.B(_0206_),
    .C(_0208_),
    .A(net476),
    .Y(_0209_));
 sg13g2_mux4_1 _1711_ (.S0(net493),
    .A0(\mem[116] ),
    .A1(\mem[124] ),
    .A2(\mem[84] ),
    .A3(\mem[92] ),
    .S1(net487),
    .X(_0210_));
 sg13g2_nand2_1 _1712_ (.Y(_0211_),
    .A(\mem[252] ),
    .B(net493));
 sg13g2_a21oi_1 _1713_ (.A1(\mem[244] ),
    .A2(net502),
    .Y(_0212_),
    .B1(net546));
 sg13g2_nand2_1 _1714_ (.Y(_0213_),
    .A(\mem[188] ),
    .B(net493));
 sg13g2_a21oi_1 _1715_ (.A1(\mem[180] ),
    .A2(net502),
    .Y(_0214_),
    .B1(net472));
 sg13g2_a221oi_1 _1716_ (.B2(_0214_),
    .C1(net487),
    .B1(_0213_),
    .A1(_0211_),
    .Y(_0215_),
    .A2(_0212_));
 sg13g2_a221oi_1 _1717_ (.B2(\mem[212] ),
    .C1(net548),
    .B1(net500),
    .A1(\mem[220] ),
    .Y(_0216_),
    .A2(net569));
 sg13g2_a221oi_1 _1718_ (.B2(\mem[148] ),
    .C1(net471),
    .B1(net501),
    .A1(\mem[156] ),
    .Y(_0217_),
    .A2(net569));
 sg13g2_nor3_2 _1719_ (.A(net480),
    .B(_0216_),
    .C(_0217_),
    .Y(_0218_));
 sg13g2_o21ai_1 _1720_ (.B1(_0779_),
    .Y(_0219_),
    .A1(_0215_),
    .A2(_0218_));
 sg13g2_a22oi_1 _1721_ (.Y(_0220_),
    .B1(net490),
    .B2(_0462_),
    .A2(net580),
    .A1(_0461_));
 sg13g2_a22oi_1 _1722_ (.Y(_0221_),
    .B1(net492),
    .B2(_0460_),
    .A2(net579),
    .A1(_0459_));
 sg13g2_a21oi_1 _1723_ (.A1(_0463_),
    .A2(net568),
    .Y(_0222_),
    .B1(net480));
 sg13g2_o21ai_1 _1724_ (.B1(_0222_),
    .Y(_0223_),
    .A1(\mem[132] ),
    .A2(net492));
 sg13g2_a21oi_1 _1725_ (.A1(net478),
    .A2(_0220_),
    .Y(_0224_),
    .B1(net470));
 sg13g2_a21oi_1 _1726_ (.A1(_0458_),
    .A2(net579),
    .Y(_0225_),
    .B1(net484));
 sg13g2_o21ai_1 _1727_ (.B1(_0225_),
    .Y(_0226_),
    .A1(\mem[236] ),
    .A2(net499));
 sg13g2_a21oi_1 _1728_ (.A1(net484),
    .A2(_0221_),
    .Y(_0227_),
    .B1(net545));
 sg13g2_a22oi_1 _1729_ (.Y(_0228_),
    .B1(_0226_),
    .B2(_0227_),
    .A2(_0224_),
    .A1(_0223_));
 sg13g2_o21ai_1 _1730_ (.B1(_0209_),
    .Y(_0229_),
    .A1(net476),
    .A2(_0210_));
 sg13g2_a21oi_1 _1731_ (.A1(net475),
    .A2(_0228_),
    .Y(_0230_),
    .B1(net549));
 sg13g2_a22oi_1 _1732_ (.Y(\rdata_curr_b[3] ),
    .B1(_0230_),
    .B2(_0219_),
    .A2(_0229_),
    .A1(net549));
 sg13g2_a21oi_1 _1733_ (.A1(_0472_),
    .A2(net578),
    .Y(_0231_),
    .B1(net483));
 sg13g2_o21ai_1 _1734_ (.B1(_0231_),
    .Y(_0232_),
    .A1(\mem[107] ),
    .A2(net498));
 sg13g2_a21oi_1 _1735_ (.A1(_0473_),
    .A2(net578),
    .Y(_0233_),
    .B1(net480));
 sg13g2_o21ai_1 _1736_ (.B1(_0233_),
    .Y(_0234_),
    .A1(\mem[75] ),
    .A2(net498));
 sg13g2_nand3_1 _1737_ (.B(_0232_),
    .C(_0234_),
    .A(net477),
    .Y(_0235_));
 sg13g2_mux4_1 _1738_ (.S0(net492),
    .A0(\mem[115] ),
    .A1(\mem[123] ),
    .A2(\mem[83] ),
    .A3(\mem[91] ),
    .S1(net485),
    .X(_0236_));
 sg13g2_nand2_1 _1739_ (.Y(_0237_),
    .A(\mem[179] ),
    .B(net504));
 sg13g2_a21oi_1 _1740_ (.A1(\mem[187] ),
    .A2(net495),
    .Y(_0238_),
    .B1(net473));
 sg13g2_nand2_1 _1741_ (.Y(_0239_),
    .A(\mem[251] ),
    .B(net495));
 sg13g2_a21oi_1 _1742_ (.A1(\mem[243] ),
    .A2(net504),
    .Y(_0240_),
    .B1(net547));
 sg13g2_a221oi_1 _1743_ (.B2(_0240_),
    .C1(net488),
    .B1(_0239_),
    .A1(_0237_),
    .Y(_0241_),
    .A2(_0238_));
 sg13g2_a221oi_1 _1744_ (.B2(\mem[211] ),
    .C1(net547),
    .B1(net503),
    .A1(\mem[219] ),
    .Y(_0242_),
    .A2(net571));
 sg13g2_a221oi_1 _1745_ (.B2(\mem[147] ),
    .C1(net473),
    .B1(net504),
    .A1(\mem[155] ),
    .Y(_0243_),
    .A2(net570));
 sg13g2_nor3_1 _1746_ (.A(net481),
    .B(_0242_),
    .C(_0243_),
    .Y(_0244_));
 sg13g2_o21ai_1 _1747_ (.B1(_0779_),
    .Y(_0245_),
    .A1(_0241_),
    .A2(_0244_));
 sg13g2_a22oi_1 _1748_ (.Y(_0246_),
    .B1(net491),
    .B2(_0470_),
    .A2(net581),
    .A1(_0469_));
 sg13g2_a22oi_1 _1749_ (.Y(_0247_),
    .B1(net494),
    .B2(_0468_),
    .A2(net582),
    .A1(_0467_));
 sg13g2_a21oi_1 _1750_ (.A1(_0471_),
    .A2(net570),
    .Y(_0248_),
    .B1(net482));
 sg13g2_o21ai_1 _1751_ (.B1(_0248_),
    .Y(_0249_),
    .A1(\mem[131] ),
    .A2(net494));
 sg13g2_a21oi_1 _1752_ (.A1(net482),
    .A2(_0246_),
    .Y(_0250_),
    .B1(net471));
 sg13g2_a21oi_1 _1753_ (.A1(_0466_),
    .A2(net584),
    .Y(_0251_),
    .B1(net489));
 sg13g2_o21ai_1 _1754_ (.B1(_0251_),
    .Y(_0252_),
    .A1(\mem[235] ),
    .A2(net506));
 sg13g2_a21oi_1 _1755_ (.A1(net486),
    .A2(_0247_),
    .Y(_0253_),
    .B1(net546));
 sg13g2_a22oi_1 _1756_ (.Y(_0254_),
    .B1(_0252_),
    .B2(_0253_),
    .A2(_0250_),
    .A1(_0249_));
 sg13g2_o21ai_1 _1757_ (.B1(_0235_),
    .Y(_0255_),
    .A1(net477),
    .A2(_0236_));
 sg13g2_a21oi_1 _1758_ (.A1(net475),
    .A2(_0254_),
    .Y(_0256_),
    .B1(net549));
 sg13g2_a22oi_1 _1759_ (.Y(\rdata_curr_b[4] ),
    .B1(_0256_),
    .B2(_0245_),
    .A2(_0255_),
    .A1(net549));
 sg13g2_a21oi_1 _1760_ (.A1(_0480_),
    .A2(net578),
    .Y(_0257_),
    .B1(net483));
 sg13g2_o21ai_1 _1761_ (.B1(_0257_),
    .Y(_0258_),
    .A1(\mem[106] ),
    .A2(net498));
 sg13g2_a21oi_1 _1762_ (.A1(_0481_),
    .A2(net578),
    .Y(_0259_),
    .B1(net480));
 sg13g2_o21ai_1 _1763_ (.B1(_0259_),
    .Y(_0260_),
    .A1(\mem[74] ),
    .A2(net498));
 sg13g2_nand3_1 _1764_ (.B(_0258_),
    .C(_0260_),
    .A(net477),
    .Y(_0261_));
 sg13g2_mux4_1 _1765_ (.S0(net492),
    .A0(\mem[114] ),
    .A1(\mem[122] ),
    .A2(\mem[82] ),
    .A3(\mem[90] ),
    .S1(net485),
    .X(_0262_));
 sg13g2_nand2_1 _1766_ (.Y(_0263_),
    .A(\mem[250] ),
    .B(net495));
 sg13g2_a21oi_1 _1767_ (.A1(\mem[242] ),
    .A2(net505),
    .Y(_0264_),
    .B1(net547));
 sg13g2_nand2_1 _1768_ (.Y(_0265_),
    .A(\mem[186] ),
    .B(net495));
 sg13g2_a21oi_1 _1769_ (.A1(\mem[178] ),
    .A2(net505),
    .Y(_0266_),
    .B1(net473));
 sg13g2_a221oi_1 _1770_ (.B2(_0266_),
    .C1(net488),
    .B1(_0265_),
    .A1(_0263_),
    .Y(_0267_),
    .A2(_0264_));
 sg13g2_a221oi_1 _1771_ (.B2(\mem[210] ),
    .C1(net547),
    .B1(net503),
    .A1(\mem[218] ),
    .Y(_0268_),
    .A2(net570));
 sg13g2_a221oi_1 _1772_ (.B2(\mem[146] ),
    .C1(net472),
    .B1(net504),
    .A1(\mem[154] ),
    .Y(_0269_),
    .A2(net570));
 sg13g2_nor3_1 _1773_ (.A(net481),
    .B(_0268_),
    .C(_0269_),
    .Y(_0270_));
 sg13g2_o21ai_1 _1774_ (.B1(_0779_),
    .Y(_0271_),
    .A1(_0267_),
    .A2(_0270_));
 sg13g2_a22oi_1 _1775_ (.Y(_0272_),
    .B1(net491),
    .B2(_0478_),
    .A2(net581),
    .A1(_0477_));
 sg13g2_a22oi_1 _1776_ (.Y(_0273_),
    .B1(net497),
    .B2(_0476_),
    .A2(net581),
    .A1(_0475_));
 sg13g2_a21oi_1 _1777_ (.A1(_0479_),
    .A2(net568),
    .Y(_0274_),
    .B1(net479));
 sg13g2_o21ai_1 _1778_ (.B1(_0274_),
    .Y(_0275_),
    .A1(\mem[130] ),
    .A2(net497));
 sg13g2_a21oi_1 _1779_ (.A1(net479),
    .A2(_0272_),
    .Y(_0276_),
    .B1(net471));
 sg13g2_a21oi_1 _1780_ (.A1(_0474_),
    .A2(net581),
    .Y(_0277_),
    .B1(net486));
 sg13g2_o21ai_1 _1781_ (.B1(_0277_),
    .Y(_0278_),
    .A1(\mem[234] ),
    .A2(net501));
 sg13g2_a21oi_1 _1782_ (.A1(net486),
    .A2(_0273_),
    .Y(_0279_),
    .B1(net545));
 sg13g2_a22oi_1 _1783_ (.Y(_0280_),
    .B1(_0278_),
    .B2(_0279_),
    .A2(_0276_),
    .A1(_0275_));
 sg13g2_o21ai_1 _1784_ (.B1(_0261_),
    .Y(_0281_),
    .A1(net477),
    .A2(_0262_));
 sg13g2_a21oi_1 _1785_ (.A1(net475),
    .A2(_0280_),
    .Y(_0282_),
    .B1(net549));
 sg13g2_a22oi_1 _1786_ (.Y(\rdata_curr_b[5] ),
    .B1(_0282_),
    .B2(_0271_),
    .A2(_0281_),
    .A1(net550));
 sg13g2_a21oi_1 _1787_ (.A1(_0488_),
    .A2(net578),
    .Y(_0283_),
    .B1(net483));
 sg13g2_o21ai_1 _1788_ (.B1(_0283_),
    .Y(_0284_),
    .A1(\mem[105] ),
    .A2(net498));
 sg13g2_a21oi_1 _1789_ (.A1(_0489_),
    .A2(net578),
    .Y(_0285_),
    .B1(net480));
 sg13g2_o21ai_1 _1790_ (.B1(_0285_),
    .Y(_0286_),
    .A1(\mem[73] ),
    .A2(net498));
 sg13g2_nand3_1 _1791_ (.B(_0284_),
    .C(_0286_),
    .A(net477),
    .Y(_0287_));
 sg13g2_mux4_1 _1792_ (.S0(net492),
    .A0(\mem[113] ),
    .A1(\mem[121] ),
    .A2(\mem[81] ),
    .A3(\mem[89] ),
    .S1(net485),
    .X(_0288_));
 sg13g2_nand2_1 _1793_ (.Y(_0289_),
    .A(\mem[249] ),
    .B(net495));
 sg13g2_a21oi_1 _1794_ (.A1(\mem[241] ),
    .A2(net505),
    .Y(_0290_),
    .B1(net547));
 sg13g2_nand2_1 _1795_ (.Y(_0291_),
    .A(\mem[185] ),
    .B(net494));
 sg13g2_a21oi_1 _1796_ (.A1(\mem[177] ),
    .A2(net504),
    .Y(_0292_),
    .B1(net473));
 sg13g2_a221oi_1 _1797_ (.B2(_0292_),
    .C1(net488),
    .B1(_0291_),
    .A1(_0289_),
    .Y(_0293_),
    .A2(_0290_));
 sg13g2_a221oi_1 _1798_ (.B2(\mem[209] ),
    .C1(net546),
    .B1(net505),
    .A1(\mem[217] ),
    .Y(_0294_),
    .A2(net570));
 sg13g2_a221oi_1 _1799_ (.B2(\mem[145] ),
    .C1(net472),
    .B1(net505),
    .A1(\mem[153] ),
    .Y(_0295_),
    .A2(net570));
 sg13g2_nor3_1 _1800_ (.A(net481),
    .B(_0294_),
    .C(_0295_),
    .Y(_0296_));
 sg13g2_o21ai_1 _1801_ (.B1(_0779_),
    .Y(_0297_),
    .A1(_0293_),
    .A2(_0296_));
 sg13g2_a22oi_1 _1802_ (.Y(_0298_),
    .B1(net491),
    .B2(_0486_),
    .A2(net580),
    .A1(_0485_));
 sg13g2_a22oi_1 _1803_ (.Y(_0299_),
    .B1(net491),
    .B2(_0484_),
    .A2(net580),
    .A1(_0483_));
 sg13g2_a21oi_1 _1804_ (.A1(_0487_),
    .A2(net568),
    .Y(_0300_),
    .B1(net479));
 sg13g2_o21ai_1 _1805_ (.B1(_0300_),
    .Y(_0301_),
    .A1(\mem[129] ),
    .A2(net491));
 sg13g2_a21oi_1 _1806_ (.A1(net479),
    .A2(_0298_),
    .Y(_0302_),
    .B1(net470));
 sg13g2_a21oi_1 _1807_ (.A1(_0482_),
    .A2(net581),
    .Y(_0303_),
    .B1(net486));
 sg13g2_o21ai_1 _1808_ (.B1(_0303_),
    .Y(_0304_),
    .A1(\mem[233] ),
    .A2(net501));
 sg13g2_a21oi_1 _1809_ (.A1(net486),
    .A2(_0299_),
    .Y(_0305_),
    .B1(net545));
 sg13g2_a22oi_1 _1810_ (.Y(_0306_),
    .B1(_0304_),
    .B2(_0305_),
    .A2(_0302_),
    .A1(_0301_));
 sg13g2_o21ai_1 _1811_ (.B1(_0287_),
    .Y(_0307_),
    .A1(net477),
    .A2(_0288_));
 sg13g2_a21oi_1 _1812_ (.A1(net475),
    .A2(_0306_),
    .Y(_0308_),
    .B1(net549));
 sg13g2_a22oi_1 _1813_ (.Y(\rdata_curr_b[6] ),
    .B1(_0308_),
    .B2(_0297_),
    .A2(_0307_),
    .A1(net550));
 sg13g2_a21oi_1 _1814_ (.A1(_0496_),
    .A2(net578),
    .Y(_0309_),
    .B1(net483));
 sg13g2_o21ai_1 _1815_ (.B1(_0309_),
    .Y(_0310_),
    .A1(\mem[104] ),
    .A2(net498));
 sg13g2_a21oi_1 _1816_ (.A1(_0497_),
    .A2(net578),
    .Y(_0311_),
    .B1(net480));
 sg13g2_o21ai_1 _1817_ (.B1(_0311_),
    .Y(_0312_),
    .A1(\mem[72] ),
    .A2(net498));
 sg13g2_nand3_1 _1818_ (.B(_0310_),
    .C(_0312_),
    .A(net477),
    .Y(_0313_));
 sg13g2_mux4_1 _1819_ (.S0(net493),
    .A0(\mem[112] ),
    .A1(\mem[120] ),
    .A2(\mem[80] ),
    .A3(\mem[88] ),
    .S1(net487),
    .X(_0314_));
 sg13g2_nand2_1 _1820_ (.Y(_0315_),
    .A(\mem[248] ),
    .B(net494));
 sg13g2_a21oi_1 _1821_ (.A1(\mem[240] ),
    .A2(net504),
    .Y(_0316_),
    .B1(net546));
 sg13g2_nand2_1 _1822_ (.Y(_0317_),
    .A(\mem[184] ),
    .B(net494));
 sg13g2_a21oi_1 _1823_ (.A1(\mem[176] ),
    .A2(net504),
    .Y(_0318_),
    .B1(net472));
 sg13g2_a221oi_1 _1824_ (.B2(_0318_),
    .C1(net488),
    .B1(_0317_),
    .A1(_0315_),
    .Y(_0319_),
    .A2(_0316_));
 sg13g2_a221oi_1 _1825_ (.B2(\mem[208] ),
    .C1(net546),
    .B1(net503),
    .A1(\mem[216] ),
    .Y(_0320_),
    .A2(net570));
 sg13g2_a221oi_1 _1826_ (.B2(\mem[144] ),
    .C1(net472),
    .B1(net504),
    .A1(\mem[152] ),
    .Y(_0321_),
    .A2(net570));
 sg13g2_nor3_1 _1827_ (.A(net481),
    .B(_0320_),
    .C(_0321_),
    .Y(_0322_));
 sg13g2_o21ai_1 _1828_ (.B1(_0779_),
    .Y(_0323_),
    .A1(_0319_),
    .A2(_0322_));
 sg13g2_a22oi_1 _1829_ (.Y(_0324_),
    .B1(net491),
    .B2(_0494_),
    .A2(net581),
    .A1(_0493_));
 sg13g2_a22oi_1 _1830_ (.Y(_0325_),
    .B1(net490),
    .B2(_0492_),
    .A2(net580),
    .A1(_0491_));
 sg13g2_a21oi_1 _1831_ (.A1(_0495_),
    .A2(net568),
    .Y(_0326_),
    .B1(net478));
 sg13g2_o21ai_1 _1832_ (.B1(_0326_),
    .Y(_0327_),
    .A1(\mem[128] ),
    .A2(net491));
 sg13g2_a21oi_1 _1833_ (.A1(net479),
    .A2(_0324_),
    .Y(_0328_),
    .B1(net470));
 sg13g2_a21oi_1 _1834_ (.A1(_0490_),
    .A2(net581),
    .Y(_0329_),
    .B1(net486));
 sg13g2_o21ai_1 _1835_ (.B1(_0329_),
    .Y(_0330_),
    .A1(\mem[232] ),
    .A2(net501));
 sg13g2_a21oi_1 _1836_ (.A1(net486),
    .A2(_0325_),
    .Y(_0331_),
    .B1(net545));
 sg13g2_a22oi_1 _1837_ (.Y(_0332_),
    .B1(_0330_),
    .B2(_0331_),
    .A2(_0328_),
    .A1(_0327_));
 sg13g2_o21ai_1 _1838_ (.B1(_0313_),
    .Y(_0333_),
    .A1(net477),
    .A2(_0314_));
 sg13g2_a21oi_1 _1839_ (.A1(net475),
    .A2(_0332_),
    .Y(_0334_),
    .B1(net549));
 sg13g2_a22oi_1 _1840_ (.Y(\rdata_curr_b[7] ),
    .B1(_0334_),
    .B2(_0323_),
    .A2(_0333_),
    .A1(net549));
 sg13g2_mux4_1 _1841_ (.S0(net9),
    .A0(\rdata_curr_b[0] ),
    .A1(\rdata_curr_b[4] ),
    .A2(\rdata_buff_b[0] ),
    .A3(\rdata_buff_b[4] ),
    .S1(read_buffer_b),
    .X(uo_out[4]));
 sg13g2_mux4_1 _1842_ (.S0(net9),
    .A0(\rdata_curr_b[1] ),
    .A1(\rdata_curr_b[5] ),
    .A2(\rdata_buff_b[1] ),
    .A3(\rdata_buff_b[5] ),
    .S1(read_buffer_b),
    .X(uo_out[5]));
 sg13g2_mux4_1 _1843_ (.S0(net9),
    .A0(\rdata_curr_b[2] ),
    .A1(\rdata_curr_b[6] ),
    .A2(\rdata_buff_b[2] ),
    .A3(\rdata_buff_b[6] ),
    .S1(read_buffer_b),
    .X(uo_out[6]));
 sg13g2_mux4_1 _1844_ (.S0(net9),
    .A0(\rdata_curr_b[3] ),
    .A1(\rdata_curr_b[7] ),
    .A2(\rdata_buff_b[3] ),
    .A3(\rdata_buff_b[7] ),
    .S1(read_buffer_b),
    .X(uo_out[7]));
 sg13g2_nand2_2 _1845_ (.Y(_0335_),
    .A(net11),
    .B(net577));
 sg13g2_nor2_1 _1846_ (.A(_0508_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_nand2_2 _1847_ (.Y(_0337_),
    .A(net4),
    .B(net513));
 sg13g2_nand3_1 _1848_ (.B(net512),
    .C(net469),
    .A(net585),
    .Y(_0338_));
 sg13g2_mux2_1 _1849_ (.A0(net613),
    .A1(net326),
    .S(_0338_),
    .X(_0000_));
 sg13g2_nand2_2 _1850_ (.Y(_0339_),
    .A(net11),
    .B(_0335_));
 sg13g2_nor2_2 _1851_ (.A(_0508_),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_nand2b_2 _1852_ (.Y(_0341_),
    .B(net537),
    .A_N(_0339_));
 sg13g2_nand2b_2 _1853_ (.Y(_0342_),
    .B(_0340_),
    .A_N(_0337_));
 sg13g2_mux2_1 _1854_ (.A0(net626),
    .A1(net429),
    .S(_0342_),
    .X(_0001_));
 sg13g2_mux2_1 _1855_ (.A0(net604),
    .A1(net332),
    .S(_0338_),
    .X(_0002_));
 sg13g2_mux2_1 _1856_ (.A0(net594),
    .A1(net413),
    .S(_0338_),
    .X(_0003_));
 sg13g2_mux2_1 _1857_ (.A0(net617),
    .A1(net404),
    .S(_0342_),
    .X(_0004_));
 sg13g2_nor2_2 _1858_ (.A(net537),
    .B(_0335_),
    .Y(_0343_));
 sg13g2_or2_2 _1859_ (.X(_0344_),
    .B(_0335_),
    .A(net537));
 sg13g2_nor2_2 _1860_ (.A(_0337_),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_mux2_1 _1861_ (.A0(net378),
    .A1(net621),
    .S(_0345_),
    .X(_0005_));
 sg13g2_mux2_1 _1862_ (.A0(net608),
    .A1(net423),
    .S(_0342_),
    .X(_0006_));
 sg13g2_mux2_1 _1863_ (.A0(net599),
    .A1(net426),
    .S(_0342_),
    .X(_0007_));
 sg13g2_mux2_1 _1864_ (.A0(net382),
    .A1(net612),
    .S(_0345_),
    .X(_0008_));
 sg13g2_nor2_2 _1865_ (.A(net536),
    .B(_0339_),
    .Y(_0346_));
 sg13g2_or2_2 _1866_ (.X(_0347_),
    .B(_0339_),
    .A(net536));
 sg13g2_nor2_2 _1867_ (.A(_0337_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_mux2_1 _1868_ (.A0(net408),
    .A1(net625),
    .S(_0348_),
    .X(_0009_));
 sg13g2_mux2_1 _1869_ (.A0(net359),
    .A1(net594),
    .S(_0345_),
    .X(_0010_));
 sg13g2_mux2_1 _1870_ (.A0(net295),
    .A1(net617),
    .S(_0348_),
    .X(_0011_));
 sg13g2_nand2_2 _1871_ (.Y(_0349_),
    .A(net585),
    .B(net522));
 sg13g2_nor3_2 _1872_ (.A(_0508_),
    .B(_0335_),
    .C(_0349_),
    .Y(_0350_));
 sg13g2_mux2_1 _1873_ (.A0(net343),
    .A1(net619),
    .S(_0350_),
    .X(_0012_));
 sg13g2_mux2_1 _1874_ (.A0(net245),
    .A1(net609),
    .S(_0348_),
    .X(_0013_));
 sg13g2_mux2_1 _1875_ (.A0(net410),
    .A1(net599),
    .S(_0348_),
    .X(_0014_));
 sg13g2_mux2_1 _1876_ (.A0(net240),
    .A1(net612),
    .S(_0350_),
    .X(_0015_));
 sg13g2_nor2_2 _1877_ (.A(_0341_),
    .B(_0349_),
    .Y(_0351_));
 sg13g2_mux2_1 _1878_ (.A0(net427),
    .A1(net621),
    .S(_0351_),
    .X(_0016_));
 sg13g2_mux2_1 _1879_ (.A0(net417),
    .A1(net603),
    .S(_0350_),
    .X(_0017_));
 sg13g2_nand3_1 _1880_ (.B(net509),
    .C(_0346_),
    .A(net513),
    .Y(_0352_));
 sg13g2_mux2_1 _1881_ (.A0(net616),
    .A1(net280),
    .S(_0352_),
    .X(_0018_));
 sg13g2_mux2_1 _1882_ (.A0(net346),
    .A1(net594),
    .S(_0350_),
    .X(_0019_));
 sg13g2_nor2_2 _1883_ (.A(_0344_),
    .B(_0349_),
    .Y(_0353_));
 sg13g2_mux2_1 _1884_ (.A0(net262),
    .A1(net619),
    .S(_0353_),
    .X(_0020_));
 sg13g2_mux2_1 _1885_ (.A0(net335),
    .A1(net603),
    .S(_0351_),
    .X(_0021_));
 sg13g2_nand3_1 _1886_ (.B(net508),
    .C(net469),
    .A(net521),
    .Y(_0354_));
 sg13g2_mux2_1 _1887_ (.A0(net620),
    .A1(net411),
    .S(_0354_),
    .X(_0022_));
 sg13g2_nor3_2 _1888_ (.A(net520),
    .B(_0530_),
    .C(_0347_),
    .Y(_0355_));
 sg13g2_mux2_1 _1889_ (.A0(net372),
    .A1(net612),
    .S(_0355_),
    .X(_0023_));
 sg13g2_nand3_1 _1890_ (.B(net509),
    .C(_0336_),
    .A(net517),
    .Y(_0356_));
 sg13g2_mux2_1 _1891_ (.A0(net623),
    .A1(net370),
    .S(_0356_),
    .X(_0024_));
 sg13g2_mux2_1 _1892_ (.A0(net407),
    .A1(net594),
    .S(_0351_),
    .X(_0025_));
 sg13g2_nand3_1 _1893_ (.B(net508),
    .C(_0343_),
    .A(net525),
    .Y(_0357_));
 sg13g2_mux2_1 _1894_ (.A0(net601),
    .A1(net303),
    .S(_0357_),
    .X(_0026_));
 sg13g2_nand3_1 _1895_ (.B(net551),
    .C(_0346_),
    .A(net518),
    .Y(_0358_));
 sg13g2_mux2_1 _1896_ (.A0(net616),
    .A1(net311),
    .S(_0358_),
    .X(_0027_));
 sg13g2_nand3_1 _1897_ (.B(net551),
    .C(_0336_),
    .A(net519),
    .Y(_0359_));
 sg13g2_mux2_1 _1898_ (.A0(net623),
    .A1(net406),
    .S(_0359_),
    .X(_0028_));
 sg13g2_mux2_1 _1899_ (.A0(net397),
    .A1(net612),
    .S(_0353_),
    .X(_0029_));
 sg13g2_mux2_1 _1900_ (.A0(net609),
    .A1(net297),
    .S(_0352_),
    .X(_0030_));
 sg13g2_mux2_1 _1901_ (.A0(net615),
    .A1(net321),
    .S(_0356_),
    .X(_0031_));
 sg13g2_mux2_1 _1902_ (.A0(net271),
    .A1(net603),
    .S(_0355_),
    .X(_0032_));
 sg13g2_nor2_2 _1903_ (.A(_0347_),
    .B(_0349_),
    .Y(_0360_));
 sg13g2_mux2_1 _1904_ (.A0(net312),
    .A1(net622),
    .S(_0360_),
    .X(_0033_));
 sg13g2_mux2_1 _1905_ (.A0(net625),
    .A1(net422),
    .S(_0358_),
    .X(_0034_));
 sg13g2_nand3_1 _1906_ (.B(net508),
    .C(_0343_),
    .A(net511),
    .Y(_0361_));
 sg13g2_mux2_1 _1907_ (.A0(net593),
    .A1(net318),
    .S(_0361_),
    .X(_0035_));
 sg13g2_nor4_2 _1908_ (.A(net544),
    .B(_0508_),
    .C(net520),
    .Y(_0362_),
    .D(_0335_));
 sg13g2_mux2_1 _1909_ (.A0(net399),
    .A1(net624),
    .S(_0362_),
    .X(_0036_));
 sg13g2_mux2_1 _1910_ (.A0(net327),
    .A1(net603),
    .S(_0353_),
    .X(_0037_));
 sg13g2_mux2_1 _1911_ (.A0(net276),
    .A1(net592),
    .S(_0353_),
    .X(_0038_));
 sg13g2_mux2_1 _1912_ (.A0(net274),
    .A1(net613),
    .S(_0360_),
    .X(_0039_));
 sg13g2_nand3_1 _1913_ (.B(net517),
    .C(net469),
    .A(_0506_),
    .Y(_0363_));
 sg13g2_nor2_1 _1914_ (.A(net623),
    .B(_0363_),
    .Y(_0364_));
 sg13g2_a21oi_1 _1915_ (.A1(_0439_),
    .A2(_0363_),
    .Y(_0040_),
    .B1(_0364_));
 sg13g2_mux2_1 _1916_ (.A0(net334),
    .A1(net594),
    .S(_0355_),
    .X(_0041_));
 sg13g2_nand3_1 _1917_ (.B(net551),
    .C(_0343_),
    .A(net516),
    .Y(_0365_));
 sg13g2_mux2_1 _1918_ (.A0(net608),
    .A1(net388),
    .S(_0365_),
    .X(_0042_));
 sg13g2_mux2_1 _1919_ (.A0(net287),
    .A1(net595),
    .S(_0360_),
    .X(_0043_));
 sg13g2_mux2_1 _1920_ (.A0(net618),
    .A1(net323),
    .S(_0363_),
    .X(_0044_));
 sg13g2_nand3_1 _1921_ (.B(net516),
    .C(_0340_),
    .A(_0506_),
    .Y(_0366_));
 sg13g2_mux2_1 _1922_ (.A0(net620),
    .A1(net390),
    .S(_0366_),
    .X(_0045_));
 sg13g2_mux2_1 _1923_ (.A0(net606),
    .A1(net338),
    .S(_0363_),
    .X(_0046_));
 sg13g2_nand2_2 _1924_ (.Y(_0367_),
    .A(net566),
    .B(net513));
 sg13g2_or2_2 _1925_ (.X(_0368_),
    .B(_0367_),
    .A(_0341_));
 sg13g2_mux2_1 _1926_ (.A0(net602),
    .A1(net356),
    .S(_0368_),
    .X(_0047_));
 sg13g2_mux2_1 _1927_ (.A0(net597),
    .A1(net355),
    .S(_0363_),
    .X(_0048_));
 sg13g2_mux2_1 _1928_ (.A0(net611),
    .A1(net401),
    .S(_0366_),
    .X(_0049_));
 sg13g2_mux2_1 _1929_ (.A0(net616),
    .A1(net322),
    .S(_0359_),
    .X(_0050_));
 sg13g2_nor3_2 _1930_ (.A(net520),
    .B(_0530_),
    .C(_0344_),
    .Y(_0369_));
 sg13g2_mux2_1 _1931_ (.A0(net288),
    .A1(net620),
    .S(_0369_),
    .X(_0051_));
 sg13g2_mux2_1 _1932_ (.A0(net598),
    .A1(net324),
    .S(_0352_),
    .X(_0052_));
 sg13g2_mux2_1 _1933_ (.A0(net602),
    .A1(net379),
    .S(_0366_),
    .X(_0053_));
 sg13g2_mux2_1 _1934_ (.A0(net598),
    .A1(net362),
    .S(_0365_),
    .X(_0054_));
 sg13g2_mux2_1 _1935_ (.A0(net596),
    .A1(net330),
    .S(_0366_),
    .X(_0055_));
 sg13g2_mux2_1 _1936_ (.A0(net602),
    .A1(net391),
    .S(_0361_),
    .X(_0056_));
 sg13g2_nand2_2 _1937_ (.Y(_0370_),
    .A(net566),
    .B(net529));
 sg13g2_nor2_2 _1938_ (.A(_0347_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_nand2_1 _1939_ (.Y(_0372_),
    .A(net610),
    .B(_0371_));
 sg13g2_o21ai_1 _1940_ (.B1(_0372_),
    .Y(_0057_),
    .A1(_0480_),
    .A2(_0371_));
 sg13g2_nand3_1 _1941_ (.B(net509),
    .C(_0340_),
    .A(net513),
    .Y(_0373_));
 sg13g2_mux2_1 _1942_ (.A0(net616),
    .A1(net331),
    .S(_0373_),
    .X(_0058_));
 sg13g2_nand3_1 _1943_ (.B(net517),
    .C(_0343_),
    .A(_0506_),
    .Y(_0374_));
 sg13g2_mux2_1 _1944_ (.A0(net618),
    .A1(net320),
    .S(_0374_),
    .X(_0059_));
 sg13g2_nand3_1 _1945_ (.B(net516),
    .C(_0346_),
    .A(_0506_),
    .Y(_0375_));
 sg13g2_mux2_1 _1946_ (.A0(net620),
    .A1(net300),
    .S(_0375_),
    .X(_0060_));
 sg13g2_nand3_1 _1947_ (.B(net509),
    .C(_0340_),
    .A(net518),
    .Y(_0376_));
 sg13g2_mux2_1 _1948_ (.A0(net608),
    .A1(net409),
    .S(_0376_),
    .X(_0061_));
 sg13g2_mux2_1 _1949_ (.A0(net606),
    .A1(net313),
    .S(_0374_),
    .X(_0062_));
 sg13g2_mux2_1 _1950_ (.A0(net597),
    .A1(net308),
    .S(_0374_),
    .X(_0063_));
 sg13g2_nand3_1 _1951_ (.B(net551),
    .C(_0340_),
    .A(net518),
    .Y(_0377_));
 sg13g2_mux2_1 _1952_ (.A0(net626),
    .A1(net430),
    .S(_0377_),
    .X(_0064_));
 sg13g2_mux2_1 _1953_ (.A0(net611),
    .A1(net316),
    .S(_0375_),
    .X(_0065_));
 sg13g2_nand3_1 _1954_ (.B(net529),
    .C(net469),
    .A(net566),
    .Y(_0378_));
 sg13g2_mux2_1 _1955_ (.A0(net624),
    .A1(net418),
    .S(_0378_),
    .X(_0066_));
 sg13g2_mux2_1 _1956_ (.A0(net606),
    .A1(net395),
    .S(_0378_),
    .X(_0067_));
 sg13g2_mux2_1 _1957_ (.A0(net610),
    .A1(net302),
    .S(_0354_),
    .X(_0068_));
 sg13g2_mux2_1 _1958_ (.A0(net602),
    .A1(net301),
    .S(_0375_),
    .X(_0069_));
 sg13g2_mux2_1 _1959_ (.A0(net596),
    .A1(net328),
    .S(_0375_),
    .X(_0070_));
 sg13g2_mux2_1 _1960_ (.A0(net615),
    .A1(net414),
    .S(_0378_),
    .X(_0071_));
 sg13g2_mux2_1 _1961_ (.A0(net420),
    .A1(net612),
    .S(_0351_),
    .X(_0072_));
 sg13g2_or2_2 _1962_ (.X(_0379_),
    .B(_0370_),
    .A(_0341_));
 sg13g2_mux2_1 _1963_ (.A0(net619),
    .A1(net412),
    .S(_0379_),
    .X(_0073_));
 sg13g2_mux2_1 _1964_ (.A0(net596),
    .A1(net363),
    .S(_0378_),
    .X(_0074_));
 sg13g2_nand2_2 _1965_ (.Y(_0380_),
    .A(net585),
    .B(net527));
 sg13g2_nand3_1 _1966_ (.B(net526),
    .C(net469),
    .A(net585),
    .Y(_0381_));
 sg13g2_nor2_1 _1967_ (.A(net621),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_a21oi_1 _1968_ (.A1(_0437_),
    .A2(_0381_),
    .Y(_0075_),
    .B1(_0382_));
 sg13g2_mux2_1 _1969_ (.A0(net610),
    .A1(net339),
    .S(_0379_),
    .X(_0076_));
 sg13g2_nand3_1 _1970_ (.B(net509),
    .C(_0340_),
    .A(net523),
    .Y(_0383_));
 sg13g2_mux2_1 _1971_ (.A0(net621),
    .A1(net358),
    .S(_0383_),
    .X(_0077_));
 sg13g2_nor2_2 _1972_ (.A(_0344_),
    .B(_0370_),
    .Y(_0384_));
 sg13g2_nand2_1 _1973_ (.Y(_0385_),
    .A(net623),
    .B(_0384_));
 sg13g2_o21ai_1 _1974_ (.B1(_0385_),
    .Y(_0078_),
    .A1(_0440_),
    .A2(_0384_));
 sg13g2_mux2_1 _1975_ (.A0(net625),
    .A1(net329),
    .S(_0352_),
    .X(_0079_));
 sg13g2_mux2_1 _1976_ (.A0(net601),
    .A1(net368),
    .S(_0379_),
    .X(_0080_));
 sg13g2_mux2_1 _1977_ (.A0(net624),
    .A1(net421),
    .S(_0374_),
    .X(_0081_));
 sg13g2_mux2_1 _1978_ (.A0(net592),
    .A1(net398),
    .S(_0379_),
    .X(_0082_));
 sg13g2_nand2_1 _1979_ (.Y(_0386_),
    .A(net615),
    .B(_0384_));
 sg13g2_o21ai_1 _1980_ (.B1(_0386_),
    .Y(_0083_),
    .A1(_0448_),
    .A2(_0384_));
 sg13g2_mux2_1 _1981_ (.A0(net608),
    .A1(net336),
    .S(_0358_),
    .X(_0084_));
 sg13g2_nand2_1 _1982_ (.Y(_0387_),
    .A(net606),
    .B(_0384_));
 sg13g2_o21ai_1 _1983_ (.B1(_0387_),
    .Y(_0085_),
    .A1(_0456_),
    .A2(_0384_));
 sg13g2_mux2_1 _1984_ (.A0(net265),
    .A1(net610),
    .S(_0369_),
    .X(_0086_));
 sg13g2_mux2_1 _1985_ (.A0(net598),
    .A1(net393),
    .S(_0359_),
    .X(_0087_));
 sg13g2_nand2_1 _1986_ (.Y(_0388_),
    .A(net596),
    .B(_0384_));
 sg13g2_o21ai_1 _1987_ (.B1(_0388_),
    .Y(_0088_),
    .A1(_0464_),
    .A2(_0384_));
 sg13g2_mux2_1 _1988_ (.A0(net255),
    .A1(net603),
    .S(_0360_),
    .X(_0089_));
 sg13g2_mux2_1 _1989_ (.A0(net601),
    .A1(net296),
    .S(_0354_),
    .X(_0090_));
 sg13g2_nand3_1 _1990_ (.B(net513),
    .C(net469),
    .A(net566),
    .Y(_0389_));
 sg13g2_mux2_1 _1991_ (.A0(net623),
    .A1(net381),
    .S(_0389_),
    .X(_0091_));
 sg13g2_nand2_1 _1992_ (.Y(_0390_),
    .A(net601),
    .B(_0371_));
 sg13g2_o21ai_1 _1993_ (.B1(_0390_),
    .Y(_0092_),
    .A1(_0488_),
    .A2(_0371_));
 sg13g2_nand2_1 _1994_ (.Y(_0391_),
    .A(net592),
    .B(_0371_));
 sg13g2_o21ai_1 _1995_ (.B1(_0391_),
    .Y(_0093_),
    .A1(_0496_),
    .A2(_0371_));
 sg13g2_mux2_1 _1996_ (.A0(net269),
    .A1(net604),
    .S(_0345_),
    .X(_0094_));
 sg13g2_mux2_1 _1997_ (.A0(net616),
    .A1(net374),
    .S(_0377_),
    .X(_0095_));
 sg13g2_mux2_1 _1998_ (.A0(net608),
    .A1(net402),
    .S(_0359_),
    .X(_0096_));
 sg13g2_mux2_1 _1999_ (.A0(net615),
    .A1(net349),
    .S(_0389_),
    .X(_0097_));
 sg13g2_nand3_1 _2000_ (.B(net508),
    .C(net469),
    .A(net525),
    .Y(_0392_));
 sg13g2_mux2_1 _2001_ (.A0(net619),
    .A1(net354),
    .S(_0392_),
    .X(_0098_));
 sg13g2_mux2_1 _2002_ (.A0(net625),
    .A1(net292),
    .S(_0365_),
    .X(_0099_));
 sg13g2_mux2_1 _2003_ (.A0(net621),
    .A1(net419),
    .S(_0338_),
    .X(_0100_));
 sg13g2_mux2_1 _2004_ (.A0(net620),
    .A1(net365),
    .S(_0368_),
    .X(_0101_));
 sg13g2_mux2_1 _2005_ (.A0(net608),
    .A1(net416),
    .S(_0377_),
    .X(_0102_));
 sg13g2_or2_2 _2006_ (.X(_0393_),
    .B(_0380_),
    .A(_0341_));
 sg13g2_nor2_1 _2007_ (.A(net604),
    .B(_0393_),
    .Y(_0394_));
 sg13g2_a21oi_1 _2008_ (.A1(_0486_),
    .A2(_0393_),
    .Y(_0103_),
    .B1(_0394_));
 sg13g2_mux2_1 _2009_ (.A0(net606),
    .A1(net369),
    .S(_0389_),
    .X(_0104_));
 sg13g2_mux2_1 _2010_ (.A0(net616),
    .A1(net383),
    .S(_0365_),
    .X(_0105_));
 sg13g2_mux2_1 _2011_ (.A0(net596),
    .A1(net341),
    .S(_0389_),
    .X(_0106_));
 sg13g2_mux2_1 _2012_ (.A0(net611),
    .A1(net367),
    .S(_0368_),
    .X(_0107_));
 sg13g2_nor2_2 _2013_ (.A(_0344_),
    .B(_0367_),
    .Y(_0395_));
 sg13g2_mux2_1 _2014_ (.A0(net281),
    .A1(net623),
    .S(_0395_),
    .X(_0108_));
 sg13g2_mux2_1 _2015_ (.A0(net593),
    .A1(net357),
    .S(_0354_),
    .X(_0109_));
 sg13g2_mux2_1 _2016_ (.A0(net593),
    .A1(net348),
    .S(_0368_),
    .X(_0110_));
 sg13g2_mux2_1 _2017_ (.A0(net243),
    .A1(net615),
    .S(_0395_),
    .X(_0111_));
 sg13g2_nor2_2 _2018_ (.A(_0347_),
    .B(_0367_),
    .Y(_0396_));
 sg13g2_mux2_1 _2019_ (.A0(net241),
    .A1(net620),
    .S(_0396_),
    .X(_0112_));
 sg13g2_mux2_1 _2020_ (.A0(net613),
    .A1(net392),
    .S(_0383_),
    .X(_0113_));
 sg13g2_mux2_1 _2021_ (.A0(net247),
    .A1(net606),
    .S(_0395_),
    .X(_0114_));
 sg13g2_mux2_1 _2022_ (.A0(net246),
    .A1(net596),
    .S(_0395_),
    .X(_0115_));
 sg13g2_mux2_1 _2023_ (.A0(net256),
    .A1(net611),
    .S(_0396_),
    .X(_0116_));
 sg13g2_mux2_1 _2024_ (.A0(net263),
    .A1(net602),
    .S(_0396_),
    .X(_0117_));
 sg13g2_mux2_1 _2025_ (.A0(net258),
    .A1(net593),
    .S(_0396_),
    .X(_0118_));
 sg13g2_mux2_1 _2026_ (.A0(net310),
    .A1(net615),
    .S(_0362_),
    .X(_0119_));
 sg13g2_nor3_2 _2027_ (.A(net543),
    .B(net520),
    .C(_0341_),
    .Y(_0397_));
 sg13g2_mux2_1 _2028_ (.A0(net352),
    .A1(net619),
    .S(_0397_),
    .X(_0120_));
 sg13g2_mux2_1 _2029_ (.A0(net604),
    .A1(net342),
    .S(_0383_),
    .X(_0121_));
 sg13g2_mux2_1 _2030_ (.A0(net351),
    .A1(net606),
    .S(_0362_),
    .X(_0122_));
 sg13g2_mux2_1 _2031_ (.A0(net291),
    .A1(net596),
    .S(_0362_),
    .X(_0123_));
 sg13g2_mux2_1 _2032_ (.A0(net594),
    .A1(net377),
    .S(_0383_),
    .X(_0124_));
 sg13g2_mux2_1 _2033_ (.A0(net415),
    .A1(net610),
    .S(_0397_),
    .X(_0125_));
 sg13g2_nor3_2 _2034_ (.A(net543),
    .B(net520),
    .C(_0344_),
    .Y(_0398_));
 sg13g2_nand2_1 _2035_ (.Y(_0399_),
    .A(net624),
    .B(_0398_));
 sg13g2_o21ai_1 _2036_ (.B1(_0399_),
    .Y(_0126_),
    .A1(_0441_),
    .A2(_0398_));
 sg13g2_mux2_1 _2037_ (.A0(net347),
    .A1(net601),
    .S(_0397_),
    .X(_0127_));
 sg13g2_mux2_1 _2038_ (.A0(net309),
    .A1(net592),
    .S(_0397_),
    .X(_0128_));
 sg13g2_nand2_1 _2039_ (.Y(_0400_),
    .A(net615),
    .B(_0398_));
 sg13g2_o21ai_1 _2040_ (.B1(_0400_),
    .Y(_0129_),
    .A1(_0449_),
    .A2(_0398_));
 sg13g2_nor3_2 _2041_ (.A(net543),
    .B(net520),
    .C(_0347_),
    .Y(_0401_));
 sg13g2_nand2_1 _2042_ (.Y(_0402_),
    .A(net619),
    .B(_0401_));
 sg13g2_o21ai_1 _2043_ (.B1(_0402_),
    .Y(_0130_),
    .A1(_0473_),
    .A2(_0401_));
 sg13g2_nand2_1 _2044_ (.Y(_0403_),
    .A(net596),
    .B(_0398_));
 sg13g2_o21ai_1 _2045_ (.B1(_0403_),
    .Y(_0131_),
    .A1(_0465_),
    .A2(_0398_));
 sg13g2_mux2_1 _2046_ (.A0(net289),
    .A1(net622),
    .S(_0355_),
    .X(_0132_));
 sg13g2_nand2_1 _2047_ (.Y(_0404_),
    .A(net610),
    .B(_0401_));
 sg13g2_o21ai_1 _2048_ (.B1(_0404_),
    .Y(_0133_),
    .A1(_0481_),
    .A2(_0401_));
 sg13g2_nand2_1 _2049_ (.Y(_0405_),
    .A(net601),
    .B(_0401_));
 sg13g2_o21ai_1 _2050_ (.B1(_0405_),
    .Y(_0134_),
    .A1(_0489_),
    .A2(_0401_));
 sg13g2_nand2_1 _2051_ (.Y(_0406_),
    .A(net592),
    .B(_0401_));
 sg13g2_o21ai_1 _2052_ (.B1(_0406_),
    .Y(_0135_),
    .A1(_0497_),
    .A2(_0401_));
 sg13g2_mux2_1 _2053_ (.A0(net250),
    .A1(net601),
    .S(_0369_),
    .X(_0136_));
 sg13g2_mux2_1 _2054_ (.A0(net599),
    .A1(net431),
    .S(_0377_),
    .X(_0137_));
 sg13g2_mux2_1 _2055_ (.A0(net273),
    .A1(net592),
    .S(_0369_),
    .X(_0138_));
 sg13g2_mux2_1 _2056_ (.A0(net598),
    .A1(net425),
    .S(_0358_),
    .X(_0139_));
 sg13g2_nor2_1 _2057_ (.A(net612),
    .B(_0381_),
    .Y(_0407_));
 sg13g2_a21oi_1 _2058_ (.A1(_0446_),
    .A2(_0381_),
    .Y(_0140_),
    .B1(_0407_));
 sg13g2_nor2_1 _2059_ (.A(net621),
    .B(_0393_),
    .Y(_0408_));
 sg13g2_a21oi_1 _2060_ (.A1(_0470_),
    .A2(_0393_),
    .Y(_0141_),
    .B1(_0408_));
 sg13g2_nor2_1 _2061_ (.A(net603),
    .B(_0381_),
    .Y(_0409_));
 sg13g2_a21oi_1 _2062_ (.A1(_0454_),
    .A2(_0381_),
    .Y(_0142_),
    .B1(_0409_));
 sg13g2_nor2_1 _2063_ (.A(net594),
    .B(_0381_),
    .Y(_0410_));
 sg13g2_a21oi_1 _2064_ (.A1(_0462_),
    .A2(_0381_),
    .Y(_0143_),
    .B1(_0410_));
 sg13g2_nor2_1 _2065_ (.A(net613),
    .B(_0393_),
    .Y(_0411_));
 sg13g2_a21oi_1 _2066_ (.A1(_0478_),
    .A2(_0393_),
    .Y(_0144_),
    .B1(_0411_));
 sg13g2_nor2_2 _2067_ (.A(_0344_),
    .B(_0380_),
    .Y(_0412_));
 sg13g2_nand2_1 _2068_ (.Y(_0413_),
    .A(net621),
    .B(_0412_));
 sg13g2_o21ai_1 _2069_ (.B1(_0413_),
    .Y(_0145_),
    .A1(_0436_),
    .A2(_0412_));
 sg13g2_nor2_1 _2070_ (.A(net595),
    .B(_0393_),
    .Y(_0414_));
 sg13g2_a21oi_1 _2071_ (.A1(_0494_),
    .A2(_0393_),
    .Y(_0146_),
    .B1(_0414_));
 sg13g2_nand2_1 _2072_ (.Y(_0415_),
    .A(net612),
    .B(_0412_));
 sg13g2_o21ai_1 _2073_ (.B1(_0415_),
    .Y(_0147_),
    .A1(_0445_),
    .A2(_0412_));
 sg13g2_nor2_2 _2074_ (.A(_0347_),
    .B(_0380_),
    .Y(_0416_));
 sg13g2_nand2_1 _2075_ (.Y(_0417_),
    .A(net621),
    .B(_0416_));
 sg13g2_o21ai_1 _2076_ (.B1(_0417_),
    .Y(_0148_),
    .A1(_0469_),
    .A2(_0416_));
 sg13g2_nand2_1 _2077_ (.Y(_0418_),
    .A(net603),
    .B(_0412_));
 sg13g2_o21ai_1 _2078_ (.B1(_0418_),
    .Y(_0149_),
    .A1(_0453_),
    .A2(_0412_));
 sg13g2_nand2_1 _2079_ (.Y(_0419_),
    .A(net594),
    .B(_0412_));
 sg13g2_o21ai_1 _2080_ (.B1(_0419_),
    .Y(_0150_),
    .A1(_0461_),
    .A2(_0412_));
 sg13g2_nand2_1 _2081_ (.Y(_0420_),
    .A(net612),
    .B(_0416_));
 sg13g2_o21ai_1 _2082_ (.B1(_0420_),
    .Y(_0151_),
    .A1(_0477_),
    .A2(_0416_));
 sg13g2_nand2_1 _2083_ (.Y(_0421_),
    .A(net604),
    .B(_0416_));
 sg13g2_o21ai_1 _2084_ (.B1(_0421_),
    .Y(_0152_),
    .A1(_0485_),
    .A2(_0416_));
 sg13g2_nand2_1 _2085_ (.Y(_0422_),
    .A(net595),
    .B(_0416_));
 sg13g2_o21ai_1 _2086_ (.B1(_0422_),
    .Y(_0153_),
    .A1(_0493_),
    .A2(_0416_));
 sg13g2_nand2_1 _2087_ (.Y(_0423_),
    .A(net606),
    .B(_0398_));
 sg13g2_o21ai_1 _2088_ (.B1(_0423_),
    .Y(_0154_),
    .A1(_0457_),
    .A2(_0398_));
 sg13g2_mux2_1 _2089_ (.A0(net611),
    .A1(net400),
    .S(_0361_),
    .X(_0155_));
 sg13g2_mux2_1 _2090_ (.A0(net598),
    .A1(net371),
    .S(_0373_),
    .X(_0156_));
 sg13g2_mux2_1 _2091_ (.A0(net608),
    .A1(net373),
    .S(_0373_),
    .X(_0157_));
 sg13g2_mux2_1 _2092_ (.A0(net620),
    .A1(net307),
    .S(_0361_),
    .X(_0158_));
 sg13g2_nand3_1 _2093_ (.B(net508),
    .C(net469),
    .A(net511),
    .Y(_0424_));
 sg13g2_mux2_1 _2094_ (.A0(net593),
    .A1(net376),
    .S(_0424_),
    .X(_0159_));
 sg13g2_mux2_1 _2095_ (.A0(net602),
    .A1(net314),
    .S(_0424_),
    .X(_0160_));
 sg13g2_mux2_1 _2096_ (.A0(net625),
    .A1(net396),
    .S(_0373_),
    .X(_0161_));
 sg13g2_mux2_1 _2097_ (.A0(net611),
    .A1(net333),
    .S(_0424_),
    .X(_0162_));
 sg13g2_nand3_1 _2098_ (.B(_0529_),
    .C(_0346_),
    .A(net529),
    .Y(_0425_));
 sg13g2_mux2_1 _2099_ (.A0(net598),
    .A1(net380),
    .S(_0425_),
    .X(_0163_));
 sg13g2_mux2_1 _2100_ (.A0(net603),
    .A1(net389),
    .S(_0425_),
    .X(_0164_));
 sg13g2_mux2_1 _2101_ (.A0(net622),
    .A1(net360),
    .S(_0424_),
    .X(_0165_));
 sg13g2_mux2_1 _2102_ (.A0(net616),
    .A1(net319),
    .S(_0425_),
    .X(_0166_));
 sg13g2_mux2_1 _2103_ (.A0(net592),
    .A1(net350),
    .S(_0357_),
    .X(_0167_));
 sg13g2_mux2_1 _2104_ (.A0(net625),
    .A1(net405),
    .S(_0425_),
    .X(_0168_));
 sg13g2_mux2_1 _2105_ (.A0(net610),
    .A1(net279),
    .S(_0357_),
    .X(_0169_));
 sg13g2_nand3_1 _2106_ (.B(net508),
    .C(_0340_),
    .A(net527),
    .Y(_0426_));
 sg13g2_mux2_1 _2107_ (.A0(net598),
    .A1(net384),
    .S(_0426_),
    .X(_0170_));
 sg13g2_mux2_1 _2108_ (.A0(net604),
    .A1(net337),
    .S(_0426_),
    .X(_0171_));
 sg13g2_mux2_1 _2109_ (.A0(net619),
    .A1(net366),
    .S(_0357_),
    .X(_0172_));
 sg13g2_mux2_1 _2110_ (.A0(net616),
    .A1(net394),
    .S(_0426_),
    .X(_0173_));
 sg13g2_mux2_1 _2111_ (.A0(net592),
    .A1(net385),
    .S(_0392_),
    .X(_0174_));
 sg13g2_mux2_1 _2112_ (.A0(net601),
    .A1(net386),
    .S(_0392_),
    .X(_0175_));
 sg13g2_mux2_1 _2113_ (.A0(net625),
    .A1(net340),
    .S(_0426_),
    .X(_0176_));
 sg13g2_mux2_1 _2114_ (.A0(net610),
    .A1(net361),
    .S(_0392_),
    .X(_0177_));
 sg13g2_nor3_2 _2115_ (.A(net515),
    .B(_0530_),
    .C(_0347_),
    .Y(_0427_));
 sg13g2_mux2_1 _2116_ (.A0(net344),
    .A1(net598),
    .S(_0427_),
    .X(_0178_));
 sg13g2_mux2_1 _2117_ (.A0(net278),
    .A1(net608),
    .S(_0427_),
    .X(_0179_));
 sg13g2_mux2_1 _2118_ (.A0(net242),
    .A1(net617),
    .S(_0427_),
    .X(_0180_));
 sg13g2_nor3_2 _2119_ (.A(net515),
    .B(_0530_),
    .C(_0344_),
    .Y(_0428_));
 sg13g2_mux2_1 _2120_ (.A0(net254),
    .A1(net597),
    .S(_0428_),
    .X(_0181_));
 sg13g2_mux2_1 _2121_ (.A0(net299),
    .A1(net607),
    .S(_0428_),
    .X(_0182_));
 sg13g2_mux2_1 _2122_ (.A0(net387),
    .A1(net625),
    .S(_0427_),
    .X(_0183_));
 sg13g2_mux2_1 _2123_ (.A0(net304),
    .A1(net615),
    .S(_0428_),
    .X(_0184_));
 sg13g2_mux2_1 _2124_ (.A0(net599),
    .A1(net424),
    .S(_0376_),
    .X(_0185_));
 sg13g2_mux2_1 _2125_ (.A0(net251),
    .A1(net623),
    .S(_0428_),
    .X(_0186_));
 sg13g2_mux2_1 _2126_ (.A0(net617),
    .A1(net375),
    .S(_0376_),
    .X(_0187_));
 sg13g2_mux2_1 _2127_ (.A0(net597),
    .A1(net345),
    .S(_0356_),
    .X(_0188_));
 sg13g2_mux2_1 _2128_ (.A0(net607),
    .A1(net403),
    .S(_0356_),
    .X(_0189_));
 sg13g2_mux2_1 _2129_ (.A0(net626),
    .A1(net428),
    .S(_0376_),
    .X(_0190_));
 sg13g2_nand2_1 _2130_ (.Y(_0429_),
    .A(net619),
    .B(_0371_));
 sg13g2_o21ai_1 _2131_ (.B1(_0429_),
    .Y(_0191_),
    .A1(_0472_),
    .A2(_0371_));
 sg13g2_dfrbp_1 _2132_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net190),
    .D(_0000_),
    .Q_N(_1035_),
    .Q(\mem[158] ));
 sg13g2_dfrbp_1 _2133_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net36),
    .D(_0001_),
    .Q_N(_1034_),
    .Q(\mem[155] ));
 sg13g2_dfrbp_1 _2134_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net35),
    .D(_0002_),
    .Q_N(_1033_),
    .Q(\mem[157] ));
 sg13g2_dfrbp_1 _2135_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net34),
    .D(_0003_),
    .Q_N(_1032_),
    .Q(\mem[156] ));
 sg13g2_dfrbp_1 _2136_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net33),
    .D(_0004_),
    .Q_N(_1031_),
    .Q(\mem[154] ));
 sg13g2_dfrbp_1 _2137_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net32),
    .D(_0005_),
    .Q_N(_1030_),
    .Q(\mem[151] ));
 sg13g2_dfrbp_1 _2138_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net31),
    .D(_0006_),
    .Q_N(_1029_),
    .Q(\mem[153] ));
 sg13g2_dfrbp_1 _2139_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net30),
    .D(_0007_),
    .Q_N(_1028_),
    .Q(\mem[152] ));
 sg13g2_dfrbp_1 _2140_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net29),
    .D(_0008_),
    .Q_N(_1027_),
    .Q(\mem[150] ));
 sg13g2_dfrbp_1 _2141_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net28),
    .D(_0009_),
    .Q_N(_1026_),
    .Q(\mem[147] ));
 sg13g2_dfrbp_1 _2142_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net239),
    .D(_0010_),
    .Q_N(_1025_),
    .Q(\mem[148] ));
 sg13g2_dfrbp_1 _2143_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net238),
    .D(_0011_),
    .Q_N(_1024_),
    .Q(\mem[146] ));
 sg13g2_dfrbp_1 _2144_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net237),
    .D(_0012_),
    .Q_N(_1023_),
    .Q(\mem[143] ));
 sg13g2_dfrbp_1 _2145_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net236),
    .D(_0013_),
    .Q_N(_1022_),
    .Q(\mem[145] ));
 sg13g2_dfrbp_1 _2146_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net235),
    .D(_0014_),
    .Q_N(_1021_),
    .Q(\mem[144] ));
 sg13g2_dfrbp_1 _2147_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net234),
    .D(_0015_),
    .Q_N(_1020_),
    .Q(\mem[142] ));
 sg13g2_dfrbp_1 _2148_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net233),
    .D(_0016_),
    .Q_N(_1019_),
    .Q(\mem[139] ));
 sg13g2_dfrbp_1 _2149_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net232),
    .D(_0017_),
    .Q_N(_1018_),
    .Q(\mem[141] ));
 sg13g2_dfrbp_1 _2150_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net231),
    .D(_0018_),
    .Q_N(_1017_),
    .Q(\mem[210] ));
 sg13g2_dfrbp_1 _2151_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net230),
    .D(_0019_),
    .Q_N(_1016_),
    .Q(\mem[140] ));
 sg13g2_dfrbp_1 _2152_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net229),
    .D(_0020_),
    .Q_N(_1015_),
    .Q(\mem[135] ));
 sg13g2_dfrbp_1 _2153_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net228),
    .D(_0021_),
    .Q_N(_1014_),
    .Q(\mem[137] ));
 sg13g2_dfrbp_1 _2154_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net227),
    .D(_0022_),
    .Q_N(_1013_),
    .Q(\mem[207] ));
 sg13g2_dfrbp_1 _2155_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net226),
    .D(_0023_),
    .Q_N(_1012_),
    .Q(\mem[194] ));
 sg13g2_dfrbp_1 _2156_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net225),
    .D(_0024_),
    .Q_N(_1011_),
    .Q(\mem[255] ));
 sg13g2_dfrbp_1 _2157_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net224),
    .D(_0025_),
    .Q_N(_1010_),
    .Q(\mem[136] ));
 sg13g2_dfrbp_1 _2158_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net223),
    .D(_0026_),
    .Q_N(_1009_),
    .Q(\mem[229] ));
 sg13g2_dfrbp_1 _2159_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net222),
    .D(_0027_),
    .Q_N(_1008_),
    .Q(\mem[178] ));
 sg13g2_dfrbp_1 _2160_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net221),
    .D(_0028_),
    .Q_N(_1007_),
    .Q(\mem[191] ));
 sg13g2_dfrbp_1 _2161_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net220),
    .D(_0029_),
    .Q_N(_1006_),
    .Q(\mem[134] ));
 sg13g2_dfrbp_1 _2162_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net219),
    .D(_0030_),
    .Q_N(_1005_),
    .Q(\mem[209] ));
 sg13g2_dfrbp_1 _2163_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net218),
    .D(_0031_),
    .Q_N(_1004_),
    .Q(\mem[254] ));
 sg13g2_dfrbp_1 _2164_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net217),
    .D(_0032_),
    .Q_N(_1003_),
    .Q(\mem[193] ));
 sg13g2_dfrbp_1 _2165_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net216),
    .D(_0033_),
    .Q_N(_1002_),
    .Q(\mem[131] ));
 sg13g2_dfrbp_1 _2166_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net215),
    .D(_0034_),
    .Q_N(_1001_),
    .Q(\mem[179] ));
 sg13g2_dfrbp_1 _2167_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net214),
    .D(_0035_),
    .Q_N(_1000_),
    .Q(\mem[212] ));
 sg13g2_dfrbp_1 _2168_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net213),
    .D(_0036_),
    .Q_N(_0999_),
    .Q(\mem[79] ));
 sg13g2_dfrbp_1 _2169_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net212),
    .D(_0037_),
    .Q_N(_0998_),
    .Q(\mem[133] ));
 sg13g2_dfrbp_1 _2170_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net211),
    .D(_0038_),
    .Q_N(_0997_),
    .Q(\mem[132] ));
 sg13g2_dfrbp_1 _2171_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net210),
    .D(_0039_),
    .Q_N(_0996_),
    .Q(\mem[130] ));
 sg13g2_dfrbp_1 _2172_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net209),
    .D(_0040_),
    .Q_N(_0995_),
    .Q(\mem[127] ));
 sg13g2_dfrbp_1 _2173_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net208),
    .D(_0041_),
    .Q_N(_0994_),
    .Q(\mem[192] ));
 sg13g2_dfrbp_1 _2174_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net207),
    .D(_0042_),
    .Q_N(_0993_),
    .Q(\mem[181] ));
 sg13g2_dfrbp_1 _2175_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net206),
    .D(_0043_),
    .Q_N(_0992_),
    .Q(\mem[128] ));
 sg13g2_dfrbp_1 _2176_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net189),
    .D(_0044_),
    .Q_N(_0991_),
    .Q(\mem[126] ));
 sg13g2_dfrbp_1 _2177_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net188),
    .D(_0045_),
    .Q_N(_0990_),
    .Q(\mem[123] ));
 sg13g2_dfrbp_1 _2178_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net187),
    .D(_0046_),
    .Q_N(_0989_),
    .Q(\mem[125] ));
 sg13g2_dfrbp_1 _2179_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net186),
    .D(_0047_),
    .Q_N(_0988_),
    .Q(\mem[89] ));
 sg13g2_dfrbp_1 _2180_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net185),
    .D(_0048_),
    .Q_N(_0987_),
    .Q(\mem[124] ));
 sg13g2_dfrbp_1 _2181_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net184),
    .D(_0049_),
    .Q_N(_0986_),
    .Q(\mem[122] ));
 sg13g2_dfrbp_1 _2182_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net183),
    .D(_0050_),
    .Q_N(_0985_),
    .Q(\mem[190] ));
 sg13g2_dfrbp_1 _2183_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net182),
    .D(_0051_),
    .Q_N(_0984_),
    .Q(\mem[199] ));
 sg13g2_dfrbp_1 _2184_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net181),
    .D(_0052_),
    .Q_N(_0983_),
    .Q(\mem[208] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net180),
    .D(_0053_),
    .Q_N(_0982_),
    .Q(\mem[121] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net179),
    .D(_0054_),
    .Q_N(_0981_),
    .Q(\mem[180] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net178),
    .D(_0055_),
    .Q_N(_0980_),
    .Q(\mem[120] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net177),
    .D(_0056_),
    .Q_N(_0979_),
    .Q(\mem[213] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net176),
    .D(_0057_),
    .Q_N(_0978_),
    .Q(\mem[98] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net173),
    .D(_0058_),
    .Q_N(_0977_),
    .Q(\mem[218] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net171),
    .D(_0059_),
    .Q_N(_0976_),
    .Q(\mem[118] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net170),
    .D(_0060_),
    .Q_N(_0975_),
    .Q(\mem[115] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net169),
    .D(_0061_),
    .Q_N(_0974_),
    .Q(\mem[249] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net167),
    .D(_0062_),
    .Q_N(_0973_),
    .Q(\mem[117] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net166),
    .D(_0063_),
    .Q_N(_0972_),
    .Q(\mem[116] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net165),
    .D(_0064_),
    .Q_N(_0971_),
    .Q(\mem[187] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net164),
    .D(_0065_),
    .Q_N(_0970_),
    .Q(\mem[114] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net163),
    .D(_0066_),
    .Q_N(_0969_),
    .Q(\mem[111] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net162),
    .D(_0067_),
    .Q_N(_0968_),
    .Q(\mem[109] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net161),
    .D(_0068_),
    .Q_N(_0967_),
    .Q(\mem[206] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net160),
    .D(_0069_),
    .Q_N(_0966_),
    .Q(\mem[113] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net159),
    .D(_0070_),
    .Q_N(_0965_),
    .Q(\mem[112] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net158),
    .D(_0071_),
    .Q_N(_0964_),
    .Q(\mem[110] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net157),
    .D(_0072_),
    .Q_N(_0963_),
    .Q(\mem[138] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net156),
    .D(_0073_),
    .Q_N(_0962_),
    .Q(\mem[107] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net155),
    .D(_0074_),
    .Q_N(_0961_),
    .Q(\mem[108] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net154),
    .D(_0075_),
    .Q_N(_0960_),
    .Q(\mem[175] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net153),
    .D(_0076_),
    .Q_N(_0959_),
    .Q(\mem[106] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net152),
    .D(_0077_),
    .Q_N(_0958_),
    .Q(\mem[203] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net151),
    .D(_0078_),
    .Q_N(_0957_),
    .Q(\mem[103] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net150),
    .D(_0079_),
    .Q_N(_0956_),
    .Q(\mem[211] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net149),
    .D(_0080_),
    .Q_N(_0955_),
    .Q(\mem[105] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net148),
    .D(_0081_),
    .Q_N(_0954_),
    .Q(\mem[119] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net147),
    .D(_0082_),
    .Q_N(_0953_),
    .Q(\mem[104] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_0083_),
    .Q_N(_0952_),
    .Q(\mem[102] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net145),
    .D(_0084_),
    .Q_N(_0951_),
    .Q(\mem[177] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net144),
    .D(_0085_),
    .Q_N(_0950_),
    .Q(\mem[101] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net143),
    .D(_0086_),
    .Q_N(_0949_),
    .Q(\mem[198] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net142),
    .D(_0087_),
    .Q_N(_0948_),
    .Q(\mem[188] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net141),
    .D(_0088_),
    .Q_N(_0947_),
    .Q(\mem[100] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net140),
    .D(_0089_),
    .Q_N(_0946_),
    .Q(\mem[129] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net139),
    .D(_0090_),
    .Q_N(_0945_),
    .Q(\mem[205] ));
 sg13g2_dfrbp_1 _2223_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net138),
    .D(_0091_),
    .Q_N(_0944_),
    .Q(\mem[95] ));
 sg13g2_dfrbp_1 _2224_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net137),
    .D(_0092_),
    .Q_N(_0943_),
    .Q(\mem[97] ));
 sg13g2_dfrbp_1 _2225_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net136),
    .D(_0093_),
    .Q_N(_0942_),
    .Q(\mem[96] ));
 sg13g2_dfrbp_1 _2226_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net135),
    .D(_0094_),
    .Q_N(_0941_),
    .Q(\mem[149] ));
 sg13g2_dfrbp_1 _2227_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net134),
    .D(_0095_),
    .Q_N(_0940_),
    .Q(\mem[186] ));
 sg13g2_dfrbp_1 _2228_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net133),
    .D(_0096_),
    .Q_N(_0939_),
    .Q(\mem[189] ));
 sg13g2_dfrbp_1 _2229_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net132),
    .D(_0097_),
    .Q_N(_0938_),
    .Q(\mem[94] ));
 sg13g2_dfrbp_1 _2230_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0098_),
    .Q_N(_0937_),
    .Q(\mem[239] ));
 sg13g2_dfrbp_1 _2231_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net130),
    .D(_0099_),
    .Q_N(_0936_),
    .Q(\mem[183] ));
 sg13g2_dfrbp_1 _2232_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net129),
    .D(_0100_),
    .Q_N(_0935_),
    .Q(\mem[159] ));
 sg13g2_dfrbp_1 _2233_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net128),
    .D(_0101_),
    .Q_N(_0934_),
    .Q(\mem[91] ));
 sg13g2_dfrbp_1 _2234_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net127),
    .D(_0102_),
    .Q_N(_0933_),
    .Q(\mem[185] ));
 sg13g2_dfrbp_1 _2235_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net126),
    .D(_0103_),
    .Q_N(_0932_),
    .Q(\mem[169] ));
 sg13g2_dfrbp_1 _2236_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net125),
    .D(_0104_),
    .Q_N(_0931_),
    .Q(\mem[93] ));
 sg13g2_dfrbp_1 _2237_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net124),
    .D(_0105_),
    .Q_N(_0930_),
    .Q(\mem[182] ));
 sg13g2_dfrbp_1 _2238_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net123),
    .D(_0106_),
    .Q_N(_0929_),
    .Q(\mem[92] ));
 sg13g2_dfrbp_1 _2239_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net122),
    .D(_0107_),
    .Q_N(_0928_),
    .Q(\mem[90] ));
 sg13g2_dfrbp_1 _2240_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net121),
    .D(_0108_),
    .Q_N(_0927_),
    .Q(\mem[87] ));
 sg13g2_dfrbp_1 _2241_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net120),
    .D(_0109_),
    .Q_N(_0926_),
    .Q(\mem[204] ));
 sg13g2_dfrbp_1 _2242_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net119),
    .D(_0110_),
    .Q_N(_0925_),
    .Q(\mem[88] ));
 sg13g2_dfrbp_1 _2243_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net118),
    .D(_0111_),
    .Q_N(_0924_),
    .Q(\mem[86] ));
 sg13g2_dfrbp_1 _2244_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net117),
    .D(_0112_),
    .Q_N(_0923_),
    .Q(\mem[83] ));
 sg13g2_dfrbp_1 _2245_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net116),
    .D(_0113_),
    .Q_N(_0922_),
    .Q(\mem[202] ));
 sg13g2_dfrbp_1 _2246_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net115),
    .D(_0114_),
    .Q_N(_0921_),
    .Q(\mem[85] ));
 sg13g2_dfrbp_1 _2247_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net114),
    .D(_0115_),
    .Q_N(_0920_),
    .Q(\mem[84] ));
 sg13g2_dfrbp_1 _2248_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net113),
    .D(_0116_),
    .Q_N(_0919_),
    .Q(\mem[82] ));
 sg13g2_dfrbp_1 _2249_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net112),
    .D(_0117_),
    .Q_N(_0918_),
    .Q(\mem[81] ));
 sg13g2_dfrbp_1 _2250_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net111),
    .D(_0118_),
    .Q_N(_0917_),
    .Q(\mem[80] ));
 sg13g2_dfrbp_1 _2251_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net110),
    .D(_0119_),
    .Q_N(_0916_),
    .Q(\mem[78] ));
 sg13g2_dfrbp_1 _2252_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net109),
    .D(_0120_),
    .Q_N(_0915_),
    .Q(\mem[75] ));
 sg13g2_dfrbp_1 _2253_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net108),
    .D(_0121_),
    .Q_N(_0914_),
    .Q(\mem[201] ));
 sg13g2_dfrbp_1 _2254_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net107),
    .D(_0122_),
    .Q_N(_0913_),
    .Q(\mem[77] ));
 sg13g2_dfrbp_1 _2255_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net106),
    .D(_0123_),
    .Q_N(_0912_),
    .Q(\mem[76] ));
 sg13g2_dfrbp_1 _2256_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net105),
    .D(_0124_),
    .Q_N(_0911_),
    .Q(\mem[200] ));
 sg13g2_dfrbp_1 _2257_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net104),
    .D(_0125_),
    .Q_N(_0910_),
    .Q(\mem[74] ));
 sg13g2_dfrbp_1 _2258_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net103),
    .D(_0126_),
    .Q_N(_0909_),
    .Q(\mem[71] ));
 sg13g2_dfrbp_1 _2259_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net102),
    .D(_0127_),
    .Q_N(_0908_),
    .Q(\mem[73] ));
 sg13g2_dfrbp_1 _2260_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net101),
    .D(_0128_),
    .Q_N(_0907_),
    .Q(\mem[72] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net100),
    .D(_0129_),
    .Q_N(_0906_),
    .Q(\mem[70] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net99),
    .D(_0130_),
    .Q_N(_0905_),
    .Q(\mem[67] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net98),
    .D(_0131_),
    .Q_N(_0904_),
    .Q(\mem[68] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net97),
    .D(_0132_),
    .Q_N(_0903_),
    .Q(\mem[195] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net96),
    .D(_0133_),
    .Q_N(_0902_),
    .Q(\mem[66] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net95),
    .D(_0134_),
    .Q_N(_0901_),
    .Q(\mem[65] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net94),
    .D(_0135_),
    .Q_N(_0900_),
    .Q(\mem[64] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net93),
    .D(_0136_),
    .Q_N(_0899_),
    .Q(\mem[197] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net92),
    .D(_0137_),
    .Q_N(_0898_),
    .Q(\mem[184] ));
 sg13g2_dllrq_1 _2270_ (.D(net584),
    .GATE_N(net1),
    .RESET_B(net168),
    .Q(addrhi));
 sg13g2_dfrbp_1 _2271_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net91),
    .D(_0138_),
    .Q_N(_0897_),
    .Q(\mem[196] ));
 sg13g2_dllrq_1 _2272_ (.D(net577),
    .GATE_N(net1),
    .RESET_B(net172),
    .Q(read_buffer_a));
 sg13g2_dfrbp_1 _2273_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net90),
    .D(_0139_),
    .Q_N(_0896_),
    .Q(\mem[176] ));
 sg13g2_dllrq_1 _2274_ (.D(net9),
    .GATE_N(net1),
    .RESET_B(net174),
    .Q(read_buffer_b));
 sg13g2_dllrq_1 _2275_ (.D(net10),
    .GATE_N(net1),
    .RESET_B(net175),
    .Q(write_through));
 sg13g2_dfrbp_1 _2276_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net89),
    .D(_0140_),
    .Q_N(_0895_),
    .Q(\mem[174] ));
 sg13g2_dfrbp_1 _2277_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net88),
    .D(_0141_),
    .Q_N(_0894_),
    .Q(\mem[171] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net87),
    .D(_0142_),
    .Q_N(_0893_),
    .Q(\mem[173] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net86),
    .D(_0143_),
    .Q_N(_0892_),
    .Q(\mem[172] ));
 sg13g2_dfrbp_1 _2280_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net85),
    .D(_0144_),
    .Q_N(_0891_),
    .Q(\mem[170] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net84),
    .D(_0145_),
    .Q_N(_0890_),
    .Q(\mem[167] ));
 sg13g2_dfrbp_1 _2282_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net83),
    .D(_0146_),
    .Q_N(_0889_),
    .Q(\mem[168] ));
 sg13g2_dfrbp_1 _2283_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net82),
    .D(_0147_),
    .Q_N(_0888_),
    .Q(\mem[166] ));
 sg13g2_dfrbp_1 _2284_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net81),
    .D(_0148_),
    .Q_N(_0887_),
    .Q(\mem[163] ));
 sg13g2_dfrbp_1 _2285_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net80),
    .D(_0149_),
    .Q_N(_0886_),
    .Q(\mem[165] ));
 sg13g2_dfrbp_1 _2286_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net79),
    .D(_0150_),
    .Q_N(_0885_),
    .Q(\mem[164] ));
 sg13g2_dfrbp_1 _2287_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net78),
    .D(_0151_),
    .Q_N(_0884_),
    .Q(\mem[162] ));
 sg13g2_dfrbp_1 _2288_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net77),
    .D(_0152_),
    .Q_N(_0883_),
    .Q(\mem[161] ));
 sg13g2_dfrbp_1 _2289_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net191),
    .D(_0153_),
    .Q_N(_1036_),
    .Q(\mem[160] ));
 sg13g2_dfrbp_1 _2290_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net192),
    .D(\rdata_curr_b[0] ),
    .Q_N(_1037_),
    .Q(\rdata_buff_b[0] ));
 sg13g2_dfrbp_1 _2291_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net193),
    .D(\rdata_curr_b[1] ),
    .Q_N(_1038_),
    .Q(\rdata_buff_b[1] ));
 sg13g2_dfrbp_1 _2292_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net194),
    .D(\rdata_curr_b[2] ),
    .Q_N(_1039_),
    .Q(\rdata_buff_b[2] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net195),
    .D(\rdata_curr_b[3] ),
    .Q_N(_1040_),
    .Q(\rdata_buff_b[3] ));
 sg13g2_dfrbp_1 _2294_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net196),
    .D(\rdata_curr_b[4] ),
    .Q_N(_1041_),
    .Q(\rdata_buff_b[4] ));
 sg13g2_dfrbp_1 _2295_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net197),
    .D(\rdata_curr_b[5] ),
    .Q_N(_1042_),
    .Q(\rdata_buff_b[5] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net198),
    .D(\rdata_curr_b[6] ),
    .Q_N(_1043_),
    .Q(\rdata_buff_b[6] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net199),
    .D(\rdata_curr_b[7] ),
    .Q_N(_1044_),
    .Q(\rdata_buff_b[7] ));
 sg13g2_dfrbp_1 _2298_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net200),
    .D(\rdata_curr_a[0] ),
    .Q_N(_1045_),
    .Q(\rdata_buff_a[0] ));
 sg13g2_dfrbp_1 _2299_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net201),
    .D(\rdata_curr_a[1] ),
    .Q_N(_1046_),
    .Q(\rdata_buff_a[1] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net202),
    .D(\rdata_curr_a[2] ),
    .Q_N(_1047_),
    .Q(\rdata_buff_a[2] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net203),
    .D(\rdata_curr_a[3] ),
    .Q_N(_1048_),
    .Q(\rdata_buff_a[3] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net204),
    .D(\rdata_curr_a[4] ),
    .Q_N(_1049_),
    .Q(\rdata_buff_a[4] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net205),
    .D(\rdata_curr_a[5] ),
    .Q_N(_1050_),
    .Q(\rdata_buff_a[5] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net37),
    .D(\rdata_curr_a[6] ),
    .Q_N(_1051_),
    .Q(\rdata_buff_a[6] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net76),
    .D(\rdata_curr_a[7] ),
    .Q_N(_0882_),
    .Q(\rdata_buff_a[7] ));
 sg13g2_dfrbp_1 _2306_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net75),
    .D(_0154_),
    .Q_N(_0881_),
    .Q(\mem[69] ));
 sg13g2_dfrbp_1 _2307_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net74),
    .D(_0155_),
    .Q_N(_0880_),
    .Q(\mem[214] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net73),
    .D(_0156_),
    .Q_N(_0879_),
    .Q(\mem[216] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net72),
    .D(_0157_),
    .Q_N(_0878_),
    .Q(\mem[217] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net71),
    .D(_0158_),
    .Q_N(_0877_),
    .Q(\mem[215] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net70),
    .D(_0159_),
    .Q_N(_0876_),
    .Q(\mem[220] ));
 sg13g2_dfrbp_1 _2312_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net69),
    .D(_0160_),
    .Q_N(_0875_),
    .Q(\mem[221] ));
 sg13g2_dfrbp_1 _2313_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net68),
    .D(_0161_),
    .Q_N(_0874_),
    .Q(\mem[219] ));
 sg13g2_dfrbp_1 _2314_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net67),
    .D(_0162_),
    .Q_N(_0873_),
    .Q(\mem[222] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net66),
    .D(_0163_),
    .Q_N(_0872_),
    .Q(\mem[224] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net65),
    .D(_0164_),
    .Q_N(_0871_),
    .Q(\mem[225] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net64),
    .D(_0165_),
    .Q_N(_0870_),
    .Q(\mem[223] ));
 sg13g2_dfrbp_1 _2318_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net63),
    .D(_0166_),
    .Q_N(_0869_),
    .Q(\mem[226] ));
 sg13g2_dfrbp_1 _2319_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net62),
    .D(_0167_),
    .Q_N(_0868_),
    .Q(\mem[228] ));
 sg13g2_dfrbp_1 _2320_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net61),
    .D(_0168_),
    .Q_N(_0867_),
    .Q(\mem[227] ));
 sg13g2_dfrbp_1 _2321_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net60),
    .D(_0169_),
    .Q_N(_0866_),
    .Q(\mem[230] ));
 sg13g2_dfrbp_1 _2322_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net59),
    .D(_0170_),
    .Q_N(_0865_),
    .Q(\mem[232] ));
 sg13g2_dfrbp_1 _2323_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net58),
    .D(_0171_),
    .Q_N(_0864_),
    .Q(\mem[233] ));
 sg13g2_dfrbp_1 _2324_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net57),
    .D(_0172_),
    .Q_N(_0863_),
    .Q(\mem[231] ));
 sg13g2_dfrbp_1 _2325_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net56),
    .D(_0173_),
    .Q_N(_0862_),
    .Q(\mem[234] ));
 sg13g2_dfrbp_1 _2326_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net55),
    .D(_0174_),
    .Q_N(_0861_),
    .Q(\mem[236] ));
 sg13g2_dfrbp_1 _2327_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net54),
    .D(_0175_),
    .Q_N(_0860_),
    .Q(\mem[237] ));
 sg13g2_dfrbp_1 _2328_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net53),
    .D(_0176_),
    .Q_N(_0859_),
    .Q(\mem[235] ));
 sg13g2_dfrbp_1 _2329_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net52),
    .D(_0177_),
    .Q_N(_0858_),
    .Q(\mem[238] ));
 sg13g2_dfrbp_1 _2330_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net51),
    .D(_0178_),
    .Q_N(_0857_),
    .Q(\mem[240] ));
 sg13g2_dfrbp_1 _2331_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net50),
    .D(_0179_),
    .Q_N(_0856_),
    .Q(\mem[241] ));
 sg13g2_dfrbp_1 _2332_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net49),
    .D(_0180_),
    .Q_N(_0855_),
    .Q(\mem[242] ));
 sg13g2_dfrbp_1 _2333_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net48),
    .D(_0181_),
    .Q_N(_0854_),
    .Q(\mem[244] ));
 sg13g2_dfrbp_1 _2334_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net47),
    .D(_0182_),
    .Q_N(_0853_),
    .Q(\mem[245] ));
 sg13g2_dfrbp_1 _2335_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net46),
    .D(_0183_),
    .Q_N(_0852_),
    .Q(\mem[243] ));
 sg13g2_dfrbp_1 _2336_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net45),
    .D(_0184_),
    .Q_N(_0851_),
    .Q(\mem[246] ));
 sg13g2_dfrbp_1 _2337_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net44),
    .D(_0185_),
    .Q_N(_0850_),
    .Q(\mem[248] ));
 sg13g2_dfrbp_1 _2338_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net43),
    .D(_0186_),
    .Q_N(_0849_),
    .Q(\mem[247] ));
 sg13g2_dfrbp_1 _2339_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net42),
    .D(_0187_),
    .Q_N(_0848_),
    .Q(\mem[250] ));
 sg13g2_dfrbp_1 _2340_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net41),
    .D(_0188_),
    .Q_N(_0847_),
    .Q(\mem[252] ));
 sg13g2_dfrbp_1 _2341_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net40),
    .D(_0189_),
    .Q_N(_0846_),
    .Q(\mem[253] ));
 sg13g2_dfrbp_1 _2342_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net39),
    .D(_0190_),
    .Q_N(_0845_),
    .Q(\mem[251] ));
 sg13g2_dfrbp_1 _2343_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net38),
    .D(_0191_),
    .Q_N(_0844_),
    .Q(\mem[99] ));
 sg13g2_tiehi _2140__29 (.L_HI(net29));
 sg13g2_tiehi _2139__30 (.L_HI(net30));
 sg13g2_tiehi _2138__31 (.L_HI(net31));
 sg13g2_tiehi _2137__32 (.L_HI(net32));
 sg13g2_tiehi _2136__33 (.L_HI(net33));
 sg13g2_tiehi _2135__34 (.L_HI(net34));
 sg13g2_tiehi _2134__35 (.L_HI(net35));
 sg13g2_tiehi _2133__36 (.L_HI(net36));
 sg13g2_tiehi _2304__37 (.L_HI(net37));
 sg13g2_tiehi _2343__38 (.L_HI(net38));
 sg13g2_tiehi _2342__39 (.L_HI(net39));
 sg13g2_tiehi _2341__40 (.L_HI(net40));
 sg13g2_tiehi _2340__41 (.L_HI(net41));
 sg13g2_tiehi _2339__42 (.L_HI(net42));
 sg13g2_tiehi _2338__43 (.L_HI(net43));
 sg13g2_tiehi _2337__44 (.L_HI(net44));
 sg13g2_tiehi _2336__45 (.L_HI(net45));
 sg13g2_tiehi _2335__46 (.L_HI(net46));
 sg13g2_tiehi _2334__47 (.L_HI(net47));
 sg13g2_tiehi _2333__48 (.L_HI(net48));
 sg13g2_tiehi _2332__49 (.L_HI(net49));
 sg13g2_tiehi _2331__50 (.L_HI(net50));
 sg13g2_tiehi _2330__51 (.L_HI(net51));
 sg13g2_tiehi _2329__52 (.L_HI(net52));
 sg13g2_tiehi _2328__53 (.L_HI(net53));
 sg13g2_tiehi _2327__54 (.L_HI(net54));
 sg13g2_tiehi _2326__55 (.L_HI(net55));
 sg13g2_tiehi _2325__56 (.L_HI(net56));
 sg13g2_tiehi _2324__57 (.L_HI(net57));
 sg13g2_tiehi _2323__58 (.L_HI(net58));
 sg13g2_tiehi _2322__59 (.L_HI(net59));
 sg13g2_tiehi _2321__60 (.L_HI(net60));
 sg13g2_tiehi _2320__61 (.L_HI(net61));
 sg13g2_tiehi _2319__62 (.L_HI(net62));
 sg13g2_tiehi _2318__63 (.L_HI(net63));
 sg13g2_tiehi _2317__64 (.L_HI(net64));
 sg13g2_tiehi _2316__65 (.L_HI(net65));
 sg13g2_tiehi _2315__66 (.L_HI(net66));
 sg13g2_tiehi _2314__67 (.L_HI(net67));
 sg13g2_tiehi _2313__68 (.L_HI(net68));
 sg13g2_tiehi _2312__69 (.L_HI(net69));
 sg13g2_tiehi _2311__70 (.L_HI(net70));
 sg13g2_tiehi _2310__71 (.L_HI(net71));
 sg13g2_tiehi _2309__72 (.L_HI(net72));
 sg13g2_tiehi _2308__73 (.L_HI(net73));
 sg13g2_tiehi _2307__74 (.L_HI(net74));
 sg13g2_tiehi _2306__75 (.L_HI(net75));
 sg13g2_tiehi _2305__76 (.L_HI(net76));
 sg13g2_tiehi _2288__77 (.L_HI(net77));
 sg13g2_tiehi _2287__78 (.L_HI(net78));
 sg13g2_tiehi _2286__79 (.L_HI(net79));
 sg13g2_tiehi _2285__80 (.L_HI(net80));
 sg13g2_tiehi _2284__81 (.L_HI(net81));
 sg13g2_tiehi _2283__82 (.L_HI(net82));
 sg13g2_tiehi _2282__83 (.L_HI(net83));
 sg13g2_tiehi _2281__84 (.L_HI(net84));
 sg13g2_tiehi _2280__85 (.L_HI(net85));
 sg13g2_tiehi _2279__86 (.L_HI(net86));
 sg13g2_tiehi _2278__87 (.L_HI(net87));
 sg13g2_tiehi _2277__88 (.L_HI(net88));
 sg13g2_tiehi _2276__89 (.L_HI(net89));
 sg13g2_tiehi _2273__90 (.L_HI(net90));
 sg13g2_tiehi _2271__91 (.L_HI(net91));
 sg13g2_tiehi _2269__92 (.L_HI(net92));
 sg13g2_tiehi _2268__93 (.L_HI(net93));
 sg13g2_tiehi _2267__94 (.L_HI(net94));
 sg13g2_tiehi _2266__95 (.L_HI(net95));
 sg13g2_tiehi _2265__96 (.L_HI(net96));
 sg13g2_tiehi _2264__97 (.L_HI(net97));
 sg13g2_tiehi _2263__98 (.L_HI(net98));
 sg13g2_tiehi _2262__99 (.L_HI(net99));
 sg13g2_tiehi _2261__100 (.L_HI(net100));
 sg13g2_tiehi _2260__101 (.L_HI(net101));
 sg13g2_tiehi _2259__102 (.L_HI(net102));
 sg13g2_tiehi _2258__103 (.L_HI(net103));
 sg13g2_tiehi _2257__104 (.L_HI(net104));
 sg13g2_tiehi _2256__105 (.L_HI(net105));
 sg13g2_tiehi _2255__106 (.L_HI(net106));
 sg13g2_tiehi _2254__107 (.L_HI(net107));
 sg13g2_tiehi _2253__108 (.L_HI(net108));
 sg13g2_tiehi _2252__109 (.L_HI(net109));
 sg13g2_tiehi _2251__110 (.L_HI(net110));
 sg13g2_tiehi _2250__111 (.L_HI(net111));
 sg13g2_tiehi _2249__112 (.L_HI(net112));
 sg13g2_tiehi _2248__113 (.L_HI(net113));
 sg13g2_tiehi _2247__114 (.L_HI(net114));
 sg13g2_tiehi _2246__115 (.L_HI(net115));
 sg13g2_tiehi _2245__116 (.L_HI(net116));
 sg13g2_tiehi _2244__117 (.L_HI(net117));
 sg13g2_tiehi _2243__118 (.L_HI(net118));
 sg13g2_tiehi _2242__119 (.L_HI(net119));
 sg13g2_tiehi _2241__120 (.L_HI(net120));
 sg13g2_tiehi _2240__121 (.L_HI(net121));
 sg13g2_tiehi _2239__122 (.L_HI(net122));
 sg13g2_tiehi _2238__123 (.L_HI(net123));
 sg13g2_tiehi _2237__124 (.L_HI(net124));
 sg13g2_tiehi _2236__125 (.L_HI(net125));
 sg13g2_tiehi _2235__126 (.L_HI(net126));
 sg13g2_tiehi _2234__127 (.L_HI(net127));
 sg13g2_tiehi _2233__128 (.L_HI(net128));
 sg13g2_tiehi _2232__129 (.L_HI(net129));
 sg13g2_tiehi _2231__130 (.L_HI(net130));
 sg13g2_tiehi _2230__131 (.L_HI(net131));
 sg13g2_tiehi _2229__132 (.L_HI(net132));
 sg13g2_tiehi _2228__133 (.L_HI(net133));
 sg13g2_tiehi _2227__134 (.L_HI(net134));
 sg13g2_tiehi _2226__135 (.L_HI(net135));
 sg13g2_tiehi _2225__136 (.L_HI(net136));
 sg13g2_tiehi _2224__137 (.L_HI(net137));
 sg13g2_tiehi _2223__138 (.L_HI(net138));
 sg13g2_tiehi _2222__139 (.L_HI(net139));
 sg13g2_tiehi _2221__140 (.L_HI(net140));
 sg13g2_tiehi _2220__141 (.L_HI(net141));
 sg13g2_tiehi _2219__142 (.L_HI(net142));
 sg13g2_tiehi _2218__143 (.L_HI(net143));
 sg13g2_tiehi _2217__144 (.L_HI(net144));
 sg13g2_tiehi _2216__145 (.L_HI(net145));
 sg13g2_tiehi _2215__146 (.L_HI(net146));
 sg13g2_tiehi _2214__147 (.L_HI(net147));
 sg13g2_tiehi _2213__148 (.L_HI(net148));
 sg13g2_tiehi _2212__149 (.L_HI(net149));
 sg13g2_tiehi _2211__150 (.L_HI(net150));
 sg13g2_tiehi _2210__151 (.L_HI(net151));
 sg13g2_tiehi _2209__152 (.L_HI(net152));
 sg13g2_tiehi _2208__153 (.L_HI(net153));
 sg13g2_tiehi _2207__154 (.L_HI(net154));
 sg13g2_tiehi _2206__155 (.L_HI(net155));
 sg13g2_tiehi _2205__156 (.L_HI(net156));
 sg13g2_tiehi _2204__157 (.L_HI(net157));
 sg13g2_tiehi _2203__158 (.L_HI(net158));
 sg13g2_tiehi _2202__159 (.L_HI(net159));
 sg13g2_tiehi _2201__160 (.L_HI(net160));
 sg13g2_tiehi _2200__161 (.L_HI(net161));
 sg13g2_tiehi _2199__162 (.L_HI(net162));
 sg13g2_tiehi _2198__163 (.L_HI(net163));
 sg13g2_tiehi _2197__164 (.L_HI(net164));
 sg13g2_tiehi _2196__165 (.L_HI(net165));
 sg13g2_tiehi _2195__166 (.L_HI(net166));
 sg13g2_tiehi _2194__167 (.L_HI(net167));
 sg13g2_tiehi _2270__168 (.L_HI(net168));
 sg13g2_tiehi _2193__169 (.L_HI(net169));
 sg13g2_tiehi _2192__170 (.L_HI(net170));
 sg13g2_tiehi _2191__171 (.L_HI(net171));
 sg13g2_tiehi _2272__172 (.L_HI(net172));
 sg13g2_tiehi _2190__173 (.L_HI(net173));
 sg13g2_tiehi _2274__174 (.L_HI(net174));
 sg13g2_tiehi _2275__175 (.L_HI(net175));
 sg13g2_tiehi _2189__176 (.L_HI(net176));
 sg13g2_tiehi _2188__177 (.L_HI(net177));
 sg13g2_tiehi _2187__178 (.L_HI(net178));
 sg13g2_tiehi _2186__179 (.L_HI(net179));
 sg13g2_tiehi _2185__180 (.L_HI(net180));
 sg13g2_tiehi _2184__181 (.L_HI(net181));
 sg13g2_tiehi _2183__182 (.L_HI(net182));
 sg13g2_tiehi _2182__183 (.L_HI(net183));
 sg13g2_tiehi _2181__184 (.L_HI(net184));
 sg13g2_tiehi _2180__185 (.L_HI(net185));
 sg13g2_tiehi _2179__186 (.L_HI(net186));
 sg13g2_tiehi _2178__187 (.L_HI(net187));
 sg13g2_tiehi _2177__188 (.L_HI(net188));
 sg13g2_tiehi _2176__189 (.L_HI(net189));
 sg13g2_tiehi _2132__190 (.L_HI(net190));
 sg13g2_tiehi _2289__191 (.L_HI(net191));
 sg13g2_tiehi _2290__192 (.L_HI(net192));
 sg13g2_tiehi _2291__193 (.L_HI(net193));
 sg13g2_tiehi _2292__194 (.L_HI(net194));
 sg13g2_tiehi _2293__195 (.L_HI(net195));
 sg13g2_tiehi _2294__196 (.L_HI(net196));
 sg13g2_tiehi _2295__197 (.L_HI(net197));
 sg13g2_tiehi _2296__198 (.L_HI(net198));
 sg13g2_tiehi _2297__199 (.L_HI(net199));
 sg13g2_tiehi _2298__200 (.L_HI(net200));
 sg13g2_tiehi _2299__201 (.L_HI(net201));
 sg13g2_tiehi _2300__202 (.L_HI(net202));
 sg13g2_tiehi _2301__203 (.L_HI(net203));
 sg13g2_tiehi _2302__204 (.L_HI(net204));
 sg13g2_tiehi _2303__205 (.L_HI(net205));
 sg13g2_tiehi _2175__206 (.L_HI(net206));
 sg13g2_tiehi _2174__207 (.L_HI(net207));
 sg13g2_tiehi _2173__208 (.L_HI(net208));
 sg13g2_tiehi _2172__209 (.L_HI(net209));
 sg13g2_tiehi _2171__210 (.L_HI(net210));
 sg13g2_tiehi _2170__211 (.L_HI(net211));
 sg13g2_tiehi _2169__212 (.L_HI(net212));
 sg13g2_tiehi _2168__213 (.L_HI(net213));
 sg13g2_tiehi _2167__214 (.L_HI(net214));
 sg13g2_tiehi _2166__215 (.L_HI(net215));
 sg13g2_tiehi _2165__216 (.L_HI(net216));
 sg13g2_tiehi _2164__217 (.L_HI(net217));
 sg13g2_tiehi _2163__218 (.L_HI(net218));
 sg13g2_tiehi _2162__219 (.L_HI(net219));
 sg13g2_tiehi _2161__220 (.L_HI(net220));
 sg13g2_tiehi _2160__221 (.L_HI(net221));
 sg13g2_tiehi _2159__222 (.L_HI(net222));
 sg13g2_tiehi _2158__223 (.L_HI(net223));
 sg13g2_tiehi _2157__224 (.L_HI(net224));
 sg13g2_tiehi _2156__225 (.L_HI(net225));
 sg13g2_tiehi _2155__226 (.L_HI(net226));
 sg13g2_tiehi _2154__227 (.L_HI(net227));
 sg13g2_tiehi _2153__228 (.L_HI(net228));
 sg13g2_tiehi _2152__229 (.L_HI(net229));
 sg13g2_tiehi _2151__230 (.L_HI(net230));
 sg13g2_tiehi _2150__231 (.L_HI(net231));
 sg13g2_tiehi _2149__232 (.L_HI(net232));
 sg13g2_tiehi _2148__233 (.L_HI(net233));
 sg13g2_tiehi _2147__234 (.L_HI(net234));
 sg13g2_tiehi _2146__235 (.L_HI(net235));
 sg13g2_tiehi _2145__236 (.L_HI(net236));
 sg13g2_tiehi _2144__237 (.L_HI(net237));
 sg13g2_tiehi _2143__238 (.L_HI(net238));
 sg13g2_tiehi _2142__239 (.L_HI(net239));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_13 (.L_LO(net13));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_14 (.L_LO(net14));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_25 (.L_LO(net25));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_26 (.L_LO(net26));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_27 (.L_LO(net27));
 sg13g2_tiehi _2141__28 (.L_HI(net28));
 sg13g2_buf_4 fanout469 (.X(net469),
    .A(_0336_));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(net474));
 sg13g2_buf_1 fanout471 (.A(net474),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(net474),
    .X(net472));
 sg13g2_buf_1 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_0785_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_0778_),
    .X(net476));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(_0778_));
 sg13g2_buf_2 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(net480));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(net482));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(net482));
 sg13g2_buf_2 fanout482 (.A(_0773_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(net485),
    .X(net483));
 sg13g2_buf_1 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_4 fanout486 (.X(net486),
    .A(net489));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(net488));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(net489));
 sg13g2_buf_2 fanout489 (.A(_0772_),
    .X(net489));
 sg13g2_buf_4 fanout490 (.X(net490),
    .A(net491));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net497));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(net497));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(net496));
 sg13g2_buf_4 fanout494 (.X(net494),
    .A(net496));
 sg13g2_buf_1 fanout495 (.A(net496),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(_0771_));
 sg13g2_buf_2 fanout498 (.A(net500),
    .X(net498));
 sg13g2_buf_1 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(_0770_));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(net507));
 sg13g2_buf_2 fanout503 (.A(net506),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(net506),
    .X(net504));
 sg13g2_buf_1 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_0770_),
    .X(net507));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(net509));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(_0529_));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(_0520_));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(net514));
 sg13g2_buf_2 fanout512 (.A(net514),
    .X(net512));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(net514));
 sg13g2_buf_2 fanout514 (.A(_0519_),
    .X(net514));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(_0515_));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(net517));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net519));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net519));
 sg13g2_buf_2 fanout519 (.A(_0514_),
    .X(net519));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(_0513_));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(net523));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net523));
 sg13g2_buf_2 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_0512_),
    .X(net524));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(net528));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(net527));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(_0510_));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(net533));
 sg13g2_buf_2 fanout531 (.A(net533),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(net533));
 sg13g2_buf_2 fanout533 (.A(net542),
    .X(net533));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(net542));
 sg13g2_buf_2 fanout535 (.A(net542),
    .X(net535));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net540));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(net540));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net540));
 sg13g2_buf_1 fanout539 (.A(net540),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net542),
    .X(net540));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(net542));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_0509_));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(_0507_));
 sg13g2_buf_2 fanout544 (.A(_0507_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net548),
    .X(net545));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(net548));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_0784_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_0781_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_0781_),
    .X(net550));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(_0527_));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net558),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(net557),
    .X(net554));
 sg13g2_buf_1 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_0505_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(net560),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_0504_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_1 fanout562 (.A(net563),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_0504_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(read_buffer_a),
    .X(net565));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(addrhi));
 sg13g2_buf_1 fanout567 (.A(addrhi),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net571),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(net571),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_0503_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_0430_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net576),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(_0430_));
 sg13g2_buf_2 fanout577 (.A(net8),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net582),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net582),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(uio_in[0]),
    .X(net582));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(uio_in[0]));
 sg13g2_buf_1 fanout584 (.A(uio_in[0]),
    .X(net584));
 sg13g2_buf_4 fanout585 (.X(net585),
    .A(net4));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net591),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(net591));
 sg13g2_buf_1 fanout591 (.A(ui_in[4]),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(net595));
 sg13g2_buf_2 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(ui_in[3]));
 sg13g2_buf_2 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(net600),
    .X(net597));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(net600));
 sg13g2_buf_2 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(ui_in[3]),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(net605),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net605),
    .X(net602));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(net605));
 sg13g2_buf_2 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(ui_in[2]),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net609),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(net609));
 sg13g2_buf_2 fanout609 (.A(ui_in[2]),
    .X(net609));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(net614));
 sg13g2_buf_2 fanout611 (.A(net614),
    .X(net611));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(net614));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(ui_in[1]),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net618),
    .X(net615));
 sg13g2_buf_4 fanout616 (.X(net616),
    .A(net618));
 sg13g2_buf_2 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_4 fanout618 (.X(net618),
    .A(ui_in[1]));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(net622));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(net622));
 sg13g2_buf_2 fanout622 (.A(ui_in[0]),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(net626),
    .X(net623));
 sg13g2_buf_1 fanout624 (.A(net626),
    .X(net624));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(net626));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(ui_in[0]));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[5]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[6]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[7]));
 sg13g2_buf_2 input5 (.A(uio_in[1]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[2]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[3]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[4]),
    .X(net8));
 sg13g2_buf_4 input9 (.X(net9),
    .A(uio_in[5]));
 sg13g2_buf_1 input10 (.A(uio_in[6]),
    .X(net10));
 sg13g2_buf_4 input11 (.X(net11),
    .A(uio_in[7]));
 sg13g2_tielo tt_um_dlmiles_dffram32x8_2r1w_12 (.L_LO(net12));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_2_3__leaf_clk));
 sg13g2_inv_2 clkload1 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_16_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mem[142] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mem[83] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mem[242] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mem[86] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mem[102] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mem[145] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mem[84] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mem[85] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mem[101] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mem[97] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mem[197] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mem[247] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mem[69] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mem[162] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mem[244] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mem[129] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mem[82] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mem[103] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mem[80] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mem[68] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mem[66] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mem[96] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mem[135] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mem[81] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mem[127] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mem[198] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mem[100] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mem[167] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mem[99] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mem[149] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mem[171] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mem[193] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mem[98] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mem[196] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mem[130] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mem[64] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mem[132] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mem[67] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mem[241] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mem[230] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mem[210] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mem[87] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mem[170] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mem[164] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mem[65] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mem[175] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mem[70] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mem[128] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mem[199] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mem[195] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mem[172] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mem[76] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mem[183] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mem[173] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mem[174] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mem[146] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mem[205] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mem[209] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mem[169] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mem[245] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mem[115] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mem[113] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mem[206] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mem[229] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mem[246] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mem[168] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mem[71] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mem[215] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mem[116] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mem[72] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mem[78] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mem[178] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mem[131] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mem[117] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mem[221] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mem[166] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mem[114] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mem[161] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mem[212] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mem[226] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mem[118] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mem[254] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mem[190] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mem[126] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mem[208] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mem[165] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mem[158] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mem[133] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mem[112] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mem[211] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mem[120] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mem[218] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mem[157] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold94 (.A(\mem[222] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mem[192] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mem[137] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mem[177] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mem[233] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold99 (.A(\mem[125] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mem[106] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mem[235] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mem[92] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mem[201] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mem[143] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mem[240] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mem[252] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mem[140] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mem[73] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mem[88] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mem[94] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mem[228] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mem[77] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mem[75] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mem[163] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mem[239] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold116 (.A(\mem[124] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mem[89] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mem[204] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mem[203] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mem[148] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold121 (.A(\mem[223] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mem[238] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mem[180] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold124 (.A(\mem[108] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mem[160] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mem[91] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mem[231] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mem[90] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mem[105] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mem[93] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mem[255] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mem[216] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mem[194] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mem[217] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mem[186] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mem[250] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mem[220] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mem[200] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mem[151] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold140 (.A(\mem[121] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mem[224] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mem[95] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mem[150] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mem[182] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold145 (.A(\mem[232] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mem[236] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mem[237] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mem[243] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mem[181] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold150 (.A(\mem[225] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mem[123] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold152 (.A(\mem[213] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mem[202] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mem[188] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mem[234] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold156 (.A(\mem[109] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mem[219] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold158 (.A(\mem[134] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mem[104] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mem[79] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold161 (.A(\mem[214] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mem[122] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold163 (.A(\mem[189] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mem[253] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold165 (.A(\mem[154] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mem[227] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold167 (.A(\mem[191] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold168 (.A(\mem[136] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold169 (.A(\mem[147] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold170 (.A(\mem[249] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold171 (.A(\mem[144] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold172 (.A(\mem[207] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mem[107] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold174 (.A(\mem[156] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mem[110] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold176 (.A(\mem[74] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mem[185] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mem[141] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mem[111] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold180 (.A(\mem[159] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mem[138] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold182 (.A(\mem[119] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mem[179] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mem[153] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold185 (.A(\mem[248] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mem[176] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mem[152] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mem[139] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold189 (.A(\mem[251] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold190 (.A(\mem[155] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mem[187] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold192 (.A(\mem[184] ),
    .X(net431));
 sg13g2_antennanp ANTENNA_1 (.A(ui_in[4]));
 sg13g2_antennanp ANTENNA_2 (.A(ui_in[4]));
 sg13g2_antennanp ANTENNA_3 (.A(ui_in[4]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_4 FILLER_2_196 ();
 sg13g2_fill_1 FILLER_2_204 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_4 FILLER_3_215 ();
 sg13g2_decap_8 FILLER_3_232 ();
 sg13g2_decap_4 FILLER_3_239 ();
 sg13g2_decap_4 FILLER_3_253 ();
 sg13g2_fill_2 FILLER_3_266 ();
 sg13g2_fill_1 FILLER_3_272 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_4 FILLER_4_182 ();
 sg13g2_fill_1 FILLER_4_186 ();
 sg13g2_fill_2 FILLER_4_237 ();
 sg13g2_fill_1 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_fill_1 FILLER_5_175 ();
 sg13g2_fill_2 FILLER_5_202 ();
 sg13g2_fill_1 FILLER_5_267 ();
 sg13g2_fill_1 FILLER_5_282 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_172 ();
 sg13g2_fill_1 FILLER_6_174 ();
 sg13g2_fill_2 FILLER_6_201 ();
 sg13g2_fill_1 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_4 FILLER_7_154 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_170 ();
 sg13g2_fill_2 FILLER_7_180 ();
 sg13g2_fill_1 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_193 ();
 sg13g2_decap_8 FILLER_7_246 ();
 sg13g2_decap_8 FILLER_7_260 ();
 sg13g2_fill_2 FILLER_7_271 ();
 sg13g2_fill_2 FILLER_7_277 ();
 sg13g2_fill_2 FILLER_7_306 ();
 sg13g2_fill_1 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_fill_2 FILLER_8_180 ();
 sg13g2_fill_1 FILLER_8_182 ();
 sg13g2_fill_1 FILLER_8_193 ();
 sg13g2_fill_2 FILLER_8_213 ();
 sg13g2_fill_1 FILLER_8_215 ();
 sg13g2_fill_2 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_233 ();
 sg13g2_decap_8 FILLER_8_240 ();
 sg13g2_fill_2 FILLER_8_247 ();
 sg13g2_decap_4 FILLER_8_275 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_294 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_fill_2 FILLER_8_305 ();
 sg13g2_fill_1 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_317 ();
 sg13g2_decap_8 FILLER_8_324 ();
 sg13g2_decap_8 FILLER_8_331 ();
 sg13g2_decap_8 FILLER_8_338 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_4 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_137 ();
 sg13g2_fill_1 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_236 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_fill_2 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_4 FILLER_9_324 ();
 sg13g2_fill_1 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_4 FILLER_10_133 ();
 sg13g2_fill_1 FILLER_10_137 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_fill_1 FILLER_10_179 ();
 sg13g2_decap_4 FILLER_10_258 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_decap_4 FILLER_11_171 ();
 sg13g2_fill_1 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_185 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_fill_2 FILLER_11_232 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_fill_1 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_344 ();
 sg13g2_decap_8 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_358 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_4 FILLER_12_133 ();
 sg13g2_fill_2 FILLER_12_137 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_213 ();
 sg13g2_decap_8 FILLER_12_219 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_fill_1 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_fill_2 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_fill_2 FILLER_14_170 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_4 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_217 ();
 sg13g2_decap_4 FILLER_14_232 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_4 FILLER_14_248 ();
 sg13g2_fill_1 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_4 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_decap_8 FILLER_15_184 ();
 sg13g2_decap_4 FILLER_15_191 ();
 sg13g2_fill_1 FILLER_15_199 ();
 sg13g2_fill_2 FILLER_15_275 ();
 sg13g2_fill_2 FILLER_15_281 ();
 sg13g2_fill_1 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_208 ();
 sg13g2_fill_2 FILLER_16_218 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_270 ();
 sg13g2_decap_4 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_4 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_237 ();
 sg13g2_fill_2 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_fill_1 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_fill_2 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_300 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_decap_4 FILLER_19_262 ();
 sg13g2_fill_1 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_272 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_decap_4 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_decap_4 FILLER_20_232 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_fill_2 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_4 FILLER_20_287 ();
 sg13g2_decap_4 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_4 FILLER_21_119 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_265 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_fill_1 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_decap_4 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_decap_4 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_fill_2 FILLER_23_150 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_decap_4 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_180 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_fill_2 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_297 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_decap_4 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_fill_2 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_126 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_decap_4 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_202 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_4 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_4 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_fill_2 FILLER_26_146 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_decap_4 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_decap_4 FILLER_26_313 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_decap_8 FILLER_27_165 ();
 sg13g2_fill_2 FILLER_27_172 ();
 sg13g2_decap_8 FILLER_27_178 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_decap_4 FILLER_27_207 ();
 sg13g2_decap_4 FILLER_27_215 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_fill_2 FILLER_27_235 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_340 ();
 sg13g2_decap_4 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_decap_4 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_157 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_4 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_fill_2 FILLER_28_282 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_332 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_4 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_decap_4 FILLER_29_170 ();
 sg13g2_fill_1 FILLER_29_174 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_246 ();
 sg13g2_fill_2 FILLER_29_262 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_166 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_184 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_206 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_decap_4 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_172 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_256 ();
 sg13g2_decap_8 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_283 ();
 sg13g2_fill_1 FILLER_31_285 ();
 sg13g2_decap_4 FILLER_31_290 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_4 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_4 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_fill_1 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_246 ();
 sg13g2_decap_8 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_260 ();
 sg13g2_decap_4 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_290 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_decap_4 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_decap_4 FILLER_32_336 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_decap_4 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_229 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_decap_4 FILLER_33_243 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_decap_4 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_fill_1 FILLER_33_300 ();
 sg13g2_decap_4 FILLER_33_306 ();
 sg13g2_fill_2 FILLER_33_323 ();
 sg13g2_fill_1 FILLER_33_325 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_decap_4 FILLER_33_346 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_2 FILLER_33_375 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_383 ();
 sg13g2_decap_8 FILLER_33_390 ();
 sg13g2_decap_8 FILLER_33_397 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_304 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_decap_4 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_171 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_295 ();
 sg13g2_fill_2 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_342 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_4 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_decap_4 FILLER_36_163 ();
 sg13g2_fill_1 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_fill_1 FILLER_36_180 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_2 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_291 ();
 sg13g2_fill_1 FILLER_36_293 ();
 sg13g2_decap_4 FILLER_36_304 ();
 sg13g2_decap_4 FILLER_36_317 ();
 sg13g2_fill_2 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_145 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_decap_4 FILLER_37_261 ();
 sg13g2_decap_4 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_fill_2 FILLER_37_318 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_fill_1 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_370 ();
 sg13g2_decap_8 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_4 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_130 ();
 sg13g2_decap_8 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_143 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_decap_4 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_267 ();
 sg13g2_decap_8 FILLER_38_274 ();
 sg13g2_decap_4 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_336 ();
 sg13g2_decap_4 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_4 FILLER_39_140 ();
 sg13g2_fill_1 FILLER_39_144 ();
 sg13g2_fill_2 FILLER_39_155 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_fill_1 FILLER_39_202 ();
 sg13g2_decap_8 FILLER_39_208 ();
 sg13g2_decap_8 FILLER_39_215 ();
 sg13g2_decap_8 FILLER_39_222 ();
 sg13g2_decap_4 FILLER_39_229 ();
 sg13g2_fill_2 FILLER_39_233 ();
 sg13g2_decap_8 FILLER_39_243 ();
 sg13g2_decap_8 FILLER_39_250 ();
 sg13g2_decap_4 FILLER_39_257 ();
 sg13g2_decap_4 FILLER_39_290 ();
 sg13g2_fill_2 FILLER_39_294 ();
 sg13g2_fill_1 FILLER_39_310 ();
 sg13g2_fill_1 FILLER_39_325 ();
 sg13g2_fill_1 FILLER_39_336 ();
 sg13g2_fill_2 FILLER_39_342 ();
 sg13g2_fill_1 FILLER_39_344 ();
 sg13g2_fill_2 FILLER_39_359 ();
 sg13g2_decap_8 FILLER_39_387 ();
 sg13g2_decap_8 FILLER_39_394 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_decap_4 FILLER_40_179 ();
 sg13g2_fill_1 FILLER_40_183 ();
 sg13g2_decap_8 FILLER_40_192 ();
 sg13g2_fill_1 FILLER_40_199 ();
 sg13g2_decap_8 FILLER_40_208 ();
 sg13g2_fill_2 FILLER_40_215 ();
 sg13g2_decap_8 FILLER_40_233 ();
 sg13g2_decap_4 FILLER_40_254 ();
 sg13g2_fill_2 FILLER_40_258 ();
 sg13g2_decap_4 FILLER_40_276 ();
 sg13g2_decap_8 FILLER_40_285 ();
 sg13g2_decap_8 FILLER_40_292 ();
 sg13g2_decap_8 FILLER_40_299 ();
 sg13g2_decap_8 FILLER_40_306 ();
 sg13g2_decap_8 FILLER_40_313 ();
 sg13g2_fill_2 FILLER_40_320 ();
 sg13g2_fill_2 FILLER_40_325 ();
 sg13g2_decap_8 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_396 ();
 sg13g2_decap_4 FILLER_40_403 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_4 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_195 ();
 sg13g2_decap_4 FILLER_41_207 ();
 sg13g2_fill_1 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_218 ();
 sg13g2_fill_1 FILLER_41_236 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_fill_1 FILLER_41_331 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_4 FILLER_42_119 ();
 sg13g2_fill_2 FILLER_42_149 ();
 sg13g2_fill_1 FILLER_42_151 ();
 sg13g2_fill_1 FILLER_42_156 ();
 sg13g2_decap_8 FILLER_42_167 ();
 sg13g2_decap_8 FILLER_42_174 ();
 sg13g2_fill_2 FILLER_42_181 ();
 sg13g2_fill_1 FILLER_42_183 ();
 sg13g2_fill_1 FILLER_42_190 ();
 sg13g2_fill_1 FILLER_42_217 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_246 ();
 sg13g2_fill_1 FILLER_42_262 ();
 sg13g2_fill_1 FILLER_42_268 ();
 sg13g2_fill_2 FILLER_42_290 ();
 sg13g2_fill_1 FILLER_42_292 ();
 sg13g2_fill_1 FILLER_42_342 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_4 FILLER_43_119 ();
 sg13g2_fill_1 FILLER_43_123 ();
 sg13g2_fill_2 FILLER_43_171 ();
 sg13g2_fill_1 FILLER_43_173 ();
 sg13g2_fill_1 FILLER_43_211 ();
 sg13g2_fill_2 FILLER_43_232 ();
 sg13g2_fill_2 FILLER_43_240 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_fill_1 FILLER_43_284 ();
 sg13g2_fill_1 FILLER_43_288 ();
 sg13g2_fill_2 FILLER_43_302 ();
 sg13g2_fill_2 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_342 ();
 sg13g2_fill_1 FILLER_43_362 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_decap_4 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_4 FILLER_44_119 ();
 sg13g2_fill_1 FILLER_44_123 ();
 sg13g2_fill_2 FILLER_44_147 ();
 sg13g2_fill_1 FILLER_44_149 ();
 sg13g2_decap_8 FILLER_44_173 ();
 sg13g2_fill_2 FILLER_44_180 ();
 sg13g2_fill_2 FILLER_44_194 ();
 sg13g2_fill_1 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_205 ();
 sg13g2_decap_4 FILLER_44_212 ();
 sg13g2_decap_4 FILLER_44_222 ();
 sg13g2_fill_2 FILLER_44_246 ();
 sg13g2_decap_4 FILLER_44_268 ();
 sg13g2_decap_8 FILLER_44_276 ();
 sg13g2_decap_8 FILLER_44_283 ();
 sg13g2_decap_8 FILLER_44_290 ();
 sg13g2_fill_1 FILLER_44_297 ();
 sg13g2_fill_2 FILLER_44_312 ();
 sg13g2_fill_1 FILLER_44_314 ();
 sg13g2_decap_4 FILLER_44_320 ();
 sg13g2_fill_2 FILLER_44_339 ();
 sg13g2_fill_1 FILLER_44_341 ();
 sg13g2_fill_2 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_147 ();
 sg13g2_fill_2 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_fill_2 FILLER_45_192 ();
 sg13g2_fill_1 FILLER_45_194 ();
 sg13g2_decap_8 FILLER_45_200 ();
 sg13g2_fill_1 FILLER_45_207 ();
 sg13g2_fill_1 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_234 ();
 sg13g2_decap_8 FILLER_45_241 ();
 sg13g2_decap_8 FILLER_45_248 ();
 sg13g2_fill_1 FILLER_45_255 ();
 sg13g2_decap_8 FILLER_45_283 ();
 sg13g2_decap_8 FILLER_45_290 ();
 sg13g2_decap_8 FILLER_45_307 ();
 sg13g2_decap_4 FILLER_45_314 ();
 sg13g2_fill_2 FILLER_45_318 ();
 sg13g2_fill_1 FILLER_45_325 ();
 sg13g2_fill_2 FILLER_45_336 ();
 sg13g2_fill_1 FILLER_45_338 ();
 sg13g2_fill_2 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_351 ();
 sg13g2_decap_8 FILLER_45_379 ();
 sg13g2_decap_8 FILLER_45_386 ();
 sg13g2_decap_8 FILLER_45_393 ();
 sg13g2_decap_8 FILLER_45_400 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_fill_2 FILLER_46_126 ();
 sg13g2_fill_1 FILLER_46_128 ();
 sg13g2_fill_2 FILLER_46_190 ();
 sg13g2_fill_2 FILLER_46_227 ();
 sg13g2_decap_4 FILLER_46_237 ();
 sg13g2_decap_8 FILLER_46_255 ();
 sg13g2_fill_2 FILLER_46_262 ();
 sg13g2_fill_2 FILLER_46_318 ();
 sg13g2_fill_1 FILLER_46_320 ();
 sg13g2_fill_2 FILLER_46_326 ();
 sg13g2_decap_8 FILLER_46_347 ();
 sg13g2_decap_4 FILLER_46_354 ();
 sg13g2_fill_2 FILLER_46_358 ();
 sg13g2_decap_8 FILLER_46_369 ();
 sg13g2_fill_2 FILLER_46_376 ();
 sg13g2_decap_8 FILLER_46_387 ();
 sg13g2_decap_8 FILLER_46_394 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_4 FILLER_47_126 ();
 sg13g2_fill_2 FILLER_47_161 ();
 sg13g2_fill_2 FILLER_47_229 ();
 sg13g2_decap_4 FILLER_47_261 ();
 sg13g2_fill_1 FILLER_47_265 ();
 sg13g2_fill_2 FILLER_47_275 ();
 sg13g2_fill_1 FILLER_47_277 ();
 sg13g2_fill_1 FILLER_47_283 ();
 sg13g2_fill_1 FILLER_47_311 ();
 sg13g2_fill_2 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_365 ();
 sg13g2_decap_8 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_379 ();
 sg13g2_decap_8 FILLER_47_386 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_4 FILLER_48_133 ();
 sg13g2_fill_2 FILLER_48_145 ();
 sg13g2_fill_1 FILLER_48_147 ();
 sg13g2_fill_1 FILLER_48_201 ();
 sg13g2_fill_2 FILLER_48_253 ();
 sg13g2_fill_2 FILLER_48_277 ();
 sg13g2_fill_2 FILLER_48_287 ();
 sg13g2_fill_2 FILLER_48_302 ();
 sg13g2_fill_1 FILLER_48_310 ();
 sg13g2_fill_2 FILLER_48_324 ();
 sg13g2_decap_8 FILLER_48_376 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_fill_2 FILLER_49_133 ();
 sg13g2_fill_2 FILLER_49_140 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_decap_8 FILLER_49_180 ();
 sg13g2_decap_4 FILLER_49_187 ();
 sg13g2_fill_1 FILLER_49_191 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_4 FILLER_49_218 ();
 sg13g2_fill_2 FILLER_49_227 ();
 sg13g2_fill_1 FILLER_49_229 ();
 sg13g2_fill_1 FILLER_49_235 ();
 sg13g2_fill_2 FILLER_49_241 ();
 sg13g2_fill_1 FILLER_49_243 ();
 sg13g2_fill_1 FILLER_49_249 ();
 sg13g2_fill_2 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_262 ();
 sg13g2_decap_8 FILLER_49_272 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_4 FILLER_49_294 ();
 sg13g2_fill_1 FILLER_49_298 ();
 sg13g2_fill_2 FILLER_49_324 ();
 sg13g2_fill_1 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_388 ();
 sg13g2_decap_8 FILLER_49_395 ();
 sg13g2_decap_8 FILLER_49_402 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_fill_2 FILLER_50_152 ();
 sg13g2_fill_1 FILLER_50_190 ();
 sg13g2_fill_1 FILLER_50_201 ();
 sg13g2_decap_8 FILLER_50_207 ();
 sg13g2_fill_1 FILLER_50_214 ();
 sg13g2_fill_2 FILLER_50_249 ();
 sg13g2_decap_8 FILLER_50_293 ();
 sg13g2_decap_4 FILLER_50_300 ();
 sg13g2_fill_1 FILLER_50_319 ();
 sg13g2_fill_1 FILLER_50_333 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_fill_1 FILLER_51_208 ();
 sg13g2_fill_1 FILLER_51_244 ();
 sg13g2_fill_2 FILLER_51_307 ();
 sg13g2_fill_2 FILLER_51_334 ();
 sg13g2_fill_1 FILLER_51_336 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_fill_2 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_4 FILLER_52_133 ();
 sg13g2_decap_4 FILLER_52_145 ();
 sg13g2_fill_2 FILLER_52_232 ();
 sg13g2_fill_1 FILLER_52_234 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_306 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_2 FILLER_52_324 ();
 sg13g2_decap_4 FILLER_52_339 ();
 sg13g2_fill_2 FILLER_52_370 ();
 sg13g2_decap_8 FILLER_52_376 ();
 sg13g2_decap_8 FILLER_52_383 ();
 sg13g2_decap_8 FILLER_52_390 ();
 sg13g2_decap_8 FILLER_52_397 ();
 sg13g2_decap_4 FILLER_52_404 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_4 FILLER_53_133 ();
 sg13g2_fill_1 FILLER_53_137 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_fill_2 FILLER_53_203 ();
 sg13g2_fill_1 FILLER_53_205 ();
 sg13g2_decap_4 FILLER_53_219 ();
 sg13g2_decap_8 FILLER_53_231 ();
 sg13g2_decap_4 FILLER_53_238 ();
 sg13g2_fill_1 FILLER_53_242 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_decap_8 FILLER_53_254 ();
 sg13g2_decap_4 FILLER_53_261 ();
 sg13g2_fill_2 FILLER_53_265 ();
 sg13g2_decap_8 FILLER_53_276 ();
 sg13g2_decap_4 FILLER_53_283 ();
 sg13g2_fill_1 FILLER_53_331 ();
 sg13g2_fill_2 FILLER_53_347 ();
 sg13g2_fill_2 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_387 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_decap_8 FILLER_53_401 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_fill_2 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_153 ();
 sg13g2_decap_8 FILLER_54_160 ();
 sg13g2_decap_8 FILLER_54_167 ();
 sg13g2_fill_2 FILLER_54_174 ();
 sg13g2_decap_4 FILLER_54_181 ();
 sg13g2_fill_1 FILLER_54_185 ();
 sg13g2_fill_1 FILLER_54_212 ();
 sg13g2_decap_8 FILLER_54_227 ();
 sg13g2_fill_1 FILLER_54_247 ();
 sg13g2_decap_4 FILLER_54_253 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_fill_2 FILLER_54_287 ();
 sg13g2_fill_1 FILLER_54_301 ();
 sg13g2_fill_2 FILLER_54_326 ();
 sg13g2_fill_1 FILLER_54_328 ();
 sg13g2_decap_4 FILLER_54_339 ();
 sg13g2_decap_8 FILLER_54_382 ();
 sg13g2_decap_8 FILLER_54_389 ();
 sg13g2_decap_8 FILLER_54_396 ();
 sg13g2_decap_4 FILLER_54_403 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_decap_4 FILLER_55_152 ();
 sg13g2_decap_4 FILLER_55_166 ();
 sg13g2_fill_2 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_221 ();
 sg13g2_decap_4 FILLER_55_247 ();
 sg13g2_fill_2 FILLER_55_259 ();
 sg13g2_decap_4 FILLER_55_287 ();
 sg13g2_fill_1 FILLER_55_291 ();
 sg13g2_decap_8 FILLER_55_300 ();
 sg13g2_fill_2 FILLER_55_316 ();
 sg13g2_fill_1 FILLER_55_347 ();
 sg13g2_fill_2 FILLER_55_358 ();
 sg13g2_decap_8 FILLER_55_386 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_4 FILLER_56_133 ();
 sg13g2_fill_2 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_241 ();
 sg13g2_decap_8 FILLER_56_291 ();
 sg13g2_decap_8 FILLER_56_298 ();
 sg13g2_decap_8 FILLER_56_305 ();
 sg13g2_fill_2 FILLER_56_341 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_fill_1 FILLER_56_358 ();
 sg13g2_decap_4 FILLER_56_403 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_4 FILLER_57_140 ();
 sg13g2_fill_1 FILLER_57_144 ();
 sg13g2_fill_1 FILLER_57_167 ();
 sg13g2_fill_2 FILLER_57_178 ();
 sg13g2_fill_1 FILLER_57_180 ();
 sg13g2_fill_2 FILLER_57_248 ();
 sg13g2_decap_4 FILLER_57_283 ();
 sg13g2_fill_2 FILLER_57_302 ();
 sg13g2_fill_1 FILLER_57_304 ();
 sg13g2_fill_1 FILLER_57_310 ();
 sg13g2_fill_1 FILLER_57_316 ();
 sg13g2_fill_1 FILLER_57_322 ();
 sg13g2_fill_1 FILLER_57_344 ();
 sg13g2_fill_2 FILLER_57_355 ();
 sg13g2_decap_8 FILLER_57_383 ();
 sg13g2_decap_8 FILLER_57_390 ();
 sg13g2_decap_8 FILLER_57_397 ();
 sg13g2_decap_4 FILLER_57_404 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_fill_2 FILLER_58_242 ();
 sg13g2_fill_1 FILLER_58_244 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_fill_1 FILLER_58_263 ();
 sg13g2_decap_8 FILLER_58_274 ();
 sg13g2_fill_2 FILLER_58_281 ();
 sg13g2_decap_8 FILLER_58_342 ();
 sg13g2_decap_8 FILLER_58_381 ();
 sg13g2_decap_8 FILLER_58_388 ();
 sg13g2_decap_8 FILLER_58_395 ();
 sg13g2_decap_8 FILLER_58_402 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_fill_1 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_153 ();
 sg13g2_decap_8 FILLER_59_216 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_fill_2 FILLER_59_235 ();
 sg13g2_fill_2 FILLER_59_295 ();
 sg13g2_fill_2 FILLER_59_335 ();
 sg13g2_fill_1 FILLER_59_345 ();
 sg13g2_decap_4 FILLER_59_356 ();
 sg13g2_fill_1 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_59_387 ();
 sg13g2_decap_8 FILLER_59_394 ();
 sg13g2_decap_8 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_fill_2 FILLER_60_152 ();
 sg13g2_fill_1 FILLER_60_154 ();
 sg13g2_fill_2 FILLER_60_181 ();
 sg13g2_fill_2 FILLER_60_215 ();
 sg13g2_fill_2 FILLER_60_253 ();
 sg13g2_fill_2 FILLER_60_302 ();
 sg13g2_fill_1 FILLER_60_323 ();
 sg13g2_decap_8 FILLER_60_384 ();
 sg13g2_decap_8 FILLER_60_391 ();
 sg13g2_decap_8 FILLER_60_398 ();
 sg13g2_decap_4 FILLER_60_405 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_fill_1 FILLER_61_119 ();
 sg13g2_fill_2 FILLER_61_183 ();
 sg13g2_fill_2 FILLER_61_190 ();
 sg13g2_fill_1 FILLER_61_192 ();
 sg13g2_fill_1 FILLER_61_210 ();
 sg13g2_decap_4 FILLER_61_220 ();
 sg13g2_fill_2 FILLER_61_224 ();
 sg13g2_fill_2 FILLER_61_252 ();
 sg13g2_fill_2 FILLER_61_269 ();
 sg13g2_fill_1 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_289 ();
 sg13g2_decap_8 FILLER_61_304 ();
 sg13g2_fill_1 FILLER_61_311 ();
 sg13g2_fill_2 FILLER_61_321 ();
 sg13g2_fill_2 FILLER_61_332 ();
 sg13g2_fill_1 FILLER_61_334 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_fill_2 FILLER_62_126 ();
 sg13g2_fill_1 FILLER_62_128 ();
 sg13g2_decap_4 FILLER_62_155 ();
 sg13g2_fill_1 FILLER_62_169 ();
 sg13g2_fill_1 FILLER_62_183 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_fill_1 FILLER_62_232 ();
 sg13g2_decap_4 FILLER_62_259 ();
 sg13g2_fill_1 FILLER_62_263 ();
 sg13g2_fill_2 FILLER_62_290 ();
 sg13g2_decap_4 FILLER_62_318 ();
 sg13g2_decap_8 FILLER_62_326 ();
 sg13g2_decap_4 FILLER_62_333 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_fill_2 FILLER_62_356 ();
 sg13g2_fill_1 FILLER_62_358 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_4 FILLER_63_133 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_fill_2 FILLER_63_143 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_fill_1 FILLER_63_191 ();
 sg13g2_decap_8 FILLER_63_199 ();
 sg13g2_decap_8 FILLER_63_214 ();
 sg13g2_decap_4 FILLER_63_221 ();
 sg13g2_decap_8 FILLER_63_233 ();
 sg13g2_fill_1 FILLER_63_240 ();
 sg13g2_decap_8 FILLER_63_249 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_324 ();
 sg13g2_decap_4 FILLER_63_340 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_decap_8 FILLER_63_369 ();
 sg13g2_decap_8 FILLER_63_376 ();
 sg13g2_decap_8 FILLER_63_383 ();
 sg13g2_decap_8 FILLER_63_390 ();
 sg13g2_decap_8 FILLER_63_397 ();
 sg13g2_decap_4 FILLER_63_404 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_4 FILLER_64_147 ();
 sg13g2_fill_1 FILLER_64_151 ();
 sg13g2_fill_1 FILLER_64_199 ();
 sg13g2_fill_2 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_212 ();
 sg13g2_decap_4 FILLER_64_223 ();
 sg13g2_decap_8 FILLER_64_231 ();
 sg13g2_decap_4 FILLER_64_238 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_decap_4 FILLER_64_259 ();
 sg13g2_fill_1 FILLER_64_263 ();
 sg13g2_decap_4 FILLER_64_287 ();
 sg13g2_fill_1 FILLER_64_311 ();
 sg13g2_decap_4 FILLER_64_364 ();
 sg13g2_decap_8 FILLER_64_377 ();
 sg13g2_decap_8 FILLER_64_384 ();
 sg13g2_decap_8 FILLER_64_391 ();
 sg13g2_decap_8 FILLER_64_398 ();
 sg13g2_decap_4 FILLER_64_405 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_fill_2 FILLER_65_140 ();
 sg13g2_fill_1 FILLER_65_178 ();
 sg13g2_fill_2 FILLER_65_203 ();
 sg13g2_fill_1 FILLER_65_205 ();
 sg13g2_fill_1 FILLER_65_237 ();
 sg13g2_fill_1 FILLER_65_260 ();
 sg13g2_fill_2 FILLER_65_266 ();
 sg13g2_fill_1 FILLER_65_268 ();
 sg13g2_decap_4 FILLER_65_277 ();
 sg13g2_fill_2 FILLER_65_321 ();
 sg13g2_fill_2 FILLER_65_333 ();
 sg13g2_decap_8 FILLER_65_387 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_fill_2 FILLER_66_133 ();
 sg13g2_fill_2 FILLER_66_161 ();
 sg13g2_fill_1 FILLER_66_163 ();
 sg13g2_fill_2 FILLER_66_209 ();
 sg13g2_decap_4 FILLER_66_277 ();
 sg13g2_fill_2 FILLER_66_281 ();
 sg13g2_fill_2 FILLER_66_291 ();
 sg13g2_fill_1 FILLER_66_293 ();
 sg13g2_fill_2 FILLER_66_304 ();
 sg13g2_fill_2 FILLER_66_316 ();
 sg13g2_fill_1 FILLER_66_318 ();
 sg13g2_fill_1 FILLER_66_338 ();
 sg13g2_fill_1 FILLER_66_349 ();
 sg13g2_decap_8 FILLER_66_376 ();
 sg13g2_decap_8 FILLER_66_383 ();
 sg13g2_decap_8 FILLER_66_390 ();
 sg13g2_decap_8 FILLER_66_397 ();
 sg13g2_decap_4 FILLER_66_404 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_fill_2 FILLER_67_140 ();
 sg13g2_fill_2 FILLER_67_184 ();
 sg13g2_fill_2 FILLER_67_222 ();
 sg13g2_fill_1 FILLER_67_224 ();
 sg13g2_fill_2 FILLER_67_265 ();
 sg13g2_decap_8 FILLER_67_380 ();
 sg13g2_decap_8 FILLER_67_387 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_4 FILLER_68_161 ();
 sg13g2_fill_1 FILLER_68_169 ();
 sg13g2_fill_2 FILLER_68_205 ();
 sg13g2_fill_1 FILLER_68_207 ();
 sg13g2_fill_1 FILLER_68_217 ();
 sg13g2_fill_2 FILLER_68_227 ();
 sg13g2_fill_1 FILLER_68_229 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_fill_2 FILLER_68_261 ();
 sg13g2_fill_1 FILLER_68_263 ();
 sg13g2_fill_1 FILLER_68_290 ();
 sg13g2_fill_2 FILLER_68_296 ();
 sg13g2_fill_1 FILLER_68_298 ();
 sg13g2_decap_4 FILLER_68_303 ();
 sg13g2_fill_2 FILLER_68_307 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_fill_1 FILLER_68_320 ();
 sg13g2_fill_2 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_367 ();
 sg13g2_decap_8 FILLER_68_374 ();
 sg13g2_decap_8 FILLER_68_381 ();
 sg13g2_decap_8 FILLER_68_388 ();
 sg13g2_decap_8 FILLER_68_395 ();
 sg13g2_decap_8 FILLER_68_402 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_192 ();
 sg13g2_decap_8 FILLER_69_199 ();
 sg13g2_decap_8 FILLER_69_206 ();
 sg13g2_decap_8 FILLER_69_216 ();
 sg13g2_decap_4 FILLER_69_223 ();
 sg13g2_fill_2 FILLER_69_238 ();
 sg13g2_fill_1 FILLER_69_240 ();
 sg13g2_decap_8 FILLER_69_252 ();
 sg13g2_fill_1 FILLER_69_274 ();
 sg13g2_decap_4 FILLER_69_286 ();
 sg13g2_fill_2 FILLER_69_290 ();
 sg13g2_decap_4 FILLER_69_311 ();
 sg13g2_fill_2 FILLER_69_315 ();
 sg13g2_decap_4 FILLER_69_322 ();
 sg13g2_fill_1 FILLER_69_326 ();
 sg13g2_fill_1 FILLER_69_336 ();
 sg13g2_decap_8 FILLER_69_363 ();
 sg13g2_decap_8 FILLER_69_370 ();
 sg13g2_decap_8 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_fill_2 FILLER_70_147 ();
 sg13g2_fill_2 FILLER_70_194 ();
 sg13g2_decap_8 FILLER_70_262 ();
 sg13g2_decap_4 FILLER_70_269 ();
 sg13g2_fill_1 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_277 ();
 sg13g2_decap_4 FILLER_70_284 ();
 sg13g2_fill_1 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_315 ();
 sg13g2_fill_1 FILLER_70_317 ();
 sg13g2_decap_8 FILLER_70_363 ();
 sg13g2_decap_8 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_398 ();
 sg13g2_decap_4 FILLER_70_405 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_4 FILLER_71_140 ();
 sg13g2_fill_1 FILLER_71_144 ();
 sg13g2_decap_8 FILLER_71_269 ();
 sg13g2_decap_8 FILLER_71_276 ();
 sg13g2_decap_8 FILLER_71_283 ();
 sg13g2_decap_4 FILLER_71_290 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_4 FILLER_72_147 ();
 sg13g2_fill_2 FILLER_72_151 ();
 sg13g2_fill_2 FILLER_72_176 ();
 sg13g2_fill_1 FILLER_72_187 ();
 sg13g2_fill_1 FILLER_72_258 ();
 sg13g2_fill_1 FILLER_72_263 ();
 sg13g2_decap_4 FILLER_72_268 ();
 sg13g2_fill_2 FILLER_72_298 ();
 sg13g2_fill_1 FILLER_72_304 ();
 sg13g2_decap_8 FILLER_72_348 ();
 sg13g2_decap_8 FILLER_72_355 ();
 sg13g2_decap_8 FILLER_72_362 ();
 sg13g2_decap_8 FILLER_72_369 ();
 sg13g2_decap_8 FILLER_72_376 ();
 sg13g2_decap_8 FILLER_72_383 ();
 sg13g2_decap_8 FILLER_72_390 ();
 sg13g2_decap_8 FILLER_72_397 ();
 sg13g2_decap_4 FILLER_72_404 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_4 FILLER_73_161 ();
 sg13g2_decap_4 FILLER_73_202 ();
 sg13g2_fill_1 FILLER_73_206 ();
 sg13g2_decap_8 FILLER_73_219 ();
 sg13g2_decap_8 FILLER_73_226 ();
 sg13g2_fill_1 FILLER_73_236 ();
 sg13g2_decap_8 FILLER_73_241 ();
 sg13g2_decap_4 FILLER_73_248 ();
 sg13g2_fill_1 FILLER_73_252 ();
 sg13g2_decap_4 FILLER_73_279 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_fill_1 FILLER_73_311 ();
 sg13g2_decap_8 FILLER_73_348 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_73_376 ();
 sg13g2_decap_8 FILLER_73_383 ();
 sg13g2_decap_8 FILLER_73_390 ();
 sg13g2_decap_8 FILLER_73_397 ();
 sg13g2_decap_4 FILLER_73_404 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_fill_2 FILLER_74_168 ();
 sg13g2_fill_1 FILLER_74_170 ();
 sg13g2_fill_2 FILLER_74_207 ();
 sg13g2_decap_8 FILLER_74_244 ();
 sg13g2_fill_2 FILLER_74_267 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_311 ();
 sg13g2_decap_8 FILLER_74_340 ();
 sg13g2_decap_8 FILLER_74_347 ();
 sg13g2_decap_8 FILLER_74_354 ();
 sg13g2_decap_8 FILLER_74_361 ();
 sg13g2_decap_8 FILLER_74_368 ();
 sg13g2_decap_8 FILLER_74_375 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_330 ();
 sg13g2_decap_8 FILLER_75_337 ();
 sg13g2_decap_8 FILLER_75_344 ();
 sg13g2_decap_8 FILLER_75_351 ();
 sg13g2_decap_8 FILLER_75_358 ();
 sg13g2_decap_8 FILLER_75_365 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_4 FILLER_76_182 ();
 sg13g2_decap_4 FILLER_76_244 ();
 sg13g2_fill_2 FILLER_76_248 ();
 sg13g2_decap_8 FILLER_76_253 ();
 sg13g2_fill_1 FILLER_76_268 ();
 sg13g2_decap_4 FILLER_76_290 ();
 sg13g2_decap_8 FILLER_76_327 ();
 sg13g2_decap_8 FILLER_76_334 ();
 sg13g2_decap_8 FILLER_76_341 ();
 sg13g2_decap_8 FILLER_76_348 ();
 sg13g2_decap_8 FILLER_76_355 ();
 sg13g2_decap_8 FILLER_76_362 ();
 sg13g2_decap_8 FILLER_76_369 ();
 sg13g2_decap_8 FILLER_76_376 ();
 sg13g2_decap_8 FILLER_76_383 ();
 sg13g2_decap_8 FILLER_76_390 ();
 sg13g2_decap_8 FILLER_76_397 ();
 sg13g2_decap_4 FILLER_76_404 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_4 FILLER_77_189 ();
 sg13g2_fill_2 FILLER_77_193 ();
 sg13g2_fill_2 FILLER_77_230 ();
 sg13g2_fill_1 FILLER_77_232 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_4 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_335 ();
 sg13g2_decap_8 FILLER_77_342 ();
 sg13g2_decap_8 FILLER_77_349 ();
 sg13g2_decap_8 FILLER_77_356 ();
 sg13g2_decap_8 FILLER_77_363 ();
 sg13g2_decap_8 FILLER_77_370 ();
 sg13g2_decap_8 FILLER_77_377 ();
 sg13g2_decap_8 FILLER_77_384 ();
 sg13g2_decap_8 FILLER_77_391 ();
 sg13g2_decap_8 FILLER_77_398 ();
 sg13g2_decap_4 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_fill_1 FILLER_78_210 ();
 sg13g2_fill_1 FILLER_78_219 ();
 sg13g2_fill_2 FILLER_78_246 ();
 sg13g2_fill_2 FILLER_78_269 ();
 sg13g2_decap_8 FILLER_78_332 ();
 sg13g2_decap_8 FILLER_78_339 ();
 sg13g2_decap_8 FILLER_78_346 ();
 sg13g2_decap_8 FILLER_78_353 ();
 sg13g2_decap_8 FILLER_78_360 ();
 sg13g2_decap_8 FILLER_78_367 ();
 sg13g2_decap_8 FILLER_78_374 ();
 sg13g2_decap_8 FILLER_78_381 ();
 sg13g2_decap_8 FILLER_78_388 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_291 ();
 sg13g2_decap_8 FILLER_79_298 ();
 sg13g2_decap_8 FILLER_79_309 ();
 sg13g2_decap_8 FILLER_79_316 ();
 sg13g2_decap_8 FILLER_79_323 ();
 sg13g2_decap_8 FILLER_79_330 ();
 sg13g2_decap_8 FILLER_79_337 ();
 sg13g2_decap_8 FILLER_79_344 ();
 sg13g2_decap_8 FILLER_79_351 ();
 sg13g2_decap_8 FILLER_79_358 ();
 sg13g2_decap_8 FILLER_79_365 ();
 sg13g2_decap_8 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_379 ();
 sg13g2_decap_8 FILLER_79_386 ();
 sg13g2_decap_8 FILLER_79_393 ();
 sg13g2_decap_8 FILLER_79_400 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_fill_2 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_238 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_decap_4 FILLER_80_260 ();
 sg13g2_fill_2 FILLER_80_285 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_295 ();
 sg13g2_decap_8 FILLER_80_301 ();
 sg13g2_decap_4 FILLER_80_308 ();
 sg13g2_decap_8 FILLER_80_336 ();
 sg13g2_decap_8 FILLER_80_343 ();
 sg13g2_decap_8 FILLER_80_350 ();
 sg13g2_decap_8 FILLER_80_357 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_4 FILLER_80_371 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_384 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_4 FILLER_80_405 ();
 assign uio_oe[0] = net12;
 assign uio_oe[1] = net13;
 assign uio_oe[2] = net14;
 assign uio_oe[3] = net15;
 assign uio_oe[4] = net16;
 assign uio_oe[5] = net17;
 assign uio_oe[6] = net18;
 assign uio_oe[7] = net19;
 assign uio_out[0] = net20;
 assign uio_out[1] = net21;
 assign uio_out[2] = net22;
 assign uio_out[3] = net23;
 assign uio_out[4] = net24;
 assign uio_out[5] = net25;
 assign uio_out[6] = net26;
 assign uio_out[7] = net27;
endmodule

module tt_um_rebeccargb_vga_timing_experiments (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire clknet_0_clk;
 wire net33;
 wire \color_in[0] ;
 wire \color_in[1] ;
 wire \color_in[2] ;
 wire \color_in[3] ;
 wire \color_in[4] ;
 wire \color_in[5] ;
 wire \hbackporch[0] ;
 wire \hbackporch[1] ;
 wire \hbackporch[2] ;
 wire \hbackporch[3] ;
 wire \hbackporch[4] ;
 wire \hbackporch[5] ;
 wire \hbackporch[6] ;
 wire \hbackporch[7] ;
 wire \hbackporch[8] ;
 wire \hbackporch[9] ;
 wire \hdisplay[0] ;
 wire \hdisplay[10] ;
 wire \hdisplay[1] ;
 wire \hdisplay[2] ;
 wire \hdisplay[3] ;
 wire \hdisplay[4] ;
 wire \hdisplay[5] ;
 wire \hdisplay[6] ;
 wire \hdisplay[7] ;
 wire \hdisplay[8] ;
 wire \hdisplay[9] ;
 wire \hfrontporch[0] ;
 wire \hfrontporch[1] ;
 wire \hfrontporch[2] ;
 wire \hfrontporch[3] ;
 wire \hfrontporch[4] ;
 wire \hfrontporch[5] ;
 wire \hfrontporch[6] ;
 wire \hfrontporch[7] ;
 wire \hfrontporch[8] ;
 wire \hfrontporch[9] ;
 wire \hpos[0] ;
 wire \hpos[10] ;
 wire \hpos[11] ;
 wire \hpos[1] ;
 wire \hpos[2] ;
 wire \hpos[3] ;
 wire \hpos[4] ;
 wire \hpos[5] ;
 wire \hpos[6] ;
 wire \hpos[7] ;
 wire \hpos[8] ;
 wire \hpos[9] ;
 wire hsync;
 wire \hsynclength[0] ;
 wire \hsynclength[1] ;
 wire \hsynclength[2] ;
 wire \hsynclength[3] ;
 wire \hsynclength[4] ;
 wire \hsynclength[5] ;
 wire \hsynclength[6] ;
 wire \hsynclength[7] ;
 wire \hsynclength[8] ;
 wire \hsynclength[9] ;
 wire hsyncpolarity;
 wire \hvsync_gen.vbackporch[0] ;
 wire \hvsync_gen.vbackporch[1] ;
 wire \hvsync_gen.vbackporch[2] ;
 wire \hvsync_gen.vbackporch[3] ;
 wire \hvsync_gen.vbackporch[4] ;
 wire \hvsync_gen.vbackporch[5] ;
 wire \hvsync_gen.vbackporch[6] ;
 wire \hvsync_gen.vbackporch[7] ;
 wire \hvsync_gen.vdisplay[0] ;
 wire \hvsync_gen.vdisplay[10] ;
 wire \hvsync_gen.vdisplay[1] ;
 wire \hvsync_gen.vdisplay[2] ;
 wire \hvsync_gen.vdisplay[3] ;
 wire \hvsync_gen.vdisplay[4] ;
 wire \hvsync_gen.vdisplay[5] ;
 wire \hvsync_gen.vdisplay[6] ;
 wire \hvsync_gen.vdisplay[7] ;
 wire \hvsync_gen.vdisplay[8] ;
 wire \hvsync_gen.vdisplay[9] ;
 wire \hvsync_gen.vfrontporch[0] ;
 wire \hvsync_gen.vfrontporch[1] ;
 wire \hvsync_gen.vfrontporch[2] ;
 wire \hvsync_gen.vfrontporch[3] ;
 wire \hvsync_gen.vfrontporch[4] ;
 wire \hvsync_gen.vfrontporch[5] ;
 wire \hvsync_gen.vfrontporch[6] ;
 wire \hvsync_gen.vfrontporch[7] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[10] ;
 wire \hvsync_gen.vpos[11] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \hvsync_gen.vsynclength[0] ;
 wire \hvsync_gen.vsynclength[1] ;
 wire \hvsync_gen.vsynclength[2] ;
 wire \hvsync_gen.vsynclength[3] ;
 wire \hvsync_gen.vsynclength[4] ;
 wire \hvsync_gen.vsynclength[5] ;
 wire \hvsync_gen.vsynclength[6] ;
 wire \hvsync_gen.vsynclength[7] ;
 wire \hvsync_gen.vsyncpolarity ;
 wire \pat.pattern[0] ;
 wire \pat.pattern[1] ;
 wire \pat.pattern[2] ;
 wire \pat.pattern[3] ;
 wire \pat.pattern[4] ;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;

 sg13g2_inv_1 _1700_ (.Y(_0789_),
    .A(net5));
 sg13g2_inv_2 _1701_ (.Y(_0790_),
    .A(net14));
 sg13g2_inv_1 _1702_ (.Y(_0791_),
    .A(net13));
 sg13g2_inv_1 _1703_ (.Y(_0792_),
    .A(net12));
 sg13g2_inv_1 _1704_ (.Y(_0793_),
    .A(net148));
 sg13g2_inv_1 _1705_ (.Y(_0794_),
    .A(net336));
 sg13g2_inv_2 _1706_ (.Y(_0795_),
    .A(\hpos[0] ));
 sg13g2_inv_1 _1707_ (.Y(_0796_),
    .A(net1));
 sg13g2_inv_1 _1708_ (.Y(_0797_),
    .A(net335));
 sg13g2_inv_1 _1709_ (.Y(_0798_),
    .A(\hvsync_gen.vfrontporch[1] ));
 sg13g2_inv_1 _1710_ (.Y(_0799_),
    .A(\hvsync_gen.vsynclength[1] ));
 sg13g2_inv_1 _1711_ (.Y(_0800_),
    .A(net333));
 sg13g2_inv_1 _1712_ (.Y(_0801_),
    .A(_0004_));
 sg13g2_inv_1 _1713_ (.Y(_0802_),
    .A(net330));
 sg13g2_inv_1 _1714_ (.Y(_0803_),
    .A(_0005_));
 sg13g2_inv_4 _1715_ (.A(net329),
    .Y(_0804_));
 sg13g2_inv_1 _1716_ (.Y(_0805_),
    .A(\hvsync_gen.vbackporch[4] ));
 sg13g2_inv_1 _1717_ (.Y(_0806_),
    .A(_0006_));
 sg13g2_inv_2 _1718_ (.Y(_0807_),
    .A(\hvsync_gen.vpos[5] ));
 sg13g2_inv_1 _1719_ (.Y(_0808_),
    .A(\hvsync_gen.vdisplay[5] ));
 sg13g2_inv_2 _1720_ (.Y(_0809_),
    .A(_0007_));
 sg13g2_inv_2 _1721_ (.Y(_0810_),
    .A(net323));
 sg13g2_inv_1 _1722_ (.Y(_0811_),
    .A(\hvsync_gen.vdisplay[6] ));
 sg13g2_inv_1 _1723_ (.Y(_0812_),
    .A(\hvsync_gen.vbackporch[6] ));
 sg13g2_inv_1 _1724_ (.Y(_0813_),
    .A(_0008_));
 sg13g2_inv_1 _1725_ (.Y(_0814_),
    .A(net320));
 sg13g2_inv_1 _1726_ (.Y(_0815_),
    .A(net319));
 sg13g2_inv_1 _1727_ (.Y(_0816_),
    .A(\hvsync_gen.vdisplay[8] ));
 sg13g2_inv_2 _1728_ (.Y(_0817_),
    .A(_0010_));
 sg13g2_inv_1 _1729_ (.Y(_0818_),
    .A(\hvsync_gen.vdisplay[9] ));
 sg13g2_inv_2 _1730_ (.Y(_0819_),
    .A(net359));
 sg13g2_inv_4 _1731_ (.A(net356),
    .Y(_0820_));
 sg13g2_inv_4 _1732_ (.A(net354),
    .Y(_0821_));
 sg13g2_inv_1 _1733_ (.Y(_0822_),
    .A(\hfrontporch[4] ));
 sg13g2_inv_1 _1734_ (.Y(_0823_),
    .A(\hdisplay[4] ));
 sg13g2_inv_1 _1735_ (.Y(_0824_),
    .A(\hbackporch[4] ));
 sg13g2_inv_4 _1736_ (.A(net352),
    .Y(_0825_));
 sg13g2_inv_1 _1737_ (.Y(_0826_),
    .A(\hsynclength[5] ));
 sg13g2_inv_1 _1738_ (.Y(_0827_),
    .A(\hbackporch[5] ));
 sg13g2_inv_2 _1739_ (.Y(_0828_),
    .A(net349));
 sg13g2_inv_1 _1740_ (.Y(_0829_),
    .A(\hsynclength[6] ));
 sg13g2_inv_2 _1741_ (.Y(_0830_),
    .A(net347));
 sg13g2_inv_1 _1742_ (.Y(_0831_),
    .A(_0021_));
 sg13g2_inv_1 _1743_ (.Y(_0832_),
    .A(net346));
 sg13g2_inv_1 _1744_ (.Y(_0833_),
    .A(\hfrontporch[8] ));
 sg13g2_inv_1 _1745_ (.Y(_0834_),
    .A(\hdisplay[8] ));
 sg13g2_inv_1 _1746_ (.Y(_0835_),
    .A(\hdisplay[9] ));
 sg13g2_inv_1 _1747_ (.Y(_0836_),
    .A(net171));
 sg13g2_inv_1 _1748_ (.Y(_0837_),
    .A(\hdisplay[10] ));
 sg13g2_inv_1 _1749_ (.Y(_0838_),
    .A(net339));
 sg13g2_inv_1 _1750_ (.Y(_0839_),
    .A(net338));
 sg13g2_inv_1 _1751_ (.Y(_0840_),
    .A(\color_in[0] ));
 sg13g2_inv_1 _1752_ (.Y(_0841_),
    .A(\color_in[2] ));
 sg13g2_inv_1 _1753_ (.Y(_0842_),
    .A(\color_in[4] ));
 sg13g2_inv_2 _1754_ (.Y(_0843_),
    .A(\color_in[5] ));
 sg13g2_nand2b_1 _1755_ (.Y(_0844_),
    .B(\pat.pattern[0] ),
    .A_N(\pat.pattern[1] ));
 sg13g2_nor2_2 _1756_ (.A(net341),
    .B(_0838_),
    .Y(_0845_));
 sg13g2_nand2_2 _1757_ (.Y(_0846_),
    .A(\pat.pattern[4] ),
    .B(_0845_));
 sg13g2_nor2_1 _1758_ (.A(net317),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_nand2_1 _1759_ (.Y(_0848_),
    .A(_0006_),
    .B(_0847_));
 sg13g2_nor2_2 _1760_ (.A(net335),
    .B(net333),
    .Y(_0849_));
 sg13g2_nand2_1 _1761_ (.Y(_0850_),
    .A(_0005_),
    .B(_0849_));
 sg13g2_xnor2_1 _1762_ (.Y(_0851_),
    .A(_0804_),
    .B(_0850_));
 sg13g2_o21ai_1 _1763_ (.B1(_0848_),
    .Y(_0852_),
    .A1(net295),
    .A2(_0851_));
 sg13g2_nand2_1 _1764_ (.Y(_0853_),
    .A(net353),
    .B(_0852_));
 sg13g2_nand2_1 _1765_ (.Y(_0854_),
    .A(net335),
    .B(net334));
 sg13g2_nor2_1 _1766_ (.A(net295),
    .B(_0849_),
    .Y(_0855_));
 sg13g2_a22oi_1 _1767_ (.Y(_0856_),
    .B1(_0854_),
    .B2(_0855_),
    .A2(net295),
    .A1(_0801_));
 sg13g2_nand2_1 _1768_ (.Y(_0857_),
    .A(net357),
    .B(_0856_));
 sg13g2_nand2_1 _1769_ (.Y(_0858_),
    .A(\hvsync_gen.vpos[1] ),
    .B(_0819_));
 sg13g2_xor2_1 _1770_ (.B(_0856_),
    .A(net357),
    .X(_0859_));
 sg13g2_nand2_1 _1771_ (.Y(_0860_),
    .A(_0858_),
    .B(_0859_));
 sg13g2_xnor2_1 _1772_ (.Y(_0861_),
    .A(_0803_),
    .B(_0855_));
 sg13g2_xor2_1 _1773_ (.B(_0861_),
    .A(_0017_),
    .X(_0862_));
 sg13g2_a21o_1 _1774_ (.A2(_0860_),
    .A1(_0857_),
    .B1(_0862_),
    .X(_0863_));
 sg13g2_nand2_1 _1775_ (.Y(_0864_),
    .A(net355),
    .B(_0861_));
 sg13g2_xnor2_1 _1776_ (.Y(_0865_),
    .A(net354),
    .B(_0852_));
 sg13g2_a21o_1 _1777_ (.A2(_0864_),
    .A1(_0863_),
    .B1(_0865_),
    .X(_0866_));
 sg13g2_nor2_2 _1778_ (.A(net332),
    .B(net328),
    .Y(_0867_));
 sg13g2_and2_1 _1779_ (.A(_0849_),
    .B(_0867_),
    .X(_0868_));
 sg13g2_xnor2_1 _1780_ (.Y(_0869_),
    .A(_0807_),
    .B(_0868_));
 sg13g2_nor2_1 _1781_ (.A(net295),
    .B(_0869_),
    .Y(_0870_));
 sg13g2_a21oi_2 _1782_ (.B1(_0870_),
    .Y(_0871_),
    .A2(net295),
    .A1(_0809_));
 sg13g2_nand2_1 _1783_ (.Y(_0872_),
    .A(net351),
    .B(_0871_));
 sg13g2_xnor2_1 _1784_ (.Y(_0873_),
    .A(net351),
    .B(_0871_));
 sg13g2_a21o_1 _1785_ (.A2(_0866_),
    .A1(_0853_),
    .B1(_0873_),
    .X(_0874_));
 sg13g2_nand2_2 _1786_ (.Y(_0875_),
    .A(\pat.pattern[0] ),
    .B(\pat.pattern[1] ));
 sg13g2_nor3_2 _1787_ (.A(net342),
    .B(net340),
    .C(_0875_),
    .Y(_0876_));
 sg13g2_a21o_2 _1788_ (.A2(_0876_),
    .A1(\pat.pattern[4] ),
    .B1(net295),
    .X(_0877_));
 sg13g2_nand3_1 _1789_ (.B(_0866_),
    .C(_0873_),
    .A(_0853_),
    .Y(_0878_));
 sg13g2_nand3_1 _1790_ (.B(_0877_),
    .C(_0878_),
    .A(_0874_),
    .Y(_0879_));
 sg13g2_nand2_2 _1791_ (.Y(_0880_),
    .A(net337),
    .B(_0845_));
 sg13g2_nor2_1 _1792_ (.A(net317),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_nor2_1 _1793_ (.A(net155),
    .B(net359),
    .Y(_0882_));
 sg13g2_nor3_2 _1794_ (.A(\hpos[0] ),
    .B(\hpos[1] ),
    .C(net357),
    .Y(_0883_));
 sg13g2_nand2_1 _1795_ (.Y(_0884_),
    .A(_0820_),
    .B(_0883_));
 sg13g2_nor2_2 _1796_ (.A(net333),
    .B(net332),
    .Y(_0885_));
 sg13g2_nor2_2 _1797_ (.A(net336),
    .B(net335),
    .Y(_0886_));
 sg13g2_and2_1 _1798_ (.A(_0885_),
    .B(_0886_),
    .X(_0887_));
 sg13g2_nand2_1 _1799_ (.Y(_0888_),
    .A(_0885_),
    .B(_0886_));
 sg13g2_nor2_1 _1800_ (.A(_0795_),
    .B(_0819_),
    .Y(_0889_));
 sg13g2_and2_2 _1801_ (.A(net357),
    .B(_0889_),
    .X(_0890_));
 sg13g2_and2_1 _1802_ (.A(net355),
    .B(_0890_),
    .X(_0891_));
 sg13g2_nand2_2 _1803_ (.Y(_0892_),
    .A(net355),
    .B(_0890_));
 sg13g2_nand2_1 _1804_ (.Y(_0893_),
    .A(net333),
    .B(net331));
 sg13g2_nand2_2 _1805_ (.Y(_0894_),
    .A(net336),
    .B(net335));
 sg13g2_or2_2 _1806_ (.X(_0895_),
    .B(_0894_),
    .A(_0893_));
 sg13g2_nand4_1 _1807_ (.B(_0888_),
    .C(_0892_),
    .A(_0884_),
    .Y(_0896_),
    .D(_0895_));
 sg13g2_nor3_1 _1808_ (.A(net317),
    .B(_0880_),
    .C(_0896_),
    .Y(_0897_));
 sg13g2_nand2b_2 _1809_ (.Y(_0898_),
    .B(\pat.pattern[1] ),
    .A_N(\pat.pattern[0] ));
 sg13g2_nor3_1 _1810_ (.A(net342),
    .B(net340),
    .C(_0898_),
    .Y(_0899_));
 sg13g2_nand2_1 _1811_ (.Y(_0900_),
    .A(net337),
    .B(_0899_));
 sg13g2_xnor2_1 _1812_ (.Y(_0901_),
    .A(\hvsync_gen.vpos[1] ),
    .B(net359));
 sg13g2_inv_1 _1813_ (.Y(_0902_),
    .A(_0901_));
 sg13g2_nor2_1 _1814_ (.A(_0900_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_nor3_1 _1815_ (.A(net342),
    .B(net340),
    .C(net317),
    .Y(_0904_));
 sg13g2_inv_1 _1816_ (.Y(_0905_),
    .A(_0904_));
 sg13g2_nand2_1 _1817_ (.Y(_0906_),
    .A(\hvsync_gen.vpos[0] ),
    .B(_0795_));
 sg13g2_xor2_1 _1818_ (.B(\hpos[0] ),
    .A(net336),
    .X(_0907_));
 sg13g2_nor3_1 _1819_ (.A(_0839_),
    .B(_0905_),
    .C(_0907_),
    .Y(_0908_));
 sg13g2_nor3_2 _1820_ (.A(_0897_),
    .B(_0903_),
    .C(_0908_),
    .Y(_0909_));
 sg13g2_nand2_1 _1821_ (.Y(_0910_),
    .A(net337),
    .B(_0876_));
 sg13g2_nor2_1 _1822_ (.A(_0800_),
    .B(net358),
    .Y(_0911_));
 sg13g2_xor2_1 _1823_ (.B(net358),
    .A(net334),
    .X(_0912_));
 sg13g2_nor2_1 _1824_ (.A(_0910_),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_nor2_1 _1825_ (.A(_0875_),
    .B(_0880_),
    .Y(_0914_));
 sg13g2_nor2_2 _1826_ (.A(_0821_),
    .B(_0892_),
    .Y(_0915_));
 sg13g2_nand2_2 _1827_ (.Y(_0916_),
    .A(net350),
    .B(_0915_));
 sg13g2_nor2_1 _1828_ (.A(net353),
    .B(_0884_),
    .Y(_0917_));
 sg13g2_nor2_2 _1829_ (.A(net329),
    .B(net326),
    .Y(_0918_));
 sg13g2_and2_1 _1830_ (.A(_0885_),
    .B(_0918_),
    .X(_0919_));
 sg13g2_nand2_2 _1831_ (.Y(_0920_),
    .A(_0887_),
    .B(_0918_));
 sg13g2_nand2_2 _1832_ (.Y(_0921_),
    .A(net328),
    .B(net326));
 sg13g2_nor2_2 _1833_ (.A(_0895_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_a21oi_1 _1834_ (.A1(_0825_),
    .A2(_0917_),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_nand3_1 _1835_ (.B(_0920_),
    .C(_0923_),
    .A(_0916_),
    .Y(_0924_));
 sg13g2_nand4_1 _1836_ (.B(_0916_),
    .C(_0920_),
    .A(_0914_),
    .Y(_0925_),
    .D(_0923_));
 sg13g2_nor2_1 _1837_ (.A(_0880_),
    .B(_0898_),
    .Y(_0926_));
 sg13g2_nor2_1 _1838_ (.A(net328),
    .B(_0888_),
    .Y(_0927_));
 sg13g2_inv_1 _1839_ (.Y(_0928_),
    .A(_0927_));
 sg13g2_nor2_1 _1840_ (.A(net172),
    .B(_0895_),
    .Y(_0929_));
 sg13g2_nor4_1 _1841_ (.A(_0915_),
    .B(_0917_),
    .C(_0927_),
    .D(_0929_),
    .Y(_0930_));
 sg13g2_or2_1 _1842_ (.X(_0931_),
    .B(\pat.pattern[1] ),
    .A(\pat.pattern[0] ));
 sg13g2_nor2_1 _1843_ (.A(_0880_),
    .B(net316),
    .Y(_0932_));
 sg13g2_nand2_1 _1844_ (.Y(_0933_),
    .A(_0004_),
    .B(_0886_));
 sg13g2_nor2_1 _1845_ (.A(net170),
    .B(_0894_),
    .Y(_0934_));
 sg13g2_nor2_1 _1846_ (.A(_0883_),
    .B(_0934_),
    .Y(_0935_));
 sg13g2_nand3b_1 _1847_ (.B(_0933_),
    .C(_0935_),
    .Y(_0936_),
    .A_N(_0890_));
 sg13g2_nor3_1 _1848_ (.A(_0880_),
    .B(net316),
    .C(_0936_),
    .Y(_0937_));
 sg13g2_nor2b_1 _1849_ (.A(net339),
    .B_N(net341),
    .Y(_0938_));
 sg13g2_nand2_1 _1850_ (.Y(_0939_),
    .A(net337),
    .B(_0938_));
 sg13g2_nor2_1 _1851_ (.A(_0875_),
    .B(net306),
    .Y(_0940_));
 sg13g2_xor2_1 _1852_ (.B(net349),
    .A(net325),
    .X(_0941_));
 sg13g2_nor3_1 _1853_ (.A(_0875_),
    .B(net306),
    .C(_0941_),
    .Y(_0942_));
 sg13g2_nor2_1 _1854_ (.A(_0804_),
    .B(net354),
    .Y(_0943_));
 sg13g2_xor2_1 _1855_ (.B(net353),
    .A(net328),
    .X(_0944_));
 sg13g2_inv_1 _1856_ (.Y(_0945_),
    .A(_0944_));
 sg13g2_nor3_1 _1857_ (.A(net317),
    .B(net306),
    .C(_0944_),
    .Y(_0946_));
 sg13g2_nor2_1 _1858_ (.A(_0898_),
    .B(net306),
    .Y(_0947_));
 sg13g2_nor2_1 _1859_ (.A(_0807_),
    .B(net351),
    .Y(_0948_));
 sg13g2_xor2_1 _1860_ (.B(net350),
    .A(net327),
    .X(_0949_));
 sg13g2_nor3_1 _1861_ (.A(_0898_),
    .B(net306),
    .C(_0949_),
    .Y(_0950_));
 sg13g2_nor2_1 _1862_ (.A(net316),
    .B(net306),
    .Y(_0951_));
 sg13g2_nand2_1 _1863_ (.Y(_0952_),
    .A(net332),
    .B(_0820_));
 sg13g2_xnor2_1 _1864_ (.Y(_0953_),
    .A(net331),
    .B(net355));
 sg13g2_nor2_1 _1865_ (.A(_0942_),
    .B(_0950_),
    .Y(_0954_));
 sg13g2_nor2_1 _1866_ (.A(_0937_),
    .B(_0946_),
    .Y(_0955_));
 sg13g2_a22oi_1 _1867_ (.Y(_0956_),
    .B1(_0951_),
    .B2(_0953_),
    .A2(_0930_),
    .A1(_0926_));
 sg13g2_nand4_1 _1868_ (.B(_0954_),
    .C(_0955_),
    .A(_0925_),
    .Y(_0957_),
    .D(_0956_));
 sg13g2_nor2_1 _1869_ (.A(_0913_),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_nand2_1 _1870_ (.Y(_0959_),
    .A(_0909_),
    .B(_0958_));
 sg13g2_nand3_1 _1871_ (.B(net339),
    .C(\pat.pattern[4] ),
    .A(net342),
    .Y(_0960_));
 sg13g2_nor2_2 _1872_ (.A(_0931_),
    .B(_0960_),
    .Y(_0961_));
 sg13g2_inv_1 _1873_ (.Y(_0962_),
    .A(_0961_));
 sg13g2_nand2_2 _1874_ (.Y(_0963_),
    .A(\pat.pattern[4] ),
    .B(_0938_));
 sg13g2_o21ai_1 _1875_ (.B1(_0962_),
    .Y(_0964_),
    .A1(_0898_),
    .A2(_0963_));
 sg13g2_nor2_1 _1876_ (.A(_0846_),
    .B(net316),
    .Y(_0965_));
 sg13g2_a21o_2 _1877_ (.A2(_0899_),
    .A1(\pat.pattern[4] ),
    .B1(net294),
    .X(_0966_));
 sg13g2_nor2_1 _1878_ (.A(_0846_),
    .B(_0875_),
    .Y(_0967_));
 sg13g2_nor2_1 _1879_ (.A(net317),
    .B(_0963_),
    .Y(_0968_));
 sg13g2_nor2_2 _1880_ (.A(net293),
    .B(_0968_),
    .Y(_0969_));
 sg13g2_or2_1 _1881_ (.X(_0970_),
    .B(_0968_),
    .A(net293));
 sg13g2_nor4_2 _1882_ (.A(net341),
    .B(net339),
    .C(net337),
    .Y(_0971_),
    .D(net316));
 sg13g2_a21oi_1 _1883_ (.A1(net337),
    .A2(_0876_),
    .Y(_0972_),
    .B1(_0971_));
 sg13g2_nand3_1 _1884_ (.B(net341),
    .C(net340),
    .A(\pat.pattern[1] ),
    .Y(_0973_));
 sg13g2_nor2_1 _1885_ (.A(net338),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_inv_1 _1886_ (.Y(_0975_),
    .A(_0974_));
 sg13g2_nand3b_1 _1887_ (.B(net339),
    .C(net341),
    .Y(_0976_),
    .A_N(\pat.pattern[4] ));
 sg13g2_nor2_2 _1888_ (.A(net317),
    .B(_0960_),
    .Y(_0977_));
 sg13g2_inv_1 _1889_ (.Y(_0978_),
    .A(_0977_));
 sg13g2_o21ai_1 _1890_ (.B1(_0978_),
    .Y(_0979_),
    .A1(_0875_),
    .A2(_0963_));
 sg13g2_nor2_2 _1891_ (.A(_0846_),
    .B(_0898_),
    .Y(_0980_));
 sg13g2_nor2_1 _1892_ (.A(net316),
    .B(_0963_),
    .Y(_0981_));
 sg13g2_or2_2 _1893_ (.X(_0982_),
    .B(_0981_),
    .A(_0980_));
 sg13g2_nand4_1 _1894_ (.B(_0905_),
    .C(_0972_),
    .A(_0900_),
    .Y(_0983_),
    .D(_0976_));
 sg13g2_nor3_1 _1895_ (.A(_0964_),
    .B(_0966_),
    .C(_0982_),
    .Y(_0984_));
 sg13g2_nand4_1 _1896_ (.B(_0939_),
    .C(_0969_),
    .A(_0880_),
    .Y(_0985_),
    .D(_0975_));
 sg13g2_nor4_1 _1897_ (.A(_0877_),
    .B(_0979_),
    .C(_0983_),
    .D(_0985_),
    .Y(_0986_));
 sg13g2_and2_1 _1898_ (.A(_0984_),
    .B(_0986_),
    .X(_0987_));
 sg13g2_nor2_2 _1899_ (.A(net317),
    .B(_0976_),
    .Y(_0988_));
 sg13g2_nor2_2 _1900_ (.A(net337),
    .B(_0905_),
    .Y(_0989_));
 sg13g2_a22oi_1 _1901_ (.Y(_0990_),
    .B1(_0989_),
    .B2(net347),
    .A2(_0988_),
    .A1(net356));
 sg13g2_nor2_2 _1902_ (.A(net316),
    .B(_0976_),
    .Y(_0991_));
 sg13g2_nor2_2 _1903_ (.A(_0875_),
    .B(_0976_),
    .Y(_0992_));
 sg13g2_a22oi_1 _1904_ (.Y(_0993_),
    .B1(_0992_),
    .B2(net350),
    .A2(_0991_),
    .A1(net358));
 sg13g2_and2_1 _1905_ (.A(\pat.pattern[0] ),
    .B(_0974_),
    .X(_0994_));
 sg13g2_nor2_2 _1906_ (.A(\pat.pattern[0] ),
    .B(_0975_),
    .Y(_0995_));
 sg13g2_a22oi_1 _1907_ (.Y(_0996_),
    .B1(_0995_),
    .B2(_0008_),
    .A2(_0994_),
    .A1(_0020_));
 sg13g2_nor3_2 _1908_ (.A(_0844_),
    .B(net306),
    .C(_0945_),
    .Y(_0997_));
 sg13g2_nor2_2 _1909_ (.A(_0898_),
    .B(_0976_),
    .Y(_0998_));
 sg13g2_nor3_1 _1910_ (.A(_0821_),
    .B(_0898_),
    .C(_0976_),
    .Y(_0999_));
 sg13g2_a221oi_1 _1911_ (.B2(_0842_),
    .C1(_0999_),
    .B1(_0997_),
    .A1(net349),
    .Y(_1000_),
    .A2(_0971_));
 sg13g2_nand4_1 _1912_ (.B(_0993_),
    .C(_0996_),
    .A(_0990_),
    .Y(_1001_),
    .D(_1000_));
 sg13g2_nor2_1 _1913_ (.A(net289),
    .B(_1001_),
    .Y(_1002_));
 sg13g2_nand2b_1 _1914_ (.Y(_1003_),
    .B(_0926_),
    .A_N(_0930_));
 sg13g2_nor3_1 _1915_ (.A(net316),
    .B(net306),
    .C(_0953_),
    .Y(_1004_));
 sg13g2_a221oi_1 _1916_ (.B2(_0949_),
    .C1(_1004_),
    .B1(_0947_),
    .A1(_0940_),
    .Y(_1005_),
    .A2(_0941_));
 sg13g2_a22oi_1 _1917_ (.Y(_1006_),
    .B1(_0932_),
    .B2(_0936_),
    .A2(_0924_),
    .A1(_0914_));
 sg13g2_nand3_1 _1918_ (.B(_1005_),
    .C(_1006_),
    .A(_1003_),
    .Y(_1007_));
 sg13g2_nor2b_1 _1919_ (.A(_0910_),
    .B_N(_0912_),
    .Y(_1008_));
 sg13g2_nand3_1 _1920_ (.B(_0904_),
    .C(_0907_),
    .A(net337),
    .Y(_1009_));
 sg13g2_o21ai_1 _1921_ (.B1(_1009_),
    .Y(_1010_),
    .A1(_0900_),
    .A2(_0901_));
 sg13g2_a21o_1 _1922_ (.A2(_0896_),
    .A1(_0881_),
    .B1(_1010_),
    .X(_1011_));
 sg13g2_nor3_1 _1923_ (.A(_1007_),
    .B(_1008_),
    .C(_1011_),
    .Y(_1012_));
 sg13g2_o21ai_1 _1924_ (.B1(_1002_),
    .Y(_1013_),
    .A1(\color_in[4] ),
    .A2(_1012_));
 sg13g2_a21oi_1 _1925_ (.A1(\color_in[4] ),
    .A2(_0959_),
    .Y(_1014_),
    .B1(_1013_));
 sg13g2_xnor2_1 _1926_ (.Y(_1015_),
    .A(net331),
    .B(_0933_));
 sg13g2_nor2_1 _1927_ (.A(net294),
    .B(_1015_),
    .Y(_1016_));
 sg13g2_a21oi_2 _1928_ (.B1(_1016_),
    .Y(_1017_),
    .A2(net294),
    .A1(_0803_));
 sg13g2_nand2b_1 _1929_ (.Y(_1018_),
    .B(_0894_),
    .A_N(_0886_));
 sg13g2_mux2_1 _1930_ (.A0(_1018_),
    .A1(_0003_),
    .S(net294),
    .X(_1019_));
 sg13g2_nand2_1 _1931_ (.Y(_1020_),
    .A(net359),
    .B(_1019_));
 sg13g2_xnor2_1 _1932_ (.Y(_1021_),
    .A(net359),
    .B(_1019_));
 sg13g2_nand2b_1 _1933_ (.Y(_1022_),
    .B(_0906_),
    .A_N(_1021_));
 sg13g2_nor2_1 _1934_ (.A(_0886_),
    .B(net294),
    .Y(_1023_));
 sg13g2_xnor2_1 _1935_ (.Y(_1024_),
    .A(_0801_),
    .B(_1023_));
 sg13g2_xor2_1 _1936_ (.B(_1024_),
    .A(_0016_),
    .X(_1025_));
 sg13g2_a21o_1 _1937_ (.A2(_1022_),
    .A1(_1020_),
    .B1(_1025_),
    .X(_1026_));
 sg13g2_nand2_1 _1938_ (.Y(_1027_),
    .A(net357),
    .B(_1024_));
 sg13g2_xnor2_1 _1939_ (.Y(_1028_),
    .A(net355),
    .B(_1017_));
 sg13g2_a21oi_1 _1940_ (.A1(_1026_),
    .A2(_1027_),
    .Y(_1029_),
    .B1(_1028_));
 sg13g2_a21oi_1 _1941_ (.A1(net355),
    .A2(_1017_),
    .Y(_1030_),
    .B1(_1029_));
 sg13g2_nor2_1 _1942_ (.A(_0804_),
    .B(_0887_),
    .Y(_1031_));
 sg13g2_nor3_1 _1943_ (.A(_0927_),
    .B(_0965_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_a21oi_2 _1944_ (.B1(_1032_),
    .Y(_1033_),
    .A2(net294),
    .A1(_0806_));
 sg13g2_nand2_1 _1945_ (.Y(_1034_),
    .A(net354),
    .B(_1033_));
 sg13g2_xnor2_1 _1946_ (.Y(_1035_),
    .A(_0821_),
    .B(_1033_));
 sg13g2_nand2b_1 _1947_ (.Y(_1036_),
    .B(_1030_),
    .A_N(_1035_));
 sg13g2_nand2b_1 _1948_ (.Y(_1037_),
    .B(_1035_),
    .A_N(_1030_));
 sg13g2_nand3_1 _1949_ (.B(_1036_),
    .C(_1037_),
    .A(_0966_),
    .Y(_1038_));
 sg13g2_nand2_1 _1950_ (.Y(_1039_),
    .A(_0010_),
    .B(_0977_));
 sg13g2_nor2_2 _1951_ (.A(net327),
    .B(net323),
    .Y(_1040_));
 sg13g2_nand2_1 _1952_ (.Y(_1041_),
    .A(_0009_),
    .B(_1040_));
 sg13g2_xnor2_1 _1953_ (.Y(_1042_),
    .A(_0815_),
    .B(_1041_));
 sg13g2_o21ai_1 _1954_ (.B1(_1039_),
    .Y(_1043_),
    .A1(_0977_),
    .A2(_1042_));
 sg13g2_and2_1 _1955_ (.A(net345),
    .B(_1043_),
    .X(_1044_));
 sg13g2_nor2_1 _1956_ (.A(_0977_),
    .B(_1040_),
    .Y(_1045_));
 sg13g2_nand2_1 _1957_ (.Y(_1046_),
    .A(\hvsync_gen.vpos[5] ),
    .B(net323));
 sg13g2_a22oi_1 _1958_ (.Y(_1047_),
    .B1(_1045_),
    .B2(_1046_),
    .A2(_0977_),
    .A1(_0813_));
 sg13g2_nand2_1 _1959_ (.Y(_1048_),
    .A(net348),
    .B(_1047_));
 sg13g2_xnor2_1 _1960_ (.Y(_1049_),
    .A(net348),
    .B(_1047_));
 sg13g2_or2_1 _1961_ (.X(_1050_),
    .B(_1049_),
    .A(_0948_));
 sg13g2_xnor2_1 _1962_ (.Y(_1051_),
    .A(_0009_),
    .B(_1045_));
 sg13g2_xnor2_1 _1963_ (.Y(_1052_),
    .A(_0021_),
    .B(_1051_));
 sg13g2_a21o_1 _1964_ (.A2(_1050_),
    .A1(_1048_),
    .B1(_1052_),
    .X(_1053_));
 sg13g2_nand2b_1 _1965_ (.Y(_1054_),
    .B(\hpos[7] ),
    .A_N(_1051_));
 sg13g2_xnor2_1 _1966_ (.Y(_1055_),
    .A(net345),
    .B(_1043_));
 sg13g2_a21oi_1 _1967_ (.A1(_1053_),
    .A2(_1054_),
    .Y(_1056_),
    .B1(_1055_));
 sg13g2_nand2_1 _1968_ (.Y(_1057_),
    .A(_0012_),
    .B(_0977_));
 sg13g2_nor4_2 _1969_ (.A(\hvsync_gen.vpos[5] ),
    .B(net323),
    .C(net320),
    .Y(_1058_),
    .D(net319));
 sg13g2_nand2b_1 _1970_ (.Y(_1059_),
    .B(_1058_),
    .A_N(\hvsync_gen.vpos[9] ));
 sg13g2_xnor2_1 _1971_ (.Y(_1060_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_1058_));
 sg13g2_o21ai_1 _1972_ (.B1(_1057_),
    .Y(_1061_),
    .A1(_0977_),
    .A2(_1060_));
 sg13g2_nand2_1 _1973_ (.Y(_1062_),
    .A(net343),
    .B(_1061_));
 sg13g2_xor2_1 _1974_ (.B(_1061_),
    .A(net343),
    .X(_1063_));
 sg13g2_nor3_1 _1975_ (.A(_1044_),
    .B(_1056_),
    .C(_1063_),
    .Y(_1064_));
 sg13g2_o21ai_1 _1976_ (.B1(_1063_),
    .Y(_1065_),
    .A1(_1044_),
    .A2(_1056_));
 sg13g2_nand2_1 _1977_ (.Y(_1066_),
    .A(_0979_),
    .B(_1065_));
 sg13g2_nor2_1 _1978_ (.A(_1064_),
    .B(_1066_),
    .Y(_1067_));
 sg13g2_nand2_1 _1979_ (.Y(_1068_),
    .A(_0007_),
    .B(_0980_));
 sg13g2_nand2_1 _1980_ (.Y(_1069_),
    .A(_0006_),
    .B(_0885_));
 sg13g2_xnor2_1 _1981_ (.Y(_1070_),
    .A(_0807_),
    .B(_1069_));
 sg13g2_o21ai_1 _1982_ (.B1(_1068_),
    .Y(_1071_),
    .A1(_0980_),
    .A2(_1070_));
 sg13g2_nand2_1 _1983_ (.Y(_1072_),
    .A(net351),
    .B(_1071_));
 sg13g2_nor2_1 _1984_ (.A(_0885_),
    .B(_0980_),
    .Y(_1073_));
 sg13g2_a22oi_1 _1985_ (.Y(_1074_),
    .B1(_1073_),
    .B2(_0893_),
    .A2(_0980_),
    .A1(_0803_));
 sg13g2_nand2_1 _1986_ (.Y(_1075_),
    .A(net356),
    .B(_1074_));
 sg13g2_xnor2_1 _1987_ (.Y(_1076_),
    .A(_0820_),
    .B(_1074_));
 sg13g2_nand2b_1 _1988_ (.Y(_1077_),
    .B(_1076_),
    .A_N(_0911_));
 sg13g2_xnor2_1 _1989_ (.Y(_1078_),
    .A(_0806_),
    .B(_1073_));
 sg13g2_xor2_1 _1990_ (.B(_1078_),
    .A(_0018_),
    .X(_1079_));
 sg13g2_a21oi_1 _1991_ (.A1(_1075_),
    .A2(_1077_),
    .Y(_1080_),
    .B1(_1079_));
 sg13g2_a21oi_1 _1992_ (.A1(net353),
    .A2(_1078_),
    .Y(_1081_),
    .B1(_1080_));
 sg13g2_xnor2_1 _1993_ (.Y(_1082_),
    .A(_0825_),
    .B(_1071_));
 sg13g2_nand2b_1 _1994_ (.Y(_1083_),
    .B(_1082_),
    .A_N(_1081_));
 sg13g2_nand2_1 _1995_ (.Y(_1084_),
    .A(_0810_),
    .B(_0919_));
 sg13g2_xnor2_1 _1996_ (.Y(_1085_),
    .A(_0810_),
    .B(_0919_));
 sg13g2_nor2_1 _1997_ (.A(_0980_),
    .B(_1085_),
    .Y(_1086_));
 sg13g2_a21oi_1 _1998_ (.A1(_0813_),
    .A2(_0980_),
    .Y(_1087_),
    .B1(_1086_));
 sg13g2_xnor2_1 _1999_ (.Y(_1088_),
    .A(net348),
    .B(_1087_));
 sg13g2_and3_1 _2000_ (.X(_1089_),
    .A(_1072_),
    .B(_1083_),
    .C(_1088_));
 sg13g2_a21oi_1 _2001_ (.A1(_1072_),
    .A2(_1083_),
    .Y(_1090_),
    .B1(_1088_));
 sg13g2_nor2_1 _2002_ (.A(_1089_),
    .B(_1090_),
    .Y(_1091_));
 sg13g2_nand2_1 _2003_ (.Y(_1092_),
    .A(net322),
    .B(_0918_));
 sg13g2_xnor2_1 _2004_ (.Y(_1093_),
    .A(net321),
    .B(_1092_));
 sg13g2_mux2_1 _2005_ (.A0(_0009_),
    .A1(_1093_),
    .S(_0962_),
    .X(_1094_));
 sg13g2_nand2_1 _2006_ (.Y(_1095_),
    .A(net347),
    .B(_1094_));
 sg13g2_nor2_1 _2007_ (.A(_0918_),
    .B(_0961_),
    .Y(_1096_));
 sg13g2_a22oi_1 _2008_ (.Y(_1097_),
    .B1(_1096_),
    .B2(_0921_),
    .A2(_0961_),
    .A1(_0809_));
 sg13g2_and2_1 _2009_ (.A(net351),
    .B(_1097_),
    .X(_1098_));
 sg13g2_xnor2_1 _2010_ (.Y(_1099_),
    .A(net351),
    .B(_1097_));
 sg13g2_nor2_1 _2011_ (.A(_0943_),
    .B(_1099_),
    .Y(_1100_));
 sg13g2_xnor2_1 _2012_ (.Y(_1101_),
    .A(net322),
    .B(_1096_));
 sg13g2_xor2_1 _2013_ (.B(_1101_),
    .A(_0020_),
    .X(_1102_));
 sg13g2_o21ai_1 _2014_ (.B1(_1102_),
    .Y(_1103_),
    .A1(_1098_),
    .A2(_1100_));
 sg13g2_nand2b_1 _2015_ (.Y(_1104_),
    .B(net348),
    .A_N(_1101_));
 sg13g2_xnor2_1 _2016_ (.Y(_1105_),
    .A(net347),
    .B(_1094_));
 sg13g2_a21o_1 _2017_ (.A2(_1104_),
    .A1(_1103_),
    .B1(_1105_),
    .X(_1106_));
 sg13g2_nand3_1 _2018_ (.B(_0814_),
    .C(_1040_),
    .A(_0804_),
    .Y(_1107_));
 sg13g2_nand2_1 _2019_ (.Y(_1108_),
    .A(_0804_),
    .B(_1058_));
 sg13g2_a21oi_1 _2020_ (.A1(net319),
    .A2(_1107_),
    .Y(_1109_),
    .B1(_0961_));
 sg13g2_a22oi_1 _2021_ (.Y(_1110_),
    .B1(_1108_),
    .B2(_1109_),
    .A2(_0961_),
    .A1(_0817_));
 sg13g2_xnor2_1 _2022_ (.Y(_1111_),
    .A(net345),
    .B(_1110_));
 sg13g2_a21oi_1 _2023_ (.A1(_1095_),
    .A2(_1106_),
    .Y(_1112_),
    .B1(_1111_));
 sg13g2_nand3_1 _2024_ (.B(_1106_),
    .C(_1111_),
    .A(_1095_),
    .Y(_1113_));
 sg13g2_nor2b_1 _2025_ (.A(_1112_),
    .B_N(_1113_),
    .Y(_1114_));
 sg13g2_nand2_1 _2026_ (.Y(_1115_),
    .A(net322),
    .B(_0967_));
 sg13g2_nand2_1 _2027_ (.Y(_1116_),
    .A(_0007_),
    .B(_0867_));
 sg13g2_xnor2_1 _2028_ (.Y(_1117_),
    .A(_0810_),
    .B(_1116_));
 sg13g2_o21ai_1 _2029_ (.B1(_1115_),
    .Y(_1118_),
    .A1(net293),
    .A2(_1117_));
 sg13g2_nand2_1 _2030_ (.Y(_1119_),
    .A(net348),
    .B(_1118_));
 sg13g2_nor2_1 _2031_ (.A(_0867_),
    .B(net293),
    .Y(_1120_));
 sg13g2_nand2_1 _2032_ (.Y(_1121_),
    .A(net332),
    .B(net328));
 sg13g2_a22oi_1 _2033_ (.Y(_1122_),
    .B1(_1120_),
    .B2(_1121_),
    .A2(net293),
    .A1(_0806_));
 sg13g2_nand2_1 _2034_ (.Y(_1123_),
    .A(net353),
    .B(_1122_));
 sg13g2_xnor2_1 _2035_ (.Y(_1124_),
    .A(_0821_),
    .B(_1122_));
 sg13g2_nand2_1 _2036_ (.Y(_1125_),
    .A(_0952_),
    .B(_1124_));
 sg13g2_xnor2_1 _2037_ (.Y(_1126_),
    .A(_0809_),
    .B(_1120_));
 sg13g2_xor2_1 _2038_ (.B(_1126_),
    .A(_0019_),
    .X(_1127_));
 sg13g2_a21o_1 _2039_ (.A2(_1125_),
    .A1(_1123_),
    .B1(_1127_),
    .X(_1128_));
 sg13g2_nand2_1 _2040_ (.Y(_1129_),
    .A(net351),
    .B(_1126_));
 sg13g2_xnor2_1 _2041_ (.Y(_1130_),
    .A(net348),
    .B(_1118_));
 sg13g2_a21o_1 _2042_ (.A2(_1129_),
    .A1(_1128_),
    .B1(_1130_),
    .X(_1131_));
 sg13g2_a21oi_1 _2043_ (.A1(_0867_),
    .A2(_1040_),
    .Y(_1132_),
    .B1(_0814_));
 sg13g2_nand3_1 _2044_ (.B(_0867_),
    .C(_1040_),
    .A(_0814_),
    .Y(_1133_));
 sg13g2_nor2_1 _2045_ (.A(net293),
    .B(_1132_),
    .Y(_1134_));
 sg13g2_nor3_1 _2046_ (.A(_0009_),
    .B(_0846_),
    .C(_0875_),
    .Y(_1135_));
 sg13g2_a21o_1 _2047_ (.A2(_1134_),
    .A1(_1133_),
    .B1(_1135_),
    .X(_1136_));
 sg13g2_xnor2_1 _2048_ (.Y(_1137_),
    .A(_0830_),
    .B(_1136_));
 sg13g2_nand3_1 _2049_ (.B(_1131_),
    .C(_1137_),
    .A(_1119_),
    .Y(_1138_));
 sg13g2_a21o_1 _2050_ (.A2(_1131_),
    .A1(_1119_),
    .B1(_1137_),
    .X(_1139_));
 sg13g2_nand3_1 _2051_ (.B(_1138_),
    .C(_1139_),
    .A(_0970_),
    .Y(_1140_));
 sg13g2_a221oi_1 _2052_ (.B2(_0964_),
    .C1(_1067_),
    .B1(_1114_),
    .A1(_0982_),
    .Y(_1141_),
    .A2(_1091_));
 sg13g2_and4_1 _2053_ (.A(_0879_),
    .B(_1014_),
    .C(_1038_),
    .D(_1140_),
    .X(_1142_));
 sg13g2_nand2b_1 _2054_ (.Y(_1143_),
    .B(net358),
    .A_N(\hdisplay[2] ));
 sg13g2_a22oi_1 _2055_ (.Y(_1144_),
    .B1(_0819_),
    .B2(\hdisplay[1] ),
    .A2(\hdisplay[0] ),
    .A1(_0795_));
 sg13g2_o21ai_1 _2056_ (.B1(_1143_),
    .Y(_1145_),
    .A1(_0819_),
    .A2(\hdisplay[1] ));
 sg13g2_nand2b_1 _2057_ (.Y(_1146_),
    .B(\hdisplay[2] ),
    .A_N(net358));
 sg13g2_o21ai_1 _2058_ (.B1(_1146_),
    .Y(_1147_),
    .A1(_1144_),
    .A2(_1145_));
 sg13g2_o21ai_1 _2059_ (.B1(_1147_),
    .Y(_1148_),
    .A1(_0820_),
    .A2(\hdisplay[3] ));
 sg13g2_a22oi_1 _2060_ (.Y(_1149_),
    .B1(_0821_),
    .B2(\hdisplay[4] ),
    .A2(\hdisplay[3] ),
    .A1(_0820_));
 sg13g2_nor2_1 _2061_ (.A(_0825_),
    .B(\hdisplay[5] ),
    .Y(_1150_));
 sg13g2_a221oi_1 _2062_ (.B2(_1149_),
    .C1(_1150_),
    .B1(_1148_),
    .A1(net354),
    .Y(_1151_),
    .A2(_0823_));
 sg13g2_a221oi_1 _2063_ (.B2(\hdisplay[6] ),
    .C1(_1151_),
    .B1(_0828_),
    .A1(_0825_),
    .Y(_1152_),
    .A2(\hdisplay[5] ));
 sg13g2_nand2b_1 _2064_ (.Y(_1153_),
    .B(net347),
    .A_N(\hdisplay[7] ));
 sg13g2_o21ai_1 _2065_ (.B1(_1153_),
    .Y(_1154_),
    .A1(_0828_),
    .A2(\hdisplay[6] ));
 sg13g2_a22oi_1 _2066_ (.Y(_1155_),
    .B1(_0832_),
    .B2(\hdisplay[8] ),
    .A2(\hdisplay[7] ),
    .A1(_0830_));
 sg13g2_o21ai_1 _2067_ (.B1(_1155_),
    .Y(_1156_),
    .A1(_1152_),
    .A2(_1154_));
 sg13g2_a22oi_1 _2068_ (.Y(_1157_),
    .B1(_0835_),
    .B2(net344),
    .A2(_0834_),
    .A1(net346));
 sg13g2_a22oi_1 _2069_ (.Y(_1158_),
    .B1(_1156_),
    .B2(_1157_),
    .A2(\hdisplay[10] ),
    .A1(_0836_));
 sg13g2_o21ai_1 _2070_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_0835_),
    .A2(net344));
 sg13g2_nor2_1 _2071_ (.A(_0814_),
    .B(\hvsync_gen.vdisplay[7] ),
    .Y(_1160_));
 sg13g2_a22oi_1 _2072_ (.Y(_1161_),
    .B1(_0797_),
    .B2(\hvsync_gen.vdisplay[1] ),
    .A2(\hvsync_gen.vdisplay[0] ),
    .A1(_0794_));
 sg13g2_nand2b_1 _2073_ (.Y(_1162_),
    .B(net333),
    .A_N(\hvsync_gen.vdisplay[2] ));
 sg13g2_o21ai_1 _2074_ (.B1(_1162_),
    .Y(_1163_),
    .A1(_0797_),
    .A2(\hvsync_gen.vdisplay[1] ));
 sg13g2_nor2_1 _2075_ (.A(_1161_),
    .B(_1163_),
    .Y(_1164_));
 sg13g2_a221oi_1 _2076_ (.B2(\hvsync_gen.vdisplay[3] ),
    .C1(_1164_),
    .B1(_0802_),
    .A1(_0800_),
    .Y(_1165_),
    .A2(\hvsync_gen.vdisplay[2] ));
 sg13g2_nand2b_1 _2077_ (.Y(_1166_),
    .B(net329),
    .A_N(\hvsync_gen.vdisplay[4] ));
 sg13g2_o21ai_1 _2078_ (.B1(_1166_),
    .Y(_1167_),
    .A1(_0802_),
    .A2(\hvsync_gen.vdisplay[3] ));
 sg13g2_a22oi_1 _2079_ (.Y(_1168_),
    .B1(_0807_),
    .B2(\hvsync_gen.vdisplay[5] ),
    .A2(\hvsync_gen.vdisplay[4] ),
    .A1(_0804_));
 sg13g2_o21ai_1 _2080_ (.B1(_1168_),
    .Y(_1169_),
    .A1(_1165_),
    .A2(_1167_));
 sg13g2_a22oi_1 _2081_ (.Y(_1170_),
    .B1(net323),
    .B2(_0811_),
    .A2(_0808_),
    .A1(net327));
 sg13g2_a22oi_1 _2082_ (.Y(_1171_),
    .B1(_1169_),
    .B2(_1170_),
    .A2(\hvsync_gen.vdisplay[6] ),
    .A1(_0810_));
 sg13g2_a22oi_1 _2083_ (.Y(_1172_),
    .B1(_0815_),
    .B2(\hvsync_gen.vdisplay[8] ),
    .A2(\hvsync_gen.vdisplay[7] ),
    .A1(_0814_));
 sg13g2_o21ai_1 _2084_ (.B1(_1172_),
    .Y(_1173_),
    .A1(_1160_),
    .A2(_1171_));
 sg13g2_a22oi_1 _2085_ (.Y(_1174_),
    .B1(net318),
    .B2(_0818_),
    .A2(_0816_),
    .A1(\hvsync_gen.vpos[8] ));
 sg13g2_and2_1 _2086_ (.A(_1173_),
    .B(_1174_),
    .X(_1175_));
 sg13g2_nor2b_1 _2087_ (.A(\hvsync_gen.vdisplay[10] ),
    .B_N(\hvsync_gen.vpos[10] ),
    .Y(_1176_));
 sg13g2_nor2b_1 _2088_ (.A(\hvsync_gen.vpos[10] ),
    .B_N(\hvsync_gen.vdisplay[10] ),
    .Y(_1177_));
 sg13g2_o21ai_1 _2089_ (.B1(_0014_),
    .Y(_1178_),
    .A1(net318),
    .A2(_0818_));
 sg13g2_nor4_1 _2090_ (.A(_1175_),
    .B(_1176_),
    .C(_1177_),
    .D(_1178_),
    .Y(_1179_));
 sg13g2_o21ai_1 _2091_ (.B1(_0024_),
    .Y(_1180_),
    .A1(_0836_),
    .A2(\hdisplay[10] ));
 sg13g2_nor4_2 _2092_ (.A(\hvsync_gen.vpos[11] ),
    .B(_1176_),
    .C(_1179_),
    .Y(_1181_),
    .D(_1180_));
 sg13g2_nand2_2 _2093_ (.Y(_1182_),
    .A(_1159_),
    .B(_1181_));
 sg13g2_a221oi_1 _2094_ (.B2(_1142_),
    .C1(_1182_),
    .B1(_1141_),
    .A1(_0842_),
    .Y(uo_out[4]),
    .A2(net289));
 sg13g2_nor3_1 _2095_ (.A(_0997_),
    .B(_1007_),
    .C(_1008_),
    .Y(_1183_));
 sg13g2_nor2b_2 _2096_ (.A(_1011_),
    .B_N(_1183_),
    .Y(_1184_));
 sg13g2_a21oi_1 _2097_ (.A1(_0909_),
    .A2(_0958_),
    .Y(_1185_),
    .B1(_0843_));
 sg13g2_a22oi_1 _2098_ (.Y(_1186_),
    .B1(_0998_),
    .B2(net328),
    .A2(_0992_),
    .A1(net327));
 sg13g2_a22oi_1 _2099_ (.Y(_1187_),
    .B1(_0989_),
    .B2(net321),
    .A2(_0971_),
    .A1(net325));
 sg13g2_a22oi_1 _2100_ (.Y(_1188_),
    .B1(_0991_),
    .B2(net334),
    .A2(_0988_),
    .A1(net331));
 sg13g2_nand4_1 _2101_ (.B(_1186_),
    .C(_1187_),
    .A(_0996_),
    .Y(_1189_),
    .D(_1188_));
 sg13g2_nor3_1 _2102_ (.A(net289),
    .B(_1185_),
    .C(_1189_),
    .Y(_1190_));
 sg13g2_o21ai_1 _2103_ (.B1(_1190_),
    .Y(_1191_),
    .A1(\color_in[5] ),
    .A2(_1184_));
 sg13g2_nand2_1 _2104_ (.Y(_1192_),
    .A(_1034_),
    .B(_1037_));
 sg13g2_a21oi_1 _2105_ (.A1(net326),
    .A2(_0928_),
    .Y(_1193_),
    .B1(net294));
 sg13g2_a22oi_1 _2106_ (.Y(_1194_),
    .B1(_1193_),
    .B2(_0920_),
    .A2(net294),
    .A1(_0809_));
 sg13g2_xnor2_1 _2107_ (.Y(_1195_),
    .A(net351),
    .B(_1194_));
 sg13g2_xnor2_1 _2108_ (.Y(_1196_),
    .A(_1192_),
    .B(_1195_));
 sg13g2_a21oi_1 _2109_ (.A1(net345),
    .A2(_1110_),
    .Y(_1197_),
    .B1(_1112_));
 sg13g2_xnor2_1 _2110_ (.Y(_1198_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_1108_));
 sg13g2_mux2_1 _2111_ (.A0(_0012_),
    .A1(_1198_),
    .S(_0962_),
    .X(_1199_));
 sg13g2_xor2_1 _2112_ (.B(_1199_),
    .A(net343),
    .X(_1200_));
 sg13g2_xnor2_1 _2113_ (.Y(_1201_),
    .A(_1197_),
    .B(_1200_));
 sg13g2_a21oi_1 _2114_ (.A1(net348),
    .A2(_1087_),
    .Y(_1202_),
    .B1(_1090_));
 sg13g2_xnor2_1 _2115_ (.Y(_1203_),
    .A(net321),
    .B(_1084_));
 sg13g2_mux2_1 _2116_ (.A0(_1203_),
    .A1(_0009_),
    .S(_0980_),
    .X(_1204_));
 sg13g2_xnor2_1 _2117_ (.Y(_1205_),
    .A(_0830_),
    .B(_1204_));
 sg13g2_xnor2_1 _2118_ (.Y(_1206_),
    .A(_1202_),
    .B(_1205_));
 sg13g2_o21ai_1 _2119_ (.B1(_1139_),
    .Y(_1207_),
    .A1(_0830_),
    .A2(_1136_));
 sg13g2_nand2_1 _2120_ (.Y(_1208_),
    .A(net319),
    .B(_1133_));
 sg13g2_a21oi_1 _2121_ (.A1(_0867_),
    .A2(_1058_),
    .Y(_1209_),
    .B1(net293));
 sg13g2_a22oi_1 _2122_ (.Y(_1210_),
    .B1(_1208_),
    .B2(_1209_),
    .A2(net293),
    .A1(_0817_));
 sg13g2_xnor2_1 _2123_ (.Y(_1211_),
    .A(net345),
    .B(_1210_));
 sg13g2_xnor2_1 _2124_ (.Y(_1212_),
    .A(_1207_),
    .B(_1211_));
 sg13g2_nand2_1 _2125_ (.Y(_1213_),
    .A(_0872_),
    .B(_0874_));
 sg13g2_nand3_1 _2126_ (.B(net324),
    .C(_0868_),
    .A(_0807_),
    .Y(_1214_));
 sg13g2_a21o_1 _2127_ (.A2(_0868_),
    .A1(_0807_),
    .B1(net324),
    .X(_1215_));
 sg13g2_a21oi_1 _2128_ (.A1(_1214_),
    .A2(_1215_),
    .Y(_1216_),
    .B1(net295));
 sg13g2_a21oi_1 _2129_ (.A1(_0813_),
    .A2(net295),
    .Y(_1217_),
    .B1(_1216_));
 sg13g2_xnor2_1 _2130_ (.Y(_1218_),
    .A(net348),
    .B(_1217_));
 sg13g2_xnor2_1 _2131_ (.Y(_1219_),
    .A(_1213_),
    .B(_1218_));
 sg13g2_nand2_1 _2132_ (.Y(_1220_),
    .A(_1062_),
    .B(_1065_));
 sg13g2_xnor2_1 _2133_ (.Y(_1221_),
    .A(\hvsync_gen.vpos[10] ),
    .B(_1059_));
 sg13g2_mux2_1 _2134_ (.A0(_0013_),
    .A1(_1221_),
    .S(_0978_),
    .X(_1222_));
 sg13g2_xnor2_1 _2135_ (.Y(_1223_),
    .A(\hpos[10] ),
    .B(_1222_));
 sg13g2_xnor2_1 _2136_ (.Y(_1224_),
    .A(_1220_),
    .B(_1223_));
 sg13g2_a22oi_1 _2137_ (.Y(_1225_),
    .B1(_1219_),
    .B2(_0877_),
    .A2(_1212_),
    .A1(_0970_));
 sg13g2_a221oi_1 _2138_ (.B2(_0982_),
    .C1(_1191_),
    .B1(_1206_),
    .A1(_0966_),
    .Y(_1226_),
    .A2(_1196_));
 sg13g2_a22oi_1 _2139_ (.Y(_1227_),
    .B1(_1224_),
    .B2(_0979_),
    .A2(_1201_),
    .A1(_0964_));
 sg13g2_and2_1 _2140_ (.A(_1225_),
    .B(_1227_),
    .X(_1228_));
 sg13g2_a221oi_1 _2141_ (.B2(_1228_),
    .C1(_1182_),
    .B1(_1226_),
    .A1(_0843_),
    .Y(uo_out[0]),
    .A2(net289));
 sg13g2_nand3_1 _2142_ (.B(_1125_),
    .C(_1127_),
    .A(_1123_),
    .Y(_1229_));
 sg13g2_and2_1 _2143_ (.A(_1128_),
    .B(_1229_),
    .X(_1230_));
 sg13g2_nand3_1 _2144_ (.B(_1077_),
    .C(_1079_),
    .A(_1075_),
    .Y(_1231_));
 sg13g2_nor2b_1 _2145_ (.A(_1080_),
    .B_N(_1231_),
    .Y(_1232_));
 sg13g2_nand3_1 _2146_ (.B(_1050_),
    .C(_1052_),
    .A(_1048_),
    .Y(_1233_));
 sg13g2_and2_1 _2147_ (.A(_1053_),
    .B(_1233_),
    .X(_1234_));
 sg13g2_a22oi_1 _2148_ (.Y(_1235_),
    .B1(_1234_),
    .B2(_0979_),
    .A2(_1232_),
    .A1(_0982_));
 sg13g2_nand3_1 _2149_ (.B(_1022_),
    .C(_1025_),
    .A(_1020_),
    .Y(_1236_));
 sg13g2_and2_1 _2150_ (.A(_1026_),
    .B(_1236_),
    .X(_1237_));
 sg13g2_a221oi_1 _2151_ (.B2(_0009_),
    .C1(_0987_),
    .B1(_0995_),
    .A1(_0830_),
    .Y(_1238_),
    .A2(_0994_));
 sg13g2_a22oi_1 _2152_ (.Y(_1239_),
    .B1(_0992_),
    .B2(net332),
    .A2(_0989_),
    .A1(net326));
 sg13g2_a22oi_1 _2153_ (.Y(_1240_),
    .B1(_0998_),
    .B2(net334),
    .A2(_0971_),
    .A1(net328));
 sg13g2_a22oi_1 _2154_ (.Y(_1241_),
    .B1(_0991_),
    .B2(net336),
    .A2(_0988_),
    .A1(\hvsync_gen.vpos[1] ));
 sg13g2_nand4_1 _2155_ (.B(_1239_),
    .C(_1240_),
    .A(_1238_),
    .Y(_1242_),
    .D(_1241_));
 sg13g2_nand3_1 _2156_ (.B(_0860_),
    .C(_0862_),
    .A(_0857_),
    .Y(_1243_));
 sg13g2_and2_1 _2157_ (.A(_0863_),
    .B(_0877_),
    .X(_1244_));
 sg13g2_or3_1 _2158_ (.A(_1098_),
    .B(_1100_),
    .C(_1102_),
    .X(_1245_));
 sg13g2_nand3_1 _2159_ (.B(_1103_),
    .C(_1245_),
    .A(_0964_),
    .Y(_1246_));
 sg13g2_o21ai_1 _2160_ (.B1(_1246_),
    .Y(_1247_),
    .A1(\color_in[2] ),
    .A2(_1184_));
 sg13g2_a221oi_1 _2161_ (.B2(_1244_),
    .C1(_1247_),
    .B1(_1243_),
    .A1(_0970_),
    .Y(_1248_),
    .A2(_1230_));
 sg13g2_a221oi_1 _2162_ (.B2(_1237_),
    .C1(_1242_),
    .B1(_0966_),
    .A1(\color_in[2] ),
    .Y(_1249_),
    .A2(_0959_));
 sg13g2_and2_1 _2163_ (.A(_1235_),
    .B(_1249_),
    .X(_1250_));
 sg13g2_a221oi_1 _2164_ (.B2(_1250_),
    .C1(_1182_),
    .B1(_1248_),
    .A1(_0029_),
    .Y(uo_out[5]),
    .A2(_0987_));
 sg13g2_nand3_1 _2165_ (.B(_1104_),
    .C(_1105_),
    .A(_1103_),
    .Y(_1251_));
 sg13g2_nand3_1 _2166_ (.B(_1106_),
    .C(_1251_),
    .A(_0964_),
    .Y(_1252_));
 sg13g2_nand3_1 _2167_ (.B(_1027_),
    .C(_1028_),
    .A(_1026_),
    .Y(_1253_));
 sg13g2_nand2_1 _2168_ (.Y(_1254_),
    .A(_0966_),
    .B(_1253_));
 sg13g2_or2_1 _2169_ (.X(_1255_),
    .B(_1254_),
    .A(_1029_));
 sg13g2_or2_1 _2170_ (.X(_1256_),
    .B(_1184_),
    .A(\color_in[3] ));
 sg13g2_a22oi_1 _2171_ (.Y(_1257_),
    .B1(_0992_),
    .B2(net328),
    .A2(_0989_),
    .A1(net325));
 sg13g2_a22oi_1 _2172_ (.Y(_1258_),
    .B1(_0991_),
    .B2(net335),
    .A2(_0988_),
    .A1(net334));
 sg13g2_a22oi_1 _2173_ (.Y(_1259_),
    .B1(_0998_),
    .B2(net332),
    .A2(_0971_),
    .A1(net326));
 sg13g2_nand4_1 _2174_ (.B(_1257_),
    .C(_1258_),
    .A(_1238_),
    .Y(_1260_),
    .D(_1259_));
 sg13g2_a21oi_1 _2175_ (.A1(\color_in[3] ),
    .A2(_0959_),
    .Y(_1261_),
    .B1(_1260_));
 sg13g2_nand4_1 _2176_ (.B(_1255_),
    .C(_1256_),
    .A(_1252_),
    .Y(_1262_),
    .D(_1261_));
 sg13g2_nand2b_1 _2177_ (.Y(_1263_),
    .B(_1081_),
    .A_N(_1082_));
 sg13g2_nand3_1 _2178_ (.B(_1083_),
    .C(_1263_),
    .A(_0982_),
    .Y(_1264_));
 sg13g2_nand3_1 _2179_ (.B(_1054_),
    .C(_1055_),
    .A(_1053_),
    .Y(_1265_));
 sg13g2_nand2_1 _2180_ (.Y(_1266_),
    .A(_0979_),
    .B(_1265_));
 sg13g2_o21ai_1 _2181_ (.B1(_1264_),
    .Y(_1267_),
    .A1(_1056_),
    .A2(_1266_));
 sg13g2_nand3_1 _2182_ (.B(_1129_),
    .C(_1130_),
    .A(_1128_),
    .Y(_1268_));
 sg13g2_nand3_1 _2183_ (.B(_1131_),
    .C(_1268_),
    .A(_0970_),
    .Y(_1269_));
 sg13g2_nand3_1 _2184_ (.B(_0864_),
    .C(_0865_),
    .A(_0863_),
    .Y(_1270_));
 sg13g2_and3_1 _2185_ (.X(_1271_),
    .A(_0866_),
    .B(_0877_),
    .C(_1270_));
 sg13g2_nor3_1 _2186_ (.A(_1262_),
    .B(_1267_),
    .C(_1271_),
    .Y(_1272_));
 sg13g2_a221oi_1 _2187_ (.B2(_1272_),
    .C1(_1182_),
    .B1(_1269_),
    .A1(_0030_),
    .Y(uo_out[1]),
    .A2(net289));
 sg13g2_a22oi_1 _2188_ (.Y(_1273_),
    .B1(_0995_),
    .B2(_0007_),
    .A2(_0994_),
    .A1(_0825_));
 sg13g2_o21ai_1 _2189_ (.B1(_1273_),
    .Y(_1274_),
    .A1(_0953_),
    .A2(_0969_));
 sg13g2_nand2_1 _2190_ (.Y(_1275_),
    .A(_0944_),
    .B(_0964_));
 sg13g2_a22oi_1 _2191_ (.Y(_1276_),
    .B1(_0998_),
    .B2(net357),
    .A2(_0991_),
    .A1(\hpos[0] ));
 sg13g2_a22oi_1 _2192_ (.Y(_1277_),
    .B1(_0982_),
    .B2(_0912_),
    .A2(_0913_),
    .A1(\color_in[0] ));
 sg13g2_a22oi_1 _2193_ (.Y(_1278_),
    .B1(_0992_),
    .B2(net355),
    .A2(_0971_),
    .A1(net353));
 sg13g2_a21oi_1 _2194_ (.A1(_0877_),
    .A2(_0902_),
    .Y(_1279_),
    .B1(_1274_));
 sg13g2_a22oi_1 _2195_ (.Y(_1280_),
    .B1(_0989_),
    .B2(net350),
    .A2(_0988_),
    .A1(\hpos[1] ));
 sg13g2_and4_1 _2196_ (.A(_1275_),
    .B(_1276_),
    .C(_1278_),
    .D(_1280_),
    .X(_1281_));
 sg13g2_a22oi_1 _2197_ (.Y(_1282_),
    .B1(_0979_),
    .B2(_0949_),
    .A2(_0966_),
    .A1(_0907_));
 sg13g2_nand4_1 _2198_ (.B(_1279_),
    .C(_1281_),
    .A(_1277_),
    .Y(_1283_),
    .D(_1282_));
 sg13g2_nand2b_1 _2199_ (.Y(_1284_),
    .B(_0909_),
    .A_N(net289));
 sg13g2_o21ai_1 _2200_ (.B1(\color_in[0] ),
    .Y(_1285_),
    .A1(_0957_),
    .A2(_1284_));
 sg13g2_o21ai_1 _2201_ (.B1(_1285_),
    .Y(_1286_),
    .A1(\color_in[0] ),
    .A2(_1184_));
 sg13g2_nor2_1 _2202_ (.A(_1283_),
    .B(_1286_),
    .Y(_1287_));
 sg13g2_nor2_2 _2203_ (.A(_1182_),
    .B(_1287_),
    .Y(uo_out[6]));
 sg13g2_or2_1 _2204_ (.X(_1288_),
    .B(_0859_),
    .A(_0858_));
 sg13g2_nand3_1 _2205_ (.B(_0877_),
    .C(_1288_),
    .A(_0860_),
    .Y(_1289_));
 sg13g2_xnor2_1 _2206_ (.Y(_1290_),
    .A(_0952_),
    .B(_1124_));
 sg13g2_o21ai_1 _2207_ (.B1(_1289_),
    .Y(_1291_),
    .A1(_0969_),
    .A2(_1290_));
 sg13g2_xor2_1 _2208_ (.B(_1049_),
    .A(_0948_),
    .X(_1292_));
 sg13g2_nor2_1 _2209_ (.A(\color_in[1] ),
    .B(_1011_),
    .Y(_1293_));
 sg13g2_a21oi_1 _2210_ (.A1(\color_in[1] ),
    .A2(_0909_),
    .Y(_1294_),
    .B1(_1293_));
 sg13g2_a22oi_1 _2211_ (.Y(_1295_),
    .B1(_0998_),
    .B2(net355),
    .A2(_0992_),
    .A1(net353));
 sg13g2_a22oi_1 _2212_ (.Y(_1296_),
    .B1(_0991_),
    .B2(net359),
    .A2(_0989_),
    .A1(net349));
 sg13g2_a22oi_1 _2213_ (.Y(_1297_),
    .B1(_0988_),
    .B2(net357),
    .A2(_0971_),
    .A1(net350));
 sg13g2_nand4_1 _2214_ (.B(_1295_),
    .C(_1296_),
    .A(_1273_),
    .Y(_1298_),
    .D(_1297_));
 sg13g2_nor3_1 _2215_ (.A(net289),
    .B(_1294_),
    .C(_1298_),
    .Y(_1299_));
 sg13g2_nand2b_1 _2216_ (.Y(_1300_),
    .B(_1021_),
    .A_N(_0906_));
 sg13g2_nand3_1 _2217_ (.B(_1022_),
    .C(_1300_),
    .A(_0966_),
    .Y(_1301_));
 sg13g2_xor2_1 _2218_ (.B(_1099_),
    .A(_0943_),
    .X(_1302_));
 sg13g2_xnor2_1 _2219_ (.Y(_1303_),
    .A(_0911_),
    .B(_1076_));
 sg13g2_mux2_1 _2220_ (.A0(_1183_),
    .A1(_0958_),
    .S(\color_in[1] ),
    .X(_1304_));
 sg13g2_a21oi_1 _2221_ (.A1(_0964_),
    .A2(_1302_),
    .Y(_1305_),
    .B1(_1291_));
 sg13g2_a22oi_1 _2222_ (.Y(_1306_),
    .B1(_1303_),
    .B2(_0982_),
    .A2(_1292_),
    .A1(_0979_));
 sg13g2_and4_1 _2223_ (.A(_1299_),
    .B(_1301_),
    .C(_1304_),
    .D(_1306_),
    .X(_1307_));
 sg13g2_a221oi_1 _2224_ (.B2(_1307_),
    .C1(_1182_),
    .B1(_1305_),
    .A1(_0028_),
    .Y(uo_out[2]),
    .A2(net289));
 sg13g2_o21ai_1 _2225_ (.B1(_0011_),
    .Y(_1308_),
    .A1(\hvsync_gen.vfrontporch[7] ),
    .A2(\hvsync_gen.vdisplay[7] ));
 sg13g2_nand2_1 _2226_ (.Y(_1309_),
    .A(\hvsync_gen.vdisplay[8] ),
    .B(\hvsync_gen.vdisplay[9] ));
 sg13g2_xor2_1 _2227_ (.B(\hvsync_gen.vdisplay[9] ),
    .A(\hvsync_gen.vdisplay[8] ),
    .X(_1310_));
 sg13g2_nor2_1 _2228_ (.A(_1308_),
    .B(_1310_),
    .Y(_1311_));
 sg13g2_inv_1 _2229_ (.Y(_1312_),
    .A(_1311_));
 sg13g2_xor2_1 _2230_ (.B(_1310_),
    .A(_1308_),
    .X(_1313_));
 sg13g2_or3_1 _2231_ (.A(\hvsync_gen.vfrontporch[7] ),
    .B(\hvsync_gen.vdisplay[7] ),
    .C(_0011_),
    .X(_1314_));
 sg13g2_and2_1 _2232_ (.A(_1308_),
    .B(_1314_),
    .X(_1315_));
 sg13g2_and2_1 _2233_ (.A(\hvsync_gen.vfrontporch[7] ),
    .B(\hvsync_gen.vdisplay[7] ),
    .X(_1316_));
 sg13g2_xor2_1 _2234_ (.B(\hvsync_gen.vdisplay[7] ),
    .A(\hvsync_gen.vfrontporch[7] ),
    .X(_1317_));
 sg13g2_nor2_1 _2235_ (.A(\hvsync_gen.vfrontporch[6] ),
    .B(\hvsync_gen.vdisplay[6] ),
    .Y(_1318_));
 sg13g2_nor2_1 _2236_ (.A(_1317_),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_xor2_1 _2237_ (.B(_1318_),
    .A(_1317_),
    .X(_1320_));
 sg13g2_a21oi_1 _2238_ (.A1(\hvsync_gen.vsynclength[7] ),
    .A2(_1320_),
    .Y(_1321_),
    .B1(_1319_));
 sg13g2_nor2b_1 _2239_ (.A(_1321_),
    .B_N(_1315_),
    .Y(_1322_));
 sg13g2_xnor2_1 _2240_ (.Y(_1323_),
    .A(_1315_),
    .B(_1321_));
 sg13g2_xnor2_1 _2241_ (.Y(_1324_),
    .A(\hvsync_gen.vsynclength[7] ),
    .B(_1320_));
 sg13g2_xnor2_1 _2242_ (.Y(_1325_),
    .A(\hvsync_gen.vfrontporch[6] ),
    .B(\hvsync_gen.vdisplay[6] ));
 sg13g2_nor2_1 _2243_ (.A(\hvsync_gen.vfrontporch[5] ),
    .B(\hvsync_gen.vdisplay[5] ),
    .Y(_1326_));
 sg13g2_o21ai_1 _2244_ (.B1(_1325_),
    .Y(_1327_),
    .A1(\hvsync_gen.vfrontporch[5] ),
    .A2(\hvsync_gen.vdisplay[5] ));
 sg13g2_xnor2_1 _2245_ (.Y(_1328_),
    .A(_1325_),
    .B(_1326_));
 sg13g2_nand2_1 _2246_ (.Y(_1329_),
    .A(\hvsync_gen.vsynclength[6] ),
    .B(_1328_));
 sg13g2_a21oi_1 _2247_ (.A1(_1327_),
    .A2(_1329_),
    .Y(_1330_),
    .B1(_1324_));
 sg13g2_nand3_1 _2248_ (.B(_1327_),
    .C(_1329_),
    .A(_1324_),
    .Y(_1331_));
 sg13g2_xnor2_1 _2249_ (.Y(_1332_),
    .A(\hvsync_gen.vsynclength[6] ),
    .B(_1328_));
 sg13g2_or2_1 _2250_ (.X(_1333_),
    .B(\hvsync_gen.vdisplay[4] ),
    .A(\hvsync_gen.vfrontporch[4] ));
 sg13g2_xnor2_1 _2251_ (.Y(_1334_),
    .A(\hvsync_gen.vfrontporch[5] ),
    .B(\hvsync_gen.vdisplay[5] ));
 sg13g2_and2_1 _2252_ (.A(_1333_),
    .B(_1334_),
    .X(_1335_));
 sg13g2_xor2_1 _2253_ (.B(_1334_),
    .A(_1333_),
    .X(_1336_));
 sg13g2_a21oi_1 _2254_ (.A1(\hvsync_gen.vsynclength[5] ),
    .A2(_1336_),
    .Y(_1337_),
    .B1(_1335_));
 sg13g2_or2_1 _2255_ (.X(_1338_),
    .B(_1337_),
    .A(_1332_));
 sg13g2_inv_1 _2256_ (.Y(_1339_),
    .A(_1338_));
 sg13g2_xnor2_1 _2257_ (.Y(_1340_),
    .A(_1332_),
    .B(_1337_));
 sg13g2_and2_1 _2258_ (.A(\hvsync_gen.vfrontporch[4] ),
    .B(\hvsync_gen.vdisplay[4] ),
    .X(_1341_));
 sg13g2_xnor2_1 _2259_ (.Y(_1342_),
    .A(\hvsync_gen.vfrontporch[4] ),
    .B(\hvsync_gen.vdisplay[4] ));
 sg13g2_nor2_1 _2260_ (.A(\hvsync_gen.vfrontporch[3] ),
    .B(\hvsync_gen.vdisplay[3] ),
    .Y(_1343_));
 sg13g2_o21ai_1 _2261_ (.B1(_1342_),
    .Y(_1344_),
    .A1(\hvsync_gen.vfrontporch[3] ),
    .A2(\hvsync_gen.vdisplay[3] ));
 sg13g2_xnor2_1 _2262_ (.Y(_1345_),
    .A(_1342_),
    .B(_1343_));
 sg13g2_nand2_1 _2263_ (.Y(_1346_),
    .A(\hvsync_gen.vsynclength[4] ),
    .B(_1345_));
 sg13g2_xnor2_1 _2264_ (.Y(_1347_),
    .A(\hvsync_gen.vsynclength[5] ),
    .B(_1336_));
 sg13g2_a21oi_2 _2265_ (.B1(_1347_),
    .Y(_1348_),
    .A2(_1346_),
    .A1(_1344_));
 sg13g2_inv_1 _2266_ (.Y(_1349_),
    .A(_1348_));
 sg13g2_nand3_1 _2267_ (.B(_1346_),
    .C(_1347_),
    .A(_1344_),
    .Y(_1350_));
 sg13g2_inv_1 _2268_ (.Y(_1351_),
    .A(_1350_));
 sg13g2_nor2b_2 _2269_ (.A(_1348_),
    .B_N(_1350_),
    .Y(_1352_));
 sg13g2_xnor2_1 _2270_ (.Y(_1353_),
    .A(\hvsync_gen.vsynclength[4] ),
    .B(_1345_));
 sg13g2_nand2_1 _2271_ (.Y(_1354_),
    .A(\hvsync_gen.vfrontporch[3] ),
    .B(\hvsync_gen.vdisplay[3] ));
 sg13g2_nand2b_2 _2272_ (.Y(_1355_),
    .B(_1354_),
    .A_N(_1343_));
 sg13g2_or2_1 _2273_ (.X(_1356_),
    .B(\hvsync_gen.vdisplay[2] ),
    .A(\hvsync_gen.vfrontporch[2] ));
 sg13g2_and2_1 _2274_ (.A(_1355_),
    .B(_1356_),
    .X(_1357_));
 sg13g2_xor2_1 _2275_ (.B(_1356_),
    .A(_1355_),
    .X(_1358_));
 sg13g2_a21oi_1 _2276_ (.A1(\hvsync_gen.vsynclength[3] ),
    .A2(_1358_),
    .Y(_1359_),
    .B1(_1357_));
 sg13g2_or2_1 _2277_ (.X(_1360_),
    .B(_1359_),
    .A(_1353_));
 sg13g2_xnor2_1 _2278_ (.Y(_1361_),
    .A(_1353_),
    .B(_1359_));
 sg13g2_xnor2_1 _2279_ (.Y(_1362_),
    .A(\hvsync_gen.vsynclength[3] ),
    .B(_1358_));
 sg13g2_and2_1 _2280_ (.A(\hvsync_gen.vfrontporch[2] ),
    .B(\hvsync_gen.vdisplay[2] ),
    .X(_1363_));
 sg13g2_xnor2_1 _2281_ (.Y(_1364_),
    .A(\hvsync_gen.vfrontporch[2] ),
    .B(\hvsync_gen.vdisplay[2] ));
 sg13g2_nor2_1 _2282_ (.A(\hvsync_gen.vfrontporch[1] ),
    .B(\hvsync_gen.vdisplay[1] ),
    .Y(_1365_));
 sg13g2_o21ai_1 _2283_ (.B1(_1364_),
    .Y(_1366_),
    .A1(\hvsync_gen.vfrontporch[1] ),
    .A2(\hvsync_gen.vdisplay[1] ));
 sg13g2_xnor2_1 _2284_ (.Y(_1367_),
    .A(_1364_),
    .B(_1365_));
 sg13g2_nand2_1 _2285_ (.Y(_1368_),
    .A(\hvsync_gen.vsynclength[2] ),
    .B(_1367_));
 sg13g2_and2_1 _2286_ (.A(_1366_),
    .B(_1368_),
    .X(_1369_));
 sg13g2_nor2_1 _2287_ (.A(_1362_),
    .B(_1369_),
    .Y(_1370_));
 sg13g2_xor2_1 _2288_ (.B(_1369_),
    .A(_1362_),
    .X(_1371_));
 sg13g2_xnor2_1 _2289_ (.Y(_1372_),
    .A(\hvsync_gen.vsynclength[2] ),
    .B(_1367_));
 sg13g2_nand2_1 _2290_ (.Y(_1373_),
    .A(\hvsync_gen.vfrontporch[1] ),
    .B(\hvsync_gen.vdisplay[1] ));
 sg13g2_xor2_1 _2291_ (.B(\hvsync_gen.vdisplay[1] ),
    .A(\hvsync_gen.vfrontporch[1] ),
    .X(_1374_));
 sg13g2_nor2_1 _2292_ (.A(\hvsync_gen.vfrontporch[0] ),
    .B(\hvsync_gen.vdisplay[0] ),
    .Y(_1375_));
 sg13g2_nor2_1 _2293_ (.A(_1374_),
    .B(_1375_),
    .Y(_1376_));
 sg13g2_xor2_1 _2294_ (.B(_1375_),
    .A(_1374_),
    .X(_1377_));
 sg13g2_a21oi_1 _2295_ (.A1(\hvsync_gen.vsynclength[1] ),
    .A2(_1377_),
    .Y(_1378_),
    .B1(_1376_));
 sg13g2_nor2_1 _2296_ (.A(_1372_),
    .B(_1378_),
    .Y(_1379_));
 sg13g2_xor2_1 _2297_ (.B(_1378_),
    .A(_1372_),
    .X(_1380_));
 sg13g2_nand2_1 _2298_ (.Y(_1381_),
    .A(\hvsync_gen.vfrontporch[0] ),
    .B(\hvsync_gen.vdisplay[0] ));
 sg13g2_xnor2_1 _2299_ (.Y(_1382_),
    .A(\hvsync_gen.vfrontporch[0] ),
    .B(\hvsync_gen.vdisplay[0] ));
 sg13g2_nand2_1 _2300_ (.Y(_1383_),
    .A(\hvsync_gen.vsynclength[0] ),
    .B(_1382_));
 sg13g2_xnor2_1 _2301_ (.Y(_1384_),
    .A(\hvsync_gen.vsynclength[1] ),
    .B(_1377_));
 sg13g2_nor2_1 _2302_ (.A(_1383_),
    .B(_1384_),
    .Y(_1385_));
 sg13g2_a21o_1 _2303_ (.A2(_1385_),
    .A1(_1380_),
    .B1(_1379_),
    .X(_1386_));
 sg13g2_a21oi_2 _2304_ (.B1(_1370_),
    .Y(_1387_),
    .A2(_1386_),
    .A1(_1371_));
 sg13g2_or4_1 _2305_ (.A(_1348_),
    .B(_1351_),
    .C(_1361_),
    .D(_1387_),
    .X(_1388_));
 sg13g2_o21ai_1 _2306_ (.B1(_1349_),
    .Y(_1389_),
    .A1(_1351_),
    .A2(_1360_));
 sg13g2_inv_1 _2307_ (.Y(_1390_),
    .A(_1389_));
 sg13g2_a21oi_2 _2308_ (.B1(_1340_),
    .Y(_1391_),
    .A2(_1390_),
    .A1(_1388_));
 sg13g2_nor2_1 _2309_ (.A(_1339_),
    .B(_1391_),
    .Y(_1392_));
 sg13g2_nand2b_1 _2310_ (.Y(_1393_),
    .B(_1338_),
    .A_N(_1330_));
 sg13g2_o21ai_1 _2311_ (.B1(_1331_),
    .Y(_1394_),
    .A1(_1391_),
    .A2(_1393_));
 sg13g2_nor2b_1 _2312_ (.A(_1394_),
    .B_N(_1323_),
    .Y(_1395_));
 sg13g2_nor2b_1 _2313_ (.A(_1310_),
    .B_N(_1322_),
    .Y(_1396_));
 sg13g2_or2_1 _2314_ (.X(_1397_),
    .B(_1396_),
    .A(_1311_));
 sg13g2_a21oi_2 _2315_ (.B1(_1397_),
    .Y(_1398_),
    .A2(_1395_),
    .A1(_1313_));
 sg13g2_nor3_2 _2316_ (.A(\hvsync_gen.vdisplay[8] ),
    .B(\hvsync_gen.vdisplay[9] ),
    .C(\hvsync_gen.vdisplay[10] ),
    .Y(_1399_));
 sg13g2_o21ai_1 _2317_ (.B1(\hvsync_gen.vdisplay[10] ),
    .Y(_1400_),
    .A1(\hvsync_gen.vdisplay[8] ),
    .A2(\hvsync_gen.vdisplay[9] ));
 sg13g2_inv_1 _2318_ (.Y(_1401_),
    .A(_1400_));
 sg13g2_nand2_1 _2319_ (.Y(_1402_),
    .A(_1398_),
    .B(_1399_));
 sg13g2_o21ai_1 _2320_ (.B1(_1402_),
    .Y(_1403_),
    .A1(_1398_),
    .A2(_1400_));
 sg13g2_nand2_1 _2321_ (.Y(_1404_),
    .A(net174),
    .B(_1403_));
 sg13g2_nor2_2 _2322_ (.A(_1399_),
    .B(_1401_),
    .Y(_1405_));
 sg13g2_xnor2_1 _2323_ (.Y(_1406_),
    .A(_1398_),
    .B(_1405_));
 sg13g2_nor2_1 _2324_ (.A(\hvsync_gen.vpos[10] ),
    .B(_1406_),
    .Y(_1407_));
 sg13g2_xor2_1 _2325_ (.B(_1406_),
    .A(_0013_),
    .X(_1408_));
 sg13g2_nor2_1 _2326_ (.A(_1313_),
    .B(_1322_),
    .Y(_1409_));
 sg13g2_or2_1 _2327_ (.X(_1410_),
    .B(_1409_),
    .A(_1396_));
 sg13g2_mux2_1 _2328_ (.A0(_1410_),
    .A1(_1313_),
    .S(_1395_),
    .X(_1411_));
 sg13g2_nand3_1 _2329_ (.B(_1388_),
    .C(_1390_),
    .A(_1340_),
    .Y(_1412_));
 sg13g2_nand2b_1 _2330_ (.Y(_1413_),
    .B(_1412_),
    .A_N(_1391_));
 sg13g2_xnor2_1 _2331_ (.Y(_1414_),
    .A(net322),
    .B(_1413_));
 sg13g2_o21ai_1 _2332_ (.B1(_1360_),
    .Y(_1415_),
    .A1(_1361_),
    .A2(_1387_));
 sg13g2_xnor2_1 _2333_ (.Y(_1416_),
    .A(_1352_),
    .B(_1415_));
 sg13g2_nor2_1 _2334_ (.A(net326),
    .B(_1416_),
    .Y(_1417_));
 sg13g2_xnor2_1 _2335_ (.Y(_1418_),
    .A(_1361_),
    .B(_1387_));
 sg13g2_xnor2_1 _2336_ (.Y(_1419_),
    .A(_1371_),
    .B(_1386_));
 sg13g2_xnor2_1 _2337_ (.Y(_1420_),
    .A(_1380_),
    .B(_1385_));
 sg13g2_xor2_1 _2338_ (.B(_1384_),
    .A(_1383_),
    .X(_1421_));
 sg13g2_xor2_1 _2339_ (.B(_1382_),
    .A(\hvsync_gen.vsynclength[0] ),
    .X(_1422_));
 sg13g2_nor3_1 _2340_ (.A(_0031_),
    .B(_0794_),
    .C(_1422_),
    .Y(_1423_));
 sg13g2_nand2b_1 _2341_ (.Y(_1424_),
    .B(_0003_),
    .A_N(_1423_));
 sg13g2_o21ai_1 _2342_ (.B1(net335),
    .Y(_1425_),
    .A1(_0003_),
    .A2(_1423_));
 sg13g2_nand2_1 _2343_ (.Y(_1426_),
    .A(_1421_),
    .B(_1425_));
 sg13g2_o21ai_1 _2344_ (.B1(_1426_),
    .Y(_1427_),
    .A1(_1421_),
    .A2(_1424_));
 sg13g2_xnor2_1 _2345_ (.Y(_1428_),
    .A(_0004_),
    .B(_1420_));
 sg13g2_nor2_1 _2346_ (.A(net333),
    .B(_1420_),
    .Y(_1429_));
 sg13g2_a21oi_1 _2347_ (.A1(_1427_),
    .A2(_1428_),
    .Y(_1430_),
    .B1(_1429_));
 sg13g2_a21oi_1 _2348_ (.A1(net330),
    .A2(_1419_),
    .Y(_1431_),
    .B1(_1430_));
 sg13g2_nor2_1 _2349_ (.A(net329),
    .B(_1418_),
    .Y(_1432_));
 sg13g2_nor2_1 _2350_ (.A(net330),
    .B(_1419_),
    .Y(_1433_));
 sg13g2_nor3_1 _2351_ (.A(_1431_),
    .B(_1432_),
    .C(_1433_),
    .Y(_1434_));
 sg13g2_a221oi_1 _2352_ (.B2(net329),
    .C1(_1434_),
    .B1(_1418_),
    .A1(net326),
    .Y(_1435_),
    .A2(_1416_));
 sg13g2_o21ai_1 _2353_ (.B1(_1414_),
    .Y(_1436_),
    .A1(_1417_),
    .A2(_1435_));
 sg13g2_nor2_1 _2354_ (.A(net323),
    .B(_1413_),
    .Y(_1437_));
 sg13g2_nand2b_1 _2355_ (.Y(_1438_),
    .B(_1331_),
    .A_N(_1330_));
 sg13g2_xor2_1 _2356_ (.B(_1438_),
    .A(_1392_),
    .X(_1439_));
 sg13g2_inv_1 _2357_ (.Y(_1440_),
    .A(_1439_));
 sg13g2_o21ai_1 _2358_ (.B1(_1436_),
    .Y(_1441_),
    .A1(net320),
    .A2(_1440_));
 sg13g2_xor2_1 _2359_ (.B(_1394_),
    .A(_1323_),
    .X(_1442_));
 sg13g2_a22oi_1 _2360_ (.Y(_1443_),
    .B1(_1442_),
    .B2(net319),
    .A2(_1440_),
    .A1(net320));
 sg13g2_o21ai_1 _2361_ (.B1(_1443_),
    .Y(_1444_),
    .A1(_1437_),
    .A2(_1441_));
 sg13g2_nor2_1 _2362_ (.A(net319),
    .B(_1442_),
    .Y(_1445_));
 sg13g2_nor2_1 _2363_ (.A(net318),
    .B(_1411_),
    .Y(_1446_));
 sg13g2_nor2_1 _2364_ (.A(_1445_),
    .B(_1446_),
    .Y(_1447_));
 sg13g2_a221oi_1 _2365_ (.B2(_1447_),
    .C1(_1408_),
    .B1(_1444_),
    .A1(net318),
    .Y(_1448_),
    .A2(_1411_));
 sg13g2_xnor2_1 _2366_ (.Y(_1449_),
    .A(\hvsync_gen.vpos[11] ),
    .B(_1403_));
 sg13g2_o21ai_1 _2367_ (.B1(_1449_),
    .Y(_1450_),
    .A1(_1407_),
    .A2(_1448_));
 sg13g2_o21ai_1 _2368_ (.B1(_1373_),
    .Y(_1451_),
    .A1(_1365_),
    .A2(_1381_));
 sg13g2_a21oi_1 _2369_ (.A1(_1356_),
    .A2(_1451_),
    .Y(_1452_),
    .B1(_1363_));
 sg13g2_o21ai_1 _2370_ (.B1(_1354_),
    .Y(_1453_),
    .A1(_1343_),
    .A2(_1452_));
 sg13g2_a21oi_1 _2371_ (.A1(_1333_),
    .A2(_1453_),
    .Y(_1454_),
    .B1(_1341_));
 sg13g2_a221oi_1 _2372_ (.B2(_1453_),
    .C1(_1341_),
    .B1(_1333_),
    .A1(\hvsync_gen.vfrontporch[5] ),
    .Y(_1455_),
    .A2(\hvsync_gen.vdisplay[5] ));
 sg13g2_nor3_1 _2373_ (.A(_1325_),
    .B(_1326_),
    .C(_1455_),
    .Y(_1456_));
 sg13g2_a21o_1 _2374_ (.A2(\hvsync_gen.vdisplay[6] ),
    .A1(\hvsync_gen.vfrontporch[6] ),
    .B1(_1456_),
    .X(_1457_));
 sg13g2_a21oi_2 _2375_ (.B1(_1316_),
    .Y(_1458_),
    .A2(_1457_),
    .A1(_1317_));
 sg13g2_nor2_1 _2376_ (.A(_1309_),
    .B(_1458_),
    .Y(_1459_));
 sg13g2_nor3_1 _2377_ (.A(_0002_),
    .B(_1309_),
    .C(_1458_),
    .Y(_1460_));
 sg13g2_xnor2_1 _2378_ (.Y(_1461_),
    .A(_0002_),
    .B(_1459_));
 sg13g2_nand2b_1 _2379_ (.Y(_1462_),
    .B(_1461_),
    .A_N(\hvsync_gen.vpos[10] ));
 sg13g2_nor2_1 _2380_ (.A(_0011_),
    .B(_1458_),
    .Y(_1463_));
 sg13g2_xnor2_1 _2381_ (.Y(_1464_),
    .A(\hvsync_gen.vdisplay[9] ),
    .B(_1463_));
 sg13g2_nor2_1 _2382_ (.A(net318),
    .B(_1464_),
    .Y(_1465_));
 sg13g2_xnor2_1 _2383_ (.Y(_1466_),
    .A(\hvsync_gen.vdisplay[8] ),
    .B(_1458_));
 sg13g2_nor2_1 _2384_ (.A(_0010_),
    .B(_1466_),
    .Y(_1467_));
 sg13g2_xnor2_1 _2385_ (.Y(_1468_),
    .A(_0012_),
    .B(_1464_));
 sg13g2_nor2b_1 _2386_ (.A(_1467_),
    .B_N(_1468_),
    .Y(_1469_));
 sg13g2_nand2b_1 _2387_ (.Y(_1470_),
    .B(_1468_),
    .A_N(_1467_));
 sg13g2_xnor2_1 _2388_ (.Y(_1471_),
    .A(_1317_),
    .B(_1457_));
 sg13g2_nor2_1 _2389_ (.A(net320),
    .B(_1471_),
    .Y(_1472_));
 sg13g2_xnor2_1 _2390_ (.Y(_1473_),
    .A(_1334_),
    .B(_1454_));
 sg13g2_o21ai_1 _2391_ (.B1(_1325_),
    .Y(_1474_),
    .A1(_1326_),
    .A2(_1455_));
 sg13g2_nor2b_1 _2392_ (.A(_1456_),
    .B_N(_1474_),
    .Y(_1475_));
 sg13g2_xnor2_1 _2393_ (.Y(_1476_),
    .A(net322),
    .B(_1475_));
 sg13g2_a221oi_1 _2394_ (.B2(net327),
    .C1(_1476_),
    .B1(_1473_),
    .A1(net320),
    .Y(_1477_),
    .A2(_1471_));
 sg13g2_nor2b_1 _2395_ (.A(_1472_),
    .B_N(_1477_),
    .Y(_1478_));
 sg13g2_xnor2_1 _2396_ (.Y(_1479_),
    .A(_1342_),
    .B(_1453_));
 sg13g2_nand2b_1 _2397_ (.Y(_1480_),
    .B(net329),
    .A_N(_1479_));
 sg13g2_nor2_1 _2398_ (.A(net327),
    .B(_1473_),
    .Y(_1481_));
 sg13g2_a21oi_1 _2399_ (.A1(_0804_),
    .A2(_1479_),
    .Y(_1482_),
    .B1(_1481_));
 sg13g2_nand3_1 _2400_ (.B(_1480_),
    .C(_1482_),
    .A(_1478_),
    .Y(_1483_));
 sg13g2_xnor2_1 _2401_ (.Y(_1484_),
    .A(_1355_),
    .B(_1452_));
 sg13g2_nor2_1 _2402_ (.A(net330),
    .B(_1484_),
    .Y(_1485_));
 sg13g2_nand2_1 _2403_ (.Y(_1486_),
    .A(net330),
    .B(_1484_));
 sg13g2_xor2_1 _2404_ (.B(_1451_),
    .A(_1364_),
    .X(_1487_));
 sg13g2_nand2_1 _2405_ (.Y(_1488_),
    .A(_0004_),
    .B(_1487_));
 sg13g2_nand2b_1 _2406_ (.Y(_1489_),
    .B(_0801_),
    .A_N(_1487_));
 sg13g2_a221oi_1 _2407_ (.B2(_1489_),
    .C1(_1485_),
    .B1(_1488_),
    .A1(net330),
    .Y(_1490_),
    .A2(_1484_));
 sg13g2_xnor2_1 _2408_ (.Y(_1491_),
    .A(_1374_),
    .B(_1381_));
 sg13g2_nor2_1 _2409_ (.A(net333),
    .B(_1487_),
    .Y(_1492_));
 sg13g2_o21ai_1 _2410_ (.B1(_1486_),
    .Y(_1493_),
    .A1(_1485_),
    .A2(_1492_));
 sg13g2_xnor2_1 _2411_ (.Y(_1494_),
    .A(_0003_),
    .B(_1491_));
 sg13g2_a21oi_1 _2412_ (.A1(net336),
    .A2(_1382_),
    .Y(_1495_),
    .B1(_1494_));
 sg13g2_a21oi_1 _2413_ (.A1(_0797_),
    .A2(_1491_),
    .Y(_1496_),
    .B1(_1495_));
 sg13g2_nand2b_1 _2414_ (.Y(_1497_),
    .B(_1490_),
    .A_N(_1496_));
 sg13g2_a21o_1 _2415_ (.A2(_1497_),
    .A1(_1493_),
    .B1(_1483_),
    .X(_1498_));
 sg13g2_nand2b_1 _2416_ (.Y(_1499_),
    .B(_1478_),
    .A_N(_1482_));
 sg13g2_nand2_2 _2417_ (.Y(_1500_),
    .A(_0010_),
    .B(_1466_));
 sg13g2_nand2_1 _2418_ (.Y(_0146_),
    .A(_0810_),
    .B(_1475_));
 sg13g2_a21oi_1 _2419_ (.A1(net320),
    .A2(_1471_),
    .Y(_0147_),
    .B1(_0146_));
 sg13g2_nor2_1 _2420_ (.A(_1472_),
    .B(_0147_),
    .Y(_0148_));
 sg13g2_nand4_1 _2421_ (.B(_1499_),
    .C(_1500_),
    .A(_1498_),
    .Y(_0149_),
    .D(_0148_));
 sg13g2_a21oi_1 _2422_ (.A1(_1469_),
    .A2(_0149_),
    .Y(_0150_),
    .B1(_1465_));
 sg13g2_xnor2_1 _2423_ (.Y(_0151_),
    .A(_0013_),
    .B(_1461_));
 sg13g2_o21ai_1 _2424_ (.B1(_1462_),
    .Y(_0152_),
    .A1(_0150_),
    .A2(_0151_));
 sg13g2_nand2b_1 _2425_ (.Y(_0153_),
    .B(_0794_),
    .A_N(_1382_));
 sg13g2_nand4_1 _2426_ (.B(_1495_),
    .C(_1500_),
    .A(_1490_),
    .Y(_0154_),
    .D(_0153_));
 sg13g2_and2_1 _2427_ (.A(net174),
    .B(_1460_),
    .X(_0155_));
 sg13g2_nor4_1 _2428_ (.A(_1470_),
    .B(_1483_),
    .C(_0151_),
    .D(_0154_),
    .Y(_0156_));
 sg13g2_nor2_1 _2429_ (.A(_0014_),
    .B(_1460_),
    .Y(_0157_));
 sg13g2_nor2_1 _2430_ (.A(_0156_),
    .B(_0157_),
    .Y(_0158_));
 sg13g2_a221oi_1 _2431_ (.B2(_0158_),
    .C1(_0155_),
    .B1(_0152_),
    .A1(_1404_),
    .Y(_0159_),
    .A2(_1450_));
 sg13g2_xor2_1 _2432_ (.B(_0159_),
    .A(\hvsync_gen.vsyncpolarity ),
    .X(_0001_));
 sg13g2_nand2_1 _2433_ (.Y(_0160_),
    .A(\hfrontporch[9] ),
    .B(\hdisplay[9] ));
 sg13g2_nor2_1 _2434_ (.A(_0833_),
    .B(_0834_),
    .Y(_0161_));
 sg13g2_nand2_2 _2435_ (.Y(_0162_),
    .A(_0833_),
    .B(_0834_));
 sg13g2_nand2b_2 _2436_ (.Y(_0163_),
    .B(_0162_),
    .A_N(_0161_));
 sg13g2_and2_1 _2437_ (.A(\hfrontporch[7] ),
    .B(\hdisplay[7] ),
    .X(_0164_));
 sg13g2_or2_2 _2438_ (.X(_0165_),
    .B(\hdisplay[7] ),
    .A(\hfrontporch[7] ));
 sg13g2_nand2b_2 _2439_ (.Y(_0166_),
    .B(_0165_),
    .A_N(_0164_));
 sg13g2_and2_1 _2440_ (.A(\hfrontporch[6] ),
    .B(\hdisplay[6] ),
    .X(_0167_));
 sg13g2_or2_2 _2441_ (.X(_0168_),
    .B(\hdisplay[6] ),
    .A(\hfrontporch[6] ));
 sg13g2_nand2b_2 _2442_ (.Y(_0169_),
    .B(_0168_),
    .A_N(_0167_));
 sg13g2_and2_1 _2443_ (.A(\hfrontporch[5] ),
    .B(\hdisplay[5] ),
    .X(_0170_));
 sg13g2_or2_1 _2444_ (.X(_0171_),
    .B(\hdisplay[5] ),
    .A(\hfrontporch[5] ));
 sg13g2_xnor2_1 _2445_ (.Y(_0172_),
    .A(\hfrontporch[5] ),
    .B(\hdisplay[5] ));
 sg13g2_nor2_1 _2446_ (.A(_0822_),
    .B(_0823_),
    .Y(_0173_));
 sg13g2_or2_1 _2447_ (.X(_0174_),
    .B(\hdisplay[4] ),
    .A(\hfrontporch[4] ));
 sg13g2_xnor2_1 _2448_ (.Y(_0175_),
    .A(\hfrontporch[4] ),
    .B(\hdisplay[4] ));
 sg13g2_nand2_1 _2449_ (.Y(_0176_),
    .A(\hfrontporch[3] ),
    .B(\hdisplay[3] ));
 sg13g2_nor2_1 _2450_ (.A(\hfrontporch[3] ),
    .B(\hdisplay[3] ),
    .Y(_0177_));
 sg13g2_xnor2_1 _2451_ (.Y(_0178_),
    .A(\hfrontporch[3] ),
    .B(\hdisplay[3] ));
 sg13g2_and2_1 _2452_ (.A(\hfrontporch[2] ),
    .B(\hdisplay[2] ),
    .X(_0179_));
 sg13g2_nor2_1 _2453_ (.A(\hfrontporch[2] ),
    .B(\hdisplay[2] ),
    .Y(_0180_));
 sg13g2_xor2_1 _2454_ (.B(\hdisplay[2] ),
    .A(\hfrontporch[2] ),
    .X(_0181_));
 sg13g2_nand2_1 _2455_ (.Y(_0182_),
    .A(\hfrontporch[1] ),
    .B(\hdisplay[1] ));
 sg13g2_nor2_1 _2456_ (.A(\hfrontporch[1] ),
    .B(\hdisplay[1] ),
    .Y(_0183_));
 sg13g2_xnor2_1 _2457_ (.Y(_0184_),
    .A(\hfrontporch[1] ),
    .B(\hdisplay[1] ));
 sg13g2_nand2_2 _2458_ (.Y(_0185_),
    .A(\hfrontporch[0] ),
    .B(\hdisplay[0] ));
 sg13g2_o21ai_1 _2459_ (.B1(_0182_),
    .Y(_0186_),
    .A1(_0184_),
    .A2(_0185_));
 sg13g2_a21oi_2 _2460_ (.B1(_0179_),
    .Y(_0187_),
    .A2(_0186_),
    .A1(_0181_));
 sg13g2_o21ai_1 _2461_ (.B1(_0176_),
    .Y(_0188_),
    .A1(_0177_),
    .A2(_0187_));
 sg13g2_a21o_1 _2462_ (.A2(_0188_),
    .A1(_0174_),
    .B1(_0173_),
    .X(_0189_));
 sg13g2_a21o_1 _2463_ (.A2(_0189_),
    .A1(_0171_),
    .B1(_0170_),
    .X(_0190_));
 sg13g2_a21o_1 _2464_ (.A2(_0190_),
    .A1(_0168_),
    .B1(_0167_),
    .X(_0191_));
 sg13g2_a21o_1 _2465_ (.A2(_0191_),
    .A1(_0165_),
    .B1(_0164_),
    .X(_0192_));
 sg13g2_a21oi_1 _2466_ (.A1(_0162_),
    .A2(_0192_),
    .Y(_0193_),
    .B1(_0161_));
 sg13g2_nor2_1 _2467_ (.A(\hfrontporch[9] ),
    .B(\hdisplay[9] ),
    .Y(_0194_));
 sg13g2_xor2_1 _2468_ (.B(\hdisplay[9] ),
    .A(\hfrontporch[9] ),
    .X(_0195_));
 sg13g2_o21ai_1 _2469_ (.B1(_0160_),
    .Y(_0196_),
    .A1(_0193_),
    .A2(_0194_));
 sg13g2_nand2_1 _2470_ (.Y(_0197_),
    .A(\hdisplay[10] ),
    .B(_0196_));
 sg13g2_xnor2_1 _2471_ (.Y(_0198_),
    .A(_0837_),
    .B(_0196_));
 sg13g2_nand2b_1 _2472_ (.Y(_0199_),
    .B(\hpos[10] ),
    .A_N(_0198_));
 sg13g2_xnor2_1 _2473_ (.Y(_0200_),
    .A(_0023_),
    .B(_0198_));
 sg13g2_xor2_1 _2474_ (.B(_0195_),
    .A(_0193_),
    .X(_0201_));
 sg13g2_xor2_1 _2475_ (.B(_0192_),
    .A(_0163_),
    .X(_0202_));
 sg13g2_xor2_1 _2476_ (.B(_0191_),
    .A(_0166_),
    .X(_0203_));
 sg13g2_nand2_1 _2477_ (.Y(_0204_),
    .A(_0831_),
    .B(_0203_));
 sg13g2_nor2_1 _2478_ (.A(_0831_),
    .B(_0203_),
    .Y(_0205_));
 sg13g2_xor2_1 _2479_ (.B(_0190_),
    .A(_0169_),
    .X(_0206_));
 sg13g2_xor2_1 _2480_ (.B(_0189_),
    .A(_0172_),
    .X(_0207_));
 sg13g2_nand2_1 _2481_ (.Y(_0208_),
    .A(net352),
    .B(_0207_));
 sg13g2_xnor2_1 _2482_ (.Y(_0209_),
    .A(_0184_),
    .B(_0185_));
 sg13g2_or2_1 _2483_ (.X(_0210_),
    .B(\hdisplay[0] ),
    .A(\hfrontporch[0] ));
 sg13g2_nand2_1 _2484_ (.Y(_0211_),
    .A(_0185_),
    .B(_0210_));
 sg13g2_nand3_1 _2485_ (.B(_0185_),
    .C(_0210_),
    .A(_0795_),
    .Y(_0212_));
 sg13g2_xnor2_1 _2486_ (.Y(_0213_),
    .A(_0015_),
    .B(_0209_));
 sg13g2_a22oi_1 _2487_ (.Y(_0214_),
    .B1(_0212_),
    .B2(_0213_),
    .A2(_0209_),
    .A1(net359));
 sg13g2_xnor2_1 _2488_ (.Y(_0215_),
    .A(_0181_),
    .B(_0186_));
 sg13g2_xor2_1 _2489_ (.B(_0215_),
    .A(_0016_),
    .X(_0216_));
 sg13g2_xnor2_1 _2490_ (.Y(_0217_),
    .A(_0178_),
    .B(_0187_));
 sg13g2_a22oi_1 _2491_ (.Y(_0218_),
    .B1(_0217_),
    .B2(net356),
    .A2(_0215_),
    .A1(net358));
 sg13g2_o21ai_1 _2492_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0214_),
    .A2(_0216_));
 sg13g2_nand2b_1 _2493_ (.Y(_0220_),
    .B(_0820_),
    .A_N(_0217_));
 sg13g2_xor2_1 _2494_ (.B(_0188_),
    .A(_0175_),
    .X(_0221_));
 sg13g2_a22oi_1 _2495_ (.Y(_0222_),
    .B1(_0221_),
    .B2(net354),
    .A2(_0220_),
    .A1(_0219_));
 sg13g2_nand2b_1 _2496_ (.Y(_0223_),
    .B(_0821_),
    .A_N(_0221_));
 sg13g2_o21ai_1 _2497_ (.B1(_0223_),
    .Y(_0224_),
    .A1(net350),
    .A2(_0207_));
 sg13g2_o21ai_1 _2498_ (.B1(_0208_),
    .Y(_0225_),
    .A1(_0222_),
    .A2(_0224_));
 sg13g2_xnor2_1 _2499_ (.Y(_0226_),
    .A(_0020_),
    .B(_0206_));
 sg13g2_a22oi_1 _2500_ (.Y(_0227_),
    .B1(_0225_),
    .B2(_0226_),
    .A2(_0206_),
    .A1(net349));
 sg13g2_a21oi_1 _2501_ (.A1(_0204_),
    .A2(_0227_),
    .Y(_0228_),
    .B1(_0205_));
 sg13g2_o21ai_1 _2502_ (.B1(_0228_),
    .Y(_0229_),
    .A1(net346),
    .A2(_0202_));
 sg13g2_a22oi_1 _2503_ (.Y(_0230_),
    .B1(_0202_),
    .B2(net346),
    .A2(_0201_),
    .A1(net344));
 sg13g2_nand2_1 _2504_ (.Y(_0231_),
    .A(_0229_),
    .B(_0230_));
 sg13g2_o21ai_1 _2505_ (.B1(_0231_),
    .Y(_0232_),
    .A1(net344),
    .A2(_0201_));
 sg13g2_o21ai_1 _2506_ (.B1(_0199_),
    .Y(_0233_),
    .A1(_0200_),
    .A2(_0232_));
 sg13g2_xnor2_1 _2507_ (.Y(_0234_),
    .A(_0024_),
    .B(_0197_));
 sg13g2_a22oi_1 _2508_ (.Y(_0235_),
    .B1(_0233_),
    .B2(_0234_),
    .A2(_0197_),
    .A1(net152));
 sg13g2_nand2_1 _2509_ (.Y(_0236_),
    .A(_0837_),
    .B(_0194_));
 sg13g2_a21oi_1 _2510_ (.A1(_0833_),
    .A2(_0834_),
    .Y(_0237_),
    .B1(_0195_));
 sg13g2_xnor2_1 _2511_ (.Y(_0238_),
    .A(_0162_),
    .B(_0195_));
 sg13g2_a21oi_2 _2512_ (.B1(_0237_),
    .Y(_0239_),
    .A2(_0238_),
    .A1(\hsynclength[9] ));
 sg13g2_o21ai_1 _2513_ (.B1(\hdisplay[10] ),
    .Y(_0240_),
    .A1(\hfrontporch[9] ),
    .A2(\hdisplay[9] ));
 sg13g2_nand2_1 _2514_ (.Y(_0241_),
    .A(_0236_),
    .B(_0240_));
 sg13g2_nor2b_1 _2515_ (.A(_0239_),
    .B_N(_0241_),
    .Y(_0242_));
 sg13g2_xor2_1 _2516_ (.B(_0241_),
    .A(_0239_),
    .X(_0243_));
 sg13g2_inv_1 _2517_ (.Y(_0244_),
    .A(_0243_));
 sg13g2_xnor2_1 _2518_ (.Y(_0245_),
    .A(\hsynclength[9] ),
    .B(_0238_));
 sg13g2_and2_1 _2519_ (.A(_0163_),
    .B(_0165_),
    .X(_0246_));
 sg13g2_xor2_1 _2520_ (.B(_0165_),
    .A(_0163_),
    .X(_0247_));
 sg13g2_a21oi_2 _2521_ (.B1(_0246_),
    .Y(_0248_),
    .A2(_0247_),
    .A1(\hsynclength[8] ));
 sg13g2_nor2_1 _2522_ (.A(_0245_),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_or2_1 _2523_ (.X(_0250_),
    .B(_0248_),
    .A(_0245_));
 sg13g2_xnor2_1 _2524_ (.Y(_0251_),
    .A(_0245_),
    .B(_0248_));
 sg13g2_inv_1 _2525_ (.Y(_0252_),
    .A(_0251_));
 sg13g2_xnor2_1 _2526_ (.Y(_0253_),
    .A(\hsynclength[8] ),
    .B(_0247_));
 sg13g2_and2_1 _2527_ (.A(_0166_),
    .B(_0168_),
    .X(_0254_));
 sg13g2_xor2_1 _2528_ (.B(_0168_),
    .A(_0166_),
    .X(_0255_));
 sg13g2_a21oi_1 _2529_ (.A1(\hsynclength[7] ),
    .A2(_0255_),
    .Y(_0256_),
    .B1(_0254_));
 sg13g2_nor2_1 _2530_ (.A(_0253_),
    .B(_0256_),
    .Y(_0257_));
 sg13g2_inv_1 _2531_ (.Y(_0258_),
    .A(_0257_));
 sg13g2_xor2_1 _2532_ (.B(_0256_),
    .A(_0253_),
    .X(_0259_));
 sg13g2_nand2_1 _2533_ (.Y(_0260_),
    .A(_0169_),
    .B(_0171_));
 sg13g2_xor2_1 _2534_ (.B(_0171_),
    .A(_0169_),
    .X(_0261_));
 sg13g2_nand2_1 _2535_ (.Y(_0262_),
    .A(\hsynclength[6] ),
    .B(_0261_));
 sg13g2_xnor2_1 _2536_ (.Y(_0263_),
    .A(\hsynclength[7] ),
    .B(_0255_));
 sg13g2_a21oi_2 _2537_ (.B1(_0263_),
    .Y(_0264_),
    .A2(_0262_),
    .A1(_0260_));
 sg13g2_nand3_1 _2538_ (.B(_0262_),
    .C(_0263_),
    .A(_0260_),
    .Y(_0265_));
 sg13g2_nor2b_2 _2539_ (.A(_0264_),
    .B_N(_0265_),
    .Y(_0266_));
 sg13g2_o21ai_1 _2540_ (.B1(_0175_),
    .Y(_0267_),
    .A1(\hfrontporch[3] ),
    .A2(\hdisplay[3] ));
 sg13g2_xnor2_1 _2541_ (.Y(_0268_),
    .A(_0175_),
    .B(_0177_));
 sg13g2_nand2_1 _2542_ (.Y(_0269_),
    .A(\hsynclength[4] ),
    .B(_0268_));
 sg13g2_and2_1 _2543_ (.A(_0172_),
    .B(_0174_),
    .X(_0270_));
 sg13g2_xor2_1 _2544_ (.B(_0174_),
    .A(_0172_),
    .X(_0271_));
 sg13g2_xnor2_1 _2545_ (.Y(_0272_),
    .A(\hsynclength[5] ),
    .B(_0271_));
 sg13g2_a21oi_2 _2546_ (.B1(_0272_),
    .Y(_0273_),
    .A2(_0269_),
    .A1(_0267_));
 sg13g2_nand3_1 _2547_ (.B(_0269_),
    .C(_0272_),
    .A(_0267_),
    .Y(_0274_));
 sg13g2_nor2b_2 _2548_ (.A(_0273_),
    .B_N(_0274_),
    .Y(_0275_));
 sg13g2_xnor2_1 _2549_ (.Y(_0276_),
    .A(\hsynclength[4] ),
    .B(_0268_));
 sg13g2_o21ai_1 _2550_ (.B1(_0178_),
    .Y(_0277_),
    .A1(\hfrontporch[2] ),
    .A2(\hdisplay[2] ));
 sg13g2_xnor2_1 _2551_ (.Y(_0278_),
    .A(_0178_),
    .B(_0180_));
 sg13g2_nand2_1 _2552_ (.Y(_0279_),
    .A(\hsynclength[3] ),
    .B(_0278_));
 sg13g2_and2_1 _2553_ (.A(_0277_),
    .B(_0279_),
    .X(_0280_));
 sg13g2_nor2_1 _2554_ (.A(_0276_),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_or2_1 _2555_ (.X(_0282_),
    .B(_0280_),
    .A(_0276_));
 sg13g2_xor2_1 _2556_ (.B(_0280_),
    .A(_0276_),
    .X(_0283_));
 sg13g2_xnor2_1 _2557_ (.Y(_0284_),
    .A(\hsynclength[3] ),
    .B(_0278_));
 sg13g2_nor2_1 _2558_ (.A(_0181_),
    .B(_0183_),
    .Y(_0285_));
 sg13g2_xor2_1 _2559_ (.B(_0183_),
    .A(_0181_),
    .X(_0286_));
 sg13g2_a21oi_1 _2560_ (.A1(\hsynclength[2] ),
    .A2(_0286_),
    .Y(_0287_),
    .B1(_0285_));
 sg13g2_nor2_1 _2561_ (.A(_0284_),
    .B(_0287_),
    .Y(_0288_));
 sg13g2_inv_1 _2562_ (.Y(_0289_),
    .A(_0288_));
 sg13g2_xnor2_1 _2563_ (.Y(_0290_),
    .A(_0284_),
    .B(_0287_));
 sg13g2_inv_1 _2564_ (.Y(_0291_),
    .A(_0290_));
 sg13g2_xnor2_1 _2565_ (.Y(_0292_),
    .A(\hsynclength[2] ),
    .B(_0286_));
 sg13g2_and2_1 _2566_ (.A(_0184_),
    .B(_0210_),
    .X(_0293_));
 sg13g2_xor2_1 _2567_ (.B(_0210_),
    .A(_0184_),
    .X(_0294_));
 sg13g2_a21oi_1 _2568_ (.A1(\hsynclength[1] ),
    .A2(_0294_),
    .Y(_0295_),
    .B1(_0293_));
 sg13g2_nor2_1 _2569_ (.A(_0292_),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_xor2_1 _2570_ (.B(_0295_),
    .A(_0292_),
    .X(_0297_));
 sg13g2_nand2_1 _2571_ (.Y(_0298_),
    .A(\hsynclength[0] ),
    .B(_0211_));
 sg13g2_xnor2_1 _2572_ (.Y(_0299_),
    .A(\hsynclength[1] ),
    .B(_0294_));
 sg13g2_nor2_2 _2573_ (.A(_0298_),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_a21oi_1 _2574_ (.A1(_0297_),
    .A2(_0300_),
    .Y(_0301_),
    .B1(_0296_));
 sg13g2_o21ai_1 _2575_ (.B1(_0289_),
    .Y(_0302_),
    .A1(_0290_),
    .A2(_0301_));
 sg13g2_nand3_1 _2576_ (.B(_0283_),
    .C(_0302_),
    .A(_0275_),
    .Y(_0303_));
 sg13g2_a21oi_1 _2577_ (.A1(_0274_),
    .A2(_0281_),
    .Y(_0304_),
    .B1(_0273_));
 sg13g2_xnor2_1 _2578_ (.Y(_0305_),
    .A(\hsynclength[6] ),
    .B(_0261_));
 sg13g2_a21oi_2 _2579_ (.B1(_0270_),
    .Y(_0306_),
    .A2(_0271_),
    .A1(\hsynclength[5] ));
 sg13g2_nor2_1 _2580_ (.A(_0305_),
    .B(_0306_),
    .Y(_0307_));
 sg13g2_xnor2_1 _2581_ (.Y(_0308_),
    .A(_0305_),
    .B(_0306_));
 sg13g2_inv_1 _2582_ (.Y(_0309_),
    .A(_0308_));
 sg13g2_a21oi_2 _2583_ (.B1(_0308_),
    .Y(_0310_),
    .A2(_0304_),
    .A1(_0303_));
 sg13g2_a21o_1 _2584_ (.A2(_0307_),
    .A1(_0265_),
    .B1(_0264_),
    .X(_0311_));
 sg13g2_a21o_1 _2585_ (.A2(_0310_),
    .A1(_0266_),
    .B1(_0311_),
    .X(_0312_));
 sg13g2_a21oi_1 _2586_ (.A1(_0259_),
    .A2(_0312_),
    .Y(_0313_),
    .B1(_0257_));
 sg13g2_o21ai_1 _2587_ (.B1(_0250_),
    .Y(_0314_),
    .A1(_0251_),
    .A2(_0313_));
 sg13g2_a21o_1 _2588_ (.A2(_0314_),
    .A1(_0244_),
    .B1(_0242_),
    .X(_0315_));
 sg13g2_nand2b_1 _2589_ (.Y(_0316_),
    .B(_0239_),
    .A_N(_0236_));
 sg13g2_nor2_1 _2590_ (.A(_0314_),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_a21o_1 _2591_ (.A2(_0315_),
    .A1(_0236_),
    .B1(_0317_),
    .X(_0318_));
 sg13g2_nand2_1 _2592_ (.Y(_0319_),
    .A(net169),
    .B(_0318_));
 sg13g2_xnor2_1 _2593_ (.Y(_0320_),
    .A(_0244_),
    .B(_0314_));
 sg13g2_nor2_1 _2594_ (.A(\hpos[10] ),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_xnor2_1 _2595_ (.Y(_0322_),
    .A(_0251_),
    .B(_0313_));
 sg13g2_nand3_1 _2596_ (.B(_0304_),
    .C(_0308_),
    .A(_0303_),
    .Y(_0323_));
 sg13g2_nor2b_2 _2597_ (.A(_0310_),
    .B_N(_0323_),
    .Y(_0324_));
 sg13g2_xnor2_1 _2598_ (.Y(_0325_),
    .A(_0020_),
    .B(_0324_));
 sg13g2_a21oi_1 _2599_ (.A1(_0283_),
    .A2(_0302_),
    .Y(_0326_),
    .B1(_0281_));
 sg13g2_xnor2_1 _2600_ (.Y(_0327_),
    .A(_0275_),
    .B(_0326_));
 sg13g2_inv_1 _2601_ (.Y(_0328_),
    .A(_0327_));
 sg13g2_xnor2_1 _2602_ (.Y(_0329_),
    .A(_0283_),
    .B(_0302_));
 sg13g2_nand2b_1 _2603_ (.Y(_0330_),
    .B(_0821_),
    .A_N(_0329_));
 sg13g2_xnor2_1 _2604_ (.Y(_0331_),
    .A(_0297_),
    .B(_0300_));
 sg13g2_xor2_1 _2605_ (.B(_0299_),
    .A(_0298_),
    .X(_0332_));
 sg13g2_xor2_1 _2606_ (.B(_0211_),
    .A(\hsynclength[0] ),
    .X(_0333_));
 sg13g2_nor3_1 _2607_ (.A(_0795_),
    .B(_0032_),
    .C(_0333_),
    .Y(_0334_));
 sg13g2_nand2b_1 _2608_ (.Y(_0335_),
    .B(_0015_),
    .A_N(_0334_));
 sg13g2_o21ai_1 _2609_ (.B1(net359),
    .Y(_0336_),
    .A1(_0015_),
    .A2(_0334_));
 sg13g2_nand2_1 _2610_ (.Y(_0337_),
    .A(_0332_),
    .B(_0336_));
 sg13g2_o21ai_1 _2611_ (.B1(_0337_),
    .Y(_0338_),
    .A1(_0332_),
    .A2(_0335_));
 sg13g2_xnor2_1 _2612_ (.Y(_0339_),
    .A(_0016_),
    .B(_0331_));
 sg13g2_xnor2_1 _2613_ (.Y(_0340_),
    .A(_0290_),
    .B(_0301_));
 sg13g2_nor2_1 _2614_ (.A(net358),
    .B(_0331_),
    .Y(_0341_));
 sg13g2_a21oi_1 _2615_ (.A1(_0338_),
    .A2(_0339_),
    .Y(_0342_),
    .B1(_0341_));
 sg13g2_o21ai_1 _2616_ (.B1(_0342_),
    .Y(_0343_),
    .A1(net356),
    .A2(_0340_));
 sg13g2_a22oi_1 _2617_ (.Y(_0344_),
    .B1(_0340_),
    .B2(net356),
    .A2(_0329_),
    .A1(net354));
 sg13g2_a22oi_1 _2618_ (.Y(_0345_),
    .B1(_0343_),
    .B2(_0344_),
    .A2(_0327_),
    .A1(_0825_));
 sg13g2_a221oi_1 _2619_ (.B2(_0345_),
    .C1(_0325_),
    .B1(_0330_),
    .A1(net350),
    .Y(_0346_),
    .A2(_0328_));
 sg13g2_nor2_1 _2620_ (.A(_0307_),
    .B(_0310_),
    .Y(_0347_));
 sg13g2_xor2_1 _2621_ (.B(_0347_),
    .A(_0266_),
    .X(_0348_));
 sg13g2_nand2_1 _2622_ (.Y(_0349_),
    .A(_0828_),
    .B(_0324_));
 sg13g2_o21ai_1 _2623_ (.B1(_0349_),
    .Y(_0350_),
    .A1(net347),
    .A2(_0348_));
 sg13g2_xnor2_1 _2624_ (.Y(_0351_),
    .A(_0259_),
    .B(_0312_));
 sg13g2_a22oi_1 _2625_ (.Y(_0352_),
    .B1(_0351_),
    .B2(net346),
    .A2(_0348_),
    .A1(net347));
 sg13g2_o21ai_1 _2626_ (.B1(_0352_),
    .Y(_0353_),
    .A1(_0346_),
    .A2(_0350_));
 sg13g2_nor2_1 _2627_ (.A(net343),
    .B(_0322_),
    .Y(_0354_));
 sg13g2_nor2_1 _2628_ (.A(net346),
    .B(_0351_),
    .Y(_0355_));
 sg13g2_nor2_1 _2629_ (.A(_0354_),
    .B(_0355_),
    .Y(_0356_));
 sg13g2_xor2_1 _2630_ (.B(_0320_),
    .A(_0023_),
    .X(_0357_));
 sg13g2_a221oi_1 _2631_ (.B2(_0356_),
    .C1(_0357_),
    .B1(_0353_),
    .A1(net343),
    .Y(_0358_),
    .A2(_0322_));
 sg13g2_xnor2_1 _2632_ (.Y(_0359_),
    .A(\hpos[11] ),
    .B(_0318_));
 sg13g2_o21ai_1 _2633_ (.B1(_0359_),
    .Y(_0360_),
    .A1(_0321_),
    .A2(_0358_));
 sg13g2_a21oi_1 _2634_ (.A1(_0319_),
    .A2(_0360_),
    .Y(_0361_),
    .B1(_0235_));
 sg13g2_xor2_1 _2635_ (.B(_0361_),
    .A(hsyncpolarity),
    .X(_0000_));
 sg13g2_nand2_1 _2636_ (.Y(_0362_),
    .A(\hbackporch[4] ),
    .B(_0283_));
 sg13g2_xnor2_1 _2637_ (.Y(_0363_),
    .A(\hbackporch[5] ),
    .B(_0275_));
 sg13g2_a21oi_1 _2638_ (.A1(_0282_),
    .A2(_0362_),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_and3_2 _2639_ (.X(_0365_),
    .A(_0282_),
    .B(_0362_),
    .C(_0363_));
 sg13g2_xnor2_1 _2640_ (.Y(_0366_),
    .A(\hbackporch[4] ),
    .B(_0283_));
 sg13g2_a21oi_1 _2641_ (.A1(\hbackporch[3] ),
    .A2(_0291_),
    .Y(_0367_),
    .B1(_0288_));
 sg13g2_nor2_1 _2642_ (.A(_0366_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_a21oi_1 _2643_ (.A1(\hbackporch[2] ),
    .A2(_0297_),
    .Y(_0369_),
    .B1(_0296_));
 sg13g2_xor2_1 _2644_ (.B(_0290_),
    .A(\hbackporch[3] ),
    .X(_0370_));
 sg13g2_nor2_1 _2645_ (.A(_0369_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_a21oi_1 _2646_ (.A1(\hbackporch[1] ),
    .A2(_0332_),
    .Y(_0372_),
    .B1(_0300_));
 sg13g2_xnor2_1 _2647_ (.Y(_0373_),
    .A(\hbackporch[2] ),
    .B(_0297_));
 sg13g2_nor2_1 _2648_ (.A(_0372_),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_nand2_1 _2649_ (.Y(_0375_),
    .A(\hbackporch[0] ),
    .B(_0333_));
 sg13g2_xnor2_1 _2650_ (.Y(_0376_),
    .A(\hbackporch[1] ),
    .B(_0332_));
 sg13g2_nor2_1 _2651_ (.A(_0375_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_xor2_1 _2652_ (.B(_0373_),
    .A(_0372_),
    .X(_0378_));
 sg13g2_a21o_1 _2653_ (.A2(_0378_),
    .A1(_0377_),
    .B1(_0374_),
    .X(_0379_));
 sg13g2_xor2_1 _2654_ (.B(_0370_),
    .A(_0369_),
    .X(_0380_));
 sg13g2_a21oi_2 _2655_ (.B1(_0371_),
    .Y(_0381_),
    .A2(_0380_),
    .A1(_0379_));
 sg13g2_xnor2_1 _2656_ (.Y(_0382_),
    .A(_0366_),
    .B(_0367_));
 sg13g2_nor2_1 _2657_ (.A(_0381_),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_nor2_1 _2658_ (.A(_0364_),
    .B(_0368_),
    .Y(_0384_));
 sg13g2_o21ai_1 _2659_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_nor2b_1 _2660_ (.A(_0365_),
    .B_N(_0385_),
    .Y(_0386_));
 sg13g2_xor2_1 _2661_ (.B(_0308_),
    .A(\hbackporch[6] ),
    .X(_0387_));
 sg13g2_a21oi_2 _2662_ (.B1(_0273_),
    .Y(_0388_),
    .A2(_0274_),
    .A1(\hbackporch[5] ));
 sg13g2_nor2_1 _2663_ (.A(_0387_),
    .B(_0388_),
    .Y(_0389_));
 sg13g2_inv_1 _2664_ (.Y(_0390_),
    .A(_0389_));
 sg13g2_xnor2_1 _2665_ (.Y(_0391_),
    .A(_0387_),
    .B(_0388_));
 sg13g2_inv_1 _2666_ (.Y(_0392_),
    .A(_0391_));
 sg13g2_a21oi_2 _2667_ (.B1(_0307_),
    .Y(_0393_),
    .A2(_0309_),
    .A1(\hbackporch[6] ));
 sg13g2_xnor2_1 _2668_ (.Y(_0394_),
    .A(\hbackporch[7] ),
    .B(_0266_));
 sg13g2_nand2_1 _2669_ (.Y(_0395_),
    .A(_0393_),
    .B(_0394_));
 sg13g2_nor2_1 _2670_ (.A(_0393_),
    .B(_0394_),
    .Y(_0396_));
 sg13g2_xor2_1 _2671_ (.B(_0394_),
    .A(_0393_),
    .X(_0397_));
 sg13g2_and2_1 _2672_ (.A(_0392_),
    .B(_0397_),
    .X(_0398_));
 sg13g2_nand3b_1 _2673_ (.B(_0385_),
    .C(_0398_),
    .Y(_0399_),
    .A_N(_0365_));
 sg13g2_a21oi_2 _2674_ (.B1(_0396_),
    .Y(_0400_),
    .A2(_0395_),
    .A1(_0389_));
 sg13g2_nand2_1 _2675_ (.Y(_0401_),
    .A(\hbackporch[8] ),
    .B(_0259_));
 sg13g2_xnor2_1 _2676_ (.Y(_0402_),
    .A(\hbackporch[8] ),
    .B(_0259_));
 sg13g2_a21oi_2 _2677_ (.B1(_0264_),
    .Y(_0403_),
    .A2(_0265_),
    .A1(\hbackporch[7] ));
 sg13g2_nor2_1 _2678_ (.A(_0402_),
    .B(_0403_),
    .Y(_0404_));
 sg13g2_xnor2_1 _2679_ (.Y(_0405_),
    .A(_0402_),
    .B(_0403_));
 sg13g2_a21o_1 _2680_ (.A2(_0400_),
    .A1(_0399_),
    .B1(_0405_),
    .X(_0406_));
 sg13g2_nand3_1 _2681_ (.B(_0400_),
    .C(_0405_),
    .A(_0399_),
    .Y(_0407_));
 sg13g2_nand3_1 _2682_ (.B(_0406_),
    .C(_0407_),
    .A(_0022_),
    .Y(_0408_));
 sg13g2_a21o_1 _2683_ (.A2(_0407_),
    .A1(_0406_),
    .B1(_0022_),
    .X(_0409_));
 sg13g2_nor2b_1 _2684_ (.A(_0404_),
    .B_N(_0406_),
    .Y(_0410_));
 sg13g2_xor2_1 _2685_ (.B(_0251_),
    .A(\hbackporch[9] ),
    .X(_0411_));
 sg13g2_and3_1 _2686_ (.X(_0412_),
    .A(_0258_),
    .B(_0401_),
    .C(_0411_));
 sg13g2_nand3_1 _2687_ (.B(_0401_),
    .C(_0411_),
    .A(_0258_),
    .Y(_0413_));
 sg13g2_a21oi_1 _2688_ (.A1(_0258_),
    .A2(_0401_),
    .Y(_0414_),
    .B1(_0411_));
 sg13g2_nor2_1 _2689_ (.A(_0412_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_xor2_1 _2690_ (.B(_0415_),
    .A(net343),
    .X(_0416_));
 sg13g2_xnor2_1 _2691_ (.Y(_0417_),
    .A(_0410_),
    .B(_0416_));
 sg13g2_nand3b_1 _2692_ (.B(_0385_),
    .C(_0392_),
    .Y(_0418_),
    .A_N(_0365_));
 sg13g2_xnor2_1 _2693_ (.Y(_0419_),
    .A(_0021_),
    .B(_0397_));
 sg13g2_xnor2_1 _2694_ (.Y(_0420_),
    .A(_0386_),
    .B(_0392_));
 sg13g2_xnor2_1 _2695_ (.Y(_0421_),
    .A(_0381_),
    .B(_0382_));
 sg13g2_xnor2_1 _2696_ (.Y(_0422_),
    .A(_0018_),
    .B(_0421_));
 sg13g2_nor2_1 _2697_ (.A(_0364_),
    .B(_0365_),
    .Y(_0423_));
 sg13g2_xor2_1 _2698_ (.B(_0423_),
    .A(_0019_),
    .X(_0424_));
 sg13g2_or3_1 _2699_ (.A(_0368_),
    .B(_0383_),
    .C(_0424_),
    .X(_0425_));
 sg13g2_o21ai_1 _2700_ (.B1(_0424_),
    .Y(_0426_),
    .A1(_0368_),
    .A2(_0383_));
 sg13g2_xor2_1 _2701_ (.B(_0380_),
    .A(_0379_),
    .X(_0427_));
 sg13g2_nor2_1 _2702_ (.A(_0017_),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_and2_1 _2703_ (.A(_0017_),
    .B(_0427_),
    .X(_0429_));
 sg13g2_xor2_1 _2704_ (.B(_0378_),
    .A(_0377_),
    .X(_0430_));
 sg13g2_xor2_1 _2705_ (.B(_0376_),
    .A(_0375_),
    .X(_0431_));
 sg13g2_xnor2_1 _2706_ (.Y(_0432_),
    .A(_0795_),
    .B(_0333_));
 sg13g2_xnor2_1 _2707_ (.Y(_0433_),
    .A(\hbackporch[0] ),
    .B(_0432_));
 sg13g2_o21ai_1 _2708_ (.B1(_0433_),
    .Y(_0434_),
    .A1(_0015_),
    .A2(_0431_));
 sg13g2_a221oi_1 _2709_ (.B2(_0015_),
    .C1(_0434_),
    .B1(_0431_),
    .A1(_0016_),
    .Y(_0435_),
    .A2(_0430_));
 sg13g2_o21ai_1 _2710_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0016_),
    .A2(_0430_));
 sg13g2_nor3_1 _2711_ (.A(_0428_),
    .B(_0429_),
    .C(_0436_),
    .Y(_0437_));
 sg13g2_nand4_1 _2712_ (.B(_0425_),
    .C(_0426_),
    .A(_0422_),
    .Y(_0438_),
    .D(_0437_));
 sg13g2_nand2b_1 _2713_ (.Y(_0439_),
    .B(_0415_),
    .A_N(_0405_));
 sg13g2_a21o_1 _2714_ (.A2(_0400_),
    .A1(_0399_),
    .B1(_0439_),
    .X(_0440_));
 sg13g2_a21oi_1 _2715_ (.A1(_0404_),
    .A2(_0413_),
    .Y(_0441_),
    .B1(_0414_));
 sg13g2_a21oi_1 _2716_ (.A1(\hbackporch[9] ),
    .A2(_0252_),
    .Y(_0442_),
    .B1(_0249_));
 sg13g2_nor2_1 _2717_ (.A(_0243_),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_inv_1 _2718_ (.Y(_0444_),
    .A(_0443_));
 sg13g2_xnor2_1 _2719_ (.Y(_0445_),
    .A(_0243_),
    .B(_0442_));
 sg13g2_a21o_1 _2720_ (.A2(_0441_),
    .A1(_0440_),
    .B1(_0445_),
    .X(_0446_));
 sg13g2_nand3_1 _2721_ (.B(_0441_),
    .C(_0445_),
    .A(_0440_),
    .Y(_0447_));
 sg13g2_a21oi_1 _2722_ (.A1(_0446_),
    .A2(_0447_),
    .Y(_0448_),
    .B1(_0023_));
 sg13g2_nand3_1 _2723_ (.B(_0446_),
    .C(_0447_),
    .A(_0023_),
    .Y(_0449_));
 sg13g2_nor2b_1 _2724_ (.A(_0448_),
    .B_N(_0449_),
    .Y(_0450_));
 sg13g2_mux2_1 _2725_ (.A0(_0240_),
    .A1(_0236_),
    .S(_0239_),
    .X(_0451_));
 sg13g2_xnor2_1 _2726_ (.Y(_0452_),
    .A(_0024_),
    .B(_0451_));
 sg13g2_inv_1 _2727_ (.Y(_0453_),
    .A(_0452_));
 sg13g2_a21oi_1 _2728_ (.A1(_0444_),
    .A2(_0446_),
    .Y(_0454_),
    .B1(_0453_));
 sg13g2_and3_1 _2729_ (.X(_0455_),
    .A(_0444_),
    .B(_0446_),
    .C(_0453_));
 sg13g2_xnor2_1 _2730_ (.Y(_0456_),
    .A(_0020_),
    .B(_0420_));
 sg13g2_and3_1 _2731_ (.X(_0457_),
    .A(_0390_),
    .B(_0418_),
    .C(_0419_));
 sg13g2_a21oi_1 _2732_ (.A1(_0390_),
    .A2(_0418_),
    .Y(_0458_),
    .B1(_0419_));
 sg13g2_nor3_1 _2733_ (.A(_0438_),
    .B(_0457_),
    .C(_0458_),
    .Y(_0459_));
 sg13g2_nand4_1 _2734_ (.B(_0409_),
    .C(_0456_),
    .A(_0408_),
    .Y(_0460_),
    .D(_0459_));
 sg13g2_nor4_2 _2735_ (.A(_0417_),
    .B(_0454_),
    .C(_0455_),
    .Y(_0461_),
    .D(_0460_));
 sg13g2_nand2_1 _2736_ (.Y(_0462_),
    .A(_0450_),
    .B(_0461_));
 sg13g2_a21oi_2 _2737_ (.B1(_0796_),
    .Y(_0463_),
    .A2(_0461_),
    .A1(_0450_));
 sg13g2_nand2_2 _2738_ (.Y(_0464_),
    .A(net1),
    .B(_0462_));
 sg13g2_and2_1 _2739_ (.A(net147),
    .B(net287),
    .X(_0033_));
 sg13g2_nor3_1 _2740_ (.A(net156),
    .B(_0889_),
    .C(_0464_),
    .Y(_0034_));
 sg13g2_o21ai_1 _2741_ (.B1(net287),
    .Y(_0465_),
    .A1(net357),
    .A2(_0889_));
 sg13g2_nor2_1 _2742_ (.A(_0890_),
    .B(_0465_),
    .Y(_0035_));
 sg13g2_nand2b_1 _2743_ (.Y(_0466_),
    .B(_0889_),
    .A_N(_0016_));
 sg13g2_xnor2_1 _2744_ (.Y(_0467_),
    .A(_0820_),
    .B(_0466_));
 sg13g2_nor2_1 _2745_ (.A(_0464_),
    .B(_0467_),
    .Y(_0036_));
 sg13g2_o21ai_1 _2746_ (.B1(net287),
    .Y(_0468_),
    .A1(net353),
    .A2(_0891_));
 sg13g2_nor2_1 _2747_ (.A(_0915_),
    .B(_0468_),
    .Y(_0037_));
 sg13g2_nor2_1 _2748_ (.A(net161),
    .B(_0892_),
    .Y(_0469_));
 sg13g2_xnor2_1 _2749_ (.Y(_0470_),
    .A(net350),
    .B(_0469_));
 sg13g2_nor2_1 _2750_ (.A(_0464_),
    .B(_0470_),
    .Y(_0038_));
 sg13g2_xnor2_1 _2751_ (.Y(_0471_),
    .A(_0828_),
    .B(_0916_));
 sg13g2_nor2_1 _2752_ (.A(_0464_),
    .B(_0471_),
    .Y(_0039_));
 sg13g2_nor2_1 _2753_ (.A(_0020_),
    .B(_0916_),
    .Y(_0472_));
 sg13g2_xnor2_1 _2754_ (.Y(_0473_),
    .A(net347),
    .B(_0472_));
 sg13g2_nor2_1 _2755_ (.A(_0464_),
    .B(_0473_),
    .Y(_0040_));
 sg13g2_nor3_2 _2756_ (.A(_0828_),
    .B(_0830_),
    .C(_0916_),
    .Y(_0474_));
 sg13g2_o21ai_1 _2757_ (.B1(_0463_),
    .Y(_0475_),
    .A1(net345),
    .A2(_0474_));
 sg13g2_a21oi_1 _2758_ (.A1(net345),
    .A2(_0474_),
    .Y(_0041_),
    .B1(_0475_));
 sg13g2_nand2b_1 _2759_ (.Y(_0476_),
    .B(_0474_),
    .A_N(net163));
 sg13g2_xnor2_1 _2760_ (.Y(_0477_),
    .A(net343),
    .B(_0476_));
 sg13g2_and2_1 _2761_ (.A(net288),
    .B(net164),
    .X(_0042_));
 sg13g2_nand3_1 _2762_ (.B(net343),
    .C(_0474_),
    .A(net345),
    .Y(_0478_));
 sg13g2_xnor2_1 _2763_ (.Y(_0479_),
    .A(_0836_),
    .B(_0478_));
 sg13g2_nor2_1 _2764_ (.A(_0464_),
    .B(_0479_),
    .Y(_0043_));
 sg13g2_nor2_1 _2765_ (.A(_0023_),
    .B(_0478_),
    .Y(_0480_));
 sg13g2_xnor2_1 _2766_ (.Y(_0481_),
    .A(net152),
    .B(_0480_));
 sg13g2_nor2_1 _2767_ (.A(_0464_),
    .B(net153),
    .Y(_0044_));
 sg13g2_nand2b_1 _2768_ (.Y(_0482_),
    .B(net377),
    .A_N(net375));
 sg13g2_nand2b_1 _2769_ (.Y(_0483_),
    .B(net2),
    .A_N(net3));
 sg13g2_nor2_2 _2770_ (.A(_0482_),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_nor2_2 _2771_ (.A(net2),
    .B(net3),
    .Y(_0485_));
 sg13g2_nor2_2 _2772_ (.A(net377),
    .B(net375),
    .Y(_0486_));
 sg13g2_nand2b_1 _2773_ (.Y(_0487_),
    .B(_0485_),
    .A_N(net375));
 sg13g2_inv_1 _2774_ (.Y(_0488_),
    .A(net313));
 sg13g2_nor2_2 _2775_ (.A(net4),
    .B(net313),
    .Y(_0489_));
 sg13g2_and2_2 _2776_ (.A(net2),
    .B(net3),
    .X(_0490_));
 sg13g2_nand2_2 _2777_ (.Y(_0491_),
    .A(net377),
    .B(net375));
 sg13g2_and2_2 _2778_ (.A(net377),
    .B(_0490_),
    .X(_0492_));
 sg13g2_nand2_2 _2779_ (.Y(_0493_),
    .A(net377),
    .B(_0490_));
 sg13g2_nor2_1 _2780_ (.A(_0489_),
    .B(_0492_),
    .Y(_0494_));
 sg13g2_a21oi_1 _2781_ (.A1(net376),
    .A2(_0492_),
    .Y(_0495_),
    .B1(_0489_));
 sg13g2_a21o_1 _2782_ (.A2(_0492_),
    .A1(net376),
    .B1(_0489_),
    .X(_0496_));
 sg13g2_nor2_2 _2783_ (.A(net315),
    .B(net299),
    .Y(_0497_));
 sg13g2_a22oi_1 _2784_ (.Y(_0498_),
    .B1(net292),
    .B2(\hfrontporch[0] ),
    .A2(net315),
    .A1(net8));
 sg13g2_inv_1 _2785_ (.Y(_0045_),
    .A(_0498_));
 sg13g2_nand2_2 _2786_ (.Y(_0499_),
    .A(net9),
    .B(net300));
 sg13g2_a22oi_1 _2787_ (.Y(_0500_),
    .B1(net292),
    .B2(\hfrontporch[1] ),
    .A2(net315),
    .A1(net9));
 sg13g2_inv_1 _2788_ (.Y(_0046_),
    .A(_0500_));
 sg13g2_a22oi_1 _2789_ (.Y(_0501_),
    .B1(net292),
    .B2(\hfrontporch[2] ),
    .A2(net315),
    .A1(net10));
 sg13g2_inv_1 _2790_ (.Y(_0047_),
    .A(_0501_));
 sg13g2_a22oi_1 _2791_ (.Y(_0502_),
    .B1(net292),
    .B2(\hfrontporch[3] ),
    .A2(net315),
    .A1(net11));
 sg13g2_inv_1 _2792_ (.Y(_0048_),
    .A(_0502_));
 sg13g2_a22oi_1 _2793_ (.Y(_0049_),
    .B1(net292),
    .B2(_0822_),
    .A2(net315),
    .A1(_0792_));
 sg13g2_a22oi_1 _2794_ (.Y(_0503_),
    .B1(_0497_),
    .B2(\hfrontporch[5] ),
    .A2(net315),
    .A1(net13));
 sg13g2_inv_1 _2795_ (.Y(_0050_),
    .A(_0503_));
 sg13g2_a22oi_1 _2796_ (.Y(_0504_),
    .B1(_0497_),
    .B2(\hfrontporch[6] ),
    .A2(_0484_),
    .A1(net14));
 sg13g2_inv_1 _2797_ (.Y(_0051_),
    .A(_0504_));
 sg13g2_a22oi_1 _2798_ (.Y(_0505_),
    .B1(net292),
    .B2(\hfrontporch[7] ),
    .A2(_0484_),
    .A1(net15));
 sg13g2_inv_1 _2799_ (.Y(_0052_),
    .A(_0505_));
 sg13g2_a22oi_1 _2800_ (.Y(_0506_),
    .B1(net292),
    .B2(\hfrontporch[8] ),
    .A2(net315),
    .A1(net5));
 sg13g2_inv_1 _2801_ (.Y(_0053_),
    .A(_0506_));
 sg13g2_a22oi_1 _2802_ (.Y(_0507_),
    .B1(net292),
    .B2(\hfrontporch[9] ),
    .A2(_0484_),
    .A1(net6));
 sg13g2_inv_1 _2803_ (.Y(_0054_),
    .A(_0507_));
 sg13g2_nor2b_2 _2804_ (.A(net2),
    .B_N(net3),
    .Y(_0508_));
 sg13g2_nand2b_1 _2805_ (.Y(_0509_),
    .B(net3),
    .A_N(net2));
 sg13g2_nor2_1 _2806_ (.A(_0482_),
    .B(_0509_),
    .Y(_0510_));
 sg13g2_nor2_2 _2807_ (.A(net299),
    .B(net311),
    .Y(_0511_));
 sg13g2_a22oi_1 _2808_ (.Y(_0512_),
    .B1(net291),
    .B2(\hsynclength[0] ),
    .A2(net311),
    .A1(net8));
 sg13g2_inv_1 _2809_ (.Y(_0055_),
    .A(_0512_));
 sg13g2_a22oi_1 _2810_ (.Y(_0513_),
    .B1(net291),
    .B2(\hsynclength[1] ),
    .A2(net311),
    .A1(net9));
 sg13g2_inv_1 _2811_ (.Y(_0056_),
    .A(_0513_));
 sg13g2_a22oi_1 _2812_ (.Y(_0514_),
    .B1(net291),
    .B2(\hsynclength[2] ),
    .A2(net311),
    .A1(net10));
 sg13g2_inv_1 _2813_ (.Y(_0057_),
    .A(_0514_));
 sg13g2_a22oi_1 _2814_ (.Y(_0515_),
    .B1(net291),
    .B2(\hsynclength[3] ),
    .A2(net311),
    .A1(net11));
 sg13g2_inv_1 _2815_ (.Y(_0058_),
    .A(_0515_));
 sg13g2_nand2_2 _2816_ (.Y(_0516_),
    .A(net12),
    .B(net300));
 sg13g2_a22oi_1 _2817_ (.Y(_0517_),
    .B1(net291),
    .B2(\hsynclength[4] ),
    .A2(net311),
    .A1(net12));
 sg13g2_inv_1 _2818_ (.Y(_0059_),
    .A(_0517_));
 sg13g2_a22oi_1 _2819_ (.Y(_0060_),
    .B1(net291),
    .B2(_0826_),
    .A2(net311),
    .A1(_0791_));
 sg13g2_a22oi_1 _2820_ (.Y(_0061_),
    .B1(_0511_),
    .B2(_0829_),
    .A2(net312),
    .A1(_0790_));
 sg13g2_a22oi_1 _2821_ (.Y(_0518_),
    .B1(_0511_),
    .B2(\hsynclength[7] ),
    .A2(net312),
    .A1(net15));
 sg13g2_inv_1 _2822_ (.Y(_0062_),
    .A(_0518_));
 sg13g2_a22oi_1 _2823_ (.Y(_0519_),
    .B1(_0511_),
    .B2(\hsynclength[8] ),
    .A2(net312),
    .A1(net5));
 sg13g2_inv_1 _2824_ (.Y(_0063_),
    .A(_0519_));
 sg13g2_a22oi_1 _2825_ (.Y(_0520_),
    .B1(net291),
    .B2(\hsynclength[9] ),
    .A2(net311),
    .A1(net6));
 sg13g2_inv_1 _2826_ (.Y(_0064_),
    .A(_0520_));
 sg13g2_nand2_1 _2827_ (.Y(_0521_),
    .A(\hbackporch[0] ),
    .B(net302));
 sg13g2_nand2_2 _2828_ (.Y(_0522_),
    .A(net8),
    .B(net300));
 sg13g2_o21ai_1 _2829_ (.B1(_0521_),
    .Y(_0065_),
    .A1(_0493_),
    .A2(_0522_));
 sg13g2_nand2_1 _2830_ (.Y(_0523_),
    .A(\hbackporch[1] ),
    .B(net302));
 sg13g2_o21ai_1 _2831_ (.B1(_0523_),
    .Y(_0066_),
    .A1(_0493_),
    .A2(_0499_));
 sg13g2_nand2_1 _2832_ (.Y(_0524_),
    .A(\hbackporch[2] ),
    .B(net302));
 sg13g2_nand2_2 _2833_ (.Y(_0525_),
    .A(net10),
    .B(net300));
 sg13g2_o21ai_1 _2834_ (.B1(_0524_),
    .Y(_0067_),
    .A1(_0493_),
    .A2(_0525_));
 sg13g2_nand2_1 _2835_ (.Y(_0526_),
    .A(\hbackporch[3] ),
    .B(net302));
 sg13g2_nand2_2 _2836_ (.Y(_0527_),
    .A(net11),
    .B(net300));
 sg13g2_o21ai_1 _2837_ (.B1(_0526_),
    .Y(_0068_),
    .A1(_0493_),
    .A2(_0527_));
 sg13g2_nor2_2 _2838_ (.A(net12),
    .B(net299),
    .Y(_0528_));
 sg13g2_a22oi_1 _2839_ (.Y(_0069_),
    .B1(_0528_),
    .B2(_0492_),
    .A2(net302),
    .A1(_0824_));
 sg13g2_nor2_2 _2840_ (.A(net13),
    .B(_0496_),
    .Y(_0529_));
 sg13g2_a22oi_1 _2841_ (.Y(_0070_),
    .B1(_0529_),
    .B2(_0492_),
    .A2(_0494_),
    .A1(_0827_));
 sg13g2_nand2_1 _2842_ (.Y(_0530_),
    .A(\hbackporch[6] ),
    .B(_0494_));
 sg13g2_nand2_2 _2843_ (.Y(_0531_),
    .A(net14),
    .B(net301));
 sg13g2_o21ai_1 _2844_ (.B1(_0530_),
    .Y(_0071_),
    .A1(_0493_),
    .A2(_0531_));
 sg13g2_nand2_1 _2845_ (.Y(_0532_),
    .A(\hbackporch[7] ),
    .B(net302));
 sg13g2_nand2_2 _2846_ (.Y(_0533_),
    .A(net15),
    .B(net301));
 sg13g2_o21ai_1 _2847_ (.B1(_0532_),
    .Y(_0072_),
    .A1(_0493_),
    .A2(_0533_));
 sg13g2_nand2_1 _2848_ (.Y(_0534_),
    .A(\hbackporch[8] ),
    .B(net302));
 sg13g2_nand2_1 _2849_ (.Y(_0535_),
    .A(net5),
    .B(net301));
 sg13g2_o21ai_1 _2850_ (.B1(_0534_),
    .Y(_0073_),
    .A1(_0493_),
    .A2(_0535_));
 sg13g2_nand2_1 _2851_ (.Y(_0536_),
    .A(\hbackporch[9] ),
    .B(net302));
 sg13g2_nand2_1 _2852_ (.Y(_0537_),
    .A(net6),
    .B(net301));
 sg13g2_o21ai_1 _2853_ (.B1(_0536_),
    .Y(_0074_),
    .A1(_0493_),
    .A2(_0537_));
 sg13g2_nor3_1 _2854_ (.A(net2),
    .B(net3),
    .C(net4),
    .Y(_0538_));
 sg13g2_nand2b_2 _2855_ (.Y(_0539_),
    .B(_0485_),
    .A_N(net377));
 sg13g2_a21oi_1 _2856_ (.A1(net376),
    .A2(_0492_),
    .Y(_0540_),
    .B1(_0538_));
 sg13g2_nand2_1 _2857_ (.Y(_0541_),
    .A(\hvsync_gen.vdisplay[0] ),
    .B(net304));
 sg13g2_o21ai_1 _2858_ (.B1(_0541_),
    .Y(_0075_),
    .A1(_0522_),
    .A2(_0539_));
 sg13g2_nand2_1 _2859_ (.Y(_0542_),
    .A(\hvsync_gen.vdisplay[1] ),
    .B(net304));
 sg13g2_o21ai_1 _2860_ (.B1(_0542_),
    .Y(_0076_),
    .A1(_0499_),
    .A2(_0539_));
 sg13g2_nand2_1 _2861_ (.Y(_0543_),
    .A(\hvsync_gen.vdisplay[2] ),
    .B(net304));
 sg13g2_o21ai_1 _2862_ (.B1(_0543_),
    .Y(_0077_),
    .A1(_0525_),
    .A2(_0539_));
 sg13g2_nand2_1 _2863_ (.Y(_0544_),
    .A(\hvsync_gen.vdisplay[3] ),
    .B(net304));
 sg13g2_o21ai_1 _2864_ (.B1(_0544_),
    .Y(_0078_),
    .A1(_0527_),
    .A2(_0539_));
 sg13g2_nand2_1 _2865_ (.Y(_0545_),
    .A(\hvsync_gen.vdisplay[4] ),
    .B(net304));
 sg13g2_o21ai_1 _2866_ (.B1(_0545_),
    .Y(_0079_),
    .A1(_0516_),
    .A2(_0539_));
 sg13g2_nand2_1 _2867_ (.Y(_0546_),
    .A(\hvsync_gen.vdisplay[5] ),
    .B(net305));
 sg13g2_o21ai_1 _2868_ (.B1(_0546_),
    .Y(_0080_),
    .A1(_0529_),
    .A2(net305));
 sg13g2_nand2b_1 _2869_ (.Y(_0547_),
    .B(net375),
    .A_N(net377));
 sg13g2_and2_2 _2870_ (.A(net376),
    .B(_0538_),
    .X(_0548_));
 sg13g2_a22oi_1 _2871_ (.Y(_0081_),
    .B1(_0548_),
    .B2(_0790_),
    .A2(net305),
    .A1(_0811_));
 sg13g2_nor2_1 _2872_ (.A(net15),
    .B(_0496_),
    .Y(_0549_));
 sg13g2_nand2_1 _2873_ (.Y(_0550_),
    .A(\hvsync_gen.vdisplay[7] ),
    .B(net305));
 sg13g2_o21ai_1 _2874_ (.B1(_0550_),
    .Y(_0082_),
    .A1(net305),
    .A2(_0549_));
 sg13g2_a22oi_1 _2875_ (.Y(_0083_),
    .B1(_0548_),
    .B2(_0789_),
    .A2(net304),
    .A1(_0816_));
 sg13g2_nand2_1 _2876_ (.Y(_0551_),
    .A(\hvsync_gen.vdisplay[9] ),
    .B(net304));
 sg13g2_o21ai_1 _2877_ (.B1(_0551_),
    .Y(_0084_),
    .A1(_0537_),
    .A2(_0539_));
 sg13g2_nand2_1 _2878_ (.Y(_0552_),
    .A(\hvsync_gen.vdisplay[10] ),
    .B(net304));
 sg13g2_nand2_2 _2879_ (.Y(_0553_),
    .A(net7),
    .B(net301));
 sg13g2_inv_1 _2880_ (.Y(_0554_),
    .A(_0553_));
 sg13g2_o21ai_1 _2881_ (.B1(_0552_),
    .Y(_0085_),
    .A1(_0539_),
    .A2(_0553_));
 sg13g2_a22oi_1 _2882_ (.Y(_0555_),
    .B1(_0554_),
    .B2(net312),
    .A2(net291),
    .A1(hsyncpolarity));
 sg13g2_inv_1 _2883_ (.Y(_0086_),
    .A(_0555_));
 sg13g2_or2_2 _2884_ (.X(_0556_),
    .B(_0547_),
    .A(_0483_));
 sg13g2_and2_2 _2885_ (.A(net300),
    .B(net310),
    .X(_0557_));
 sg13g2_nand2_1 _2886_ (.Y(_0558_),
    .A(\hvsync_gen.vfrontporch[0] ),
    .B(_0557_));
 sg13g2_o21ai_1 _2887_ (.B1(_0558_),
    .Y(_0087_),
    .A1(_0522_),
    .A2(net310));
 sg13g2_nor3_1 _2888_ (.A(net9),
    .B(net299),
    .C(net310),
    .Y(_0559_));
 sg13g2_a21oi_1 _2889_ (.A1(_0798_),
    .A2(_0557_),
    .Y(_0088_),
    .B1(_0559_));
 sg13g2_nand2_1 _2890_ (.Y(_0560_),
    .A(\hvsync_gen.vfrontporch[2] ),
    .B(_0557_));
 sg13g2_o21ai_1 _2891_ (.B1(_0560_),
    .Y(_0089_),
    .A1(_0525_),
    .A2(net310));
 sg13g2_nand2_1 _2892_ (.Y(_0561_),
    .A(\hvsync_gen.vfrontporch[3] ),
    .B(net310));
 sg13g2_nor2_2 _2893_ (.A(net11),
    .B(net299),
    .Y(_0562_));
 sg13g2_o21ai_1 _2894_ (.B1(_0561_),
    .Y(_0090_),
    .A1(_0557_),
    .A2(_0562_));
 sg13g2_nand2_1 _2895_ (.Y(_0563_),
    .A(\hvsync_gen.vfrontporch[4] ),
    .B(_0557_));
 sg13g2_o21ai_1 _2896_ (.B1(_0563_),
    .Y(_0091_),
    .A1(_0516_),
    .A2(_0556_));
 sg13g2_nand2_1 _2897_ (.Y(_0564_),
    .A(\hvsync_gen.vfrontporch[5] ),
    .B(_0557_));
 sg13g2_nand2_2 _2898_ (.Y(_0565_),
    .A(net13),
    .B(net300));
 sg13g2_o21ai_1 _2899_ (.B1(_0564_),
    .Y(_0092_),
    .A1(net310),
    .A2(_0565_));
 sg13g2_nand2_1 _2900_ (.Y(_0566_),
    .A(\hvsync_gen.vfrontporch[6] ),
    .B(_0557_));
 sg13g2_o21ai_1 _2901_ (.B1(_0566_),
    .Y(_0093_),
    .A1(_0531_),
    .A2(net310));
 sg13g2_nand2_1 _2902_ (.Y(_0567_),
    .A(\hvsync_gen.vfrontporch[7] ),
    .B(_0557_));
 sg13g2_o21ai_1 _2903_ (.B1(_0567_),
    .Y(_0094_),
    .A1(_0533_),
    .A2(net310));
 sg13g2_or2_2 _2904_ (.X(_0568_),
    .B(_0547_),
    .A(_0509_));
 sg13g2_and2_1 _2905_ (.A(net301),
    .B(net309),
    .X(_0569_));
 sg13g2_nand2_1 _2906_ (.Y(_0570_),
    .A(\hvsync_gen.vsynclength[0] ),
    .B(net290));
 sg13g2_o21ai_1 _2907_ (.B1(_0570_),
    .Y(_0095_),
    .A1(_0522_),
    .A2(net309));
 sg13g2_nor3_1 _2908_ (.A(net9),
    .B(net299),
    .C(net309),
    .Y(_0571_));
 sg13g2_a21oi_1 _2909_ (.A1(_0799_),
    .A2(net290),
    .Y(_0096_),
    .B1(_0571_));
 sg13g2_nand2_1 _2910_ (.Y(_0572_),
    .A(\hvsync_gen.vsynclength[2] ),
    .B(net290));
 sg13g2_o21ai_1 _2911_ (.B1(_0572_),
    .Y(_0097_),
    .A1(_0525_),
    .A2(net309));
 sg13g2_nand2_1 _2912_ (.Y(_0573_),
    .A(\hvsync_gen.vsynclength[3] ),
    .B(net290));
 sg13g2_o21ai_1 _2913_ (.B1(_0573_),
    .Y(_0098_),
    .A1(_0527_),
    .A2(net309));
 sg13g2_nand2_1 _2914_ (.Y(_0574_),
    .A(\hvsync_gen.vsynclength[4] ),
    .B(net290));
 sg13g2_o21ai_1 _2915_ (.B1(_0574_),
    .Y(_0099_),
    .A1(_0516_),
    .A2(net309));
 sg13g2_nand2_1 _2916_ (.Y(_0575_),
    .A(\hvsync_gen.vsynclength[5] ),
    .B(_0569_));
 sg13g2_o21ai_1 _2917_ (.B1(_0575_),
    .Y(_0100_),
    .A1(_0565_),
    .A2(_0568_));
 sg13g2_nand2_1 _2918_ (.Y(_0576_),
    .A(\hvsync_gen.vsynclength[6] ),
    .B(net290));
 sg13g2_o21ai_1 _2919_ (.B1(_0576_),
    .Y(_0101_),
    .A1(_0531_),
    .A2(_0568_));
 sg13g2_nand2_1 _2920_ (.Y(_0577_),
    .A(\hvsync_gen.vsynclength[7] ),
    .B(net290));
 sg13g2_o21ai_1 _2921_ (.B1(_0577_),
    .Y(_0102_),
    .A1(_0533_),
    .A2(net309));
 sg13g2_nand2_2 _2922_ (.Y(_0578_),
    .A(net375),
    .B(_0490_));
 sg13g2_nor2b_2 _2923_ (.A(_0489_),
    .B_N(_0578_),
    .Y(_0579_));
 sg13g2_nor2_2 _2924_ (.A(net8),
    .B(net299),
    .Y(_0580_));
 sg13g2_nand2_1 _2925_ (.Y(_0581_),
    .A(\hvsync_gen.vbackporch[0] ),
    .B(net298));
 sg13g2_o21ai_1 _2926_ (.B1(_0581_),
    .Y(_0103_),
    .A1(net298),
    .A2(_0580_));
 sg13g2_nand2_1 _2927_ (.Y(_0582_),
    .A(\hvsync_gen.vbackporch[1] ),
    .B(net298));
 sg13g2_o21ai_1 _2928_ (.B1(_0582_),
    .Y(_0104_),
    .A1(_0499_),
    .A2(_0578_));
 sg13g2_nand2_1 _2929_ (.Y(_0583_),
    .A(\hvsync_gen.vbackporch[2] ),
    .B(net298));
 sg13g2_o21ai_1 _2930_ (.B1(_0583_),
    .Y(_0105_),
    .A1(_0525_),
    .A2(_0578_));
 sg13g2_nand2_1 _2931_ (.Y(_0584_),
    .A(\hvsync_gen.vbackporch[3] ),
    .B(net298));
 sg13g2_o21ai_1 _2932_ (.B1(_0584_),
    .Y(_0106_),
    .A1(_0527_),
    .A2(_0578_));
 sg13g2_nand2_1 _2933_ (.Y(_0585_),
    .A(\hvsync_gen.vbackporch[4] ),
    .B(_0579_));
 sg13g2_o21ai_1 _2934_ (.B1(_0585_),
    .Y(_0107_),
    .A1(_0516_),
    .A2(_0578_));
 sg13g2_nand2_1 _2935_ (.Y(_0586_),
    .A(\hvsync_gen.vbackporch[5] ),
    .B(net298));
 sg13g2_o21ai_1 _2936_ (.B1(_0586_),
    .Y(_0108_),
    .A1(_0529_),
    .A2(_0579_));
 sg13g2_nand2_1 _2937_ (.Y(_0587_),
    .A(\hvsync_gen.vbackporch[6] ),
    .B(net298));
 sg13g2_o21ai_1 _2938_ (.B1(_0587_),
    .Y(_0109_),
    .A1(_0531_),
    .A2(_0578_));
 sg13g2_nand2_1 _2939_ (.Y(_0588_),
    .A(\hvsync_gen.vbackporch[7] ),
    .B(net298));
 sg13g2_o21ai_1 _2940_ (.B1(_0588_),
    .Y(_0110_),
    .A1(_0533_),
    .A2(_0578_));
 sg13g2_nand2_1 _2941_ (.Y(_0589_),
    .A(\hvsync_gen.vsyncpolarity ),
    .B(net290));
 sg13g2_o21ai_1 _2942_ (.B1(_0589_),
    .Y(_0111_),
    .A1(_0553_),
    .A2(net309));
 sg13g2_a21oi_2 _2943_ (.B1(_0486_),
    .Y(_0590_),
    .A2(_0492_),
    .A1(net375));
 sg13g2_nand2_1 _2944_ (.Y(_0591_),
    .A(\pat.pattern[0] ),
    .B(net303));
 sg13g2_nand2_1 _2945_ (.Y(_0592_),
    .A(_0486_),
    .B(_0490_));
 sg13g2_nand2_2 _2946_ (.Y(_0593_),
    .A(net300),
    .B(_0592_));
 sg13g2_nand3_1 _2947_ (.B(_0490_),
    .C(_0580_),
    .A(_0486_),
    .Y(_0594_));
 sg13g2_o21ai_1 _2948_ (.B1(_0594_),
    .Y(_0595_),
    .A1(_0025_),
    .A2(_0593_));
 sg13g2_o21ai_1 _2949_ (.B1(_0591_),
    .Y(_0112_),
    .A1(net303),
    .A2(_0595_));
 sg13g2_nand2_1 _2950_ (.Y(_0596_),
    .A(\pat.pattern[1] ),
    .B(net303));
 sg13g2_and2_2 _2951_ (.A(_0486_),
    .B(_0508_),
    .X(_0597_));
 sg13g2_nand2_1 _2952_ (.Y(_0598_),
    .A(_0486_),
    .B(_0508_));
 sg13g2_nor2_1 _2953_ (.A(_0026_),
    .B(_0598_),
    .Y(_0599_));
 sg13g2_nand2_1 _2954_ (.Y(_0600_),
    .A(_0026_),
    .B(_0598_));
 sg13g2_nor2b_1 _2955_ (.A(_0599_),
    .B_N(_0600_),
    .Y(_0601_));
 sg13g2_xnor2_1 _2956_ (.Y(_0602_),
    .A(_0025_),
    .B(_0601_));
 sg13g2_or3_1 _2957_ (.A(net9),
    .B(net299),
    .C(_0592_),
    .X(_0603_));
 sg13g2_o21ai_1 _2958_ (.B1(_0603_),
    .Y(_0604_),
    .A1(_0593_),
    .A2(_0602_));
 sg13g2_o21ai_1 _2959_ (.B1(_0596_),
    .Y(_0113_),
    .A1(net303),
    .A2(_0604_));
 sg13g2_nand2_1 _2960_ (.Y(_0605_),
    .A(net341),
    .B(_0597_));
 sg13g2_xnor2_1 _2961_ (.Y(_0606_),
    .A(net341),
    .B(_0597_));
 sg13g2_a21oi_1 _2962_ (.A1(\pat.pattern[0] ),
    .A2(_0600_),
    .Y(_0607_),
    .B1(_0599_));
 sg13g2_xor2_1 _2963_ (.B(_0607_),
    .A(_0606_),
    .X(_0608_));
 sg13g2_or2_1 _2964_ (.X(_0609_),
    .B(_0592_),
    .A(net10));
 sg13g2_o21ai_1 _2965_ (.B1(_0609_),
    .Y(_0610_),
    .A1(_0593_),
    .A2(_0608_));
 sg13g2_nand2_1 _2966_ (.Y(_0611_),
    .A(net341),
    .B(net303));
 sg13g2_o21ai_1 _2967_ (.B1(_0611_),
    .Y(_0114_),
    .A1(net303),
    .A2(_0610_));
 sg13g2_nand2_1 _2968_ (.Y(_0612_),
    .A(net339),
    .B(net303));
 sg13g2_o21ai_1 _2969_ (.B1(_0605_),
    .Y(_0613_),
    .A1(_0606_),
    .A2(_0607_));
 sg13g2_nand2_1 _2970_ (.Y(_0614_),
    .A(net339),
    .B(_0597_));
 sg13g2_xnor2_1 _2971_ (.Y(_0615_),
    .A(net339),
    .B(_0597_));
 sg13g2_xnor2_1 _2972_ (.Y(_0616_),
    .A(_0613_),
    .B(_0615_));
 sg13g2_nand3_1 _2973_ (.B(_0490_),
    .C(_0562_),
    .A(_0486_),
    .Y(_0617_));
 sg13g2_o21ai_1 _2974_ (.B1(_0617_),
    .Y(_0618_),
    .A1(_0593_),
    .A2(_0616_));
 sg13g2_o21ai_1 _2975_ (.B1(_0612_),
    .Y(_0115_),
    .A1(net303),
    .A2(_0618_));
 sg13g2_nand2_1 _2976_ (.Y(_0619_),
    .A(\pat.pattern[4] ),
    .B(_0590_));
 sg13g2_o21ai_1 _2977_ (.B1(_0614_),
    .Y(_0620_),
    .A1(_0597_),
    .A2(_0613_));
 sg13g2_a21oi_1 _2978_ (.A1(_0838_),
    .A2(_0613_),
    .Y(_0621_),
    .B1(_0620_));
 sg13g2_xnor2_1 _2979_ (.Y(_0622_),
    .A(net338),
    .B(_0621_));
 sg13g2_nand3_1 _2980_ (.B(_0490_),
    .C(_0528_),
    .A(_0486_),
    .Y(_0623_));
 sg13g2_o21ai_1 _2981_ (.B1(_0623_),
    .Y(_0624_),
    .A1(_0593_),
    .A2(_0622_));
 sg13g2_o21ai_1 _2982_ (.B1(_0619_),
    .Y(_0116_),
    .A1(_0590_),
    .A2(_0624_));
 sg13g2_nand2_1 _2983_ (.Y(_0625_),
    .A(net336),
    .B(net287));
 sg13g2_or2_1 _2984_ (.X(_0626_),
    .B(_1340_),
    .A(_0812_));
 sg13g2_xor2_1 _2985_ (.B(_1438_),
    .A(\hvsync_gen.vbackporch[7] ),
    .X(_0627_));
 sg13g2_nand3_1 _2986_ (.B(_0626_),
    .C(_0627_),
    .A(_1338_),
    .Y(_0628_));
 sg13g2_a21o_1 _2987_ (.A2(_0626_),
    .A1(_1338_),
    .B1(_0627_),
    .X(_0629_));
 sg13g2_nand2_1 _2988_ (.Y(_0630_),
    .A(\hvsync_gen.vbackporch[5] ),
    .B(_1352_));
 sg13g2_xnor2_1 _2989_ (.Y(_0631_),
    .A(_0812_),
    .B(_1340_));
 sg13g2_a21oi_1 _2990_ (.A1(_1349_),
    .A2(_0630_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_inv_1 _2991_ (.Y(_0633_),
    .A(_0632_));
 sg13g2_nand2_1 _2992_ (.Y(_0634_),
    .A(_0628_),
    .B(_0632_));
 sg13g2_xnor2_1 _2993_ (.Y(_0635_),
    .A(\hvsync_gen.vbackporch[5] ),
    .B(_1352_));
 sg13g2_or2_1 _2994_ (.X(_0636_),
    .B(_1361_),
    .A(_0805_));
 sg13g2_nand3_1 _2995_ (.B(_0635_),
    .C(_0636_),
    .A(_1360_),
    .Y(_0637_));
 sg13g2_a21oi_2 _2996_ (.B1(_1379_),
    .Y(_0638_),
    .A2(_1380_),
    .A1(\hvsync_gen.vbackporch[2] ));
 sg13g2_xnor2_1 _2997_ (.Y(_0639_),
    .A(\hvsync_gen.vbackporch[3] ),
    .B(_1371_));
 sg13g2_or2_1 _2998_ (.X(_0640_),
    .B(_0639_),
    .A(_0638_));
 sg13g2_a21oi_1 _2999_ (.A1(\hvsync_gen.vbackporch[1] ),
    .A2(_1421_),
    .Y(_0641_),
    .B1(_1385_));
 sg13g2_xnor2_1 _3000_ (.Y(_0642_),
    .A(\hvsync_gen.vbackporch[2] ),
    .B(_1380_));
 sg13g2_nor2_1 _3001_ (.A(_0641_),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_nand2_1 _3002_ (.Y(_0644_),
    .A(\hvsync_gen.vbackporch[0] ),
    .B(_1422_));
 sg13g2_xnor2_1 _3003_ (.Y(_0645_),
    .A(\hvsync_gen.vbackporch[1] ),
    .B(_1421_));
 sg13g2_nor2_1 _3004_ (.A(_0644_),
    .B(_0645_),
    .Y(_0646_));
 sg13g2_xor2_1 _3005_ (.B(_0642_),
    .A(_0641_),
    .X(_0647_));
 sg13g2_a21oi_1 _3006_ (.A1(_0646_),
    .A2(_0647_),
    .Y(_0648_),
    .B1(_0643_));
 sg13g2_and2_1 _3007_ (.A(_0638_),
    .B(_0639_),
    .X(_0649_));
 sg13g2_xor2_1 _3008_ (.B(_0639_),
    .A(_0638_),
    .X(_0650_));
 sg13g2_o21ai_1 _3009_ (.B1(_0640_),
    .Y(_0651_),
    .A1(_0648_),
    .A2(_0649_));
 sg13g2_xnor2_1 _3010_ (.Y(_0652_),
    .A(_0805_),
    .B(_1361_));
 sg13g2_a21oi_1 _3011_ (.A1(\hvsync_gen.vbackporch[3] ),
    .A2(_1371_),
    .Y(_0653_),
    .B1(_1370_));
 sg13g2_nor2_1 _3012_ (.A(_0652_),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_xor2_1 _3013_ (.B(_0653_),
    .A(_0652_),
    .X(_0655_));
 sg13g2_a21oi_1 _3014_ (.A1(_1360_),
    .A2(_0636_),
    .Y(_0656_),
    .B1(_0635_));
 sg13g2_a21o_1 _3015_ (.A2(_0636_),
    .A1(_1360_),
    .B1(_0635_),
    .X(_0657_));
 sg13g2_nand2_1 _3016_ (.Y(_0658_),
    .A(_0637_),
    .B(_0657_));
 sg13g2_nand3b_1 _3017_ (.B(_0651_),
    .C(_0655_),
    .Y(_0659_),
    .A_N(_0658_));
 sg13g2_a21oi_1 _3018_ (.A1(_0637_),
    .A2(_0654_),
    .Y(_0660_),
    .B1(_0656_));
 sg13g2_and3_1 _3019_ (.X(_0661_),
    .A(_0629_),
    .B(_0634_),
    .C(_0660_));
 sg13g2_nand3_1 _3020_ (.B(_0630_),
    .C(_0631_),
    .A(_1349_),
    .Y(_0662_));
 sg13g2_nand2_1 _3021_ (.Y(_0663_),
    .A(_0628_),
    .B(_0662_));
 sg13g2_a22oi_1 _3022_ (.Y(_0664_),
    .B1(_0663_),
    .B2(_0629_),
    .A2(_0661_),
    .A1(_0659_));
 sg13g2_a21oi_1 _3023_ (.A1(\hvsync_gen.vbackporch[7] ),
    .A2(_1331_),
    .Y(_0665_),
    .B1(_1330_));
 sg13g2_nor2b_1 _3024_ (.A(_0665_),
    .B_N(_1323_),
    .Y(_0666_));
 sg13g2_xnor2_1 _3025_ (.Y(_0667_),
    .A(_1323_),
    .B(_0665_));
 sg13g2_nor2b_1 _3026_ (.A(_1410_),
    .B_N(_0667_),
    .Y(_0668_));
 sg13g2_nor2_1 _3027_ (.A(_1396_),
    .B(_0666_),
    .Y(_0669_));
 sg13g2_nor2_1 _3028_ (.A(_1409_),
    .B(_0669_),
    .Y(_0670_));
 sg13g2_a21oi_1 _3029_ (.A1(_0664_),
    .A2(_0668_),
    .Y(_0671_),
    .B1(_0670_));
 sg13g2_xnor2_1 _3030_ (.Y(_0672_),
    .A(_1311_),
    .B(_1405_));
 sg13g2_nand2b_1 _3031_ (.Y(_0673_),
    .B(_0672_),
    .A_N(_0671_));
 sg13g2_o21ai_1 _3032_ (.B1(_0673_),
    .Y(_0674_),
    .A1(_1312_),
    .A2(_1405_));
 sg13g2_xor2_1 _3033_ (.B(_1399_),
    .A(_0014_),
    .X(_0675_));
 sg13g2_xnor2_1 _3034_ (.Y(_0676_),
    .A(_0674_),
    .B(_0675_));
 sg13g2_xnor2_1 _3035_ (.Y(_0677_),
    .A(_0671_),
    .B(_0672_));
 sg13g2_xnor2_1 _3036_ (.Y(_0678_),
    .A(_0013_),
    .B(_0677_));
 sg13g2_xor2_1 _3037_ (.B(_0667_),
    .A(_0664_),
    .X(_0679_));
 sg13g2_xnor2_1 _3038_ (.Y(_0680_),
    .A(_0817_),
    .B(_0679_));
 sg13g2_nand2_1 _3039_ (.Y(_0681_),
    .A(_0633_),
    .B(_0662_));
 sg13g2_a21o_1 _3040_ (.A2(_0660_),
    .A1(_0659_),
    .B1(_0681_),
    .X(_0682_));
 sg13g2_nand2_1 _3041_ (.Y(_0683_),
    .A(_0628_),
    .B(_0629_));
 sg13g2_xor2_1 _3042_ (.B(_0683_),
    .A(_0009_),
    .X(_0684_));
 sg13g2_a21oi_1 _3043_ (.A1(_0633_),
    .A2(_0682_),
    .Y(_0685_),
    .B1(_0684_));
 sg13g2_xor2_1 _3044_ (.B(_0655_),
    .A(_0651_),
    .X(_0686_));
 sg13g2_xnor2_1 _3045_ (.Y(_0687_),
    .A(_0648_),
    .B(_0650_));
 sg13g2_xor2_1 _3046_ (.B(_0647_),
    .A(_0646_),
    .X(_0688_));
 sg13g2_xnor2_1 _3047_ (.Y(_0689_),
    .A(_0644_),
    .B(_0645_));
 sg13g2_xnor2_1 _3048_ (.Y(_0690_),
    .A(net336),
    .B(_1422_));
 sg13g2_xnor2_1 _3049_ (.Y(_0691_),
    .A(\hvsync_gen.vbackporch[0] ),
    .B(_0690_));
 sg13g2_a21oi_1 _3050_ (.A1(_0651_),
    .A2(_0655_),
    .Y(_0692_),
    .B1(_0654_));
 sg13g2_xnor2_1 _3051_ (.Y(_0693_),
    .A(_0809_),
    .B(_0658_));
 sg13g2_or2_1 _3052_ (.X(_0694_),
    .B(_0686_),
    .A(_0006_));
 sg13g2_a21oi_1 _3053_ (.A1(_0004_),
    .A2(_0688_),
    .Y(_0695_),
    .B1(_0691_));
 sg13g2_o21ai_1 _3054_ (.B1(_0695_),
    .Y(_0696_),
    .A1(_0005_),
    .A2(_0687_));
 sg13g2_a21oi_1 _3055_ (.A1(_0006_),
    .A2(_0686_),
    .Y(_0697_),
    .B1(_0696_));
 sg13g2_xnor2_1 _3056_ (.Y(_0698_),
    .A(_0003_),
    .B(_0689_));
 sg13g2_o21ai_1 _3057_ (.B1(_0698_),
    .Y(_0699_),
    .A1(_0004_),
    .A2(_0688_));
 sg13g2_a21oi_1 _3058_ (.A1(_0005_),
    .A2(_0687_),
    .Y(_0700_),
    .B1(_0699_));
 sg13g2_nand3_1 _3059_ (.B(_0697_),
    .C(_0700_),
    .A(_0694_),
    .Y(_0701_));
 sg13g2_xnor2_1 _3060_ (.Y(_0702_),
    .A(_0692_),
    .B(_0693_));
 sg13g2_nand3_1 _3061_ (.B(_0660_),
    .C(_0681_),
    .A(_0659_),
    .Y(_0703_));
 sg13g2_a21oi_1 _3062_ (.A1(_0682_),
    .A2(_0703_),
    .Y(_0704_),
    .B1(net322));
 sg13g2_nand3_1 _3063_ (.B(_0682_),
    .C(_0684_),
    .A(_0633_),
    .Y(_0705_));
 sg13g2_nand3_1 _3064_ (.B(_0682_),
    .C(_0703_),
    .A(net322),
    .Y(_0706_));
 sg13g2_nand3b_1 _3065_ (.B(_0705_),
    .C(_0706_),
    .Y(_0707_),
    .A_N(_0704_));
 sg13g2_nor4_2 _3066_ (.A(_0685_),
    .B(_0701_),
    .C(_0702_),
    .Y(_0708_),
    .D(_0707_));
 sg13g2_a21oi_1 _3067_ (.A1(_0664_),
    .A2(_0667_),
    .Y(_0709_),
    .B1(_0666_));
 sg13g2_xnor2_1 _3068_ (.Y(_0710_),
    .A(_0012_),
    .B(_1410_));
 sg13g2_xnor2_1 _3069_ (.Y(_0711_),
    .A(_0709_),
    .B(_0710_));
 sg13g2_nand3_1 _3070_ (.B(_0708_),
    .C(_0711_),
    .A(_0680_),
    .Y(_0712_));
 sg13g2_nor3_1 _3071_ (.A(_0676_),
    .B(_0678_),
    .C(_0712_),
    .Y(_0713_));
 sg13g2_or3_1 _3072_ (.A(_0796_),
    .B(_0462_),
    .C(_0713_),
    .X(_0714_));
 sg13g2_o21ai_1 _3073_ (.B1(_0625_),
    .Y(_0117_),
    .A1(_0793_),
    .A2(net285));
 sg13g2_nand2_1 _3074_ (.Y(_0715_),
    .A(net335),
    .B(net287));
 sg13g2_o21ai_1 _3075_ (.B1(_0715_),
    .Y(_0118_),
    .A1(_1018_),
    .A2(net285));
 sg13g2_nand2_1 _3076_ (.Y(_0716_),
    .A(net333),
    .B(net287));
 sg13g2_xnor2_1 _3077_ (.Y(_0717_),
    .A(_0800_),
    .B(_0894_));
 sg13g2_o21ai_1 _3078_ (.B1(_0716_),
    .Y(_0119_),
    .A1(net285),
    .A2(_0717_));
 sg13g2_nand2_1 _3079_ (.Y(_0718_),
    .A(net330),
    .B(net287));
 sg13g2_xnor2_1 _3080_ (.Y(_0719_),
    .A(net330),
    .B(_0934_));
 sg13g2_o21ai_1 _3081_ (.B1(_0718_),
    .Y(_0120_),
    .A1(net285),
    .A2(_0719_));
 sg13g2_nand2_1 _3082_ (.Y(_0720_),
    .A(net329),
    .B(net288));
 sg13g2_xnor2_1 _3083_ (.Y(_0721_),
    .A(_0804_),
    .B(_0895_));
 sg13g2_o21ai_1 _3084_ (.B1(_0720_),
    .Y(_0121_),
    .A1(net285),
    .A2(_0721_));
 sg13g2_nand2_1 _3085_ (.Y(_0722_),
    .A(net326),
    .B(net287));
 sg13g2_xnor2_1 _3086_ (.Y(_0723_),
    .A(net327),
    .B(_0929_));
 sg13g2_o21ai_1 _3087_ (.B1(_0722_),
    .Y(_0122_),
    .A1(net285),
    .A2(_0723_));
 sg13g2_nand2_1 _3088_ (.Y(_0724_),
    .A(net323),
    .B(net288));
 sg13g2_xnor2_1 _3089_ (.Y(_0725_),
    .A(net324),
    .B(_0922_));
 sg13g2_o21ai_1 _3090_ (.B1(_0724_),
    .Y(_0123_),
    .A1(net286),
    .A2(_0725_));
 sg13g2_nand2_1 _3091_ (.Y(_0726_),
    .A(net321),
    .B(net288));
 sg13g2_nor3_1 _3092_ (.A(net322),
    .B(_0895_),
    .C(_0921_),
    .Y(_0727_));
 sg13g2_xnor2_1 _3093_ (.Y(_0728_),
    .A(net321),
    .B(_0727_));
 sg13g2_o21ai_1 _3094_ (.B1(_0726_),
    .Y(_0124_),
    .A1(net285),
    .A2(_0728_));
 sg13g2_nand2_1 _3095_ (.Y(_0729_),
    .A(net319),
    .B(_0463_));
 sg13g2_nand3_1 _3096_ (.B(net320),
    .C(_0922_),
    .A(net323),
    .Y(_0730_));
 sg13g2_inv_1 _3097_ (.Y(_0731_),
    .A(_0730_));
 sg13g2_xnor2_1 _3098_ (.Y(_0732_),
    .A(_0815_),
    .B(_0730_));
 sg13g2_o21ai_1 _3099_ (.B1(_0729_),
    .Y(_0125_),
    .A1(net286),
    .A2(_0732_));
 sg13g2_nand2_1 _3100_ (.Y(_0733_),
    .A(net318),
    .B(net288));
 sg13g2_nor2_1 _3101_ (.A(net166),
    .B(_0730_),
    .Y(_0734_));
 sg13g2_xnor2_1 _3102_ (.Y(_0735_),
    .A(net318),
    .B(_0734_));
 sg13g2_o21ai_1 _3103_ (.B1(_0733_),
    .Y(_0126_),
    .A1(net286),
    .A2(_0735_));
 sg13g2_nand2_1 _3104_ (.Y(_0736_),
    .A(net154),
    .B(net288));
 sg13g2_nand3_1 _3105_ (.B(net318),
    .C(_0731_),
    .A(net319),
    .Y(_0737_));
 sg13g2_xor2_1 _3106_ (.B(_0737_),
    .A(net154),
    .X(_0738_));
 sg13g2_o21ai_1 _3107_ (.B1(_0736_),
    .Y(_0127_),
    .A1(net286),
    .A2(_0738_));
 sg13g2_nand2_1 _3108_ (.Y(_0739_),
    .A(net150),
    .B(net288));
 sg13g2_nor2_1 _3109_ (.A(_0013_),
    .B(_0737_),
    .Y(_0740_));
 sg13g2_xnor2_1 _3110_ (.Y(_0741_),
    .A(net150),
    .B(_0740_));
 sg13g2_o21ai_1 _3111_ (.B1(_0739_),
    .Y(_0128_),
    .A1(net285),
    .A2(_0741_));
 sg13g2_nor2b_2 _3112_ (.A(_0489_),
    .B_N(_0491_),
    .Y(_0742_));
 sg13g2_o21ai_1 _3113_ (.B1(_0491_),
    .Y(_0743_),
    .A1(net377),
    .A2(net313));
 sg13g2_nor3_2 _3114_ (.A(_0485_),
    .B(_0490_),
    .C(_0491_),
    .Y(_0744_));
 sg13g2_or2_1 _3115_ (.X(_0745_),
    .B(net308),
    .A(_0522_));
 sg13g2_a21oi_1 _3116_ (.A1(_0840_),
    .A2(net308),
    .Y(_0746_),
    .B1(_0742_));
 sg13g2_a22oi_1 _3117_ (.Y(_0129_),
    .B1(_0745_),
    .B2(_0746_),
    .A2(_0742_),
    .A1(_0840_));
 sg13g2_nor2_1 _3118_ (.A(_0491_),
    .B(_0509_),
    .Y(_0747_));
 sg13g2_inv_1 _3119_ (.Y(_0748_),
    .A(net307));
 sg13g2_xnor2_1 _3120_ (.Y(_0749_),
    .A(_0028_),
    .B(net307));
 sg13g2_or2_1 _3121_ (.X(_0750_),
    .B(_0749_),
    .A(\color_in[0] ));
 sg13g2_nand2_1 _3122_ (.Y(_0751_),
    .A(\color_in[0] ),
    .B(_0749_));
 sg13g2_nand3_1 _3123_ (.B(_0750_),
    .C(_0751_),
    .A(_0744_),
    .Y(_0752_));
 sg13g2_o21ai_1 _3124_ (.B1(_0752_),
    .Y(_0753_),
    .A1(_0499_),
    .A2(net308));
 sg13g2_mux2_1 _3125_ (.A0(\color_in[1] ),
    .A1(_0753_),
    .S(_0743_),
    .X(_0130_));
 sg13g2_o21ai_1 _3126_ (.B1(_0751_),
    .Y(_0754_),
    .A1(_0028_),
    .A2(_0748_));
 sg13g2_xnor2_1 _3127_ (.Y(_0755_),
    .A(_0029_),
    .B(net307));
 sg13g2_xor2_1 _3128_ (.B(_0755_),
    .A(_0754_),
    .X(_0756_));
 sg13g2_o21ai_1 _3129_ (.B1(_0743_),
    .Y(_0757_),
    .A1(_0525_),
    .A2(net308));
 sg13g2_a21oi_1 _3130_ (.A1(net308),
    .A2(_0756_),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_a21oi_1 _3131_ (.A1(_0841_),
    .A2(_0742_),
    .Y(_0131_),
    .B1(_0758_));
 sg13g2_a22oi_1 _3132_ (.Y(_0759_),
    .B1(_0754_),
    .B2(_0755_),
    .A2(net307),
    .A1(\color_in[2] ));
 sg13g2_xnor2_1 _3133_ (.Y(_0760_),
    .A(_0030_),
    .B(net307));
 sg13g2_nand2b_1 _3134_ (.Y(_0761_),
    .B(_0760_),
    .A_N(_0759_));
 sg13g2_xor2_1 _3135_ (.B(_0760_),
    .A(_0759_),
    .X(_0762_));
 sg13g2_mux2_1 _3136_ (.A0(_0527_),
    .A1(_0762_),
    .S(net308),
    .X(_0763_));
 sg13g2_nand2_1 _3137_ (.Y(_0764_),
    .A(\color_in[3] ),
    .B(_0742_));
 sg13g2_o21ai_1 _3138_ (.B1(_0764_),
    .Y(_0132_),
    .A1(_0742_),
    .A2(_0763_));
 sg13g2_nand2_1 _3139_ (.Y(_0765_),
    .A(\color_in[3] ),
    .B(net307));
 sg13g2_xnor2_1 _3140_ (.Y(_0766_),
    .A(\color_in[4] ),
    .B(_0747_));
 sg13g2_nand3_1 _3141_ (.B(_0765_),
    .C(_0766_),
    .A(_0761_),
    .Y(_0767_));
 sg13g2_a21oi_1 _3142_ (.A1(_0761_),
    .A2(_0765_),
    .Y(_0768_),
    .B1(_0766_));
 sg13g2_nor2b_1 _3143_ (.A(_0768_),
    .B_N(net308),
    .Y(_0769_));
 sg13g2_o21ai_1 _3144_ (.B1(_0743_),
    .Y(_0770_),
    .A1(_0516_),
    .A2(_0744_));
 sg13g2_a21oi_1 _3145_ (.A1(_0767_),
    .A2(_0769_),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_a21oi_1 _3146_ (.A1(_0842_),
    .A2(_0742_),
    .Y(_0133_),
    .B1(_0771_));
 sg13g2_a21oi_1 _3147_ (.A1(\color_in[4] ),
    .A2(net307),
    .Y(_0772_),
    .B1(_0768_));
 sg13g2_xnor2_1 _3148_ (.Y(_0773_),
    .A(_0843_),
    .B(net307));
 sg13g2_xnor2_1 _3149_ (.Y(_0774_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_o21ai_1 _3150_ (.B1(_0743_),
    .Y(_0775_),
    .A1(_0565_),
    .A2(_0744_));
 sg13g2_a21oi_1 _3151_ (.A1(net308),
    .A2(_0774_),
    .Y(_0776_),
    .B1(_0775_));
 sg13g2_a21oi_1 _3152_ (.A1(_0843_),
    .A2(_0742_),
    .Y(_0134_),
    .B1(_0776_));
 sg13g2_a21oi_1 _3153_ (.A1(net375),
    .A2(_0492_),
    .Y(_0777_),
    .B1(_0488_));
 sg13g2_nand2_1 _3154_ (.Y(_0778_),
    .A(\hdisplay[0] ),
    .B(net296));
 sg13g2_o21ai_1 _3155_ (.B1(_0778_),
    .Y(_0135_),
    .A1(net313),
    .A2(_0522_));
 sg13g2_nand2_1 _3156_ (.Y(_0779_),
    .A(\hdisplay[1] ),
    .B(net296));
 sg13g2_o21ai_1 _3157_ (.B1(_0779_),
    .Y(_0136_),
    .A1(net313),
    .A2(_0499_));
 sg13g2_nand2_1 _3158_ (.Y(_0780_),
    .A(\hdisplay[2] ),
    .B(net296));
 sg13g2_o21ai_1 _3159_ (.B1(_0780_),
    .Y(_0137_),
    .A1(net313),
    .A2(_0525_));
 sg13g2_nand2_1 _3160_ (.Y(_0781_),
    .A(\hdisplay[3] ),
    .B(net296));
 sg13g2_o21ai_1 _3161_ (.B1(_0781_),
    .Y(_0138_),
    .A1(net313),
    .A2(_0527_));
 sg13g2_nand2_1 _3162_ (.Y(_0782_),
    .A(\hdisplay[4] ),
    .B(net296));
 sg13g2_o21ai_1 _3163_ (.B1(_0782_),
    .Y(_0139_),
    .A1(net313),
    .A2(_0516_));
 sg13g2_nand2_1 _3164_ (.Y(_0783_),
    .A(\hdisplay[5] ),
    .B(net296));
 sg13g2_o21ai_1 _3165_ (.B1(_0783_),
    .Y(_0140_),
    .A1(net314),
    .A2(_0565_));
 sg13g2_nand2_1 _3166_ (.Y(_0784_),
    .A(\hdisplay[6] ),
    .B(net297));
 sg13g2_o21ai_1 _3167_ (.B1(_0784_),
    .Y(_0141_),
    .A1(net314),
    .A2(_0531_));
 sg13g2_nand2_1 _3168_ (.Y(_0785_),
    .A(\hdisplay[7] ),
    .B(net297));
 sg13g2_o21ai_1 _3169_ (.B1(_0785_),
    .Y(_0142_),
    .A1(_0549_),
    .A2(net297));
 sg13g2_nand2_1 _3170_ (.Y(_0786_),
    .A(\hdisplay[8] ),
    .B(net297));
 sg13g2_o21ai_1 _3171_ (.B1(_0786_),
    .Y(_0143_),
    .A1(net314),
    .A2(_0535_));
 sg13g2_nor2_1 _3172_ (.A(net6),
    .B(net314),
    .Y(_0787_));
 sg13g2_a22oi_1 _3173_ (.Y(_0144_),
    .B1(_0787_),
    .B2(net301),
    .A2(net296),
    .A1(_0835_));
 sg13g2_nand2_1 _3174_ (.Y(_0788_),
    .A(\hdisplay[10] ),
    .B(net296));
 sg13g2_o21ai_1 _3175_ (.B1(_0788_),
    .Y(_0145_),
    .A1(net314),
    .A2(_0553_));
 sg13g2_dfrbp_1 _3176_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net143),
    .D(_0033_),
    .Q_N(_0032_),
    .Q(\hpos[0] ));
 sg13g2_dfrbp_1 _3177_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net104),
    .D(_0034_),
    .Q_N(_0015_),
    .Q(\hpos[1] ));
 sg13g2_dfrbp_1 _3178_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net103),
    .D(_0035_),
    .Q_N(_0016_),
    .Q(\hpos[2] ));
 sg13g2_dfrbp_1 _3179_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net102),
    .D(_0036_),
    .Q_N(_0017_),
    .Q(\hpos[3] ));
 sg13g2_dfrbp_1 _3180_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net101),
    .D(_0037_),
    .Q_N(_0018_),
    .Q(\hpos[4] ));
 sg13g2_dfrbp_1 _3181_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net100),
    .D(_0038_),
    .Q_N(_0019_),
    .Q(\hpos[5] ));
 sg13g2_dfrbp_1 _3182_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net99),
    .D(_0039_),
    .Q_N(_0020_),
    .Q(\hpos[6] ));
 sg13g2_dfrbp_1 _3183_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net98),
    .D(_0040_),
    .Q_N(_0021_),
    .Q(\hpos[7] ));
 sg13g2_dfrbp_1 _3184_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net97),
    .D(_0041_),
    .Q_N(_0022_),
    .Q(\hpos[8] ));
 sg13g2_dfrbp_1 _3185_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net96),
    .D(_0042_),
    .Q_N(_1584_),
    .Q(\hpos[9] ));
 sg13g2_dfrbp_1 _3186_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net95),
    .D(_0043_),
    .Q_N(_0023_),
    .Q(\hpos[10] ));
 sg13g2_dfrbp_1 _3187_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net94),
    .D(_0044_),
    .Q_N(_0024_),
    .Q(\hpos[11] ));
 sg13g2_dfrbp_1 _3188_ (.CLK(net364),
    .RESET_B(net93),
    .D(_0045_),
    .Q_N(_1583_),
    .Q(\hfrontporch[0] ));
 sg13g2_dfrbp_1 _3189_ (.CLK(net363),
    .RESET_B(net91),
    .D(_0046_),
    .Q_N(_1582_),
    .Q(\hfrontporch[1] ));
 sg13g2_dfrbp_1 _3190_ (.CLK(net363),
    .RESET_B(net89),
    .D(_0047_),
    .Q_N(_1581_),
    .Q(\hfrontporch[2] ));
 sg13g2_dfrbp_1 _3191_ (.CLK(net367),
    .RESET_B(net87),
    .D(_0048_),
    .Q_N(_1580_),
    .Q(\hfrontporch[3] ));
 sg13g2_dfrbp_1 _3192_ (.CLK(net366),
    .RESET_B(net85),
    .D(_0049_),
    .Q_N(_1579_),
    .Q(\hfrontporch[4] ));
 sg13g2_dfrbp_1 _3193_ (.CLK(net370),
    .RESET_B(net83),
    .D(_0050_),
    .Q_N(_1578_),
    .Q(\hfrontporch[5] ));
 sg13g2_dfrbp_1 _3194_ (.CLK(net370),
    .RESET_B(net81),
    .D(_0051_),
    .Q_N(_1577_),
    .Q(\hfrontporch[6] ));
 sg13g2_dfrbp_1 _3195_ (.CLK(net371),
    .RESET_B(net79),
    .D(_0052_),
    .Q_N(_1576_),
    .Q(\hfrontporch[7] ));
 sg13g2_dfrbp_1 _3196_ (.CLK(net373),
    .RESET_B(net77),
    .D(_0053_),
    .Q_N(_1575_),
    .Q(\hfrontporch[8] ));
 sg13g2_dfrbp_1 _3197_ (.CLK(net371),
    .RESET_B(net75),
    .D(_0054_),
    .Q_N(_1574_),
    .Q(\hfrontporch[9] ));
 sg13g2_dfrbp_1 _3198_ (.CLK(net363),
    .RESET_B(net73),
    .D(_0055_),
    .Q_N(_1573_),
    .Q(\hsynclength[0] ));
 sg13g2_dfrbp_1 _3199_ (.CLK(net363),
    .RESET_B(net71),
    .D(_0056_),
    .Q_N(_1572_),
    .Q(\hsynclength[1] ));
 sg13g2_dfrbp_1 _3200_ (.CLK(net363),
    .RESET_B(net69),
    .D(_0057_),
    .Q_N(_1571_),
    .Q(\hsynclength[2] ));
 sg13g2_dfrbp_1 _3201_ (.CLK(net364),
    .RESET_B(net67),
    .D(_0058_),
    .Q_N(_1570_),
    .Q(\hsynclength[3] ));
 sg13g2_dfrbp_1 _3202_ (.CLK(net366),
    .RESET_B(net65),
    .D(_0059_),
    .Q_N(_1569_),
    .Q(\hsynclength[4] ));
 sg13g2_dfrbp_1 _3203_ (.CLK(net366),
    .RESET_B(net63),
    .D(_0060_),
    .Q_N(_1568_),
    .Q(\hsynclength[5] ));
 sg13g2_dfrbp_1 _3204_ (.CLK(net370),
    .RESET_B(net61),
    .D(_0061_),
    .Q_N(_1567_),
    .Q(\hsynclength[6] ));
 sg13g2_dfrbp_1 _3205_ (.CLK(net371),
    .RESET_B(net59),
    .D(_0062_),
    .Q_N(_1566_),
    .Q(\hsynclength[7] ));
 sg13g2_dfrbp_1 _3206_ (.CLK(net371),
    .RESET_B(net57),
    .D(_0063_),
    .Q_N(_1565_),
    .Q(\hsynclength[8] ));
 sg13g2_dfrbp_1 _3207_ (.CLK(net371),
    .RESET_B(net55),
    .D(_0064_),
    .Q_N(_1564_),
    .Q(\hsynclength[9] ));
 sg13g2_dfrbp_1 _3208_ (.CLK(net365),
    .RESET_B(net53),
    .D(_0065_),
    .Q_N(_1563_),
    .Q(\hbackporch[0] ));
 sg13g2_dfrbp_1 _3209_ (.CLK(net365),
    .RESET_B(net51),
    .D(_0066_),
    .Q_N(_1562_),
    .Q(\hbackporch[1] ));
 sg13g2_dfrbp_1 _3210_ (.CLK(net363),
    .RESET_B(net49),
    .D(_0067_),
    .Q_N(_1561_),
    .Q(\hbackporch[2] ));
 sg13g2_dfrbp_1 _3211_ (.CLK(net364),
    .RESET_B(net47),
    .D(_0068_),
    .Q_N(_1560_),
    .Q(\hbackporch[3] ));
 sg13g2_dfrbp_1 _3212_ (.CLK(net367),
    .RESET_B(net45),
    .D(_0069_),
    .Q_N(_1559_),
    .Q(\hbackporch[4] ));
 sg13g2_dfrbp_1 _3213_ (.CLK(net373),
    .RESET_B(net43),
    .D(_0070_),
    .Q_N(_1558_),
    .Q(\hbackporch[5] ));
 sg13g2_dfrbp_1 _3214_ (.CLK(net370),
    .RESET_B(net40),
    .D(_0071_),
    .Q_N(_1557_),
    .Q(\hbackporch[6] ));
 sg13g2_dfrbp_1 _3215_ (.CLK(net371),
    .RESET_B(net38),
    .D(_0072_),
    .Q_N(_1556_),
    .Q(\hbackporch[7] ));
 sg13g2_dfrbp_1 _3216_ (.CLK(net371),
    .RESET_B(net36),
    .D(_0073_),
    .Q_N(_1555_),
    .Q(\hbackporch[8] ));
 sg13g2_dfrbp_1 _3217_ (.CLK(net372),
    .RESET_B(net34),
    .D(_0074_),
    .Q_N(_1554_),
    .Q(\hbackporch[9] ));
 sg13g2_dfrbp_1 _3218_ (.CLK(net360),
    .RESET_B(net32),
    .D(_0075_),
    .Q_N(_1553_),
    .Q(\hvsync_gen.vdisplay[0] ));
 sg13g2_dfrbp_1 _3219_ (.CLK(net360),
    .RESET_B(net145),
    .D(_0076_),
    .Q_N(_1552_),
    .Q(\hvsync_gen.vdisplay[1] ));
 sg13g2_dfrbp_1 _3220_ (.CLK(net360),
    .RESET_B(net142),
    .D(_0077_),
    .Q_N(_1551_),
    .Q(\hvsync_gen.vdisplay[2] ));
 sg13g2_dfrbp_1 _3221_ (.CLK(net362),
    .RESET_B(net140),
    .D(_0078_),
    .Q_N(_1550_),
    .Q(\hvsync_gen.vdisplay[3] ));
 sg13g2_dfrbp_1 _3222_ (.CLK(net362),
    .RESET_B(net138),
    .D(_0079_),
    .Q_N(_1549_),
    .Q(\hvsync_gen.vdisplay[4] ));
 sg13g2_dfrbp_1 _3223_ (.CLK(net369),
    .RESET_B(net136),
    .D(_0080_),
    .Q_N(_1548_),
    .Q(\hvsync_gen.vdisplay[5] ));
 sg13g2_dfrbp_1 _3224_ (.CLK(net368),
    .RESET_B(net134),
    .D(_0081_),
    .Q_N(_1547_),
    .Q(\hvsync_gen.vdisplay[6] ));
 sg13g2_dfrbp_1 _3225_ (.CLK(net372),
    .RESET_B(net132),
    .D(_0082_),
    .Q_N(_1546_),
    .Q(\hvsync_gen.vdisplay[7] ));
 sg13g2_dfrbp_1 _3226_ (.CLK(net368),
    .RESET_B(net130),
    .D(_0083_),
    .Q_N(_0011_),
    .Q(\hvsync_gen.vdisplay[8] ));
 sg13g2_dfrbp_1 _3227_ (.CLK(net372),
    .RESET_B(net128),
    .D(_0084_),
    .Q_N(_1545_),
    .Q(\hvsync_gen.vdisplay[9] ));
 sg13g2_dfrbp_1 _3228_ (.CLK(net368),
    .RESET_B(net126),
    .D(_0085_),
    .Q_N(_0002_),
    .Q(\hvsync_gen.vdisplay[10] ));
 sg13g2_dfrbp_1 _3229_ (.CLK(net372),
    .RESET_B(net124),
    .D(_0086_),
    .Q_N(_1544_),
    .Q(hsyncpolarity));
 sg13g2_dfrbp_1 _3230_ (.CLK(net360),
    .RESET_B(net123),
    .D(_0087_),
    .Q_N(_1543_),
    .Q(\hvsync_gen.vfrontporch[0] ));
 sg13g2_dfrbp_1 _3231_ (.CLK(net360),
    .RESET_B(net121),
    .D(_0088_),
    .Q_N(_1542_),
    .Q(\hvsync_gen.vfrontporch[1] ));
 sg13g2_dfrbp_1 _3232_ (.CLK(net361),
    .RESET_B(net119),
    .D(_0089_),
    .Q_N(_1541_),
    .Q(\hvsync_gen.vfrontporch[2] ));
 sg13g2_dfrbp_1 _3233_ (.CLK(net360),
    .RESET_B(net117),
    .D(_0090_),
    .Q_N(_1540_),
    .Q(\hvsync_gen.vfrontporch[3] ));
 sg13g2_dfrbp_1 _3234_ (.CLK(net369),
    .RESET_B(net115),
    .D(_0091_),
    .Q_N(_1539_),
    .Q(\hvsync_gen.vfrontporch[4] ));
 sg13g2_dfrbp_1 _3235_ (.CLK(net369),
    .RESET_B(net113),
    .D(_0092_),
    .Q_N(_1538_),
    .Q(\hvsync_gen.vfrontporch[5] ));
 sg13g2_dfrbp_1 _3236_ (.CLK(net368),
    .RESET_B(net111),
    .D(_0093_),
    .Q_N(_1537_),
    .Q(\hvsync_gen.vfrontporch[6] ));
 sg13g2_dfrbp_1 _3237_ (.CLK(net368),
    .RESET_B(net109),
    .D(_0094_),
    .Q_N(_1536_),
    .Q(\hvsync_gen.vfrontporch[7] ));
 sg13g2_dfrbp_1 _3238_ (.CLK(net360),
    .RESET_B(net107),
    .D(_0095_),
    .Q_N(_1535_),
    .Q(\hvsync_gen.vsynclength[0] ));
 sg13g2_dfrbp_1 _3239_ (.CLK(net362),
    .RESET_B(net105),
    .D(_0096_),
    .Q_N(_1534_),
    .Q(\hvsync_gen.vsynclength[1] ));
 sg13g2_dfrbp_1 _3240_ (.CLK(net360),
    .RESET_B(net90),
    .D(_0097_),
    .Q_N(_1533_),
    .Q(\hvsync_gen.vsynclength[2] ));
 sg13g2_dfrbp_1 _3241_ (.CLK(net362),
    .RESET_B(net86),
    .D(_0098_),
    .Q_N(_1532_),
    .Q(\hvsync_gen.vsynclength[3] ));
 sg13g2_dfrbp_1 _3242_ (.CLK(net362),
    .RESET_B(net82),
    .D(_0099_),
    .Q_N(_1531_),
    .Q(\hvsync_gen.vsynclength[4] ));
 sg13g2_dfrbp_1 _3243_ (.CLK(net369),
    .RESET_B(net78),
    .D(_0100_),
    .Q_N(_1530_),
    .Q(\hvsync_gen.vsynclength[5] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(net368),
    .RESET_B(net74),
    .D(_0101_),
    .Q_N(_1529_),
    .Q(\hvsync_gen.vsynclength[6] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(net368),
    .RESET_B(net70),
    .D(_0102_),
    .Q_N(_1528_),
    .Q(\hvsync_gen.vsynclength[7] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(net361),
    .RESET_B(net66),
    .D(_0103_),
    .Q_N(_1527_),
    .Q(\hvsync_gen.vbackporch[0] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(net361),
    .RESET_B(net62),
    .D(_0104_),
    .Q_N(_1526_),
    .Q(\hvsync_gen.vbackporch[1] ));
 sg13g2_dfrbp_1 _3248_ (.CLK(net361),
    .RESET_B(net58),
    .D(_0105_),
    .Q_N(_1525_),
    .Q(\hvsync_gen.vbackporch[2] ));
 sg13g2_dfrbp_1 _3249_ (.CLK(net362),
    .RESET_B(net54),
    .D(_0106_),
    .Q_N(_1524_),
    .Q(\hvsync_gen.vbackporch[3] ));
 sg13g2_dfrbp_1 _3250_ (.CLK(net362),
    .RESET_B(net50),
    .D(_0107_),
    .Q_N(_1523_),
    .Q(\hvsync_gen.vbackporch[4] ));
 sg13g2_dfrbp_1 _3251_ (.CLK(net369),
    .RESET_B(net46),
    .D(_0108_),
    .Q_N(_1522_),
    .Q(\hvsync_gen.vbackporch[5] ));
 sg13g2_dfrbp_1 _3252_ (.CLK(net369),
    .RESET_B(net42),
    .D(_0109_),
    .Q_N(_1521_),
    .Q(\hvsync_gen.vbackporch[6] ));
 sg13g2_dfrbp_1 _3253_ (.CLK(net368),
    .RESET_B(net37),
    .D(_0110_),
    .Q_N(_1520_),
    .Q(\hvsync_gen.vbackporch[7] ));
 sg13g2_dfrbp_1 _3254_ (.CLK(net369),
    .RESET_B(net33),
    .D(_0111_),
    .Q_N(_1519_),
    .Q(\hvsync_gen.vsyncpolarity ));
 sg13g2_dfrbp_1 _3255_ (.CLK(net365),
    .RESET_B(net146),
    .D(_0112_),
    .Q_N(_0025_),
    .Q(\pat.pattern[0] ));
 sg13g2_dfrbp_1 _3256_ (.CLK(net365),
    .RESET_B(net144),
    .D(_0113_),
    .Q_N(_0026_),
    .Q(\pat.pattern[1] ));
 sg13g2_dfrbp_1 _3257_ (.CLK(net361),
    .RESET_B(net141),
    .D(_0114_),
    .Q_N(_1518_),
    .Q(\pat.pattern[2] ));
 sg13g2_dfrbp_1 _3258_ (.CLK(net361),
    .RESET_B(net139),
    .D(_0115_),
    .Q_N(_1517_),
    .Q(\pat.pattern[3] ));
 sg13g2_dfrbp_1 _3259_ (.CLK(net361),
    .RESET_B(net41),
    .D(_0116_),
    .Q_N(_0027_),
    .Q(\pat.pattern[4] ));
 sg13g2_dfrbp_1 _3260_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net137),
    .D(_0000_),
    .Q_N(_1516_),
    .Q(hsync));
 sg13g2_dfrbp_1 _3261_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net135),
    .D(net149),
    .Q_N(_0031_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _3262_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net131),
    .D(_0118_),
    .Q_N(_0003_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _3263_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net127),
    .D(_0119_),
    .Q_N(_0004_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _3264_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(_0120_),
    .Q_N(_0005_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _3265_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net118),
    .D(_0121_),
    .Q_N(_0006_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _3266_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net114),
    .D(_0122_),
    .Q_N(_0007_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _3267_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net110),
    .D(_0123_),
    .Q_N(_0008_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _3268_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net106),
    .D(_0124_),
    .Q_N(_0009_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _3269_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net88),
    .D(_0125_),
    .Q_N(_0010_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _3270_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net80),
    .D(net167),
    .Q_N(_0012_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _3271_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net72),
    .D(_0127_),
    .Q_N(_0013_),
    .Q(\hvsync_gen.vpos[10] ));
 sg13g2_dfrbp_1 _3272_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net92),
    .D(net151),
    .Q_N(_0014_),
    .Q(\hvsync_gen.vpos[11] ));
 sg13g2_dfrbp_1 _3273_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net64),
    .D(_0001_),
    .Q_N(_1515_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _3274_ (.CLK(net366),
    .RESET_B(net56),
    .D(_0129_),
    .Q_N(_1514_),
    .Q(\color_in[0] ));
 sg13g2_dfrbp_1 _3275_ (.CLK(net366),
    .RESET_B(net52),
    .D(_0130_),
    .Q_N(_0028_),
    .Q(\color_in[1] ));
 sg13g2_dfrbp_1 _3276_ (.CLK(net366),
    .RESET_B(net48),
    .D(_0131_),
    .Q_N(_0029_),
    .Q(\color_in[2] ));
 sg13g2_dfrbp_1 _3277_ (.CLK(net370),
    .RESET_B(net44),
    .D(_0132_),
    .Q_N(_0030_),
    .Q(\color_in[3] ));
 sg13g2_dfrbp_1 _3278_ (.CLK(net370),
    .RESET_B(net39),
    .D(_0133_),
    .Q_N(_1513_),
    .Q(\color_in[4] ));
 sg13g2_dfrbp_1 _3279_ (.CLK(net370),
    .RESET_B(net35),
    .D(_0134_),
    .Q_N(_1512_),
    .Q(\color_in[5] ));
 sg13g2_dfrbp_1 _3280_ (.CLK(net365),
    .RESET_B(net133),
    .D(_0135_),
    .Q_N(_1511_),
    .Q(\hdisplay[0] ));
 sg13g2_dfrbp_1 _3281_ (.CLK(net363),
    .RESET_B(net125),
    .D(_0136_),
    .Q_N(_1510_),
    .Q(\hdisplay[1] ));
 sg13g2_dfrbp_1 _3282_ (.CLK(net363),
    .RESET_B(net116),
    .D(_0137_),
    .Q_N(_1509_),
    .Q(\hdisplay[2] ));
 sg13g2_dfrbp_1 _3283_ (.CLK(net366),
    .RESET_B(net108),
    .D(_0138_),
    .Q_N(_1508_),
    .Q(\hdisplay[3] ));
 sg13g2_dfrbp_1 _3284_ (.CLK(net366),
    .RESET_B(net84),
    .D(_0139_),
    .Q_N(_1507_),
    .Q(\hdisplay[4] ));
 sg13g2_dfrbp_1 _3285_ (.CLK(net373),
    .RESET_B(net68),
    .D(_0140_),
    .Q_N(_1506_),
    .Q(\hdisplay[5] ));
 sg13g2_dfrbp_1 _3286_ (.CLK(net370),
    .RESET_B(net129),
    .D(_0141_),
    .Q_N(_1505_),
    .Q(\hdisplay[6] ));
 sg13g2_dfrbp_1 _3287_ (.CLK(net371),
    .RESET_B(net112),
    .D(_0142_),
    .Q_N(_1504_),
    .Q(\hdisplay[7] ));
 sg13g2_dfrbp_1 _3288_ (.CLK(net372),
    .RESET_B(net76),
    .D(_0143_),
    .Q_N(_1503_),
    .Q(\hdisplay[8] ));
 sg13g2_dfrbp_1 _3289_ (.CLK(net372),
    .RESET_B(net120),
    .D(_0144_),
    .Q_N(_1502_),
    .Q(\hdisplay[9] ));
 sg13g2_dfrbp_1 _3290_ (.CLK(net372),
    .RESET_B(net60),
    .D(_0145_),
    .Q_N(_1501_),
    .Q(\hdisplay[10] ));
 sg13g2_tiehi _3254__33 (.L_HI(net33));
 sg13g2_tiehi _3217__34 (.L_HI(net34));
 sg13g2_tiehi _3279__35 (.L_HI(net35));
 sg13g2_tiehi _3216__36 (.L_HI(net36));
 sg13g2_tiehi _3253__37 (.L_HI(net37));
 sg13g2_tiehi _3215__38 (.L_HI(net38));
 sg13g2_tiehi _3278__39 (.L_HI(net39));
 sg13g2_tiehi _3214__40 (.L_HI(net40));
 sg13g2_tiehi _3259__41 (.L_HI(net41));
 sg13g2_tiehi _3252__42 (.L_HI(net42));
 sg13g2_tiehi _3213__43 (.L_HI(net43));
 sg13g2_tiehi _3277__44 (.L_HI(net44));
 sg13g2_tiehi _3212__45 (.L_HI(net45));
 sg13g2_tiehi _3251__46 (.L_HI(net46));
 sg13g2_tiehi _3211__47 (.L_HI(net47));
 sg13g2_tiehi _3276__48 (.L_HI(net48));
 sg13g2_tiehi _3210__49 (.L_HI(net49));
 sg13g2_tiehi _3250__50 (.L_HI(net50));
 sg13g2_tiehi _3209__51 (.L_HI(net51));
 sg13g2_tiehi _3275__52 (.L_HI(net52));
 sg13g2_tiehi _3208__53 (.L_HI(net53));
 sg13g2_tiehi _3249__54 (.L_HI(net54));
 sg13g2_tiehi _3207__55 (.L_HI(net55));
 sg13g2_tiehi _3274__56 (.L_HI(net56));
 sg13g2_tiehi _3206__57 (.L_HI(net57));
 sg13g2_tiehi _3248__58 (.L_HI(net58));
 sg13g2_tiehi _3205__59 (.L_HI(net59));
 sg13g2_tiehi _3290__60 (.L_HI(net60));
 sg13g2_tiehi _3204__61 (.L_HI(net61));
 sg13g2_tiehi _3247__62 (.L_HI(net62));
 sg13g2_tiehi _3203__63 (.L_HI(net63));
 sg13g2_tiehi _3273__64 (.L_HI(net64));
 sg13g2_tiehi _3202__65 (.L_HI(net65));
 sg13g2_tiehi _3246__66 (.L_HI(net66));
 sg13g2_tiehi _3201__67 (.L_HI(net67));
 sg13g2_tiehi _3285__68 (.L_HI(net68));
 sg13g2_tiehi _3200__69 (.L_HI(net69));
 sg13g2_tiehi _3245__70 (.L_HI(net70));
 sg13g2_tiehi _3199__71 (.L_HI(net71));
 sg13g2_tiehi _3271__72 (.L_HI(net72));
 sg13g2_tiehi _3198__73 (.L_HI(net73));
 sg13g2_tiehi _3244__74 (.L_HI(net74));
 sg13g2_tiehi _3197__75 (.L_HI(net75));
 sg13g2_tiehi _3288__76 (.L_HI(net76));
 sg13g2_tiehi _3196__77 (.L_HI(net77));
 sg13g2_tiehi _3243__78 (.L_HI(net78));
 sg13g2_tiehi _3195__79 (.L_HI(net79));
 sg13g2_tiehi _3270__80 (.L_HI(net80));
 sg13g2_tiehi _3194__81 (.L_HI(net81));
 sg13g2_tiehi _3242__82 (.L_HI(net82));
 sg13g2_tiehi _3193__83 (.L_HI(net83));
 sg13g2_tiehi _3284__84 (.L_HI(net84));
 sg13g2_tiehi _3192__85 (.L_HI(net85));
 sg13g2_tiehi _3241__86 (.L_HI(net86));
 sg13g2_tiehi _3191__87 (.L_HI(net87));
 sg13g2_tiehi _3269__88 (.L_HI(net88));
 sg13g2_tiehi _3190__89 (.L_HI(net89));
 sg13g2_tiehi _3240__90 (.L_HI(net90));
 sg13g2_tiehi _3189__91 (.L_HI(net91));
 sg13g2_tiehi _3272__92 (.L_HI(net92));
 sg13g2_tiehi _3188__93 (.L_HI(net93));
 sg13g2_tiehi _3187__94 (.L_HI(net94));
 sg13g2_tiehi _3186__95 (.L_HI(net95));
 sg13g2_tiehi _3185__96 (.L_HI(net96));
 sg13g2_tiehi _3184__97 (.L_HI(net97));
 sg13g2_tiehi _3183__98 (.L_HI(net98));
 sg13g2_tiehi _3182__99 (.L_HI(net99));
 sg13g2_tiehi _3181__100 (.L_HI(net100));
 sg13g2_tiehi _3180__101 (.L_HI(net101));
 sg13g2_tiehi _3179__102 (.L_HI(net102));
 sg13g2_tiehi _3178__103 (.L_HI(net103));
 sg13g2_tiehi _3177__104 (.L_HI(net104));
 sg13g2_tiehi _3239__105 (.L_HI(net105));
 sg13g2_tiehi _3268__106 (.L_HI(net106));
 sg13g2_tiehi _3238__107 (.L_HI(net107));
 sg13g2_tiehi _3283__108 (.L_HI(net108));
 sg13g2_tiehi _3237__109 (.L_HI(net109));
 sg13g2_tiehi _3267__110 (.L_HI(net110));
 sg13g2_tiehi _3236__111 (.L_HI(net111));
 sg13g2_tiehi _3287__112 (.L_HI(net112));
 sg13g2_tiehi _3235__113 (.L_HI(net113));
 sg13g2_tiehi _3266__114 (.L_HI(net114));
 sg13g2_tiehi _3234__115 (.L_HI(net115));
 sg13g2_tiehi _3282__116 (.L_HI(net116));
 sg13g2_tiehi _3233__117 (.L_HI(net117));
 sg13g2_tiehi _3265__118 (.L_HI(net118));
 sg13g2_tiehi _3232__119 (.L_HI(net119));
 sg13g2_tiehi _3289__120 (.L_HI(net120));
 sg13g2_tiehi _3231__121 (.L_HI(net121));
 sg13g2_tiehi _3264__122 (.L_HI(net122));
 sg13g2_tiehi _3230__123 (.L_HI(net123));
 sg13g2_tiehi _3229__124 (.L_HI(net124));
 sg13g2_tiehi _3281__125 (.L_HI(net125));
 sg13g2_tiehi _3228__126 (.L_HI(net126));
 sg13g2_tiehi _3263__127 (.L_HI(net127));
 sg13g2_tiehi _3227__128 (.L_HI(net128));
 sg13g2_tiehi _3286__129 (.L_HI(net129));
 sg13g2_tiehi _3226__130 (.L_HI(net130));
 sg13g2_tiehi _3262__131 (.L_HI(net131));
 sg13g2_tiehi _3225__132 (.L_HI(net132));
 sg13g2_tiehi _3280__133 (.L_HI(net133));
 sg13g2_tiehi _3224__134 (.L_HI(net134));
 sg13g2_tiehi _3261__135 (.L_HI(net135));
 sg13g2_tiehi _3223__136 (.L_HI(net136));
 sg13g2_tiehi _3260__137 (.L_HI(net137));
 sg13g2_tiehi _3222__138 (.L_HI(net138));
 sg13g2_tiehi _3258__139 (.L_HI(net139));
 sg13g2_tiehi _3221__140 (.L_HI(net140));
 sg13g2_tiehi _3257__141 (.L_HI(net141));
 sg13g2_tiehi _3220__142 (.L_HI(net142));
 sg13g2_tiehi _3176__143 (.L_HI(net143));
 sg13g2_tiehi _3256__144 (.L_HI(net144));
 sg13g2_tiehi _3219__145 (.L_HI(net145));
 sg13g2_tiehi _3255__146 (.L_HI(net146));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_21 (.L_LO(net21));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_22 (.L_LO(net22));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_23 (.L_LO(net23));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_24 (.L_LO(net24));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_25 (.L_LO(net25));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_26 (.L_LO(net26));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_27 (.L_LO(net27));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_28 (.L_LO(net28));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_29 (.L_LO(net29));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_30 (.L_LO(net30));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_31 (.L_LO(net31));
 sg13g2_tiehi _3218__32 (.L_HI(net32));
 sg13g2_buf_4 _3422_ (.X(uo_out[3]),
    .A(\hvsync_gen.vsync ));
 sg13g2_buf_1 _3423_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_0714_));
 sg13g2_buf_1 fanout286 (.A(_0714_),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(net288));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(_0463_));
 sg13g2_buf_2 fanout289 (.A(_0987_),
    .X(net289));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(_0569_));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_0511_));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(_0497_));
 sg13g2_buf_2 fanout293 (.A(_0967_),
    .X(net293));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(_0965_));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(_0847_));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(_0777_));
 sg13g2_buf_1 fanout297 (.A(_0777_),
    .X(net297));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(_0579_));
 sg13g2_buf_4 fanout299 (.X(net299),
    .A(_0496_));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(_0495_));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(_0495_));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(_0494_));
 sg13g2_buf_2 fanout303 (.A(_0590_),
    .X(net303));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(_0540_));
 sg13g2_buf_2 fanout305 (.A(_0540_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_0939_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_0747_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_0744_),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(_0568_));
 sg13g2_buf_4 fanout310 (.X(net310),
    .A(_0556_));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_0510_));
 sg13g2_buf_1 fanout312 (.A(_0510_),
    .X(net312));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(_0487_));
 sg13g2_buf_2 fanout314 (.A(_0487_),
    .X(net314));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(_0484_));
 sg13g2_buf_2 fanout316 (.A(_0931_),
    .X(net316));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_0844_));
 sg13g2_buf_2 fanout318 (.A(\hvsync_gen.vpos[9] ),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net160),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(net158),
    .X(net321));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_0008_));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_1 fanout324 (.A(net325),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(\hvsync_gen.vpos[6] ),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(\hvsync_gen.vpos[5] ));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(net329));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(net157));
 sg13g2_buf_2 fanout330 (.A(net332),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(net332),
    .X(net331));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(\hvsync_gen.vpos[3] ));
 sg13g2_buf_2 fanout333 (.A(net162),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(\hvsync_gen.vpos[2] ),
    .X(net334));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(net168));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(\hvsync_gen.vpos[0] ));
 sg13g2_buf_2 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_1 fanout338 (.A(_0027_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(\pat.pattern[3] ),
    .X(net339));
 sg13g2_buf_1 fanout340 (.A(\pat.pattern[3] ),
    .X(net340));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(\pat.pattern[2] ));
 sg13g2_buf_1 fanout342 (.A(\pat.pattern[2] ),
    .X(net342));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(\hpos[9] ));
 sg13g2_buf_1 fanout344 (.A(\hpos[9] ),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(net159),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(\hpos[8] ),
    .X(net346));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(net165));
 sg13g2_buf_2 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(\hpos[6] ));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net352));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(net352));
 sg13g2_buf_2 fanout352 (.A(\hpos[5] ),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(net354),
    .X(net353));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(\hpos[4] ));
 sg13g2_buf_2 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(net173));
 sg13g2_buf_2 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(\hpos[2] ),
    .X(net358));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(\hpos[1] ));
 sg13g2_buf_2 fanout360 (.A(net361),
    .X(net360));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(net362));
 sg13g2_buf_2 fanout362 (.A(net374),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_1 fanout364 (.A(net365),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(net367),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(net367));
 sg13g2_buf_2 fanout367 (.A(net374),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(net374),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(net373),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(net372),
    .X(net371));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(net373));
 sg13g2_buf_2 fanout373 (.A(net374),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(ui_in[7]),
    .X(net374));
 sg13g2_buf_4 fanout375 (.X(net375),
    .A(ui_in[3]));
 sg13g2_buf_1 fanout376 (.A(ui_in[3]),
    .X(net376));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(net4));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_4 input9 (.X(net9),
    .A(uio_in[1]));
 sg13g2_buf_2 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[6]),
    .X(net14));
 sg13g2_buf_2 input15 (.A(uio_in[7]),
    .X(net15));
 sg13g2_tielo tt_um_rebeccargb_vga_timing_experiments_16 (.L_LO(net16));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0032_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0031_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0117_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.vpos[11] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0128_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold6 (.A(\hpos[11] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0481_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold8 (.A(\hvsync_gen.vpos[10] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold9 (.A(\hpos[0] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0882_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold11 (.A(\hvsync_gen.vpos[4] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold12 (.A(\hvsync_gen.vpos[7] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hpos[8] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold14 (.A(\hvsync_gen.vpos[8] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0018_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold16 (.A(\hvsync_gen.vpos[2] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0022_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0477_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hpos[7] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0010_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0126_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hvsync_gen.vpos[1] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0024_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0004_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold25 (.A(\hpos[10] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0006_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold27 (.A(\hpos[3] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0014_),
    .X(net174));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_4 FILLER_0_91 ();
 sg13g2_fill_2 FILLER_0_95 ();
 sg13g2_fill_2 FILLER_0_102 ();
 sg13g2_fill_1 FILLER_0_104 ();
 sg13g2_decap_8 FILLER_0_113 ();
 sg13g2_decap_8 FILLER_0_120 ();
 sg13g2_decap_8 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_fill_2 FILLER_0_141 ();
 sg13g2_fill_2 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_4 FILLER_0_186 ();
 sg13g2_fill_2 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_197 ();
 sg13g2_fill_2 FILLER_0_204 ();
 sg13g2_fill_2 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_fill_1 FILLER_0_239 ();
 sg13g2_fill_2 FILLER_0_256 ();
 sg13g2_fill_1 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_fill_1 FILLER_0_271 ();
 sg13g2_fill_1 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_fill_1 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_4 FILLER_0_327 ();
 sg13g2_decap_4 FILLER_0_335 ();
 sg13g2_fill_2 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_4 FILLER_1_49 ();
 sg13g2_fill_2 FILLER_1_53 ();
 sg13g2_decap_8 FILLER_1_60 ();
 sg13g2_fill_2 FILLER_1_67 ();
 sg13g2_fill_1 FILLER_1_69 ();
 sg13g2_decap_8 FILLER_1_78 ();
 sg13g2_decap_8 FILLER_1_85 ();
 sg13g2_fill_2 FILLER_1_92 ();
 sg13g2_decap_8 FILLER_1_120 ();
 sg13g2_decap_8 FILLER_1_127 ();
 sg13g2_fill_1 FILLER_1_264 ();
 sg13g2_fill_1 FILLER_1_295 ();
 sg13g2_decap_8 FILLER_1_362 ();
 sg13g2_decap_8 FILLER_1_369 ();
 sg13g2_decap_8 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_390 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_4 FILLER_1_404 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_fill_1 FILLER_2_35 ();
 sg13g2_fill_2 FILLER_2_92 ();
 sg13g2_fill_1 FILLER_2_94 ();
 sg13g2_decap_4 FILLER_2_100 ();
 sg13g2_fill_2 FILLER_2_104 ();
 sg13g2_fill_2 FILLER_2_111 ();
 sg13g2_fill_2 FILLER_2_121 ();
 sg13g2_decap_4 FILLER_2_162 ();
 sg13g2_fill_2 FILLER_2_166 ();
 sg13g2_fill_1 FILLER_2_181 ();
 sg13g2_decap_8 FILLER_2_187 ();
 sg13g2_fill_2 FILLER_2_194 ();
 sg13g2_decap_4 FILLER_2_200 ();
 sg13g2_fill_1 FILLER_2_204 ();
 sg13g2_decap_4 FILLER_2_212 ();
 sg13g2_fill_2 FILLER_2_216 ();
 sg13g2_decap_8 FILLER_2_227 ();
 sg13g2_fill_2 FILLER_2_234 ();
 sg13g2_fill_1 FILLER_2_266 ();
 sg13g2_fill_1 FILLER_2_288 ();
 sg13g2_decap_8 FILLER_2_297 ();
 sg13g2_fill_1 FILLER_2_312 ();
 sg13g2_fill_1 FILLER_2_317 ();
 sg13g2_fill_2 FILLER_2_323 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_fill_2 FILLER_2_336 ();
 sg13g2_fill_1 FILLER_2_338 ();
 sg13g2_fill_2 FILLER_2_348 ();
 sg13g2_fill_1 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_fill_2 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_fill_2 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_27 ();
 sg13g2_decap_4 FILLER_3_51 ();
 sg13g2_fill_1 FILLER_3_55 ();
 sg13g2_decap_4 FILLER_3_70 ();
 sg13g2_fill_2 FILLER_3_74 ();
 sg13g2_fill_1 FILLER_3_83 ();
 sg13g2_fill_2 FILLER_3_100 ();
 sg13g2_fill_2 FILLER_3_138 ();
 sg13g2_fill_1 FILLER_3_140 ();
 sg13g2_decap_4 FILLER_3_162 ();
 sg13g2_fill_2 FILLER_3_166 ();
 sg13g2_fill_2 FILLER_3_173 ();
 sg13g2_fill_2 FILLER_3_216 ();
 sg13g2_fill_2 FILLER_3_226 ();
 sg13g2_fill_2 FILLER_3_232 ();
 sg13g2_fill_1 FILLER_3_234 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_fill_2 FILLER_3_266 ();
 sg13g2_fill_1 FILLER_3_304 ();
 sg13g2_fill_2 FILLER_3_344 ();
 sg13g2_fill_1 FILLER_3_346 ();
 sg13g2_decap_4 FILLER_3_386 ();
 sg13g2_decap_4 FILLER_3_394 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_11 ();
 sg13g2_fill_2 FILLER_4_38 ();
 sg13g2_fill_2 FILLER_4_66 ();
 sg13g2_fill_1 FILLER_4_84 ();
 sg13g2_fill_1 FILLER_4_107 ();
 sg13g2_fill_1 FILLER_4_115 ();
 sg13g2_decap_4 FILLER_4_132 ();
 sg13g2_fill_2 FILLER_4_149 ();
 sg13g2_fill_2 FILLER_4_159 ();
 sg13g2_fill_2 FILLER_4_174 ();
 sg13g2_fill_1 FILLER_4_176 ();
 sg13g2_fill_2 FILLER_4_244 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_fill_2 FILLER_4_274 ();
 sg13g2_fill_1 FILLER_4_276 ();
 sg13g2_decap_4 FILLER_4_298 ();
 sg13g2_fill_2 FILLER_4_314 ();
 sg13g2_decap_4 FILLER_4_356 ();
 sg13g2_fill_1 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_fill_1 FILLER_4_378 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_16 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_4 FILLER_5_28 ();
 sg13g2_fill_1 FILLER_5_32 ();
 sg13g2_fill_1 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_62 ();
 sg13g2_fill_1 FILLER_5_69 ();
 sg13g2_fill_2 FILLER_5_82 ();
 sg13g2_decap_4 FILLER_5_97 ();
 sg13g2_fill_1 FILLER_5_101 ();
 sg13g2_fill_2 FILLER_5_135 ();
 sg13g2_decap_4 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_154 ();
 sg13g2_fill_2 FILLER_5_159 ();
 sg13g2_decap_4 FILLER_5_169 ();
 sg13g2_decap_4 FILLER_5_185 ();
 sg13g2_fill_2 FILLER_5_194 ();
 sg13g2_fill_1 FILLER_5_196 ();
 sg13g2_fill_2 FILLER_5_204 ();
 sg13g2_fill_2 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_fill_2 FILLER_5_230 ();
 sg13g2_fill_1 FILLER_5_232 ();
 sg13g2_fill_1 FILLER_5_240 ();
 sg13g2_decap_4 FILLER_5_249 ();
 sg13g2_fill_2 FILLER_5_253 ();
 sg13g2_decap_4 FILLER_5_272 ();
 sg13g2_decap_4 FILLER_5_332 ();
 sg13g2_fill_1 FILLER_5_336 ();
 sg13g2_fill_1 FILLER_5_350 ();
 sg13g2_fill_2 FILLER_5_375 ();
 sg13g2_fill_2 FILLER_5_400 ();
 sg13g2_fill_1 FILLER_5_402 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_fill_2 FILLER_6_32 ();
 sg13g2_fill_1 FILLER_6_34 ();
 sg13g2_decap_4 FILLER_6_61 ();
 sg13g2_fill_1 FILLER_6_65 ();
 sg13g2_decap_4 FILLER_6_86 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_fill_1 FILLER_6_109 ();
 sg13g2_fill_2 FILLER_6_118 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_decap_4 FILLER_6_158 ();
 sg13g2_fill_2 FILLER_6_162 ();
 sg13g2_fill_1 FILLER_6_181 ();
 sg13g2_decap_8 FILLER_6_187 ();
 sg13g2_decap_8 FILLER_6_194 ();
 sg13g2_decap_4 FILLER_6_201 ();
 sg13g2_fill_2 FILLER_6_213 ();
 sg13g2_fill_2 FILLER_6_227 ();
 sg13g2_decap_8 FILLER_6_258 ();
 sg13g2_fill_1 FILLER_6_275 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_fill_2 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_293 ();
 sg13g2_decap_4 FILLER_6_311 ();
 sg13g2_fill_2 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_4 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_fill_1 FILLER_6_366 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_4 FILLER_7_32 ();
 sg13g2_decap_4 FILLER_7_50 ();
 sg13g2_decap_4 FILLER_7_59 ();
 sg13g2_fill_1 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_80 ();
 sg13g2_fill_2 FILLER_7_87 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_fill_2 FILLER_7_136 ();
 sg13g2_fill_1 FILLER_7_138 ();
 sg13g2_fill_2 FILLER_7_143 ();
 sg13g2_decap_8 FILLER_7_150 ();
 sg13g2_decap_4 FILLER_7_209 ();
 sg13g2_decap_4 FILLER_7_251 ();
 sg13g2_fill_2 FILLER_7_271 ();
 sg13g2_fill_2 FILLER_7_294 ();
 sg13g2_fill_1 FILLER_7_296 ();
 sg13g2_decap_8 FILLER_7_317 ();
 sg13g2_fill_1 FILLER_7_324 ();
 sg13g2_decap_4 FILLER_7_338 ();
 sg13g2_fill_1 FILLER_7_342 ();
 sg13g2_fill_2 FILLER_7_355 ();
 sg13g2_fill_1 FILLER_7_357 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_14 ();
 sg13g2_fill_1 FILLER_8_16 ();
 sg13g2_fill_1 FILLER_8_69 ();
 sg13g2_decap_4 FILLER_8_93 ();
 sg13g2_fill_2 FILLER_8_122 ();
 sg13g2_fill_1 FILLER_8_124 ();
 sg13g2_fill_1 FILLER_8_135 ();
 sg13g2_fill_2 FILLER_8_145 ();
 sg13g2_fill_2 FILLER_8_162 ();
 sg13g2_fill_1 FILLER_8_164 ();
 sg13g2_fill_1 FILLER_8_178 ();
 sg13g2_fill_2 FILLER_8_192 ();
 sg13g2_decap_4 FILLER_8_198 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_fill_2 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_fill_2 FILLER_8_266 ();
 sg13g2_fill_1 FILLER_8_268 ();
 sg13g2_fill_2 FILLER_8_290 ();
 sg13g2_fill_1 FILLER_8_292 ();
 sg13g2_decap_4 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_334 ();
 sg13g2_fill_2 FILLER_8_341 ();
 sg13g2_decap_4 FILLER_8_355 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_fill_1 FILLER_8_394 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_fill_2 FILLER_9_32 ();
 sg13g2_fill_1 FILLER_9_34 ();
 sg13g2_decap_4 FILLER_9_48 ();
 sg13g2_fill_1 FILLER_9_52 ();
 sg13g2_fill_1 FILLER_9_57 ();
 sg13g2_fill_2 FILLER_9_62 ();
 sg13g2_fill_2 FILLER_9_86 ();
 sg13g2_fill_2 FILLER_9_108 ();
 sg13g2_decap_4 FILLER_9_118 ();
 sg13g2_fill_2 FILLER_9_122 ();
 sg13g2_decap_4 FILLER_9_170 ();
 sg13g2_fill_2 FILLER_9_179 ();
 sg13g2_decap_4 FILLER_9_204 ();
 sg13g2_fill_1 FILLER_9_208 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_fill_2 FILLER_9_227 ();
 sg13g2_fill_2 FILLER_9_246 ();
 sg13g2_fill_1 FILLER_9_248 ();
 sg13g2_fill_1 FILLER_9_254 ();
 sg13g2_fill_2 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_263 ();
 sg13g2_fill_2 FILLER_9_274 ();
 sg13g2_fill_1 FILLER_9_276 ();
 sg13g2_fill_2 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_302 ();
 sg13g2_fill_1 FILLER_9_319 ();
 sg13g2_fill_2 FILLER_9_362 ();
 sg13g2_fill_2 FILLER_9_368 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_32 ();
 sg13g2_fill_1 FILLER_10_34 ();
 sg13g2_decap_4 FILLER_10_49 ();
 sg13g2_fill_1 FILLER_10_53 ();
 sg13g2_fill_2 FILLER_10_72 ();
 sg13g2_fill_2 FILLER_10_92 ();
 sg13g2_fill_1 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_149 ();
 sg13g2_fill_2 FILLER_10_156 ();
 sg13g2_fill_1 FILLER_10_158 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_2 FILLER_10_200 ();
 sg13g2_decap_4 FILLER_10_207 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_decap_4 FILLER_10_265 ();
 sg13g2_fill_1 FILLER_10_269 ();
 sg13g2_fill_2 FILLER_10_289 ();
 sg13g2_fill_1 FILLER_10_291 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_fill_1 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_fill_1 FILLER_10_331 ();
 sg13g2_decap_4 FILLER_10_336 ();
 sg13g2_decap_4 FILLER_10_345 ();
 sg13g2_fill_1 FILLER_10_349 ();
 sg13g2_fill_2 FILLER_10_368 ();
 sg13g2_fill_1 FILLER_10_370 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_11 ();
 sg13g2_fill_1 FILLER_11_20 ();
 sg13g2_fill_2 FILLER_11_96 ();
 sg13g2_fill_2 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_fill_2 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_fill_1 FILLER_11_169 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_decap_8 FILLER_11_181 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_fill_2 FILLER_11_225 ();
 sg13g2_fill_1 FILLER_11_227 ();
 sg13g2_decap_4 FILLER_11_292 ();
 sg13g2_fill_1 FILLER_11_354 ();
 sg13g2_fill_1 FILLER_11_393 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_39 ();
 sg13g2_fill_1 FILLER_12_43 ();
 sg13g2_decap_8 FILLER_12_48 ();
 sg13g2_fill_2 FILLER_12_94 ();
 sg13g2_fill_1 FILLER_12_96 ();
 sg13g2_fill_1 FILLER_12_139 ();
 sg13g2_fill_2 FILLER_12_150 ();
 sg13g2_fill_2 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_4 FILLER_12_213 ();
 sg13g2_fill_1 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_251 ();
 sg13g2_fill_1 FILLER_12_262 ();
 sg13g2_fill_1 FILLER_12_292 ();
 sg13g2_decap_4 FILLER_12_313 ();
 sg13g2_fill_2 FILLER_12_317 ();
 sg13g2_decap_4 FILLER_12_325 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_335 ();
 sg13g2_fill_2 FILLER_12_371 ();
 sg13g2_fill_2 FILLER_12_378 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_37 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_100 ();
 sg13g2_fill_1 FILLER_13_109 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_164 ();
 sg13g2_fill_2 FILLER_13_174 ();
 sg13g2_fill_2 FILLER_13_200 ();
 sg13g2_decap_4 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_fill_1 FILLER_13_256 ();
 sg13g2_fill_2 FILLER_13_265 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_fill_2 FILLER_13_293 ();
 sg13g2_fill_2 FILLER_13_316 ();
 sg13g2_fill_1 FILLER_13_318 ();
 sg13g2_decap_4 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_45 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_fill_2 FILLER_14_65 ();
 sg13g2_fill_1 FILLER_14_67 ();
 sg13g2_fill_2 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_14_101 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_fill_1 FILLER_14_228 ();
 sg13g2_fill_2 FILLER_14_241 ();
 sg13g2_fill_1 FILLER_14_243 ();
 sg13g2_fill_2 FILLER_14_250 ();
 sg13g2_fill_1 FILLER_14_252 ();
 sg13g2_decap_4 FILLER_14_262 ();
 sg13g2_decap_4 FILLER_14_274 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_310 ();
 sg13g2_fill_1 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_16 ();
 sg13g2_decap_4 FILLER_15_25 ();
 sg13g2_fill_2 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_fill_2 FILLER_15_111 ();
 sg13g2_fill_1 FILLER_15_113 ();
 sg13g2_fill_1 FILLER_15_133 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_fill_2 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_145 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_fill_2 FILLER_15_158 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_196 ();
 sg13g2_decap_4 FILLER_15_219 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_fill_2 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_2 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_decap_8 FILLER_16_45 ();
 sg13g2_decap_4 FILLER_16_72 ();
 sg13g2_fill_2 FILLER_16_76 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_107 ();
 sg13g2_fill_2 FILLER_16_122 ();
 sg13g2_fill_1 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_131 ();
 sg13g2_decap_4 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_185 ();
 sg13g2_fill_2 FILLER_16_195 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_fill_2 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_259 ();
 sg13g2_decap_4 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_decap_4 FILLER_16_290 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_2 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_371 ();
 sg13g2_fill_1 FILLER_16_373 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_15 ();
 sg13g2_fill_2 FILLER_17_22 ();
 sg13g2_fill_2 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_54 ();
 sg13g2_fill_1 FILLER_17_66 ();
 sg13g2_decap_4 FILLER_17_79 ();
 sg13g2_fill_1 FILLER_17_83 ();
 sg13g2_fill_2 FILLER_17_96 ();
 sg13g2_fill_1 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_125 ();
 sg13g2_fill_2 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_143 ();
 sg13g2_decap_4 FILLER_17_152 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_fill_2 FILLER_17_199 ();
 sg13g2_fill_1 FILLER_17_213 ();
 sg13g2_decap_4 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_260 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_decap_4 FILLER_17_288 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_353 ();
 sg13g2_fill_2 FILLER_17_381 ();
 sg13g2_fill_2 FILLER_18_31 ();
 sg13g2_fill_2 FILLER_18_40 ();
 sg13g2_fill_1 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_109 ();
 sg13g2_fill_2 FILLER_18_116 ();
 sg13g2_fill_1 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_197 ();
 sg13g2_fill_2 FILLER_18_211 ();
 sg13g2_fill_1 FILLER_18_213 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_fill_2 FILLER_18_261 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_2 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_fill_2 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_365 ();
 sg13g2_decap_4 FILLER_18_370 ();
 sg13g2_fill_2 FILLER_18_378 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_41 ();
 sg13g2_fill_1 FILLER_19_45 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_decap_4 FILLER_19_87 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_132 ();
 sg13g2_fill_2 FILLER_19_159 ();
 sg13g2_fill_1 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_170 ();
 sg13g2_decap_4 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_220 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_decap_4 FILLER_19_244 ();
 sg13g2_fill_2 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_271 ();
 sg13g2_decap_4 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_4 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_293 ();
 sg13g2_decap_4 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_decap_4 FILLER_19_355 ();
 sg13g2_fill_2 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_2 FILLER_20_31 ();
 sg13g2_fill_1 FILLER_20_47 ();
 sg13g2_decap_8 FILLER_20_57 ();
 sg13g2_fill_1 FILLER_20_64 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_fill_1 FILLER_20_138 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_247 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_decap_4 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_fill_2 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_373 ();
 sg13g2_fill_2 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_12 ();
 sg13g2_fill_1 FILLER_21_34 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_fill_2 FILLER_21_60 ();
 sg13g2_fill_1 FILLER_21_62 ();
 sg13g2_fill_1 FILLER_21_80 ();
 sg13g2_fill_2 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_93 ();
 sg13g2_fill_1 FILLER_21_99 ();
 sg13g2_fill_2 FILLER_21_109 ();
 sg13g2_decap_4 FILLER_21_143 ();
 sg13g2_fill_2 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_fill_1 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_250 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_17 ();
 sg13g2_fill_1 FILLER_22_19 ();
 sg13g2_fill_1 FILLER_22_41 ();
 sg13g2_decap_4 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_54 ();
 sg13g2_fill_2 FILLER_22_60 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_decap_4 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_fill_2 FILLER_22_191 ();
 sg13g2_decap_4 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_202 ();
 sg13g2_fill_2 FILLER_22_217 ();
 sg13g2_decap_4 FILLER_22_233 ();
 sg13g2_fill_2 FILLER_22_237 ();
 sg13g2_decap_8 FILLER_22_243 ();
 sg13g2_decap_4 FILLER_22_250 ();
 sg13g2_fill_2 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_decap_4 FILLER_22_299 ();
 sg13g2_fill_2 FILLER_22_303 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_349 ();
 sg13g2_fill_2 FILLER_22_364 ();
 sg13g2_fill_2 FILLER_23_31 ();
 sg13g2_fill_1 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_80 ();
 sg13g2_fill_2 FILLER_23_87 ();
 sg13g2_fill_1 FILLER_23_89 ();
 sg13g2_fill_2 FILLER_23_100 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_121 ();
 sg13g2_fill_1 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_decap_8 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_decap_4 FILLER_23_223 ();
 sg13g2_fill_2 FILLER_23_253 ();
 sg13g2_fill_2 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_291 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_2 FILLER_23_397 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_20 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_fill_2 FILLER_24_43 ();
 sg13g2_fill_1 FILLER_24_45 ();
 sg13g2_fill_2 FILLER_24_51 ();
 sg13g2_fill_1 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_127 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_fill_2 FILLER_24_150 ();
 sg13g2_fill_1 FILLER_24_152 ();
 sg13g2_fill_2 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_2 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_4 FILLER_24_271 ();
 sg13g2_fill_1 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_fill_1 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_25_34 ();
 sg13g2_fill_1 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_77 ();
 sg13g2_fill_2 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_90 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_183 ();
 sg13g2_decap_4 FILLER_25_205 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_fill_2 FILLER_25_226 ();
 sg13g2_fill_1 FILLER_25_228 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_279 ();
 sg13g2_fill_2 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_fill_2 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_fill_2 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_343 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_fill_1 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_15 ();
 sg13g2_fill_1 FILLER_26_17 ();
 sg13g2_fill_2 FILLER_26_22 ();
 sg13g2_fill_1 FILLER_26_24 ();
 sg13g2_decap_4 FILLER_26_46 ();
 sg13g2_fill_1 FILLER_26_50 ();
 sg13g2_decap_8 FILLER_26_101 ();
 sg13g2_decap_4 FILLER_26_108 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_124 ();
 sg13g2_decap_4 FILLER_26_128 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_230 ();
 sg13g2_decap_4 FILLER_26_238 ();
 sg13g2_fill_2 FILLER_26_242 ();
 sg13g2_decap_4 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_fill_2 FILLER_26_327 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_2 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_392 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_33 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_decap_8 FILLER_27_50 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_85 ();
 sg13g2_decap_8 FILLER_27_136 ();
 sg13g2_decap_8 FILLER_27_143 ();
 sg13g2_decap_8 FILLER_27_181 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_decap_4 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_230 ();
 sg13g2_fill_2 FILLER_27_245 ();
 sg13g2_fill_1 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_255 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_decap_4 FILLER_27_274 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_2 FILLER_27_308 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_33 ();
 sg13g2_fill_1 FILLER_28_37 ();
 sg13g2_fill_2 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_66 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_decap_8 FILLER_28_87 ();
 sg13g2_decap_4 FILLER_28_94 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_decap_4 FILLER_28_162 ();
 sg13g2_decap_4 FILLER_28_170 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_229 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_decap_4 FILLER_28_237 ();
 sg13g2_decap_4 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_334 ();
 sg13g2_fill_2 FILLER_28_341 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_4 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_28_382 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_39 ();
 sg13g2_fill_1 FILLER_29_53 ();
 sg13g2_fill_1 FILLER_29_82 ();
 sg13g2_decap_8 FILLER_29_96 ();
 sg13g2_fill_1 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_134 ();
 sg13g2_decap_8 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_decap_4 FILLER_29_198 ();
 sg13g2_decap_4 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_decap_4 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_385 ();
 sg13g2_fill_2 FILLER_29_394 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_27 ();
 sg13g2_fill_2 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_fill_2 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_1 FILLER_30_94 ();
 sg13g2_decap_4 FILLER_30_190 ();
 sg13g2_fill_2 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_336 ();
 sg13g2_decap_4 FILLER_30_345 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_11 ();
 sg13g2_decap_4 FILLER_31_20 ();
 sg13g2_fill_2 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_44 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_95 ();
 sg13g2_fill_1 FILLER_31_97 ();
 sg13g2_decap_4 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_decap_4 FILLER_31_180 ();
 sg13g2_fill_1 FILLER_31_184 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_decap_4 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_242 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_fill_2 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_258 ();
 sg13g2_decap_4 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_269 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_decap_4 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_4 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_38 ();
 sg13g2_decap_4 FILLER_32_69 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_95 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_decap_4 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_242 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_296 ();
 sg13g2_decap_4 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_4 FILLER_32_368 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_11 ();
 sg13g2_fill_1 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_71 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_fill_2 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_208 ();
 sg13g2_decap_4 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_225 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_295 ();
 sg13g2_decap_4 FILLER_33_328 ();
 sg13g2_decap_4 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_391 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_fill_2 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_69 ();
 sg13g2_fill_2 FILLER_34_101 ();
 sg13g2_decap_8 FILLER_34_120 ();
 sg13g2_decap_8 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_134 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_decap_8 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_171 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_220 ();
 sg13g2_decap_4 FILLER_34_227 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_decap_4 FILLER_34_252 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_262 ();
 sg13g2_fill_2 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_decap_4 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_1 FILLER_35_113 ();
 sg13g2_fill_2 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_203 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_248 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_288 ();
 sg13g2_decap_4 FILLER_35_310 ();
 sg13g2_decap_4 FILLER_35_321 ();
 sg13g2_decap_4 FILLER_35_336 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_fill_2 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_30 ();
 sg13g2_fill_2 FILLER_36_50 ();
 sg13g2_fill_1 FILLER_36_52 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_fill_2 FILLER_36_96 ();
 sg13g2_fill_1 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_fill_2 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_139 ();
 sg13g2_decap_4 FILLER_36_145 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_decap_4 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_219 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_decap_4 FILLER_36_276 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_38 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_fill_1 FILLER_37_83 ();
 sg13g2_decap_8 FILLER_37_113 ();
 sg13g2_decap_8 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_218 ();
 sg13g2_decap_4 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_4 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_22 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_71 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_87 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_381 ();
 assign uio_oe[0] = net16;
 assign uio_oe[1] = net17;
 assign uio_oe[2] = net18;
 assign uio_oe[3] = net19;
 assign uio_oe[4] = net20;
 assign uio_oe[5] = net21;
 assign uio_oe[6] = net22;
 assign uio_oe[7] = net23;
 assign uio_out[0] = net24;
 assign uio_out[1] = net25;
 assign uio_out[2] = net26;
 assign uio_out[3] = net27;
 assign uio_out[4] = net28;
 assign uio_out[5] = net29;
 assign uio_out[6] = net30;
 assign uio_out[7] = net31;
endmodule
